library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    234, 234, 239, 238, 237, 225, 247, 258, 240, 209, 183, 193, 199, 202, 201, 
    236, 241, 247, 244, 249, 228, 206, 211, 169, 130, 76, 82, 128, 190, 202, 
    164, 236, 247, 248, 255, 246, 143, 100, 86, 124, 74, 72, 51, 114, 191, 
    33, 157, 235, 251, 204, 182, 120, 68, 69, 156, 82, 88, 54, 40, 179, 
    41, 137, 193, 260, 170, 123, 88, 55, 50, 137, 105, 52, 75, 36, 91, 
    48, 135, 181, 178, 199, 139, 106, 78, 25, 196, 93, 51, 92, 58, 34, 
    48, 84, 170, 172, 182, 171, 152, 95, 47, 191, 73, 47, 69, 86, 67, 
    65, 87, 74, 148, 168, 210, 90, 109, 79, 187, 99, 48, 86, 103, 132, 
    72, 110, 11, 130, 106, 124, 98, 86, 119, 116, 128, 51, 79, 138, 195, 
    127, 117, 24, 107, 70, 85, 126, 94, 69, 121, 52, 40, 92, 196, 201, 
    151, 117, 34, 188, 50, 49, 120, 101, 30, 18, 4, 3, 12, 63, 48, 
    74, 117, 91, 219, 63, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 139, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 102, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    47, 65, 51, 50, 40, 60, 57, 51, 43, 53, 67, 69, 64, 54, 45, 
    39, 64, 51, 53, 43, 50, 49, 73, 83, 44, 35, 43, 55, 55, 48, 
    82, 62, 48, 52, 41, 88, 78, 51, 35, 35, 68, 52, 43, 35, 61, 
    68, 0, 49, 45, 60, 32, 58, 43, 40, 46, 88, 67, 66, 40, 38, 
    65, 27, 50, 3, 84, 48, 106, 74, 65, 1, 64, 62, 46, 46, 17, 
    62, 86, 75, 56, 156, 118, 112, 63, 62, 0, 98, 83, 50, 45, 30, 
    53, 107, 78, 93, 64, 57, 123, 74, 88, 22, 100, 60, 33, 38, 48, 
    73, 110, 15, 67, 11, 101, 120, 90, 86, 42, 89, 71, 47, 70, 53, 
    93, 96, 76, 70, 42, 85, 76, 56, 32, 40, 93, 95, 51, 44, 35, 
    108, 84, 109, 32, 100, 44, 37, 78, 41, 106, 86, 47, 34, 39, 55, 
    92, 88, 110, 11, 64, 32, 66, 136, 102, 38, 12, 9, 10, 18, 21, 
    65, 97, 80, 43, 170, 103, 68, 69, 52, 28, 25, 27, 28, 22, 35, 
    9, 48, 41, 136, 120, 39, 42, 35, 24, 16, 12, 17, 34, 33, 14, 
    26, 22, 32, 177, 49, 27, 30, 35, 35, 31, 24, 36, 24, 12, 59, 
    36, 32, 27, 78, 27, 35, 45, 37, 25, 23, 29, 16, 0, 29, 36, 
    
    -- channel=2
    132, 151, 150, 146, 139, 154, 149, 142, 135, 114, 106, 120, 140, 133, 117, 
    134, 163, 156, 147, 153, 241, 155, 139, 103, 132, 140, 112, 96, 104, 120, 
    95, 99, 145, 146, 141, 142, 110, 80, 101, 198, 166, 149, 111, 61, 127, 
    112, 140, 138, 151, 152, 152, 185, 126, 110, 156, 171, 124, 97, 52, 104, 
    182, 234, 152, 197, 335, 292, 210, 142, 88, 168, 212, 146, 129, 91, 69, 
    178, 224, 167, 161, 213, 237, 255, 167, 113, 246, 212, 116, 124, 120, 108, 
    206, 219, 116, 137, 180, 258, 237, 204, 124, 251, 181, 131, 123, 147, 123, 
    247, 259, 147, 154, 167, 267, 193, 146, 119, 216, 178, 116, 122, 137, 121, 
    273, 275, 159, 190, 164, 139, 138, 153, 145, 159, 106, 69, 90, 133, 157, 
    257, 261, 178, 227, 150, 148, 201, 245, 146, 107, 70, 59, 119, 171, 135, 
    250, 265, 176, 327, 341, 224, 251, 215, 138, 112, 95, 131, 129, 104, 85, 
    119, 228, 232, 381, 197, 68, 96, 95, 80, 90, 96, 109, 121, 121, 113, 
    92, 119, 245, 302, 86, 119, 112, 105, 95, 99, 114, 128, 122, 121, 155, 
    92, 103, 174, 177, 95, 123, 118, 106, 111, 119, 111, 98, 103, 132, 96, 
    110, 111, 109, 66, 60, 73, 84, 111, 140, 145, 110, 107, 175, 168, 81, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 67, 0, 0, 96, 40, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 89, 0, 0, 111, 29, 42, 0, 0, 89, 19, 0, 0, 0, 0, 
    0, 77, 0, 0, 17, 73, 78, 0, 0, 112, 0, 0, 0, 0, 0, 
    45, 60, 0, 0, 0, 136, 0, 0, 0, 69, 0, 0, 0, 0, 0, 
    82, 109, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 107, 0, 50, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 
    125, 97, 0, 167, 91, 10, 92, 55, 0, 0, 0, 0, 0, 0, 0, 
    49, 91, 34, 259, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 92, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 87, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 
    
    -- channel=4
    123, 115, 120, 123, 123, 114, 126, 126, 119, 111, 97, 96, 100, 106, 103, 
    120, 117, 120, 126, 122, 137, 130, 113, 85, 73, 84, 79, 76, 95, 108, 
    101, 97, 130, 124, 131, 112, 98, 59, 63, 84, 101, 75, 79, 72, 94, 
    85, 93, 135, 122, 122, 93, 107, 82, 77, 82, 104, 82, 64, 60, 67, 
    100, 131, 142, 98, 145, 132, 108, 82, 65, 64, 108, 94, 70, 60, 61, 
    122, 134, 145, 132, 93, 109, 128, 88, 75, 93, 141, 82, 69, 68, 59, 
    117, 140, 110, 106, 79, 129, 139, 119, 78, 105, 121, 87, 72, 79, 89, 
    137, 115, 107, 111, 97, 138, 127, 95, 84, 111, 114, 84, 65, 94, 88, 
    146, 132, 128, 96, 132, 78, 89, 95, 82, 112, 91, 60, 54, 80, 118, 
    141, 140, 118, 86, 104, 84, 82, 121, 109, 84, 58, 28, 59, 114, 115, 
    126, 143, 115, 117, 171, 126, 129, 117, 90, 57, 48, 59, 71, 89, 92, 
    88, 118, 121, 185, 173, 74, 60, 56, 56, 58, 63, 61, 65, 72, 68, 
    82, 85, 114, 198, 77, 60, 59, 57, 58, 60, 60, 71, 74, 66, 75, 
    69, 64, 97, 136, 76, 63, 66, 58, 53, 59, 66, 67, 62, 74, 91, 
    76, 56, 76, 54, 64, 57, 59, 60, 65, 71, 70, 58, 75, 97, 63, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 2, 0, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 14, 0, 0, 41, 24, 44, 0, 0, 
    122, 0, 0, 0, 0, 0, 27, 35, 9, 0, 63, 7, 35, 16, 0, 
    147, 0, 20, 0, 51, 41, 72, 50, 18, 0, 43, 77, 1, 47, 0, 
    111, 0, 40, 0, 0, 34, 73, 59, 71, 0, 92, 82, 0, 34, 28, 
    112, 56, 0, 32, 0, 0, 50, 63, 90, 0, 112, 62, 0, 0, 34, 
    96, 76, 58, 34, 0, 0, 96, 10, 46, 0, 61, 65, 0, 0, 0, 
    106, 33, 135, 0, 27, 0, 36, 16, 0, 19, 0, 54, 0, 0, 0, 
    43, 31, 148, 0, 86, 2, 0, 63, 23, 5, 53, 7, 0, 0, 0, 
    0, 40, 137, 0, 179, 94, 0, 55, 113, 57, 25, 20, 13, 3, 41, 
    0, 0, 86, 0, 172, 97, 21, 22, 50, 30, 31, 29, 36, 38, 56, 
    69, 0, 0, 52, 179, 39, 43, 33, 38, 34, 35, 39, 46, 45, 43, 
    84, 38, 0, 114, 78, 31, 57, 39, 31, 35, 40, 40, 53, 25, 61, 
    90, 42, 23, 31, 45, 9, 25, 37, 31, 45, 61, 35, 11, 84, 112, 
    
    -- channel=6
    134, 134, 137, 136, 137, 139, 138, 139, 135, 123, 114, 119, 126, 124, 118, 
    133, 143, 141, 138, 143, 162, 138, 130, 109, 114, 108, 104, 108, 117, 122, 
    103, 131, 142, 139, 142, 136, 98, 98, 95, 129, 91, 88, 79, 96, 119, 
    77, 142, 139, 144, 131, 140, 119, 86, 82, 121, 90, 88, 66, 59, 119, 
    90, 149, 131, 171, 172, 161, 108, 79, 66, 132, 122, 85, 88, 63, 94, 
    99, 126, 124, 130, 125, 122, 115, 96, 67, 168, 109, 70, 91, 79, 78, 
    106, 108, 114, 104, 135, 150, 124, 112, 67, 168, 93, 80, 92, 98, 83, 
    119, 115, 113, 124, 137, 151, 97, 92, 76, 143, 93, 74, 89, 95, 90, 
    123, 136, 77, 114, 118, 106, 93, 96, 111, 130, 88, 52, 83, 102, 128, 
    122, 130, 70, 141, 83, 103, 131, 121, 103, 72, 57, 61, 98, 135, 124, 
    143, 137, 81, 184, 128, 116, 136, 100, 66, 81, 76, 82, 90, 112, 101, 
    97, 124, 114, 206, 85, 43, 70, 66, 50, 62, 58, 64, 63, 61, 53, 
    50, 93, 146, 145, 34, 59, 56, 56, 53, 55, 61, 64, 59, 61, 74, 
    38, 58, 128, 67, 51, 66, 58, 55, 56, 58, 57, 49, 50, 63, 45, 
    40, 47, 64, 54, 48, 49, 47, 55, 67, 68, 51, 55, 84, 66, 28, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 5, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 30, 5, 22, 0, 7, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 31, 15, 5, 0, 22, 3, 27, 0, 0, 
    89, 0, 0, 0, 6, 0, 10, 33, 0, 0, 29, 9, 23, 21, 0, 
    93, 0, 32, 0, 0, 19, 38, 33, 9, 0, 9, 60, 0, 30, 0, 
    89, 0, 42, 18, 0, 26, 19, 35, 39, 0, 56, 61, 0, 17, 18, 
    87, 0, 1, 44, 0, 0, 9, 26, 60, 0, 69, 41, 0, 0, 23, 
    65, 0, 42, 11, 0, 0, 58, 0, 30, 0, 32, 45, 0, 0, 0, 
    52, 0, 101, 0, 34, 0, 16, 0, 0, 0, 0, 43, 0, 0, 0, 
    0, 0, 89, 0, 67, 4, 0, 5, 19, 16, 35, 5, 0, 0, 6, 
    0, 0, 75, 0, 75, 62, 0, 6, 66, 19, 0, 0, 0, 0, 12, 
    0, 0, 34, 0, 113, 53, 0, 0, 14, 0, 0, 0, 0, 0, 4, 
    10, 0, 0, 0, 123, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 20, 37, 0, 7, 1, 0, 0, 0, 0, 0, 0, 8, 
    25, 0, 0, 0, 11, 0, 0, 0, 0, 0, 11, 0, 0, 9, 44, 
    
    -- channel=8
    293, 295, 297, 305, 299, 293, 309, 307, 294, 276, 246, 244, 255, 259, 242, 
    291, 298, 304, 313, 307, 386, 331, 291, 219, 209, 231, 197, 187, 233, 258, 
    250, 246, 309, 306, 306, 314, 249, 162, 155, 250, 286, 234, 201, 158, 236, 
    242, 216, 319, 310, 307, 257, 305, 210, 189, 239, 299, 211, 167, 119, 175, 
    339, 378, 348, 319, 510, 393, 338, 221, 155, 178, 342, 251, 193, 157, 111, 
    342, 414, 370, 247, 341, 358, 402, 274, 195, 268, 402, 233, 202, 194, 147, 
    349, 403, 299, 267, 248, 371, 456, 341, 245, 311, 363, 231, 185, 222, 226, 
    401, 413, 299, 312, 261, 445, 379, 273, 236, 296, 332, 226, 185, 239, 226, 
    453, 442, 318, 309, 294, 234, 260, 253, 255, 272, 240, 158, 119, 214, 287, 
    441, 436, 358, 282, 327, 210, 271, 385, 263, 239, 160, 80, 174, 291, 302, 
    406, 438, 352, 398, 547, 380, 381, 399, 292, 164, 134, 165, 198, 253, 245, 
    272, 386, 413, 560, 495, 210, 169, 164, 166, 159, 171, 172, 190, 202, 196, 
    204, 232, 369, 569, 265, 178, 171, 159, 156, 161, 178, 206, 216, 204, 241, 
    198, 175, 270, 439, 211, 187, 186, 164, 159, 177, 182, 190, 179, 214, 229, 
    209, 166, 178, 200, 149, 143, 170, 178, 194, 211, 191, 169, 238, 289, 186, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 136, 181, 156, 94, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 93, 134, 123, 71, 84, 118, 90, 0, 
    182, 106, 0, 0, 0, 0, 49, 94, 128, 100, 75, 75, 119, 114, 0, 
    261, 192, 0, 0, 99, 19, 45, 60, 107, 180, 114, 102, 135, 142, 109, 
    249, 212, 0, 0, 0, 33, 94, 80, 110, 202, 128, 130, 142, 160, 96, 
    249, 239, 76, 0, 0, 148, 126, 105, 75, 76, 105, 122, 165, 106, 0, 
    298, 311, 231, 133, 0, 57, 33, 100, 95, 0, 63, 85, 113, 0, 0, 
    249, 294, 241, 253, 159, 82, 91, 146, 139, 58, 98, 147, 105, 0, 0, 
    311, 240, 221, 318, 260, 270, 336, 313, 269, 207, 338, 412, 437, 334, 303, 
    612, 405, 257, 269, 331, 463, 488, 496, 537, 556, 613, 641, 678, 678, 683, 
    765, 580, 360, 298, 440, 593, 593, 578, 594, 636, 689, 713, 705, 717, 762, 
    811, 712, 571, 422, 525, 614, 607, 600, 624, 670, 725, 750, 749, 827, 793, 
    789, 774, 666, 544, 577, 629, 635, 614, 627, 666, 692, 700, 742, 806, 757, 
    
    -- channel=10
    242, 243, 248, 246, 248, 237, 252, 268, 262, 233, 210, 212, 216, 224, 231, 
    247, 253, 255, 251, 252, 193, 220, 235, 216, 149, 93, 110, 153, 203, 220, 
    201, 230, 254, 259, 264, 221, 183, 150, 129, 84, 53, 60, 73, 142, 190, 
    71, 130, 231, 259, 225, 191, 109, 93, 81, 114, 71, 102, 85, 94, 171, 
    30, 47, 188, 237, 75, 89, 69, 79, 79, 123, 68, 75, 80, 71, 135, 
    45, 34, 171, 241, 120, 118, 60, 74, 52, 116, 57, 77, 84, 71, 73, 
    42, 12, 159, 210, 143, 120, 67, 71, 56, 88, 51, 67, 78, 78, 73, 
    42, 0, 73, 134, 157, 95, 52, 90, 83, 114, 78, 67, 86, 87, 130, 
    14, 9, 30, 73, 125, 114, 97, 85, 86, 115, 130, 92, 104, 122, 188, 
    42, 23, 6, 45, 54, 107, 94, 33, 71, 126, 87, 92, 84, 168, 209, 
    33, 36, 10, 51, 0, 16, 41, 22, 23, 47, 28, 11, 3, 30, 45, 
    0, 12, 16, 37, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    168, 178, 169, 175, 174, 163, 181, 185, 174, 165, 149, 142, 143, 150, 146, 
    164, 171, 177, 183, 171, 173, 185, 173, 161, 87, 89, 86, 93, 124, 144, 
    164, 139, 173, 180, 176, 230, 162, 91, 47, 91, 137, 109, 115, 73, 126, 
    134, 43, 172, 177, 178, 112, 136, 95, 89, 104, 168, 117, 96, 60, 83, 
    155, 133, 193, 132, 203, 171, 184, 110, 96, 34, 151, 127, 83, 81, 52, 
    153, 181, 196, 164, 191, 190, 203, 137, 110, 36, 218, 134, 91, 94, 52, 
    131, 229, 146, 181, 142, 139, 249, 162, 145, 108, 198, 108, 76, 79, 100, 
    159, 203, 123, 147, 118, 201, 238, 169, 118, 142, 185, 122, 79, 120, 123, 
    204, 198, 152, 131, 121, 154, 134, 118, 88, 170, 119, 129, 54, 98, 147, 
    212, 201, 192, 107, 152, 96, 100, 172, 113, 150, 132, 40, 51, 141, 175, 
    162, 194, 198, 76, 229, 124, 159, 224, 155, 81, 11, 22, 57, 91, 85, 
    117, 165, 175, 226, 336, 114, 79, 73, 54, 44, 46, 47, 44, 58, 53, 
    56, 88, 104, 305, 162, 51, 57, 49, 42, 33, 36, 42, 71, 62, 44, 
    55, 41, 70, 283, 79, 53, 54, 47, 44, 45, 51, 58, 51, 27, 106, 
    69, 39, 55, 111, 53, 41, 62, 54, 51, 56, 57, 38, 34, 96, 66, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    77, 71, 70, 67, 66, 68, 70, 65, 58, 76, 89, 90, 73, 59, 51, 
    65, 58, 68, 67, 72, 82, 49, 70, 79, 84, 66, 66, 93, 92, 63, 
    83, 140, 70, 62, 71, 137, 75, 61, 65, 142, 114, 109, 70, 96, 95, 
    10, 117, 70, 70, 58, 86, 72, 78, 99, 182, 107, 108, 83, 60, 128, 
    77, 147, 69, 117, 108, 97, 97, 74, 88, 152, 102, 59, 93, 52, 90, 
    136, 208, 80, 80, 250, 163, 111, 76, 41, 213, 141, 89, 120, 84, 50, 
    123, 165, 125, 27, 170, 166, 179, 119, 64, 236, 120, 75, 102, 107, 84, 
    146, 153, 99, 68, 118, 235, 168, 158, 96, 195, 135, 77, 124, 135, 96, 
    170, 210, 93, 167, 88, 164, 99, 91, 136, 87, 127, 99, 110, 107, 79, 
    213, 212, 98, 175, 101, 124, 148, 101, 113, 145, 105, 72, 115, 116, 87, 
    250, 195, 111, 243, 102, 86, 224, 227, 135, 80, 78, 101, 142, 168, 134, 
    290, 272, 164, 284, 209, 172, 170, 164, 146, 146, 160, 166, 168, 173, 164, 
    175, 256, 266, 247, 144, 152, 148, 149, 145, 150, 164, 171, 188, 192, 191, 
    176, 172, 299, 243, 151, 165, 142, 143, 157, 165, 180, 192, 179, 198, 222, 
    171, 176, 182, 193, 150, 178, 188, 166, 161, 160, 155, 169, 191, 183, 147, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 6, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 23, 8, 24, 0, 6, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 51, 12, 0, 0, 8, 3, 26, 0, 0, 
    84, 0, 0, 0, 21, 0, 5, 20, 0, 0, 42, 0, 29, 14, 0, 
    84, 0, 26, 0, 0, 0, 34, 34, 13, 0, 0, 47, 0, 31, 0, 
    57, 0, 37, 4, 0, 10, 37, 26, 48, 0, 53, 62, 0, 16, 10, 
    52, 8, 0, 53, 0, 0, 6, 31, 57, 0, 68, 35, 0, 0, 11, 
    38, 13, 17, 16, 0, 0, 73, 1, 29, 0, 42, 40, 0, 0, 0, 
    43, 0, 92, 0, 17, 0, 12, 2, 0, 3, 0, 55, 0, 0, 0, 
    2, 0, 98, 0, 35, 0, 0, 4, 0, 14, 52, 0, 0, 0, 11, 
    0, 0, 82, 0, 94, 20, 0, 12, 72, 31, 0, 0, 0, 0, 15, 
    0, 0, 18, 0, 114, 60, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 72, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    
    -- channel=15
    205, 218, 219, 220, 213, 218, 218, 217, 211, 187, 164, 178, 193, 179, 171, 
    215, 220, 224, 221, 235, 365, 195, 196, 131, 207, 192, 135, 135, 183, 185, 
    144, 205, 224, 220, 223, 232, 164, 101, 137, 288, 222, 200, 132, 107, 208, 
    118, 246, 218, 235, 215, 230, 254, 152, 159, 255, 218, 160, 132, 74, 185, 
    236, 358, 197, 307, 454, 281, 229, 157, 110, 256, 283, 153, 180, 115, 71, 
    203, 379, 212, 160, 383, 277, 333, 201, 124, 413, 255, 135, 189, 157, 111, 
    230, 316, 202, 164, 277, 387, 362, 259, 154, 406, 235, 161, 171, 228, 161, 
    292, 355, 178, 226, 249, 434, 211, 209, 179, 328, 261, 146, 188, 193, 177, 
    347, 391, 169, 327, 193, 185, 207, 227, 249, 172, 213, 70, 123, 218, 227, 
    395, 382, 230, 323, 209, 143, 282, 340, 161, 176, 80, 79, 196, 259, 208, 
    452, 369, 222, 529, 444, 280, 356, 312, 184, 117, 149, 189, 193, 217, 188, 
    270, 385, 336, 586, 273, 145, 160, 155, 162, 165, 183, 188, 214, 214, 201, 
    185, 237, 411, 449, 124, 190, 170, 169, 171, 185, 210, 227, 216, 218, 277, 
    192, 186, 302, 332, 189, 201, 186, 168, 180, 197, 196, 204, 197, 263, 186, 
    186, 197, 183, 182, 137, 167, 183, 191, 220, 230, 186, 196, 309, 271, 154, 
    
    -- channel=16
    216, 226, 225, 224, 214, 228, 229, 212, 203, 199, 187, 192, 201, 188, 160, 
    205, 220, 229, 228, 234, 345, 251, 217, 177, 209, 232, 179, 158, 180, 177, 
    180, 194, 221, 219, 221, 282, 223, 136, 152, 317, 339, 278, 202, 131, 195, 
    195, 199, 235, 228, 229, 232, 305, 224, 209, 319, 336, 248, 190, 106, 165, 
    387, 420, 281, 320, 544, 453, 387, 247, 166, 265, 393, 264, 214, 150, 95, 
    438, 507, 324, 248, 490, 479, 468, 299, 179, 391, 464, 261, 237, 215, 149, 
    458, 485, 287, 191, 303, 467, 533, 392, 253, 438, 425, 257, 219, 270, 234, 
    531, 520, 324, 265, 291, 559, 441, 339, 255, 383, 402, 249, 237, 278, 223, 
    594, 591, 377, 389, 306, 315, 299, 281, 293, 267, 276, 169, 150, 230, 250, 
    582, 585, 420, 407, 370, 250, 351, 443, 297, 273, 165, 95, 192, 268, 241, 
    552, 570, 417, 578, 648, 433, 510, 524, 349, 185, 170, 228, 273, 299, 272, 
    425, 555, 524, 742, 621, 328, 291, 286, 269, 253, 276, 293, 321, 336, 326, 
    326, 381, 553, 710, 359, 296, 284, 268, 260, 271, 304, 337, 352, 351, 394, 
    337, 306, 463, 549, 307, 309, 298, 275, 283, 307, 320, 334, 322, 373, 376, 
    348, 318, 320, 301, 236, 260, 292, 296, 324, 344, 316, 304, 406, 442, 305, 
    
    -- channel=17
    186, 201, 194, 205, 197, 191, 201, 204, 203, 194, 170, 158, 167, 169, 165, 
    189, 196, 199, 211, 200, 262, 221, 208, 160, 122, 141, 106, 93, 139, 171, 
    196, 137, 199, 204, 197, 202, 182, 85, 81, 127, 193, 153, 139, 68, 141, 
    195, 67, 195, 203, 222, 146, 208, 144, 121, 107, 221, 132, 119, 77, 63, 
    253, 207, 228, 173, 362, 245, 237, 160, 108, 39, 214, 182, 119, 120, 29, 
    223, 253, 248, 163, 198, 232, 293, 185, 153, 87, 290, 173, 115, 134, 88, 
    219, 279, 169, 218, 127, 219, 324, 234, 194, 126, 260, 157, 96, 126, 147, 
    261, 279, 170, 203, 136, 285, 289, 178, 167, 145, 238, 155, 99, 143, 139, 
    311, 272, 235, 181, 187, 118, 157, 170, 133, 150, 146, 129, 47, 112, 178, 
    297, 269, 283, 119, 231, 126, 137, 263, 150, 186, 134, 42, 80, 170, 207, 
    229, 269, 261, 174, 415, 258, 246, 290, 236, 105, 62, 93, 105, 128, 137, 
    114, 225, 270, 311, 384, 135, 68, 67, 93, 85, 92, 87, 95, 102, 111, 
    113, 85, 172, 393, 217, 99, 96, 83, 82, 82, 89, 108, 125, 115, 125, 
    119, 83, 82, 352, 148, 96, 106, 87, 85, 94, 95, 102, 94, 110, 141, 
    131, 87, 77, 100, 80, 68, 99, 104, 107, 114, 107, 79, 112, 180, 123, 
    
    -- channel=18
    84, 67, 76, 80, 82, 67, 75, 75, 78, 83, 76, 72, 70, 82, 88, 
    85, 64, 78, 77, 79, 65, 76, 60, 55, 68, 89, 88, 82, 82, 88, 
    78, 76, 75, 73, 83, 71, 48, 70, 94, 102, 104, 105, 115, 111, 79, 
    95, 127, 78, 73, 63, 66, 85, 111, 116, 111, 74, 96, 92, 121, 103, 
    80, 129, 81, 75, 57, 75, 57, 86, 109, 96, 79, 95, 111, 118, 125, 
    75, 86, 63, 57, 21, 22, 48, 92, 111, 119, 69, 76, 113, 111, 115, 
    66, 81, 62, 56, 97, 56, 63, 68, 96, 114, 57, 91, 108, 105, 120, 
    50, 56, 107, 68, 114, 88, 65, 76, 87, 113, 64, 88, 109, 107, 101, 
    49, 61, 75, 78, 82, 62, 67, 93, 109, 80, 80, 83, 106, 103, 102, 
    50, 72, 66, 87, 81, 97, 74, 81, 116, 82, 93, 107, 131, 108, 85, 
    63, 56, 63, 99, 69, 120, 105, 61, 86, 100, 126, 134, 133, 103, 90, 
    131, 59, 76, 96, 36, 53, 86, 86, 111, 132, 142, 139, 138, 147, 140, 
    168, 128, 67, 57, 56, 129, 134, 136, 145, 151, 153, 154, 151, 140, 147, 
    157, 145, 125, 53, 118, 141, 137, 139, 138, 143, 151, 148, 144, 158, 153, 
    153, 147, 136, 117, 145, 145, 144, 139, 143, 143, 151, 152, 153, 158, 154, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 21, 70, 51, 3, 0, 0, 
    29, 0, 0, 0, 0, 3, 50, 51, 26, 25, 114, 93, 109, 0, 0, 
    174, 0, 0, 0, 0, 0, 75, 85, 74, 0, 132, 76, 108, 67, 0, 
    184, 20, 0, 0, 95, 87, 148, 115, 103, 0, 98, 128, 71, 110, 0, 
    148, 67, 19, 0, 30, 82, 142, 116, 150, 0, 154, 138, 58, 101, 79, 
    130, 165, 0, 58, 0, 0, 133, 113, 166, 0, 168, 118, 61, 55, 80, 
    130, 179, 64, 54, 0, 26, 181, 91, 100, 0, 123, 131, 49, 61, 23, 
    170, 128, 178, 40, 50, 68, 85, 87, 14, 82, 42, 136, 36, 0, 0, 
    126, 115, 223, 47, 135, 51, 26, 144, 72, 76, 139, 79, 11, 0, 0, 
    59, 112, 218, 0, 223, 130, 75, 169, 182, 137, 93, 99, 101, 76, 96, 
    85, 90, 136, 14, 295, 186, 143, 143, 148, 139, 143, 153, 158, 159, 174, 
    183, 72, 0, 178, 268, 155, 165, 151, 151, 147, 153, 157, 172, 172, 159, 
    209, 159, 0, 269, 167, 148, 169, 157, 155, 161, 171, 172, 182, 151, 214, 
    222, 180, 144, 173, 153, 130, 147, 153, 150, 167, 184, 156, 127, 224, 234, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 66, 0, 0, 0, 8, 0, 
    0, 73, 0, 0, 0, 0, 0, 0, 5, 89, 0, 0, 0, 0, 24, 
    0, 44, 0, 0, 0, 0, 0, 0, 0, 106, 0, 0, 5, 0, 52, 
    0, 0, 0, 0, 19, 0, 0, 0, 0, 218, 0, 0, 21, 0, 0, 
    0, 0, 0, 0, 54, 23, 0, 0, 0, 182, 0, 0, 21, 24, 0, 
    0, 0, 0, 0, 32, 69, 0, 0, 0, 97, 0, 0, 42, 9, 0, 
    0, 5, 0, 10, 0, 0, 0, 0, 14, 0, 5, 0, 40, 0, 0, 
    0, 3, 0, 88, 0, 17, 16, 0, 17, 0, 0, 13, 53, 0, 0, 
    68, 0, 0, 185, 0, 6, 109, 0, 0, 0, 65, 97, 101, 64, 27, 
    170, 51, 0, 133, 0, 0, 69, 66, 55, 95, 107, 116, 116, 116, 101, 
    114, 172, 98, 0, 0, 90, 90, 94, 96, 114, 126, 131, 116, 119, 130, 
    97, 127, 249, 0, 29, 106, 80, 99, 110, 119, 128, 124, 111, 173, 114, 
    88, 131, 132, 42, 83, 125, 104, 91, 113, 107, 100, 120, 161, 106, 52, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 17, 14, 16, 6, 11, 
    19, 0, 0, 0, 0, 14, 13, 14, 18, 21, 19, 14, 3, 7, 11, 
    21, 18, 0, 0, 10, 7, 17, 14, 16, 14, 13, 7, 19, 14, 0, 
    19, 21, 7, 0, 15, 9, 5, 14, 13, 13, 14, 17, 9, 0, 28, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 0, 0, 10, 10, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 11, 2, 0, 0, 0, 12, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 12, 14, 7, 0, 0, 5, 0, 0, 5, 0, 
    4, 11, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 12, 5, 0, 5, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 
    10, 6, 8, 0, 0, 0, 15, 27, 16, 0, 0, 0, 0, 0, 0, 
    33, 25, 17, 4, 43, 18, 8, 9, 9, 7, 11, 11, 11, 13, 14, 
    20, 23, 9, 21, 14, 8, 12, 9, 8, 7, 9, 8, 20, 20, 8, 
    22, 15, 20, 36, 12, 9, 8, 9, 12, 11, 16, 21, 18, 9, 40, 
    22, 17, 21, 20, 12, 15, 22, 14, 11, 7, 15, 13, 7, 16, 25, 
    
    -- channel=23
    295, 309, 307, 309, 306, 294, 317, 338, 315, 267, 241, 249, 262, 276, 277, 
    304, 320, 315, 318, 306, 279, 273, 285, 234, 143, 93, 106, 156, 230, 269, 
    241, 257, 319, 326, 321, 262, 210, 129, 103, 77, 70, 69, 84, 127, 233, 
    107, 135, 290, 314, 284, 194, 140, 94, 82, 84, 114, 99, 86, 91, 168, 
    49, 87, 250, 215, 160, 119, 111, 97, 86, 71, 88, 94, 83, 82, 111, 
    25, 80, 246, 255, 132, 126, 128, 92, 87, 71, 100, 88, 76, 71, 72, 
    21, 72, 184, 274, 146, 131, 116, 105, 86, 64, 81, 74, 66, 66, 93, 
    39, 43, 63, 176, 136, 116, 106, 98, 111, 119, 107, 76, 66, 103, 170, 
    32, 19, 49, 87, 131, 95, 105, 97, 81, 132, 120, 103, 88, 146, 235, 
    69, 35, 52, 16, 67, 97, 77, 78, 72, 135, 97, 56, 84, 209, 252, 
    35, 47, 48, 18, 45, 18, 37, 41, 42, 25, 0, 0, 0, 0, 0, 
    0, 0, 31, 54, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    159, 158, 156, 162, 163, 151, 165, 169, 168, 162, 146, 135, 134, 141, 139, 
    158, 151, 157, 169, 155, 159, 187, 167, 152, 105, 117, 118, 115, 120, 138, 
    176, 118, 163, 167, 169, 209, 188, 128, 74, 83, 154, 113, 126, 94, 110, 
    165, 61, 168, 161, 183, 119, 147, 113, 106, 91, 184, 134, 120, 91, 64, 
    176, 129, 194, 101, 168, 164, 199, 140, 118, 39, 166, 151, 96, 93, 72, 
    214, 194, 206, 194, 190, 194, 213, 148, 135, 20, 244, 167, 98, 104, 72, 
    191, 246, 170, 174, 112, 154, 239, 183, 158, 83, 233, 149, 103, 99, 121, 
    217, 208, 160, 160, 100, 169, 251, 178, 141, 123, 207, 165, 90, 131, 123, 
    246, 212, 225, 127, 178, 165, 168, 149, 94, 192, 156, 150, 78, 91, 132, 
    239, 222, 236, 112, 184, 114, 106, 175, 161, 151, 137, 53, 44, 123, 174, 
    175, 223, 243, 75, 240, 151, 145, 215, 172, 109, 56, 48, 87, 134, 145, 
    148, 177, 185, 207, 394, 208, 147, 140, 115, 90, 90, 94, 95, 112, 114, 
    126, 130, 131, 335, 244, 95, 96, 92, 92, 85, 86, 95, 115, 108, 99, 
    124, 96, 109, 306, 136, 96, 106, 92, 84, 90, 108, 114, 108, 94, 163, 
    133, 91, 117, 156, 117, 94, 101, 90, 86, 104, 115, 90, 77, 154, 126, 
    
    -- channel=25
    132, 159, 154, 146, 135, 161, 157, 148, 135, 119, 116, 132, 145, 133, 112, 
    137, 172, 164, 149, 156, 222, 146, 152, 113, 118, 103, 82, 88, 118, 118, 
    97, 127, 146, 150, 139, 131, 90, 55, 86, 158, 112, 100, 61, 60, 137, 
    58, 122, 137, 158, 140, 136, 150, 85, 65, 149, 108, 92, 51, 28, 124, 
    117, 196, 124, 215, 310, 229, 155, 91, 44, 149, 161, 93, 87, 52, 53, 
    93, 180, 139, 114, 225, 211, 194, 117, 48, 241, 133, 63, 94, 73, 70, 
    123, 142, 125, 118, 173, 223, 201, 136, 79, 220, 109, 73, 73, 108, 77, 
    168, 182, 101, 127, 152, 264, 99, 101, 84, 171, 118, 56, 97, 100, 91, 
    179, 205, 65, 174, 102, 104, 99, 98, 129, 76, 106, 21, 59, 117, 148, 
    179, 182, 93, 170, 129, 98, 161, 181, 83, 100, 27, 45, 120, 159, 124, 
    207, 189, 86, 285, 222, 166, 208, 165, 94, 40, 47, 79, 65, 50, 30, 
    68, 171, 176, 301, 82, 0, 20, 20, 15, 15, 15, 19, 26, 19, 16, 
    0, 57, 196, 196, 0, 37, 32, 22, 7, 9, 17, 28, 26, 26, 46, 
    0, 11, 131, 76, 12, 32, 21, 25, 31, 28, 4, 1, 0, 27, 0, 
    0, 12, 12, 0, 0, 0, 10, 27, 50, 38, 6, 6, 72, 30, 0, 
    
    -- channel=26
    14, 15, 18, 7, 9, 20, 17, 12, 10, 13, 12, 26, 15, 4, 0, 
    17, 21, 26, 6, 25, 28, 0, 13, 4, 32, 0, 0, 34, 35, 1, 
    0, 71, 14, 8, 23, 66, 0, 0, 16, 86, 0, 0, 0, 41, 42, 
    0, 117, 9, 30, 0, 35, 0, 0, 0, 131, 0, 4, 0, 0, 119, 
    0, 71, 0, 121, 0, 0, 0, 0, 0, 143, 0, 0, 0, 0, 57, 
    0, 30, 0, 16, 146, 0, 0, 0, 0, 258, 0, 0, 28, 0, 0, 
    0, 0, 6, 0, 146, 76, 0, 0, 0, 231, 0, 0, 10, 24, 0, 
    0, 0, 0, 0, 91, 132, 0, 0, 0, 147, 0, 0, 45, 9, 0, 
    0, 18, 0, 63, 0, 39, 0, 0, 47, 0, 49, 0, 34, 36, 28, 
    0, 9, 0, 113, 0, 0, 54, 0, 0, 0, 0, 7, 73, 72, 1, 
    114, 1, 0, 214, 0, 0, 82, 0, 0, 0, 4, 15, 30, 40, 0, 
    135, 58, 0, 179, 0, 0, 17, 10, 0, 0, 0, 2, 0, 0, 0, 
    0, 113, 110, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 200, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 11, 7, 0, 18, 1, 0, 1, 0, 0, 0, 39, 0, 0, 
    
    -- channel=27
    324, 349, 346, 348, 336, 339, 358, 365, 338, 295, 265, 276, 300, 298, 281, 
    329, 363, 359, 358, 355, 419, 341, 324, 256, 200, 175, 141, 163, 251, 287, 
    243, 290, 354, 359, 348, 328, 244, 133, 124, 216, 201, 176, 134, 111, 267, 
    174, 170, 337, 360, 326, 273, 270, 156, 128, 195, 244, 158, 120, 54, 188, 
    255, 288, 331, 356, 498, 356, 283, 168, 97, 158, 274, 186, 144, 108, 64, 
    206, 307, 351, 257, 320, 339, 357, 220, 129, 236, 304, 167, 148, 141, 97, 
    226, 283, 261, 315, 252, 334, 380, 280, 181, 260, 267, 152, 119, 161, 156, 
    280, 324, 183, 293, 244, 385, 295, 210, 188, 253, 263, 142, 130, 181, 211, 
    324, 325, 181, 255, 217, 194, 200, 184, 196, 218, 172, 114, 82, 197, 290, 
    342, 312, 239, 208, 222, 164, 238, 314, 148, 202, 123, 49, 141, 292, 311, 
    310, 323, 236, 320, 431, 245, 287, 305, 199, 94, 31, 63, 57, 99, 92, 
    74, 273, 312, 446, 307, 46, 17, 12, 8, 6, 3, 2, 10, 7, 6, 
    0, 45, 261, 402, 104, 25, 17, 6, 0, 0, 0, 9, 22, 19, 36, 
    0, 0, 93, 286, 58, 22, 18, 1, 6, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 4, 24, 38, 32, 0, 0, 50, 50, 0, 
    
    -- channel=28
    43, 53, 46, 53, 48, 54, 44, 32, 41, 62, 69, 59, 64, 50, 43, 
    45, 41, 43, 53, 50, 147, 87, 67, 69, 109, 165, 112, 64, 56, 57, 
    79, 44, 40, 43, 30, 65, 110, 74, 86, 164, 216, 201, 170, 54, 69, 
    208, 66, 58, 44, 84, 92, 187, 156, 154, 114, 232, 135, 155, 98, 37, 
    316, 231, 122, 76, 343, 236, 240, 176, 136, 82, 232, 196, 154, 161, 26, 
    259, 280, 153, 15, 170, 211, 294, 205, 192, 104, 284, 197, 147, 178, 139, 
    268, 306, 117, 99, 99, 194, 304, 250, 223, 154, 283, 187, 140, 165, 168, 
    291, 348, 192, 177, 100, 242, 292, 183, 183, 123, 245, 181, 134, 153, 117, 
    351, 331, 267, 215, 147, 132, 167, 177, 165, 144, 104, 149, 79, 106, 81, 
    318, 310, 333, 203, 242, 132, 178, 300, 156, 153, 167, 101, 127, 100, 96, 
    285, 299, 316, 228, 490, 300, 276, 333, 296, 194, 170, 211, 217, 222, 217, 
    235, 310, 334, 323, 392, 243, 196, 198, 231, 230, 251, 256, 279, 277, 285, 
    310, 204, 254, 381, 319, 257, 253, 241, 241, 250, 276, 291, 298, 298, 330, 
    329, 275, 172, 425, 270, 260, 272, 244, 250, 268, 280, 286, 296, 306, 321, 
    335, 290, 248, 250, 224, 217, 251, 266, 273, 294, 284, 269, 309, 376, 334, 
    
    -- channel=29
    175, 188, 182, 181, 169, 194, 181, 160, 153, 168, 165, 171, 174, 146, 121, 
    161, 180, 187, 183, 200, 344, 187, 177, 150, 220, 240, 171, 150, 166, 149, 
    146, 197, 178, 169, 178, 290, 163, 111, 160, 403, 364, 303, 205, 136, 194, 
    164, 247, 191, 190, 181, 237, 321, 232, 236, 407, 328, 263, 191, 94, 204, 
    380, 499, 218, 346, 602, 467, 376, 233, 177, 335, 412, 246, 247, 154, 104, 
    421, 564, 250, 206, 562, 462, 463, 300, 173, 544, 453, 231, 283, 237, 150, 
    431, 518, 247, 137, 388, 508, 576, 393, 246, 598, 400, 245, 248, 315, 238, 
    517, 561, 298, 257, 345, 676, 426, 353, 252, 481, 396, 232, 285, 314, 205, 
    603, 659, 326, 445, 286, 334, 285, 300, 337, 262, 298, 146, 182, 246, 234, 
    627, 642, 392, 502, 362, 256, 395, 492, 298, 283, 164, 119, 257, 293, 210, 
    675, 616, 398, 738, 654, 467, 625, 586, 352, 205, 223, 308, 346, 367, 311, 
    575, 656, 559, 905, 611, 321, 347, 338, 320, 338, 372, 395, 429, 439, 421, 
    421, 506, 645, 780, 326, 380, 369, 352, 347, 370, 416, 451, 463, 465, 520, 
    433, 407, 609, 602, 362, 407, 377, 360, 380, 411, 429, 446, 426, 509, 488, 
    440, 429, 408, 392, 312, 358, 392, 390, 429, 447, 409, 410, 550, 562, 379, 
    
    -- channel=30
    0, 4, 0, 2, 0, 0, 0, 3, 13, 24, 21, 0, 0, 13, 29, 
    0, 0, 0, 13, 0, 0, 78, 31, 89, 0, 36, 19, 0, 0, 10, 
    91, 0, 0, 8, 0, 3, 135, 65, 0, 0, 57, 27, 123, 0, 0, 
    343, 0, 0, 0, 64, 0, 54, 45, 8, 0, 166, 5, 103, 48, 0, 
    265, 0, 99, 0, 43, 0, 174, 115, 81, 0, 43, 166, 0, 126, 0, 
    116, 0, 127, 0, 0, 0, 168, 119, 226, 0, 187, 194, 0, 66, 40, 
    72, 147, 0, 213, 0, 0, 96, 106, 249, 0, 241, 121, 0, 0, 58, 
    38, 140, 20, 121, 0, 0, 262, 32, 118, 0, 130, 162, 0, 0, 12, 
    105, 0, 245, 0, 5, 0, 71, 31, 0, 109, 0, 201, 0, 0, 0, 
    10, 0, 340, 0, 141, 0, 0, 109, 0, 28, 200, 5, 0, 0, 37, 
    0, 0, 325, 0, 291, 46, 0, 79, 218, 120, 0, 0, 0, 0, 19, 
    0, 0, 64, 0, 426, 160, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 81, 387, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 345, 74, 0, 12, 0, 0, 0, 0, 0, 0, 0, 41, 
    74, 0, 0, 49, 16, 0, 0, 0, 0, 0, 7, 0, 0, 36, 146, 
    
    -- channel=31
    28, 22, 24, 22, 24, 19, 29, 30, 21, 22, 24, 26, 23, 28, 29, 
    27, 25, 26, 23, 21, 0, 14, 18, 22, 0, 0, 9, 26, 34, 28, 
    17, 47, 26, 24, 26, 8, 0, 10, 9, 0, 0, 0, 0, 37, 31, 
    0, 30, 29, 21, 5, 0, 0, 0, 0, 0, 0, 0, 0, 18, 51, 
    0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 11, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 19, 27, 19, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    187, 199, 195, 196, 195, 189, 204, 220, 206, 171, 152, 156, 167, 176, 178, 
    186, 211, 204, 203, 197, 144, 193, 187, 168, 85, 40, 63, 95, 133, 165, 
    148, 147, 204, 211, 204, 190, 150, 113, 59, 12, 23, 21, 27, 59, 125, 
    77, 17, 181, 205, 184, 134, 75, 41, 13, 18, 62, 49, 42, 19, 73, 
    36, 0, 165, 151, 75, 86, 88, 55, 31, 10, 54, 56, 24, 22, 44, 
    36, 0, 163, 179, 65, 112, 73, 65, 35, 0, 68, 67, 21, 25, 18, 
    39, 2, 111, 205, 65, 51, 61, 60, 52, 0, 66, 41, 16, 8, 27, 
    31, 24, 30, 115, 71, 21, 88, 56, 57, 28, 55, 51, 11, 33, 88, 
    21, 0, 32, 1, 79, 80, 72, 36, 12, 102, 61, 76, 29, 53, 120, 
    28, 1, 29, 0, 40, 57, 42, 26, 27, 70, 57, 23, 0, 93, 162, 
    0, 23, 42, 0, 0, 0, 0, 12, 7, 15, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 33, 0, 0, 0, 4, 0, 0, 0, 3, 0, 
    0, 12, 0, 0, 0, 31, 0, 0, 0, 37, 0, 0, 0, 0, 20, 
    0, 35, 0, 0, 1, 0, 8, 0, 0, 31, 0, 0, 0, 0, 33, 
    0, 51, 0, 0, 25, 0, 0, 0, 0, 16, 0, 0, 4, 0, 0, 
    0, 30, 0, 0, 62, 0, 1, 0, 0, 79, 0, 0, 7, 0, 0, 
    0, 41, 0, 0, 65, 17, 22, 0, 0, 96, 0, 0, 0, 7, 0, 
    0, 11, 0, 0, 14, 61, 0, 0, 0, 63, 0, 0, 7, 5, 0, 
    0, 10, 0, 39, 0, 0, 0, 12, 1, 3, 15, 0, 2, 13, 5, 
    0, 1, 0, 43, 0, 0, 0, 28, 0, 0, 0, 0, 30, 36, 0, 
    72, 0, 0, 61, 0, 0, 33, 2, 0, 0, 0, 5, 9, 6, 0, 
    43, 19, 0, 94, 0, 0, 0, 0, 0, 0, 1, 2, 2, 5, 0, 
    0, 28, 0, 46, 0, 0, 0, 0, 0, 1, 5, 3, 5, 0, 1, 
    0, 1, 25, 23, 0, 0, 0, 0, 1, 2, 1, 4, 0, 8, 5, 
    0, 5, 6, 17, 0, 5, 2, 0, 6, 3, 0, 0, 17, 4, 0, 
    
    -- channel=35
    395, 419, 419, 418, 411, 404, 436, 456, 421, 346, 299, 325, 353, 369, 364, 
    409, 449, 436, 429, 423, 445, 378, 382, 275, 206, 136, 152, 210, 304, 356, 
    288, 335, 434, 442, 433, 368, 245, 166, 137, 157, 91, 87, 83, 148, 321, 
    125, 231, 402, 437, 387, 285, 222, 97, 77, 138, 133, 111, 75, 65, 246, 
    48, 197, 330, 348, 330, 212, 166, 112, 75, 134, 166, 104, 113, 75, 123, 
    0, 145, 316, 296, 228, 174, 211, 138, 95, 203, 117, 69, 103, 74, 76, 
    1, 114, 239, 360, 243, 234, 191, 136, 96, 185, 86, 80, 81, 101, 103, 
    41, 118, 72, 267, 205, 232, 91, 111, 119, 218, 116, 77, 85, 121, 203, 
    51, 90, 0, 155, 155, 114, 141, 141, 129, 187, 162, 61, 92, 207, 331, 
    111, 81, 36, 94, 88, 97, 144, 169, 78, 134, 53, 43, 123, 313, 331, 
    126, 104, 41, 179, 100, 60, 75, 52, 0, 13, 0, 0, 0, 0, 0, 
    0, 23, 62, 212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 39, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    37, 37, 37, 37, 37, 34, 38, 42, 42, 41, 38, 38, 33, 39, 44, 
    37, 38, 37, 37, 34, 1, 32, 42, 35, 14, 2, 19, 30, 35, 42, 
    47, 28, 37, 38, 37, 12, 18, 23, 29, 0, 0, 0, 9, 34, 30, 
    16, 11, 34, 36, 36, 14, 2, 16, 7, 0, 0, 7, 9, 34, 26, 
    0, 0, 20, 12, 0, 0, 0, 9, 17, 0, 0, 5, 9, 22, 40, 
    0, 0, 11, 23, 0, 0, 0, 0, 13, 0, 0, 0, 5, 6, 19, 
    0, 0, 8, 42, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 6, 1, 0, 0, 0, 1, 0, 0, 0, 6, 0, 15, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 17, 18, 13, 8, 25, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 22, 13, 29, 13, 12, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 67, 40, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 8, 0, 0, 30, 63, 11, 8, 0, 0, 
    93, 61, 0, 0, 108, 26, 81, 16, 6, 0, 62, 12, 5, 0, 0, 
    88, 148, 0, 0, 154, 80, 106, 33, 13, 0, 111, 39, 21, 13, 0, 
    76, 161, 0, 0, 21, 38, 166, 64, 59, 62, 110, 21, 0, 16, 4, 
    103, 183, 3, 0, 0, 147, 138, 69, 38, 33, 82, 32, 16, 34, 0, 
    165, 188, 71, 79, 0, 48, 31, 20, 22, 0, 31, 27, 0, 0, 0, 
    178, 169, 138, 74, 95, 0, 28, 109, 13, 48, 32, 0, 0, 0, 0, 
    183, 151, 143, 102, 175, 76, 135, 213, 127, 17, 11, 33, 61, 75, 54, 
    202, 201, 155, 181, 262, 144, 115, 111, 109, 94, 114, 125, 140, 142, 146, 
    153, 149, 130, 251, 181, 120, 119, 107, 103, 108, 130, 145, 165, 163, 175, 
    181, 138, 134, 307, 120, 124, 118, 111, 119, 134, 147, 168, 156, 170, 212, 
    182, 160, 121, 182, 99, 115, 139, 128, 124, 140, 142, 134, 153, 212, 173, 
    
    -- channel=38
    315, 331, 324, 326, 316, 321, 341, 344, 314, 281, 256, 271, 280, 277, 258, 
    307, 339, 336, 335, 332, 372, 316, 306, 243, 200, 161, 161, 199, 250, 266, 
    252, 297, 334, 336, 335, 412, 243, 168, 118, 236, 223, 180, 129, 148, 264, 
    146, 198, 332, 337, 309, 261, 251, 140, 132, 263, 246, 190, 129, 60, 223, 
    203, 308, 315, 333, 415, 319, 300, 168, 124, 186, 289, 166, 154, 83, 105, 
    231, 372, 331, 270, 454, 355, 345, 218, 120, 281, 324, 175, 180, 132, 72, 
    228, 347, 295, 276, 315, 346, 422, 270, 180, 343, 287, 161, 146, 173, 156, 
    285, 363, 190, 277, 244, 448, 331, 269, 194, 342, 277, 174, 164, 222, 219, 
    343, 391, 182, 285, 218, 279, 242, 207, 213, 261, 255, 144, 129, 215, 277, 
    400, 384, 239, 272, 246, 170, 254, 308, 198, 233, 132, 54, 139, 294, 300, 
    399, 384, 265, 384, 324, 207, 307, 358, 184, 92, 41, 43, 90, 164, 133, 
    258, 355, 315, 530, 418, 151, 144, 135, 74, 58, 59, 69, 74, 86, 74, 
    36, 204, 330, 519, 173, 76, 69, 64, 51, 44, 54, 73, 93, 85, 100, 
    40, 46, 261, 390, 91, 86, 65, 60, 60, 67, 64, 77, 52, 72, 105, 
    54, 45, 67, 180, 48, 62, 79, 72, 80, 88, 63, 55, 108, 126, 20, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    40, 47, 50, 51, 51, 48, 50, 55, 59, 46, 31, 30, 37, 39, 38, 
    51, 55, 55, 54, 53, 83, 60, 57, 23, 12, 12, 3, 1, 17, 37, 
    39, 11, 51, 53, 53, 23, 19, 0, 0, 6, 0, 0, 0, 0, 15, 
    13, 11, 39, 59, 65, 30, 34, 6, 0, 0, 10, 0, 0, 0, 0, 
    12, 27, 41, 54, 92, 66, 20, 5, 0, 0, 19, 12, 0, 0, 0, 
    2, 4, 38, 46, 0, 15, 36, 11, 0, 18, 27, 0, 0, 0, 0, 
    7, 7, 0, 44, 7, 41, 27, 21, 0, 10, 3, 0, 0, 0, 0, 
    26, 7, 12, 29, 17, 32, 11, 0, 0, 5, 4, 0, 0, 0, 0, 
    27, 11, 7, 0, 33, 0, 0, 10, 0, 14, 0, 0, 0, 0, 32, 
    11, 6, 3, 0, 0, 14, 8, 28, 6, 0, 0, 0, 0, 39, 48, 
    0, 17, 0, 25, 69, 42, 30, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    286, 306, 310, 311, 301, 303, 316, 313, 302, 269, 229, 241, 263, 251, 233, 
    294, 316, 319, 318, 325, 476, 313, 299, 202, 221, 217, 153, 147, 220, 251, 
    226, 243, 315, 313, 314, 307, 219, 97, 128, 299, 264, 214, 154, 93, 246, 
    169, 231, 309, 329, 322, 274, 323, 181, 160, 257, 281, 180, 123, 47, 173, 
    300, 418, 310, 380, 624, 432, 323, 193, 104, 218, 345, 207, 180, 111, 52, 
    274, 438, 329, 259, 405, 372, 439, 245, 143, 407, 376, 166, 184, 164, 102, 
    296, 408, 244, 264, 295, 460, 484, 341, 191, 425, 314, 183, 156, 223, 180, 
    390, 434, 231, 297, 285, 545, 330, 248, 190, 361, 319, 160, 172, 214, 190, 
    463, 477, 244, 349, 274, 193, 219, 255, 247, 230, 216, 76, 79, 207, 296, 
    480, 461, 307, 325, 275, 188, 300, 424, 205, 221, 92, 29, 171, 325, 294, 
    489, 463, 290, 551, 612, 379, 459, 414, 246, 117, 97, 165, 179, 211, 188, 
    231, 424, 408, 718, 422, 100, 96, 90, 97, 108, 123, 127, 147, 154, 143, 
    123, 189, 424, 619, 130, 138, 121, 109, 102, 113, 137, 169, 172, 164, 218, 
    118, 116, 279, 415, 155, 146, 135, 109, 120, 138, 130, 131, 120, 191, 145, 
    133, 118, 121, 103, 65, 84, 117, 136, 173, 179, 127, 114, 245, 249, 87, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    25, 26, 0, 0, 0, 5, 8, 12, 0, 46, 83, 65, 9, 0, 1, 
    0, 0, 0, 2, 0, 0, 0, 39, 150, 0, 0, 0, 67, 46, 0, 
    114, 130, 1, 1, 16, 227, 82, 78, 0, 0, 0, 0, 0, 75, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 0, 64, 23, 1, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 59, 
    19, 0, 0, 146, 288, 97, 0, 0, 0, 0, 0, 35, 8, 0, 0, 
    0, 0, 80, 5, 104, 0, 28, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 46, 105, 131, 9, 46, 19, 5, 23, 51, 0, 
    0, 0, 0, 0, 0, 214, 29, 0, 0, 2, 164, 153, 85, 0, 0, 
    24, 0, 0, 0, 0, 18, 0, 0, 0, 171, 122, 35, 0, 0, 6, 
    10, 0, 0, 0, 0, 0, 0, 116, 0, 0, 0, 0, 0, 11, 11, 
    241, 85, 0, 0, 266, 232, 162, 154, 45, 0, 0, 0, 0, 0, 0, 
    0, 185, 0, 69, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 189, 179, 11, 0, 0, 0, 0, 0, 0, 25, 0, 0, 105, 
    0, 0, 16, 184, 48, 72, 65, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    99, 107, 105, 110, 109, 105, 110, 119, 115, 93, 84, 78, 91, 106, 99, 
    104, 115, 108, 115, 100, 80, 149, 110, 86, 31, 52, 58, 45, 56, 89, 
    90, 28, 108, 116, 101, 41, 107, 66, 40, 0, 46, 42, 62, 28, 43, 
    123, 0, 102, 107, 115, 58, 61, 65, 25, 0, 85, 37, 45, 51, 0, 
    121, 0, 145, 53, 81, 126, 104, 81, 35, 0, 61, 106, 19, 59, 30, 
    119, 0, 163, 105, 0, 101, 91, 83, 76, 0, 113, 102, 0, 46, 65, 
    139, 29, 81, 132, 0, 16, 37, 90, 83, 0, 110, 78, 17, 2, 62, 
    123, 41, 113, 78, 15, 0, 120, 33, 61, 0, 70, 76, 0, 16, 73, 
    99, 5, 147, 0, 97, 21, 58, 28, 7, 72, 0, 78, 0, 15, 73, 
    24, 15, 118, 0, 82, 77, 21, 38, 73, 34, 62, 15, 0, 35, 102, 
    0, 37, 103, 0, 144, 84, 0, 17, 87, 49, 0, 0, 0, 0, 0, 
    0, 0, 63, 0, 90, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 7, 35, 0, 0, 0, 12, 0, 0, 0, 5, 0, 
    0, 34, 0, 0, 3, 18, 0, 0, 0, 89, 0, 0, 0, 10, 22, 
    0, 121, 0, 6, 0, 18, 0, 0, 0, 113, 0, 0, 0, 0, 89, 
    0, 83, 0, 99, 0, 0, 0, 0, 0, 141, 0, 0, 0, 0, 38, 
    0, 30, 0, 0, 96, 0, 0, 0, 0, 268, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 121, 75, 0, 0, 0, 228, 0, 0, 7, 22, 0, 
    0, 0, 0, 0, 83, 113, 0, 0, 0, 147, 0, 0, 35, 2, 0, 
    0, 9, 0, 53, 0, 3, 0, 0, 43, 0, 8, 0, 23, 39, 23, 
    0, 11, 0, 108, 0, 0, 52, 0, 0, 0, 0, 0, 68, 59, 0, 
    96, 0, 0, 239, 0, 0, 83, 0, 0, 0, 0, 25, 34, 12, 0, 
    95, 47, 0, 193, 0, 0, 0, 0, 0, 0, 4, 10, 9, 13, 0, 
    0, 91, 115, 0, 0, 0, 0, 0, 0, 8, 19, 17, 4, 6, 25, 
    0, 8, 180, 0, 0, 12, 0, 0, 9, 10, 6, 3, 0, 42, 0, 
    0, 9, 17, 0, 0, 18, 4, 0, 20, 6, 0, 11, 72, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    15, 15, 16, 12, 8, 22, 11, 3, 0, 7, 16, 27, 25, 8, 0, 
    14, 13, 14, 7, 21, 82, 1, 7, 0, 70, 63, 46, 49, 40, 10, 
    0, 61, 13, 7, 7, 42, 11, 29, 54, 138, 81, 89, 30, 48, 52, 
    0, 124, 18, 19, 4, 67, 64, 42, 58, 140, 61, 56, 42, 20, 90, 
    72, 158, 11, 109, 145, 88, 66, 43, 35, 159, 106, 29, 73, 28, 41, 
    85, 179, 26, 0, 195, 115, 100, 64, 16, 237, 74, 39, 90, 58, 43, 
    108, 109, 77, 0, 122, 161, 124, 86, 32, 222, 72, 51, 80, 101, 54, 
    125, 150, 78, 49, 87, 187, 64, 85, 60, 152, 83, 43, 96, 80, 56, 
    143, 190, 43, 155, 42, 94, 76, 70, 130, 34, 79, 15, 70, 91, 42, 
    168, 178, 61, 183, 74, 67, 149, 111, 68, 56, 17, 46, 106, 75, 22, 
    231, 167, 68, 303, 133, 102, 167, 144, 73, 53, 94, 109, 123, 132, 96, 
    214, 224, 154, 269, 64, 102, 128, 127, 119, 118, 133, 141, 155, 152, 142, 
    140, 192, 261, 159, 66, 135, 123, 125, 123, 134, 155, 163, 153, 161, 199, 
    148, 152, 244, 130, 108, 147, 127, 125, 134, 146, 148, 157, 152, 193, 138, 
    136, 158, 142, 144, 102, 135, 138, 139, 148, 155, 132, 154, 211, 167, 119, 
    
    -- channel=49
    255, 266, 273, 278, 275, 255, 279, 294, 278, 223, 182, 195, 228, 244, 248, 
    278, 283, 284, 282, 284, 317, 256, 227, 155, 149, 134, 104, 110, 196, 241, 
    153, 195, 280, 287, 280, 171, 156, 94, 116, 133, 105, 118, 111, 94, 210, 
    140, 173, 264, 284, 244, 198, 187, 118, 99, 89, 126, 84, 88, 83, 151, 
    148, 187, 243, 258, 295, 182, 121, 106, 67, 114, 155, 125, 115, 120, 73, 
    39, 119, 234, 140, 58, 111, 182, 145, 118, 151, 102, 81, 97, 111, 116, 
    74, 89, 149, 239, 126, 171, 140, 137, 118, 112, 98, 97, 88, 118, 126, 
    78, 126, 110, 203, 174, 143, 66, 68, 118, 125, 117, 81, 83, 90, 175, 
    83, 82, 55, 137, 116, 43, 112, 123, 137, 117, 76, 44, 59, 173, 244, 
    94, 83, 95, 83, 96, 76, 128, 180, 63, 84, 54, 64, 128, 221, 226, 
    80, 87, 73, 158, 247, 148, 77, 41, 62, 59, 55, 64, 20, 9, 14, 
    0, 24, 128, 156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 58, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 2, 11, 
    0, 0, 0, 0, 0, 0, 32, 0, 63, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 30, 80, 54, 0, 0, 28, 11, 43, 0, 0, 
    132, 0, 0, 0, 0, 0, 0, 28, 0, 0, 73, 24, 62, 28, 0, 
    125, 0, 51, 0, 0, 0, 80, 54, 43, 0, 0, 77, 0, 42, 0, 
    135, 0, 72, 28, 0, 60, 26, 53, 70, 0, 106, 130, 0, 26, 0, 
    110, 19, 14, 86, 0, 0, 26, 41, 114, 0, 141, 61, 0, 0, 24, 
    58, 29, 31, 8, 0, 0, 177, 49, 69, 0, 77, 95, 0, 0, 32, 
    62, 0, 150, 0, 8, 58, 54, 0, 0, 45, 0, 151, 0, 0, 0, 
    13, 0, 158, 0, 80, 5, 0, 0, 17, 52, 127, 16, 0, 0, 11, 
    0, 0, 167, 0, 29, 0, 0, 48, 113, 42, 0, 0, 0, 0, 0, 
    0, 0, 41, 0, 272, 166, 32, 34, 27, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 295, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 152, 61, 0, 2, 0, 0, 0, 0, 0, 3, 0, 49, 
    49, 0, 0, 62, 37, 0, 0, 0, 0, 0, 13, 0, 0, 0, 84, 
    
    -- channel=51
    269, 260, 270, 273, 275, 250, 277, 296, 283, 246, 222, 228, 235, 247, 259, 
    276, 269, 273, 276, 275, 218, 241, 240, 210, 162, 110, 129, 173, 228, 251, 
    208, 259, 282, 284, 288, 230, 200, 169, 140, 93, 71, 89, 95, 161, 218, 
    107, 164, 265, 279, 242, 209, 125, 107, 104, 105, 100, 105, 112, 116, 188, 
    59, 69, 226, 226, 86, 73, 81, 100, 103, 118, 85, 92, 107, 103, 142, 
    45, 60, 212, 204, 95, 94, 80, 99, 93, 91, 71, 103, 104, 97, 97, 
    47, 27, 187, 238, 129, 110, 72, 94, 88, 69, 75, 92, 99, 95, 106, 
    28, 31, 85, 179, 145, 70, 84, 102, 121, 111, 93, 96, 95, 105, 176, 
    10, 12, 48, 85, 130, 112, 121, 103, 112, 138, 128, 124, 120, 155, 207, 
    51, 25, 40, 39, 66, 110, 106, 56, 80, 132, 116, 107, 101, 189, 233, 
    39, 36, 45, 42, 0, 18, 12, 25, 44, 77, 53, 21, 8, 53, 68, 
    0, 19, 38, 14, 0, 31, 9, 11, 4, 3, 0, 0, 0, 0, 0, 
    0, 0, 41, 3, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    51, 60, 52, 63, 60, 48, 58, 74, 68, 49, 48, 34, 53, 65, 71, 
    53, 56, 48, 68, 44, 0, 97, 47, 86, 2, 21, 6, 0, 20, 53, 
    44, 3, 53, 75, 41, 0, 145, 79, 0, 0, 16, 36, 54, 0, 1, 
    184, 0, 52, 42, 60, 20, 14, 36, 0, 0, 115, 0, 84, 37, 0, 
    208, 0, 119, 0, 0, 0, 104, 83, 30, 0, 27, 106, 0, 77, 0, 
    121, 0, 165, 0, 0, 90, 108, 84, 102, 0, 109, 164, 0, 45, 42, 
    143, 0, 73, 162, 0, 0, 14, 95, 139, 0, 177, 87, 0, 0, 44, 
    82, 70, 50, 91, 0, 0, 173, 24, 113, 0, 110, 106, 0, 0, 83, 
    82, 0, 177, 0, 12, 18, 87, 0, 0, 38, 0, 153, 0, 0, 0, 
    18, 0, 210, 0, 84, 0, 0, 16, 0, 30, 130, 21, 0, 0, 64, 
    0, 0, 199, 0, 180, 0, 0, 14, 146, 63, 0, 0, 0, 0, 0, 
    0, 0, 84, 0, 176, 146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 298, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 130, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 83, 63, 40, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 12, 40, 0, 31, 0, 32, 0, 0, 
    145, 48, 0, 0, 20, 0, 19, 27, 35, 0, 24, 30, 30, 52, 0, 
    122, 101, 0, 0, 0, 0, 44, 11, 75, 0, 66, 34, 22, 57, 32, 
    109, 159, 0, 0, 0, 0, 61, 35, 73, 24, 80, 53, 29, 47, 20, 
    125, 180, 5, 0, 0, 34, 69, 4, 9, 0, 39, 44, 29, 0, 0, 
    190, 190, 144, 47, 0, 0, 0, 32, 0, 0, 0, 3, 0, 0, 0, 
    131, 153, 197, 100, 90, 0, 0, 122, 21, 0, 34, 31, 8, 0, 0, 
    171, 123, 169, 101, 285, 196, 189, 206, 195, 126, 192, 257, 267, 211, 197, 
    327, 225, 161, 126, 251, 260, 260, 268, 322, 340, 383, 397, 429, 422, 433, 
    506, 293, 139, 215, 287, 368, 369, 353, 363, 393, 435, 455, 451, 455, 497, 
    540, 454, 234, 347, 327, 375, 388, 368, 382, 418, 455, 470, 479, 526, 519, 
    529, 493, 404, 328, 343, 361, 380, 380, 392, 428, 441, 429, 463, 554, 521, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, 0, 1, 0, 
    3, 0, 0, 0, 0, 0, 14, 2, 0, 0, 0, 8, 8, 0, 0, 
    10, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 2, 17, 0, 
    0, 12, 4, 0, 0, 0, 0, 9, 5, 0, 3, 2, 0, 23, 0, 
    0, 0, 25, 0, 0, 17, 0, 10, 3, 0, 0, 11, 0, 0, 31, 
    44, 0, 37, 33, 0, 14, 0, 0, 0, 0, 21, 15, 0, 0, 14, 
    48, 0, 27, 0, 0, 0, 0, 10, 0, 0, 6, 9, 0, 0, 12, 
    49, 0, 49, 0, 0, 0, 24, 0, 0, 0, 0, 2, 0, 3, 9, 
    20, 0, 58, 0, 45, 0, 0, 0, 0, 0, 0, 12, 0, 0, 3, 
    0, 0, 7, 0, 5, 44, 0, 0, 43, 4, 4, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 11, 7, 0, 21, 0, 0, 0, 9, 0, 3, 
    0, 0, 0, 0, 4, 22, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    22, 9, 18, 0, 15, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    7, 11, 27, 0, 5, 0, 2, 0, 0, 0, 1, 0, 0, 0, 13, 
    12, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    36, 36, 37, 34, 37, 38, 29, 30, 37, 41, 50, 52, 50, 43, 50, 
    37, 34, 36, 31, 40, 26, 16, 32, 59, 78, 63, 57, 60, 57, 47, 
    32, 65, 32, 32, 32, 27, 40, 68, 83, 81, 41, 70, 64, 72, 60, 
    37, 78, 23, 37, 26, 70, 39, 68, 75, 79, 33, 58, 72, 78, 86, 
    41, 33, 11, 81, 10, 28, 16, 50, 68, 111, 30, 42, 74, 78, 86, 
    25, 15, 1, 37, 33, 28, 4, 45, 52, 104, 0, 46, 75, 77, 84, 
    32, 0, 24, 30, 73, 39, 0, 32, 42, 80, 10, 47, 76, 74, 54, 
    12, 15, 39, 29, 82, 23, 7, 42, 50, 60, 29, 41, 82, 53, 60, 
    1, 11, 11, 56, 27, 58, 41, 47, 73, 34, 40, 63, 89, 73, 43, 
    11, 13, 5, 74, 13, 70, 77, 23, 33, 52, 73, 106, 92, 48, 34, 
    34, 8, 5, 72, 0, 25, 47, 20, 42, 82, 98, 102, 91, 70, 68, 
    59, 43, 28, 8, 0, 48, 69, 70, 81, 94, 93, 93, 89, 83, 81, 
    77, 67, 66, 0, 31, 88, 87, 90, 93, 96, 97, 86, 79, 90, 85, 
    82, 89, 72, 0, 77, 89, 83, 87, 97, 92, 89, 84, 93, 88, 60, 
    74, 95, 81, 63, 87, 93, 92, 93, 92, 83, 79, 97, 97, 57, 79, 
    
    -- channel=59
    193, 207, 207, 204, 193, 209, 212, 206, 187, 160, 140, 159, 171, 159, 133, 
    189, 214, 214, 207, 217, 323, 199, 188, 106, 142, 121, 95, 111, 146, 148, 
    127, 180, 211, 206, 208, 240, 133, 64, 77, 228, 178, 141, 57, 68, 164, 
    40, 186, 205, 219, 193, 191, 196, 93, 83, 228, 179, 122, 55, 0, 143, 
    168, 308, 201, 298, 419, 315, 229, 113, 44, 209, 250, 108, 106, 17, 40, 
    220, 354, 230, 185, 395, 327, 303, 156, 36, 364, 270, 100, 127, 80, 35, 
    250, 282, 207, 128, 245, 372, 350, 234, 85, 370, 219, 109, 106, 150, 102, 
    322, 319, 171, 177, 201, 434, 245, 196, 120, 311, 224, 97, 126, 159, 133, 
    365, 394, 158, 265, 190, 188, 165, 157, 191, 154, 172, 31, 68, 157, 200, 
    387, 384, 183, 281, 189, 148, 253, 269, 165, 147, 21, 0, 109, 223, 185, 
    404, 382, 189, 499, 371, 236, 344, 313, 139, 41, 37, 73, 106, 148, 108, 
    241, 373, 309, 591, 302, 99, 107, 101, 66, 59, 70, 83, 101, 106, 92, 
    65, 208, 409, 475, 95, 90, 72, 66, 53, 61, 84, 112, 113, 111, 161, 
    62, 78, 322, 281, 84, 102, 78, 67, 73, 89, 85, 92, 74, 141, 97, 
    72, 77, 93, 94, 26, 61, 76, 85, 111, 120, 75, 79, 185, 161, 21, 
    
    -- channel=60
    392, 402, 402, 403, 393, 387, 416, 414, 383, 354, 324, 339, 346, 332, 311, 
    388, 395, 409, 413, 415, 521, 372, 374, 291, 280, 242, 201, 241, 328, 336, 
    316, 404, 415, 409, 416, 461, 314, 170, 165, 359, 320, 272, 194, 194, 352, 
    169, 319, 409, 415, 385, 339, 346, 213, 224, 370, 350, 254, 191, 107, 295, 
    309, 473, 395, 436, 602, 416, 369, 231, 176, 297, 382, 226, 231, 140, 130, 
    330, 567, 422, 331, 604, 462, 483, 276, 166, 478, 447, 234, 259, 206, 121, 
    329, 503, 384, 314, 409, 526, 578, 397, 230, 531, 391, 225, 220, 275, 234, 
    425, 498, 273, 357, 340, 648, 446, 368, 276, 479, 411, 221, 246, 315, 295, 
    511, 562, 284, 446, 316, 336, 308, 301, 331, 306, 327, 180, 180, 312, 373, 
    594, 561, 355, 399, 327, 245, 369, 440, 266, 332, 188, 79, 237, 404, 379, 
    621, 545, 360, 612, 566, 334, 518, 528, 307, 144, 107, 159, 212, 307, 265, 
    412, 573, 474, 808, 561, 247, 213, 200, 180, 170, 190, 194, 212, 223, 205, 
    194, 343, 553, 738, 242, 195, 176, 172, 162, 168, 191, 218, 242, 235, 273, 
    190, 182, 428, 593, 230, 208, 183, 162, 177, 194, 202, 221, 195, 248, 266, 
    197, 183, 208, 256, 154, 182, 216, 205, 218, 226, 185, 184, 289, 294, 147, 
    
    -- channel=61
    338, 348, 340, 351, 345, 333, 357, 368, 351, 325, 288, 279, 286, 294, 288, 
    333, 346, 350, 365, 349, 366, 355, 339, 285, 199, 180, 168, 192, 260, 292, 
    305, 294, 357, 363, 362, 399, 301, 188, 123, 169, 223, 170, 161, 151, 254, 
    226, 140, 354, 357, 348, 256, 262, 159, 143, 185, 266, 188, 152, 95, 170, 
    264, 252, 357, 298, 395, 278, 298, 181, 137, 94, 273, 202, 142, 117, 83, 
    263, 329, 370, 291, 360, 325, 347, 225, 159, 127, 349, 215, 156, 144, 82, 
    243, 345, 308, 328, 235, 292, 416, 279, 221, 198, 328, 186, 132, 156, 170, 
    290, 331, 212, 303, 216, 368, 354, 260, 218, 236, 307, 203, 135, 200, 213, 
    347, 335, 249, 243, 244, 242, 248, 215, 183, 265, 252, 178, 99, 187, 281, 
    374, 339, 304, 179, 277, 148, 193, 298, 190, 248, 171, 57, 101, 262, 332, 
    317, 342, 312, 211, 376, 228, 251, 337, 231, 107, 38, 35, 77, 181, 190, 
    179, 289, 308, 394, 501, 195, 117, 110, 87, 59, 53, 50, 53, 64, 65, 
    51, 129, 230, 499, 253, 58, 55, 46, 42, 32, 34, 48, 75, 68, 63, 
    53, 32, 130, 427, 127, 58, 59, 45, 38, 42, 46, 63, 45, 40, 110, 
    61, 22, 50, 159, 64, 45, 69, 56, 52, 62, 58, 31, 51, 114, 53, 
    
    -- channel=62
    52, 66, 56, 62, 52, 63, 67, 59, 45, 42, 38, 38, 47, 44, 26, 
    48, 65, 58, 68, 56, 120, 91, 62, 32, 19, 51, 31, 13, 25, 37, 
    48, 22, 61, 62, 52, 89, 63, 4, 0, 57, 117, 75, 50, 0, 36, 
    94, 0, 77, 55, 70, 33, 105, 44, 33, 44, 138, 56, 37, 0, 0, 
    168, 145, 116, 34, 248, 171, 173, 76, 28, 0, 149, 96, 36, 25, 0, 
    162, 200, 152, 36, 156, 173, 216, 108, 67, 12, 211, 94, 39, 45, 10, 
    165, 223, 100, 79, 48, 131, 238, 156, 109, 70, 195, 82, 29, 50, 68, 
    204, 236, 99, 113, 30, 189, 211, 110, 89, 76, 156, 87, 26, 77, 57, 
    251, 236, 163, 113, 91, 81, 99, 78, 60, 93, 64, 47, 0, 37, 60, 
    231, 225, 212, 93, 161, 39, 75, 191, 87, 73, 42, 0, 12, 65, 73, 
    185, 225, 209, 125, 318, 164, 154, 220, 145, 32, 0, 12, 28, 56, 51, 
    101, 190, 215, 256, 324, 104, 59, 55, 47, 28, 42, 47, 64, 72, 74, 
    76, 74, 139, 331, 160, 57, 56, 44, 36, 36, 48, 69, 84, 73, 94, 
    84, 57, 67, 286, 73, 58, 66, 49, 43, 55, 59, 69, 63, 69, 116, 
    100, 60, 57, 88, 30, 24, 47, 57, 62, 80, 73, 49, 79, 148, 90, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    156, 158, 158, 158, 159, 159, 159, 158, 160, 156, 154, 160, 159, 158, 159, 
    157, 159, 159, 158, 158, 158, 159, 159, 154, 118, 157, 163, 157, 158, 159, 
    159, 160, 161, 159, 159, 156, 160, 136, 123, 90, 140, 177, 159, 161, 160, 
    149, 148, 161, 163, 159, 135, 172, 122, 107, 82, 82, 149, 157, 159, 162, 
    95, 133, 185, 165, 160, 144, 163, 151, 146, 128, 120, 119, 118, 181, 166, 
    89, 105, 144, 147, 156, 135, 158, 164, 172, 126, 99, 93, 57, 145, 163, 
    66, 108, 126, 141, 101, 0, 31, 62, 131, 146, 139, 130, 145, 128, 158, 
    58, 73, 70, 151, 130, 82, 113, 96, 102, 73, 41, 49, 67, 79, 103, 
    123, 119, 104, 132, 141, 134, 146, 103, 97, 92, 97, 79, 92, 91, 78, 
    100, 63, 58, 51, 48, 48, 25, 20, 31, 2, 17, 5, 17, 39, 66, 
    0, 7, 0, 0, 12, 20, 0, 0, 0, 0, 0, 0, 12, 33, 80, 
    7, 63, 17, 0, 0, 2, 24, 0, 0, 0, 0, 25, 63, 73, 110, 
    0, 21, 33, 9, 4, 8, 149, 97, 89, 82, 78, 80, 86, 111, 137, 
    0, 9, 14, 5, 8, 10, 77, 98, 70, 68, 84, 108, 110, 125, 147, 
    15, 24, 21, 16, 15, 14, 40, 69, 71, 120, 118, 114, 124, 132, 147, 
    
    -- channel=65
    107, 106, 106, 106, 106, 107, 106, 110, 107, 105, 109, 105, 106, 106, 106, 
    107, 106, 106, 107, 106, 106, 106, 105, 106, 133, 106, 105, 107, 105, 106, 
    112, 111, 107, 105, 107, 112, 103, 117, 115, 117, 89, 101, 107, 105, 106, 
    93, 97, 100, 107, 112, 130, 95, 107, 61, 51, 31, 38, 95, 96, 99, 
    106, 102, 104, 110, 109, 108, 77, 104, 89, 110, 121, 118, 128, 89, 95, 
    44, 40, 83, 120, 129, 151, 156, 148, 116, 95, 50, 39, 52, 27, 89, 
    138, 121, 127, 78, 95, 56, 8, 0, 33, 121, 144, 153, 150, 136, 107, 
    38, 22, 53, 75, 88, 47, 19, 84, 111, 100, 64, 41, 21, 33, 38, 
    0, 93, 58, 78, 102, 118, 121, 128, 83, 100, 110, 119, 118, 107, 101, 
    87, 150, 139, 147, 138, 125, 118, 93, 101, 97, 93, 95, 72, 70, 71, 
    70, 75, 105, 119, 124, 131, 152, 150, 139, 132, 108, 87, 60, 60, 60, 
    48, 19, 65, 44, 37, 37, 4, 0, 8, 18, 20, 56, 98, 85, 41, 
    21, 21, 79, 73, 37, 29, 82, 277, 254, 236, 196, 131, 66, 36, 28, 
    49, 24, 33, 39, 27, 26, 78, 351, 314, 163, 55, 30, 41, 31, 37, 
    38, 0, 0, 1, 7, 2, 11, 116, 54, 22, 45, 34, 30, 26, 33, 
    
    -- channel=66
    342, 342, 342, 342, 342, 342, 343, 343, 344, 339, 342, 340, 341, 342, 343, 
    342, 342, 342, 342, 341, 341, 341, 341, 333, 281, 285, 332, 343, 342, 343, 
    337, 341, 345, 342, 346, 343, 335, 306, 243, 220, 245, 317, 341, 342, 344, 
    328, 336, 335, 345, 351, 319, 315, 309, 306, 304, 310, 329, 329, 333, 339, 
    131, 160, 293, 337, 342, 322, 344, 334, 348, 321, 257, 203, 179, 244, 328, 
    324, 358, 336, 266, 282, 182, 188, 216, 271, 305, 296, 320, 311, 337, 327, 
    112, 151, 203, 293, 288, 139, 151, 238, 316, 306, 256, 217, 215, 223, 239, 
    129, 256, 177, 253, 273, 316, 363, 283, 210, 205, 196, 210, 236, 270, 277, 
    277, 315, 320, 350, 337, 292, 262, 231, 267, 234, 244, 214, 185, 166, 173, 
    223, 167, 175, 182, 197, 201, 206, 198, 197, 178, 162, 141, 155, 161, 196, 
    16, 53, 48, 32, 27, 44, 72, 85, 91, 93, 92, 116, 163, 188, 205, 
    15, 48, 105, 68, 25, 33, 208, 196, 165, 179, 218, 238, 222, 200, 221, 
    26, 7, 31, 23, 5, 13, 155, 329, 350, 300, 211, 172, 181, 205, 236, 
    28, 8, 17, 14, 7, 9, 113, 370, 295, 203, 191, 198, 174, 191, 232, 
    15, 23, 15, 11, 20, 23, 54, 162, 173, 199, 182, 146, 174, 206, 245, 
    
    -- channel=67
    199, 201, 201, 201, 201, 202, 202, 202, 200, 200, 202, 200, 201, 201, 203, 
    201, 202, 202, 202, 201, 201, 202, 200, 195, 155, 169, 203, 202, 201, 204, 
    198, 201, 203, 203, 206, 202, 197, 177, 124, 84, 131, 192, 202, 203, 206, 
    198, 196, 204, 207, 208, 182, 190, 152, 139, 129, 130, 203, 200, 200, 206, 
    55, 82, 200, 199, 201, 173, 203, 188, 201, 185, 147, 109, 91, 143, 207, 
    120, 160, 198, 142, 165, 91, 104, 124, 156, 162, 132, 135, 104, 196, 205, 
    20, 51, 103, 130, 139, 0, 0, 63, 182, 186, 147, 109, 104, 111, 133, 
    0, 85, 16, 126, 130, 109, 168, 138, 88, 58, 29, 31, 56, 88, 128, 
    78, 147, 125, 168, 189, 168, 165, 90, 102, 91, 103, 79, 65, 55, 48, 
    94, 49, 68, 71, 76, 76, 65, 46, 55, 9, 15, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 19, 0, 37, 
    0, 0, 0, 0, 0, 0, 25, 71, 64, 28, 0, 0, 0, 15, 81, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 29, 95, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 47, 107, 
    
    -- channel=68
    189, 188, 188, 188, 188, 188, 188, 188, 186, 189, 185, 189, 188, 188, 188, 
    189, 188, 188, 188, 188, 188, 188, 189, 189, 180, 159, 178, 188, 188, 189, 
    186, 185, 188, 189, 188, 189, 185, 190, 160, 138, 148, 164, 191, 189, 190, 
    185, 190, 194, 190, 188, 190, 174, 176, 162, 159, 158, 182, 195, 194, 195, 
    121, 123, 170, 185, 187, 179, 189, 184, 187, 187, 177, 159, 142, 141, 195, 
    153, 165, 183, 167, 169, 157, 141, 148, 158, 179, 168, 164, 152, 173, 191, 
    90, 85, 126, 146, 175, 103, 77, 104, 158, 180, 167, 149, 136, 143, 138, 
    15, 132, 112, 125, 143, 156, 173, 179, 132, 114, 110, 106, 118, 131, 160, 
    62, 146, 154, 164, 172, 181, 176, 151, 144, 140, 134, 135, 123, 119, 111, 
    100, 90, 92, 91, 95, 96, 98, 93, 92, 83, 78, 65, 68, 81, 90, 
    22, 12, 15, 6, 12, 13, 13, 19, 31, 22, 24, 32, 47, 79, 93, 
    15, 17, 34, 19, 1, 0, 10, 57, 35, 33, 45, 69, 78, 72, 105, 
    32, 13, 0, 0, 0, 0, 24, 29, 21, 26, 30, 28, 72, 105, 137, 
    61, 1, 0, 0, 0, 0, 0, 0, 0, 0, 46, 97, 107, 122, 146, 
    60, 27, 20, 16, 10, 10, 21, 0, 31, 84, 103, 111, 119, 135, 156, 
    
    -- channel=69
    61, 56, 56, 56, 55, 56, 56, 57, 55, 58, 56, 55, 56, 56, 55, 
    60, 56, 56, 57, 55, 56, 55, 58, 61, 88, 10, 32, 58, 56, 55, 
    56, 54, 54, 57, 54, 60, 52, 78, 65, 82, 0, 0, 58, 55, 55, 
    52, 62, 54, 55, 57, 84, 12, 95, 67, 85, 65, 0, 60, 58, 56, 
    10, 0, 0, 49, 54, 85, 32, 71, 54, 76, 69, 46, 30, 0, 44, 
    71, 46, 32, 49, 28, 64, 5, 10, 12, 79, 85, 78, 105, 0, 41, 
    6, 0, 5, 22, 91, 151, 5, 0, 0, 51, 55, 46, 25, 29, 0, 
    0, 0, 33, 0, 41, 100, 40, 78, 38, 56, 69, 48, 30, 42, 23, 
    0, 58, 65, 38, 39, 66, 43, 100, 49, 55, 40, 58, 26, 20, 33, 
    0, 20, 12, 23, 26, 37, 61, 50, 39, 66, 31, 50, 25, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 15, 5, 0, 15, 0, 
    11, 0, 21, 27, 0, 0, 0, 69, 29, 19, 1, 5, 6, 8, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    
    -- channel=70
    164, 165, 165, 165, 165, 165, 165, 165, 164, 162, 164, 165, 165, 165, 165, 
    164, 165, 165, 165, 165, 165, 165, 165, 162, 133, 149, 164, 165, 165, 166, 
    162, 164, 166, 165, 167, 162, 164, 146, 128, 107, 136, 164, 165, 165, 166, 
    165, 166, 167, 167, 167, 147, 161, 141, 144, 141, 153, 181, 164, 166, 167, 
    96, 110, 154, 164, 164, 153, 176, 159, 165, 144, 121, 110, 104, 144, 164, 
    142, 161, 170, 138, 138, 96, 101, 112, 141, 146, 143, 150, 138, 178, 165, 
    72, 101, 109, 144, 137, 74, 106, 147, 169, 141, 118, 103, 101, 113, 132, 
    82, 126, 109, 146, 134, 133, 165, 137, 118, 114, 111, 118, 136, 140, 147, 
    166, 144, 145, 167, 161, 141, 131, 98, 121, 106, 105, 93, 90, 95, 95, 
    122, 79, 87, 87, 94, 95, 97, 95, 96, 78, 80, 65, 76, 84, 103, 
    36, 46, 33, 24, 24, 28, 27, 34, 36, 37, 42, 58, 83, 91, 109, 
    26, 63, 50, 41, 35, 40, 101, 92, 84, 86, 99, 97, 93, 98, 126, 
    42, 46, 46, 31, 32, 38, 129, 80, 88, 76, 76, 87, 103, 125, 143, 
    31, 39, 44, 38, 38, 39, 99, 123, 99, 108, 117, 127, 114, 125, 141, 
    35, 52, 49, 47, 48, 50, 76, 114, 112, 128, 113, 108, 117, 131, 146, 
    
    -- channel=71
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 10, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 20, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 10, 17, 1, 0, 0, 0, 
    1, 0, 0, 9, 0, 46, 0, 0, 0, 0, 7, 3, 22, 0, 0, 
    0, 0, 0, 0, 12, 98, 0, 0, 0, 0, 12, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 0, 21, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 41, 0, 16, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 7, 0, 0, 0, 
    10, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 13, 26, 12, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 
    51, 0, 0, 13, 7, 0, 0, 0, 3, 11, 1, 0, 0, 0, 0, 
    95, 0, 0, 2, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    79, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=72
    599, 596, 596, 596, 597, 598, 598, 598, 594, 596, 594, 599, 598, 596, 598, 
    600, 598, 598, 597, 595, 596, 596, 598, 593, 543, 506, 572, 597, 597, 599, 
    592, 592, 598, 600, 598, 599, 591, 577, 497, 453, 451, 536, 602, 599, 603, 
    586, 599, 606, 603, 602, 584, 548, 563, 512, 504, 487, 548, 609, 608, 610, 
    329, 367, 536, 589, 595, 593, 584, 596, 588, 581, 530, 460, 414, 462, 605, 
    501, 523, 563, 511, 526, 468, 438, 469, 514, 566, 532, 521, 480, 503, 596, 
    254, 274, 408, 483, 536, 279, 209, 307, 472, 563, 517, 457, 444, 439, 447, 
    102, 347, 310, 371, 481, 506, 537, 512, 399, 363, 331, 326, 355, 415, 460, 
    204, 522, 506, 537, 556, 559, 540, 498, 459, 441, 441, 419, 371, 349, 339, 
    293, 301, 305, 312, 321, 338, 335, 301, 307, 269, 249, 221, 222, 246, 280, 
    12, 17, 23, 3, 15, 36, 72, 94, 116, 96, 96, 116, 165, 241, 285, 
    6, 33, 99, 33, 0, 0, 82, 155, 107, 114, 158, 233, 251, 251, 324, 
    32, 0, 0, 0, 0, 0, 79, 216, 207, 190, 152, 148, 233, 308, 399, 
    114, 0, 0, 0, 0, 0, 0, 56, 19, 55, 172, 267, 300, 339, 426, 
    132, 18, 0, 0, 0, 0, 5, 47, 121, 230, 288, 300, 330, 380, 451, 
    
    -- channel=73
    288, 289, 289, 289, 289, 289, 289, 282, 278, 298, 308, 287, 287, 289, 289, 
    289, 289, 289, 289, 288, 288, 289, 281, 289, 315, 330, 302, 287, 289, 290, 
    287, 285, 286, 286, 286, 291, 302, 310, 356, 386, 376, 334, 290, 289, 293, 
    347, 330, 302, 282, 284, 277, 301, 308, 381, 406, 393, 381, 330, 319, 307, 
    393, 383, 345, 273, 288, 286, 292, 301, 343, 388, 419, 400, 367, 365, 330, 
    409, 387, 324, 266, 307, 339, 375, 371, 372, 375, 390, 380, 351, 373, 344, 
    418, 388, 372, 339, 351, 343, 376, 360, 372, 352, 360, 350, 353, 349, 372, 
    361, 375, 273, 273, 337, 359, 386, 353, 330, 330, 336, 339, 341, 365, 397, 
    370, 369, 348, 328, 374, 370, 403, 417, 443, 474, 495, 478, 462, 430, 403, 
    456, 488, 526, 536, 532, 527, 524, 502, 499, 487, 501, 475, 467, 427, 383, 
    281, 333, 361, 376, 373, 420, 515, 516, 504, 481, 472, 448, 434, 366, 304, 
    155, 215, 193, 165, 150, 189, 343, 377, 391, 381, 345, 331, 262, 219, 230, 
    94, 123, 80, 82, 108, 113, 125, 0, 0, 0, 0, 41, 119, 191, 265, 
    102, 98, 90, 90, 97, 98, 0, 0, 0, 0, 0, 92, 157, 221, 294, 
    99, 69, 94, 102, 91, 106, 47, 0, 0, 18, 89, 157, 190, 240, 303, 
    
    -- channel=74
    12, 12, 12, 12, 13, 13, 12, 12, 16, 12, 7, 12, 13, 12, 12, 
    12, 12, 12, 12, 13, 12, 13, 13, 15, 7, 25, 17, 12, 12, 12, 
    16, 15, 13, 12, 13, 12, 13, 10, 16, 0, 23, 23, 11, 14, 12, 
    2, 1, 8, 15, 13, 5, 30, 0, 0, 0, 0, 0, 2, 6, 7, 
    38, 47, 26, 21, 15, 0, 14, 5, 0, 0, 0, 15, 34, 45, 6, 
    0, 0, 0, 43, 30, 49, 51, 44, 29, 0, 0, 0, 0, 11, 3, 
    37, 56, 31, 21, 0, 0, 9, 0, 13, 5, 22, 35, 39, 27, 41, 
    47, 1, 26, 61, 5, 0, 0, 0, 27, 18, 3, 4, 3, 0, 0, 
    64, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 9, 15, 12, 
    20, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 
    66, 60, 45, 53, 65, 61, 25, 15, 8, 8, 9, 9, 0, 6, 32, 
    89, 96, 56, 63, 85, 93, 18, 0, 0, 0, 0, 5, 41, 46, 52, 
    83, 114, 118, 110, 105, 106, 135, 114, 118, 121, 127, 110, 88, 64, 47, 
    64, 105, 112, 106, 107, 107, 158, 232, 241, 170, 117, 90, 71, 65, 41, 
    68, 102, 102, 99, 101, 99, 122, 154, 127, 110, 92, 77, 68, 53, 34, 
    
    -- channel=75
    272, 271, 271, 271, 270, 272, 272, 272, 271, 271, 269, 271, 271, 271, 271, 
    273, 271, 271, 272, 270, 271, 270, 272, 272, 283, 234, 250, 271, 270, 271, 
    274, 272, 272, 273, 270, 275, 268, 284, 253, 221, 209, 243, 273, 273, 273, 
    249, 262, 270, 274, 275, 291, 239, 264, 201, 196, 170, 197, 271, 269, 273, 
    187, 184, 231, 274, 273, 276, 249, 266, 253, 262, 276, 257, 235, 206, 269, 
    176, 185, 262, 259, 261, 283, 263, 266, 260, 262, 196, 183, 186, 164, 265, 
    169, 165, 196, 192, 263, 127, 57, 55, 131, 274, 281, 269, 249, 265, 219, 
    27, 93, 150, 166, 206, 163, 172, 263, 223, 178, 132, 102, 108, 126, 164, 
    0, 244, 179, 219, 252, 275, 263, 239, 195, 215, 209, 222, 207, 204, 173, 
    176, 187, 182, 177, 174, 170, 165, 127, 139, 116, 124, 105, 87, 103, 120, 
    35, 29, 49, 52, 68, 82, 93, 98, 98, 84, 65, 59, 52, 81, 119, 
    21, 1, 55, 27, 0, 0, 0, 3, 0, 0, 7, 56, 140, 131, 120, 
    24, 0, 23, 16, 0, 0, 33, 188, 180, 184, 175, 117, 85, 125, 148, 
    74, 0, 0, 0, 0, 0, 0, 143, 147, 71, 45, 100, 135, 132, 173, 
    80, 0, 0, 0, 0, 0, 0, 52, 17, 79, 138, 132, 134, 150, 179, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 20, 19, 36, 41, 38, 33, 21, 12, 8, 4, 0, 0, 0, 0, 
    22, 19, 0, 1, 22, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 27, 24, 31, 30, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 28, 27, 30, 29, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 13, 17, 16, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=77
    255, 257, 257, 257, 258, 259, 259, 256, 256, 257, 263, 259, 257, 257, 258, 
    257, 258, 258, 257, 258, 257, 258, 257, 253, 242, 280, 263, 256, 257, 258, 
    263, 260, 259, 257, 257, 255, 266, 251, 262, 231, 274, 304, 259, 260, 261, 
    262, 262, 266, 259, 259, 239, 273, 222, 211, 188, 182, 252, 270, 268, 267, 
    260, 287, 306, 262, 261, 240, 252, 247, 254, 255, 283, 291, 278, 319, 279, 
    187, 200, 252, 253, 280, 286, 339, 334, 327, 255, 198, 177, 142, 233, 278, 
    254, 280, 267, 247, 212, 90, 129, 136, 205, 268, 290, 291, 295, 288, 308, 
    164, 152, 168, 237, 229, 150, 189, 222, 246, 199, 144, 133, 147, 158, 209, 
    183, 227, 191, 227, 272, 278, 296, 251, 239, 254, 272, 258, 276, 272, 231, 
    269, 264, 267, 262, 256, 242, 212, 185, 198, 165, 187, 162, 162, 174, 189, 
    89, 124, 110, 142, 168, 193, 206, 211, 195, 168, 157, 149, 144, 128, 169, 
    44, 107, 61, 22, 20, 40, 83, 0, 22, 32, 45, 77, 144, 151, 166, 
    0, 46, 59, 27, 20, 21, 195, 91, 64, 79, 117, 120, 103, 155, 204, 
    0, 16, 22, 18, 17, 19, 59, 0, 0, 34, 49, 112, 148, 179, 228, 
    32, 12, 16, 18, 12, 14, 34, 29, 16, 90, 128, 152, 166, 192, 229, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 6, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 12, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 0, 0, 0, 6, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 17, 95, 0, 0, 0, 0, 4, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 8, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 11, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    94, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 
    82, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    504, 506, 506, 506, 507, 507, 508, 505, 506, 505, 507, 508, 507, 506, 509, 
    505, 508, 508, 506, 506, 506, 507, 508, 496, 414, 472, 511, 505, 507, 509, 
    499, 502, 510, 508, 510, 504, 504, 456, 393, 364, 397, 506, 509, 510, 513, 
    513, 508, 515, 512, 510, 465, 505, 457, 463, 442, 445, 511, 516, 517, 520, 
    268, 333, 534, 500, 506, 496, 513, 506, 512, 482, 410, 357, 321, 457, 528, 
    451, 487, 470, 399, 453, 311, 354, 390, 461, 490, 474, 464, 404, 509, 519, 
    202, 261, 373, 468, 427, 148, 232, 358, 484, 460, 397, 342, 371, 341, 414, 
    188, 384, 237, 387, 456, 469, 512, 372, 321, 311, 287, 313, 345, 407, 412, 
    403, 454, 460, 473, 480, 454, 455, 400, 398, 353, 389, 325, 304, 283, 297, 
    283, 248, 261, 265, 280, 300, 288, 270, 278, 227, 219, 195, 214, 230, 276, 
    0, 64, 15, 7, 20, 49, 76, 89, 108, 85, 101, 131, 205, 239, 277, 
    0, 83, 95, 14, 0, 0, 263, 153, 140, 157, 212, 245, 212, 233, 330, 
    0, 0, 0, 0, 0, 0, 162, 184, 163, 130, 89, 146, 238, 298, 393, 
    11, 0, 0, 0, 0, 0, 26, 20, 0, 67, 195, 255, 268, 324, 410, 
    38, 20, 14, 5, 3, 8, 26, 56, 145, 238, 254, 262, 307, 355, 428, 
    
    -- channel=80
    782, 779, 779, 779, 780, 781, 782, 780, 778, 778, 781, 780, 779, 779, 782, 
    784, 782, 782, 781, 779, 780, 780, 780, 769, 704, 698, 764, 781, 781, 783, 
    777, 778, 783, 783, 785, 782, 777, 744, 662, 596, 615, 739, 785, 783, 789, 
    771, 780, 784, 788, 791, 748, 738, 719, 677, 657, 640, 726, 788, 787, 792, 
    491, 545, 732, 774, 782, 753, 756, 769, 774, 762, 703, 626, 576, 666, 789, 
    638, 681, 725, 674, 699, 619, 614, 653, 716, 739, 677, 660, 605, 682, 783, 
    418, 471, 584, 656, 666, 354, 320, 442, 649, 741, 694, 629, 616, 606, 648, 
    238, 459, 409, 545, 648, 639, 685, 651, 561, 517, 457, 442, 474, 543, 603, 
    370, 663, 642, 690, 742, 733, 715, 645, 607, 596, 609, 570, 532, 508, 493, 
    464, 496, 510, 525, 535, 542, 520, 475, 479, 422, 403, 358, 351, 370, 418, 
    70, 117, 127, 120, 137, 185, 246, 268, 275, 247, 231, 246, 304, 356, 404, 
    0, 57, 123, 29, 0, 0, 200, 223, 192, 209, 267, 345, 375, 362, 431, 
    0, 0, 0, 0, 0, 0, 200, 413, 392, 352, 286, 257, 306, 389, 508, 
    53, 0, 0, 0, 0, 0, 40, 197, 143, 126, 204, 309, 358, 424, 547, 
    77, 0, 0, 0, 0, 0, 0, 77, 129, 259, 335, 345, 392, 466, 574, 
    
    -- channel=81
    382, 379, 379, 379, 379, 380, 380, 380, 378, 382, 378, 380, 380, 379, 380, 
    382, 379, 379, 379, 376, 378, 376, 378, 380, 367, 300, 348, 378, 377, 378, 
    378, 375, 378, 380, 377, 385, 372, 382, 319, 304, 270, 321, 381, 380, 382, 
    362, 375, 379, 383, 382, 391, 330, 374, 321, 314, 283, 299, 385, 384, 385, 
    169, 187, 319, 372, 377, 389, 355, 384, 371, 390, 364, 300, 257, 252, 378, 
    338, 337, 343, 326, 346, 335, 305, 322, 327, 367, 332, 328, 312, 273, 368, 
    142, 122, 242, 304, 363, 184, 60, 98, 235, 372, 360, 321, 312, 296, 261, 
    8, 202, 167, 179, 291, 339, 343, 342, 236, 200, 172, 165, 176, 232, 271, 
    21, 347, 344, 351, 360, 369, 360, 372, 321, 316, 316, 308, 258, 216, 199, 
    171, 191, 179, 180, 180, 192, 191, 157, 169, 161, 136, 129, 125, 143, 154, 
    0, 0, 0, 0, 0, 2, 36, 49, 68, 52, 46, 50, 62, 129, 157, 
    16, 0, 88, 34, 0, 0, 3, 56, 15, 19, 47, 132, 167, 150, 178, 
    28, 0, 0, 0, 0, 0, 0, 171, 168, 167, 119, 73, 133, 177, 227, 
    119, 0, 0, 0, 0, 0, 0, 42, 45, 20, 85, 153, 180, 194, 248, 
    114, 4, 0, 0, 0, 0, 0, 0, 48, 119, 182, 184, 197, 225, 266, 
    
    -- channel=82
    40, 41, 41, 41, 41, 40, 40, 39, 40, 43, 40, 41, 41, 41, 41, 
    38, 39, 39, 39, 39, 39, 39, 39, 40, 38, 40, 36, 38, 39, 39, 
    37, 36, 38, 39, 37, 38, 42, 43, 48, 58, 83, 46, 40, 40, 40, 
    46, 46, 46, 37, 34, 35, 46, 46, 74, 84, 85, 87, 49, 48, 45, 
    49, 53, 45, 35, 37, 45, 60, 45, 57, 58, 73, 65, 49, 53, 50, 
    113, 102, 80, 44, 43, 65, 58, 56, 53, 53, 80, 93, 84, 95, 57, 
    45, 35, 48, 57, 76, 71, 95, 80, 82, 61, 59, 52, 58, 60, 52, 
    105, 123, 93, 63, 54, 89, 124, 98, 45, 30, 52, 72, 87, 87, 105, 
    124, 93, 90, 81, 64, 55, 62, 66, 97, 104, 93, 97, 88, 77, 59, 
    119, 40, 42, 30, 30, 36, 40, 53, 62, 63, 81, 75, 98, 102, 89, 
    99, 88, 78, 80, 82, 74, 61, 63, 67, 64, 82, 86, 90, 97, 99, 
    129, 157, 118, 135, 137, 134, 108, 123, 111, 104, 101, 108, 93, 76, 97, 
    145, 138, 92, 101, 130, 135, 96, 0, 0, 0, 9, 25, 77, 106, 106, 
    127, 141, 130, 127, 137, 139, 67, 0, 0, 0, 68, 112, 106, 108, 106, 
    133, 157, 158, 154, 147, 149, 121, 6, 63, 115, 109, 114, 114, 114, 106, 
    
    -- channel=83
    133, 130, 130, 130, 129, 130, 130, 131, 128, 133, 133, 128, 130, 130, 129, 
    133, 130, 130, 131, 129, 130, 128, 129, 135, 184, 99, 108, 132, 129, 129, 
    132, 131, 128, 130, 128, 137, 125, 162, 154, 173, 92, 86, 130, 129, 129, 
    120, 131, 122, 128, 133, 174, 86, 174, 134, 157, 127, 64, 128, 126, 126, 
    116, 76, 65, 125, 130, 158, 103, 141, 129, 159, 170, 151, 136, 50, 115, 
    138, 119, 132, 127, 124, 162, 122, 120, 108, 164, 138, 134, 177, 41, 116, 
    139, 92, 101, 89, 192, 211, 86, 51, 33, 148, 159, 158, 133, 156, 83, 
    49, 66, 112, 46, 121, 137, 95, 177, 143, 147, 143, 112, 94, 102, 92, 
    0, 173, 119, 123, 138, 160, 139, 181, 146, 162, 155, 180, 150, 142, 138, 
    109, 171, 171, 176, 176, 176, 202, 170, 167, 181, 169, 172, 139, 124, 109, 
    111, 93, 143, 131, 119, 127, 167, 170, 175, 180, 158, 140, 117, 112, 87, 
    91, 15, 119, 119, 88, 64, 55, 157, 133, 122, 103, 109, 127, 111, 55, 
    106, 36, 65, 94, 67, 59, 0, 177, 177, 177, 151, 100, 58, 59, 44, 
    159, 57, 54, 67, 58, 56, 0, 129, 165, 87, 34, 39, 68, 45, 56, 
    131, 48, 44, 46, 48, 48, 0, 52, 31, 8, 63, 57, 50, 53, 59, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 18, 83, 0, 0, 0, 
    23, 42, 30, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 51, 0, 
    24, 49, 23, 0, 0, 0, 14, 10, 13, 0, 0, 1, 0, 121, 0, 
    33, 60, 19, 11, 0, 0, 69, 87, 116, 0, 0, 0, 0, 0, 41, 
    105, 106, 5, 87, 0, 0, 62, 0, 0, 0, 0, 16, 45, 34, 78, 
    291, 0, 12, 41, 32, 0, 8, 0, 34, 38, 38, 23, 41, 29, 6, 
    172, 36, 59, 48, 49, 36, 22, 39, 51, 25, 61, 27, 67, 65, 62, 
    42, 76, 54, 66, 73, 85, 82, 77, 64, 54, 64, 74, 82, 55, 57, 
    3, 114, 2, 8, 33, 77, 125, 51, 72, 78, 82, 77, 43, 3, 46, 
    0, 72, 31, 0, 25, 47, 224, 0, 0, 0, 0, 0, 10, 41, 61, 
    0, 37, 44, 29, 38, 41, 90, 0, 0, 0, 7, 49, 11, 43, 53, 
    0, 17, 34, 34, 36, 41, 61, 0, 7, 53, 10, 2, 23, 37, 49, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 16, 32, 45, 50, 48, 51, 48, 43, 41, 28, 0, 0, 0, 0, 
    42, 40, 17, 33, 51, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 50, 47, 49, 52, 51, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 47, 49, 51, 51, 51, 34, 0, 19, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    17, 16, 16, 16, 16, 17, 17, 17, 15, 16, 17, 17, 16, 16, 16, 
    17, 16, 16, 16, 16, 16, 16, 16, 14, 26, 22, 15, 16, 16, 16, 
    19, 18, 16, 16, 15, 16, 19, 20, 27, 20, 26, 26, 18, 16, 17, 
    15, 17, 17, 16, 17, 20, 16, 11, 7, 3, 0, 1, 19, 18, 18, 
    28, 27, 21, 18, 17, 15, 11, 16, 14, 19, 40, 40, 34, 29, 20, 
    5, 4, 19, 26, 21, 51, 54, 50, 43, 20, 0, 0, 0, 0, 21, 
    34, 36, 25, 10, 19, 0, 0, 0, 0, 27, 41, 45, 42, 41, 34, 
    10, 0, 4, 8, 7, 0, 0, 26, 23, 8, 0, 0, 0, 0, 2, 
    0, 16, 3, 10, 23, 30, 30, 32, 18, 37, 35, 40, 44, 37, 21, 
    39, 39, 36, 37, 31, 26, 20, 11, 16, 11, 18, 13, 9, 15, 11, 
    2, 0, 7, 17, 23, 27, 31, 35, 29, 24, 18, 11, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 8, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 
    
    -- channel=87
    44, 44, 44, 44, 44, 44, 44, 46, 48, 42, 38, 44, 45, 44, 44, 
    43, 43, 43, 43, 43, 43, 43, 44, 43, 42, 28, 36, 43, 42, 42, 
    47, 46, 45, 44, 43, 45, 37, 41, 16, 5, 14, 32, 42, 44, 42, 
    15, 23, 37, 46, 45, 56, 41, 33, 0, 0, 0, 0, 27, 32, 37, 
    0, 0, 38, 50, 43, 38, 35, 36, 24, 20, 19, 18, 22, 12, 32, 
    0, 6, 23, 52, 56, 49, 51, 49, 29, 11, 0, 0, 0, 3, 21, 
    0, 0, 14, 26, 18, 0, 0, 0, 0, 36, 47, 51, 50, 41, 17, 
    0, 12, 17, 36, 14, 9, 5, 20, 14, 0, 0, 0, 0, 0, 0, 
    0, 5, 19, 27, 19, 23, 23, 22, 4, 0, 0, 1, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    69, 45, 68, 58, 57, 45, 0, 0, 0, 0, 0, 7, 51, 47, 41, 
    72, 72, 85, 85, 74, 72, 84, 209, 209, 192, 153, 97, 74, 55, 38, 
    86, 75, 76, 75, 75, 74, 128, 299, 264, 153, 100, 90, 71, 52, 34, 
    78, 84, 74, 70, 73, 66, 78, 125, 111, 113, 102, 73, 64, 49, 32, 
    
    -- channel=88
    302, 299, 299, 299, 299, 300, 299, 300, 298, 302, 296, 299, 300, 299, 299, 
    304, 301, 301, 302, 300, 301, 300, 302, 308, 328, 266, 282, 302, 301, 301, 
    301, 299, 301, 303, 300, 306, 297, 326, 301, 263, 228, 251, 304, 302, 303, 
    289, 300, 302, 303, 303, 329, 270, 302, 237, 235, 217, 244, 308, 305, 305, 
    271, 250, 259, 299, 303, 301, 276, 295, 282, 300, 305, 299, 290, 235, 302, 
    170, 178, 274, 292, 291, 309, 269, 270, 264, 296, 246, 213, 215, 196, 295, 
    230, 209, 238, 209, 287, 221, 123, 137, 189, 295, 299, 288, 253, 275, 245, 
    15, 129, 193, 195, 245, 194, 173, 284, 271, 248, 216, 173, 167, 173, 208, 
    0, 221, 184, 206, 256, 304, 299, 257, 198, 211, 201, 225, 215, 236, 223, 
    134, 215, 220, 222, 220, 221, 218, 193, 188, 172, 167, 148, 122, 128, 140, 
    96, 74, 102, 95, 102, 107, 118, 117, 126, 114, 96, 84, 80, 113, 130, 
    31, 0, 35, 26, 1, 0, 0, 59, 38, 27, 26, 62, 109, 134, 137, 
    48, 9, 26, 28, 0, 0, 0, 101, 88, 110, 135, 119, 108, 132, 171, 
    112, 0, 0, 0, 0, 0, 0, 17, 56, 36, 42, 97, 152, 159, 197, 
    119, 13, 5, 0, 0, 0, 4, 7, 8, 57, 144, 158, 155, 175, 208, 
    
    -- channel=89
    246, 247, 247, 247, 248, 248, 248, 250, 249, 242, 248, 245, 246, 247, 249, 
    245, 247, 247, 246, 246, 245, 246, 244, 235, 181, 207, 249, 247, 246, 247, 
    245, 249, 248, 246, 252, 245, 241, 201, 151, 137, 178, 241, 244, 245, 248, 
    234, 233, 238, 250, 257, 214, 233, 198, 200, 186, 189, 225, 226, 231, 238, 
    47, 97, 225, 246, 246, 225, 246, 239, 244, 217, 162, 109, 99, 182, 227, 
    233, 263, 228, 193, 202, 128, 143, 167, 200, 187, 183, 212, 193, 246, 228, 
    53, 100, 159, 219, 175, 13, 60, 132, 239, 220, 183, 150, 170, 145, 176, 
    110, 167, 84, 185, 184, 219, 262, 164, 118, 113, 97, 121, 139, 178, 181, 
    254, 232, 249, 275, 252, 195, 180, 168, 187, 167, 178, 142, 121, 83, 93, 
    171, 113, 112, 121, 127, 128, 120, 111, 123, 100, 88, 76, 95, 103, 129, 
    0, 11, 6, 3, 3, 21, 49, 60, 56, 55, 53, 72, 105, 127, 144, 
    0, 47, 79, 35, 7, 23, 164, 90, 84, 110, 156, 195, 185, 144, 163, 
    0, 0, 38, 20, 0, 2, 209, 385, 399, 330, 217, 153, 155, 147, 163, 
    0, 0, 14, 11, 2, 1, 191, 514, 408, 248, 189, 160, 112, 125, 152, 
    0, 0, 0, 0, 1, 0, 55, 201, 186, 176, 130, 85, 111, 129, 156, 
    
    -- channel=90
    0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 
    0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 52, 33, 0, 1, 2, 
    0, 3, 2, 0, 3, 0, 7, 0, 0, 0, 64, 71, 0, 1, 1, 
    17, 0, 4, 1, 2, 0, 48, 0, 0, 0, 0, 80, 0, 0, 1, 
    30, 70, 80, 7, 3, 0, 34, 0, 5, 0, 0, 0, 4, 100, 11, 
    0, 4, 31, 4, 14, 0, 36, 35, 46, 0, 0, 0, 0, 106, 22, 
    27, 95, 49, 24, 0, 0, 36, 68, 108, 1, 0, 0, 13, 6, 76, 
    104, 44, 0, 123, 4, 0, 14, 0, 7, 0, 0, 0, 22, 12, 32, 
    266, 5, 0, 31, 32, 0, 12, 0, 0, 0, 0, 0, 7, 10, 0, 
    137, 18, 36, 29, 27, 19, 0, 0, 18, 0, 10, 0, 10, 15, 35, 
    1, 54, 14, 32, 48, 61, 47, 38, 18, 8, 13, 24, 37, 11, 41, 
    0, 86, 0, 0, 0, 30, 100, 0, 0, 0, 20, 20, 23, 12, 53, 
    0, 35, 41, 0, 0, 11, 267, 2, 11, 7, 25, 38, 31, 44, 62, 
    0, 4, 21, 2, 5, 8, 161, 129, 73, 64, 49, 51, 14, 42, 57, 
    0, 0, 0, 0, 1, 3, 70, 85, 38, 70, 21, 4, 24, 31, 46, 
    
    -- channel=91
    449, 448, 448, 448, 448, 449, 450, 452, 451, 443, 444, 449, 449, 448, 449, 
    449, 448, 448, 447, 446, 446, 446, 448, 436, 379, 367, 426, 447, 446, 448, 
    447, 447, 450, 449, 450, 447, 440, 407, 328, 292, 302, 412, 449, 449, 451, 
    417, 432, 444, 454, 457, 430, 407, 405, 355, 332, 316, 357, 435, 440, 447, 
    146, 198, 392, 448, 446, 442, 430, 444, 431, 407, 350, 283, 245, 322, 435, 
    368, 396, 403, 367, 386, 306, 310, 341, 385, 398, 348, 357, 334, 345, 425, 
    113, 156, 264, 366, 369, 112, 69, 153, 302, 403, 367, 322, 329, 310, 311, 
    68, 217, 177, 265, 339, 366, 395, 340, 253, 219, 175, 180, 206, 266, 286, 
    153, 394, 385, 423, 418, 392, 362, 349, 322, 295, 307, 272, 236, 200, 192, 
    205, 174, 160, 164, 173, 180, 176, 142, 156, 128, 106, 93, 99, 130, 176, 
    0, 0, 0, 0, 0, 0, 0, 14, 26, 14, 11, 34, 77, 136, 194, 
    0, 6, 91, 15, 0, 0, 97, 40, 13, 35, 95, 165, 216, 202, 238, 
    0, 0, 0, 0, 0, 0, 114, 383, 382, 328, 236, 179, 193, 232, 276, 
    43, 0, 0, 0, 0, 0, 79, 412, 334, 218, 200, 224, 216, 229, 288, 
    49, 0, 0, 0, 0, 0, 0, 160, 174, 222, 229, 201, 226, 256, 303, 
    
    -- channel=92
    402, 399, 399, 399, 398, 400, 400, 399, 395, 400, 404, 400, 399, 399, 399, 
    401, 399, 399, 399, 397, 397, 396, 399, 395, 385, 339, 374, 398, 398, 399, 
    396, 394, 398, 400, 397, 401, 396, 395, 354, 363, 306, 362, 401, 399, 402, 
    399, 409, 402, 399, 401, 406, 351, 412, 391, 403, 379, 346, 414, 409, 407, 
    220, 231, 348, 387, 395, 425, 379, 414, 405, 417, 391, 335, 285, 297, 405, 
    421, 412, 385, 327, 352, 317, 309, 330, 365, 430, 409, 406, 404, 318, 401, 
    203, 190, 281, 357, 417, 283, 191, 225, 282, 388, 365, 329, 325, 323, 299, 
    140, 269, 232, 211, 354, 414, 406, 376, 287, 280, 268, 263, 273, 323, 321, 
    111, 424, 404, 395, 401, 404, 379, 417, 385, 371, 384, 365, 316, 283, 276, 
    237, 271, 271, 281, 287, 305, 322, 284, 283, 279, 254, 252, 240, 240, 245, 
    48, 65, 74, 62, 59, 82, 141, 165, 183, 175, 172, 178, 199, 223, 225, 
    74, 49, 158, 106, 46, 23, 169, 214, 176, 176, 188, 216, 217, 213, 228, 
    74, 0, 8, 30, 23, 15, 0, 149, 144, 136, 109, 110, 159, 215, 263, 
    158, 19, 12, 21, 17, 17, 0, 0, 0, 34, 109, 166, 207, 222, 283, 
    158, 50, 39, 37, 32, 35, 1, 23, 77, 124, 184, 204, 220, 255, 300, 
    
    -- channel=93
    838, 839, 839, 839, 840, 841, 842, 838, 836, 837, 844, 840, 840, 839, 843, 
    840, 841, 841, 839, 838, 838, 840, 837, 824, 739, 777, 833, 838, 839, 843, 
    835, 837, 843, 841, 844, 837, 841, 787, 712, 642, 712, 840, 843, 844, 849, 
    843, 845, 851, 847, 849, 786, 815, 759, 746, 723, 707, 829, 855, 854, 858, 
    530, 605, 831, 834, 840, 806, 837, 831, 850, 825, 770, 686, 621, 765, 864, 
    736, 786, 820, 716, 762, 661, 697, 738, 815, 806, 738, 734, 654, 797, 864, 
    457, 536, 645, 734, 733, 313, 376, 510, 745, 815, 756, 680, 687, 677, 733, 
    333, 552, 442, 635, 713, 692, 795, 713, 603, 539, 470, 479, 534, 615, 690, 
    531, 778, 722, 797, 843, 803, 797, 703, 703, 692, 715, 657, 620, 580, 545, 
    624, 557, 582, 587, 598, 602, 580, 523, 545, 460, 469, 405, 417, 442, 495, 
    73, 153, 142, 142, 170, 232, 300, 325, 329, 288, 280, 305, 374, 408, 473, 
    0, 138, 154, 37, 0, 0, 319, 245, 231, 252, 322, 401, 432, 399, 498, 
    0, 0, 5, 0, 0, 0, 341, 380, 358, 315, 260, 248, 325, 457, 597, 
    12, 0, 0, 0, 0, 0, 51, 93, 12, 80, 216, 368, 407, 492, 642, 
    43, 0, 0, 0, 0, 0, 0, 62, 132, 317, 377, 389, 454, 542, 668, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 116, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 56, 35, 89, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 99, 0, 97, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 61, 0, 0, 0, 6, 43, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 73, 0, 0, 0, 49, 0, 0, 95, 0, 0, 
    0, 0, 0, 0, 130, 281, 0, 0, 0, 0, 22, 36, 0, 19, 0, 
    0, 0, 0, 0, 0, 11, 0, 80, 13, 37, 43, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 19, 0, 101, 0, 0, 0, 41, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 0, 0, 41, 0, 38, 0, 0, 0, 
    25, 0, 18, 0, 0, 0, 0, 0, 1, 26, 0, 0, 0, 0, 0, 
    72, 0, 70, 100, 38, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 
    147, 0, 0, 70, 21, 0, 0, 51, 50, 83, 78, 0, 0, 0, 0, 
    327, 0, 0, 16, 0, 0, 0, 41, 168, 20, 0, 0, 0, 0, 0, 
    277, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 42, 12, 30, 49, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 55, 47, 44, 54, 58, 40, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 60, 61, 60, 61, 61, 64, 42, 38, 28, 6, 0, 0, 0, 0, 
    9, 48, 52, 54, 54, 52, 55, 52, 27, 5, 0, 0, 0, 0, 0, 
    
    -- channel=96
    18, 17, 17, 17, 17, 17, 17, 19, 22, 14, 11, 16, 17, 17, 16, 
    19, 17, 17, 18, 18, 18, 17, 18, 19, 22, 0, 9, 19, 17, 17, 
    21, 21, 18, 18, 18, 19, 13, 18, 10, 0, 0, 0, 18, 17, 16, 
    0, 1, 8, 20, 22, 28, 4, 20, 0, 0, 0, 0, 0, 3, 8, 
    0, 0, 0, 25, 20, 17, 0, 12, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 35, 17, 26, 5, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 13, 0, 0, 0, 0, 9, 19, 9, 11, 0, 
    0, 0, 5, 4, 0, 0, 0, 0, 17, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 7, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 2, 9, 12, 7, 0, 0, 0, 0, 0, 0, 2, 25, 0, 
    30, 8, 53, 55, 23, 16, 35, 192, 187, 170, 144, 110, 42, 3, 0, 
    33, 16, 24, 30, 19, 18, 78, 361, 357, 206, 80, 25, 17, 0, 0, 
    36, 14, 6, 5, 12, 8, 19, 148, 94, 37, 34, 11, 0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 23, 0, 0, 0, 
    3, 0, 1, 0, 0, 2, 11, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 37, 0, 0, 0, 14, 0, 2, 0, 0, 0, 0, 12, 7, 
    0, 12, 31, 0, 10, 0, 4, 5, 9, 1, 0, 0, 0, 39, 9, 
    0, 4, 5, 0, 15, 0, 2, 11, 25, 8, 0, 0, 0, 7, 7, 
    12, 43, 0, 42, 3, 0, 14, 1, 0, 0, 0, 0, 0, 4, 6, 
    57, 34, 0, 21, 19, 6, 11, 0, 0, 0, 8, 0, 5, 0, 0, 
    71, 0, 2, 0, 0, 0, 0, 0, 4, 0, 4, 0, 0, 2, 12, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 12, 
    0, 13, 0, 0, 0, 0, 58, 0, 0, 0, 3, 6, 12, 0, 14, 
    0, 2, 5, 0, 0, 0, 59, 1, 0, 1, 0, 0, 0, 13, 20, 
    0, 0, 0, 0, 0, 0, 3, 19, 0, 0, 0, 17, 5, 9, 22, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 21, 13, 0, 7, 9, 18, 
    
    -- channel=99
    123, 126, 126, 126, 126, 126, 126, 130, 133, 120, 118, 125, 127, 126, 127, 
    123, 126, 126, 125, 125, 125, 125, 127, 121, 73, 89, 125, 126, 125, 126, 
    122, 126, 129, 126, 129, 127, 113, 91, 30, 14, 46, 103, 125, 125, 125, 
    94, 99, 118, 130, 132, 119, 120, 93, 55, 35, 43, 89, 97, 107, 115, 
    0, 0, 115, 129, 127, 117, 131, 117, 103, 71, 12, 0, 0, 51, 105, 
    56, 84, 109, 88, 106, 6, 15, 31, 48, 60, 49, 65, 59, 107, 94, 
    0, 0, 38, 84, 67, 0, 0, 39, 107, 86, 46, 25, 44, 29, 37, 
    0, 82, 18, 113, 80, 79, 102, 39, 18, 14, 3, 25, 37, 59, 45, 
    119, 91, 87, 120, 84, 57, 46, 6, 18, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 53, 
    12, 34, 51, 31, 21, 18, 57, 0, 0, 0, 35, 74, 72, 81, 102, 
    37, 30, 75, 59, 38, 41, 169, 312, 325, 276, 185, 150, 141, 109, 100, 
    25, 47, 56, 54, 48, 49, 185, 556, 448, 288, 218, 162, 107, 92, 83, 
    21, 65, 54, 46, 57, 50, 85, 257, 231, 206, 149, 92, 98, 88, 83, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 1, 8, 12, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 45, 32, 47, 59, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 58, 52, 60, 67, 65, 18, 18, 26, 26, 8, 0, 0, 0, 0, 
    43, 67, 66, 67, 69, 68, 51, 65, 57, 28, 20, 0, 0, 0, 0, 
    31, 56, 58, 58, 60, 57, 45, 37, 43, 11, 0, 0, 0, 0, 0, 
    
    -- channel=101
    242, 242, 242, 242, 242, 243, 243, 243, 239, 243, 249, 243, 242, 242, 243, 
    244, 243, 243, 243, 242, 242, 242, 241, 239, 247, 230, 237, 242, 242, 243, 
    245, 244, 243, 243, 242, 246, 244, 245, 237, 234, 204, 242, 245, 243, 246, 
    243, 246, 246, 244, 246, 250, 221, 239, 201, 199, 168, 190, 252, 248, 249, 
    179, 192, 243, 239, 244, 255, 215, 247, 237, 258, 265, 241, 219, 220, 252, 
    188, 183, 229, 213, 242, 245, 261, 265, 261, 259, 204, 183, 169, 152, 250, 
    181, 174, 217, 196, 236, 89, 52, 64, 139, 258, 264, 249, 249, 239, 223, 
    49, 85, 98, 132, 214, 170, 164, 207, 194, 168, 123, 101, 99, 135, 153, 
    0, 255, 180, 205, 249, 265, 268, 264, 218, 231, 250, 241, 222, 205, 185, 
    169, 226, 232, 239, 233, 232, 226, 178, 187, 159, 165, 149, 125, 122, 127, 
    0, 18, 42, 54, 66, 93, 148, 156, 153, 131, 110, 93, 91, 87, 94, 
    0, 0, 2, 0, 0, 0, 0, 0, 1, 6, 16, 57, 90, 87, 77, 
    0, 0, 0, 0, 0, 0, 0, 116, 84, 75, 57, 37, 20, 59, 105, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 54, 73, 137, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 50, 65, 93, 143, 
    
    -- channel=102
    528, 529, 529, 529, 529, 531, 531, 532, 531, 525, 527, 530, 530, 529, 531, 
    531, 531, 531, 531, 530, 530, 531, 531, 523, 479, 485, 523, 531, 530, 533, 
    530, 532, 535, 532, 534, 533, 526, 503, 448, 386, 413, 510, 534, 533, 536, 
    506, 516, 532, 538, 540, 516, 508, 477, 399, 373, 356, 465, 525, 527, 535, 
    349, 392, 514, 534, 535, 513, 509, 516, 501, 487, 451, 421, 410, 468, 532, 
    334, 369, 496, 473, 499, 435, 445, 464, 489, 478, 394, 369, 329, 414, 524, 
    291, 340, 407, 411, 428, 149, 155, 247, 400, 503, 475, 439, 434, 430, 447, 
    114, 240, 262, 402, 435, 335, 368, 406, 390, 343, 270, 247, 267, 307, 349, 
    184, 439, 353, 429, 481, 487, 483, 387, 348, 338, 352, 333, 324, 332, 317, 
    293, 312, 319, 323, 324, 323, 299, 258, 269, 204, 217, 177, 164, 188, 245, 
    37, 64, 67, 72, 97, 120, 136, 144, 143, 118, 98, 104, 140, 184, 246, 
    0, 30, 44, 0, 0, 0, 51, 21, 25, 39, 91, 162, 223, 244, 276, 
    0, 0, 31, 0, 0, 0, 229, 380, 352, 319, 269, 240, 210, 257, 329, 
    0, 0, 0, 0, 0, 0, 70, 358, 281, 186, 161, 213, 250, 281, 362, 
    35, 0, 0, 0, 0, 0, 0, 141, 114, 196, 248, 238, 264, 304, 373, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 29, 13, 7, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    34, 34, 34, 34, 34, 34, 34, 34, 35, 34, 33, 34, 34, 34, 34, 
    33, 33, 33, 33, 32, 33, 33, 33, 35, 16, 0, 22, 33, 33, 33, 
    31, 31, 33, 33, 34, 35, 30, 27, 0, 0, 0, 12, 32, 34, 34, 
    28, 32, 31, 34, 35, 29, 18, 25, 21, 21, 24, 30, 29, 32, 32, 
    0, 0, 0, 30, 32, 28, 40, 33, 38, 31, 6, 0, 0, 0, 25, 
    48, 57, 33, 10, 15, 0, 0, 0, 0, 14, 20, 36, 35, 38, 24, 
    0, 0, 0, 17, 24, 0, 0, 0, 21, 21, 6, 0, 0, 0, 0, 
    0, 23, 0, 0, 0, 40, 66, 29, 0, 0, 0, 0, 1, 14, 26, 
    22, 30, 54, 60, 39, 19, 8, 6, 22, 6, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 22, 0, 0, 6, 12, 17, 
    0, 0, 0, 0, 0, 0, 0, 53, 55, 16, 24, 28, 5, 4, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 26, 18, 0, 4, 11, 14, 
    
    -- channel=105
    655, 655, 655, 655, 656, 656, 657, 655, 655, 654, 653, 656, 656, 655, 658, 
    655, 655, 655, 654, 652, 653, 653, 655, 645, 553, 553, 634, 654, 654, 657, 
    647, 649, 658, 656, 658, 657, 646, 606, 490, 437, 479, 612, 657, 657, 662, 
    641, 651, 657, 663, 664, 619, 612, 588, 558, 535, 527, 611, 657, 661, 665, 
    255, 328, 612, 645, 654, 633, 653, 650, 655, 629, 537, 435, 374, 498, 661, 
    578, 626, 617, 520, 572, 430, 443, 490, 562, 602, 561, 572, 514, 604, 651, 
    187, 238, 406, 557, 559, 167, 168, 317, 545, 605, 532, 451, 461, 439, 473, 
    101, 425, 258, 419, 512, 570, 648, 519, 373, 329, 289, 313, 362, 451, 500, 
    360, 582, 596, 635, 634, 592, 572, 512, 511, 465, 487, 427, 370, 317, 306, 
    347, 272, 277, 282, 297, 316, 304, 272, 286, 231, 211, 172, 199, 231, 288, 
    0, 0, 0, 0, 0, 0, 5, 31, 58, 33, 39, 75, 152, 236, 299, 
    0, 3, 80, 0, 0, 0, 174, 122, 73, 94, 172, 270, 278, 257, 358, 
    0, 0, 0, 0, 0, 0, 98, 303, 310, 268, 170, 142, 249, 336, 444, 
    2, 0, 0, 0, 0, 0, 0, 186, 103, 92, 210, 301, 302, 356, 464, 
    7, 0, 0, 0, 0, 0, 0, 55, 147, 275, 305, 285, 337, 401, 492, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 91, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 36, 150, 80, 109, 55, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    366, 331, 69, 2, 0, 0, 0, 0, 0, 0, 132, 250, 316, 194, 0, 
    0, 0, 0, 139, 122, 351, 390, 323, 180, 0, 0, 0, 0, 0, 0, 
    418, 409, 220, 0, 0, 0, 0, 0, 0, 52, 201, 291, 261, 262, 224, 
    59, 0, 33, 113, 0, 0, 0, 0, 208, 118, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 60, 133, 45, 0, 52, 43, 115, 216, 266, 179, 
    184, 348, 338, 325, 278, 208, 132, 70, 96, 54, 126, 95, 25, 33, 25, 
    247, 229, 289, 376, 435, 462, 435, 398, 327, 283, 206, 123, 0, 0, 0, 
    45, 57, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 4, 15, 0, 
    0, 71, 171, 106, 30, 20, 274, 207, 114, 164, 279, 177, 0, 0, 0, 
    0, 0, 24, 24, 8, 7, 76, 244, 318, 114, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    38, 32, 32, 32, 32, 32, 32, 36, 34, 32, 28, 30, 32, 32, 31, 
    37, 32, 32, 33, 31, 32, 31, 33, 34, 43, 0, 6, 34, 32, 31, 
    34, 32, 30, 33, 33, 36, 25, 41, 12, 18, 0, 0, 32, 31, 30, 
    10, 24, 22, 34, 36, 48, 0, 54, 21, 33, 23, 0, 19, 20, 24, 
    0, 0, 0, 31, 30, 41, 9, 32, 22, 30, 8, 0, 0, 0, 4, 
    35, 26, 1, 32, 0, 19, 0, 0, 0, 11, 28, 38, 68, 0, 0, 
    0, 0, 0, 0, 25, 122, 0, 0, 0, 12, 14, 11, 0, 0, 0, 
    0, 0, 34, 0, 0, 59, 18, 45, 2, 14, 30, 11, 0, 1, 0, 
    0, 0, 40, 18, 2, 9, 0, 29, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    32, 0, 42, 56, 31, 1, 0, 66, 20, 18, 18, 27, 32, 26, 0, 
    76, 0, 10, 38, 24, 12, 0, 154, 171, 152, 102, 49, 32, 0, 0, 
    114, 18, 17, 23, 17, 13, 58, 248, 241, 113, 52, 17, 9, 0, 0, 
    91, 31, 13, 15, 17, 13, 31, 74, 62, 20, 21, 6, 0, 0, 0, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 37, 26, 0, 0, 1, 
    0, 0, 1, 0, 2, 0, 4, 0, 0, 0, 51, 66, 0, 0, 1, 
    13, 0, 3, 0, 0, 0, 45, 0, 1, 0, 13, 89, 0, 0, 2, 
    0, 28, 73, 2, 0, 0, 38, 0, 15, 0, 0, 0, 0, 80, 14, 
    15, 51, 35, 0, 0, 0, 0, 6, 33, 0, 0, 0, 0, 127, 22, 
    0, 41, 13, 36, 0, 0, 34, 80, 117, 0, 0, 0, 0, 0, 51, 
    99, 80, 0, 106, 4, 0, 67, 0, 0, 0, 0, 0, 28, 27, 47, 
    296, 11, 15, 43, 33, 0, 0, 0, 3, 0, 5, 0, 0, 0, 0, 
    124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 34, 
    0, 20, 0, 0, 0, 9, 0, 0, 0, 0, 0, 4, 36, 16, 44, 
    0, 78, 0, 0, 0, 18, 135, 0, 8, 20, 50, 44, 24, 5, 57, 
    0, 21, 2, 0, 0, 0, 228, 0, 0, 0, 0, 0, 16, 47, 72, 
    0, 0, 2, 0, 0, 0, 108, 1, 0, 0, 29, 53, 14, 47, 65, 
    0, 0, 0, 0, 0, 2, 45, 15, 20, 80, 21, 4, 29, 43, 60, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 5, 1, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    220, 223, 223, 223, 223, 223, 224, 222, 221, 220, 227, 223, 222, 223, 224, 
    222, 224, 224, 223, 223, 223, 224, 223, 214, 166, 234, 239, 222, 224, 225, 
    221, 222, 225, 223, 226, 218, 227, 187, 184, 176, 205, 256, 224, 224, 227, 
    238, 230, 231, 225, 225, 183, 239, 190, 210, 199, 209, 253, 231, 230, 231, 
    162, 204, 266, 222, 224, 214, 228, 221, 228, 209, 180, 171, 166, 258, 239, 
    200, 216, 209, 178, 205, 135, 183, 197, 234, 217, 215, 206, 164, 244, 239, 
    139, 186, 206, 230, 167, 62, 149, 213, 247, 201, 176, 159, 183, 163, 227, 
    161, 174, 126, 203, 223, 197, 222, 145, 166, 168, 152, 165, 179, 200, 194, 
    276, 208, 202, 211, 221, 201, 210, 177, 188, 167, 194, 154, 158, 159, 168, 
    161, 160, 173, 180, 185, 191, 175, 169, 170, 139, 142, 131, 138, 136, 158, 
    32, 83, 54, 61, 68, 86, 108, 114, 110, 99, 104, 116, 150, 136, 148, 
    0, 75, 39, 1, 0, 18, 169, 83, 103, 114, 134, 127, 99, 124, 162, 
    0, 3, 18, 0, 0, 0, 162, 75, 53, 32, 32, 90, 113, 137, 185, 
    0, 0, 0, 0, 0, 0, 67, 14, 0, 51, 92, 102, 113, 149, 192, 
    0, 0, 0, 2, 2, 5, 31, 56, 71, 96, 89, 109, 133, 159, 196, 
    
    -- channel=113
    104, 104, 104, 104, 103, 103, 103, 104, 107, 100, 97, 104, 104, 104, 104, 
    101, 102, 102, 101, 101, 101, 100, 104, 95, 42, 51, 92, 101, 102, 102, 
    96, 98, 103, 104, 103, 99, 94, 66, 11, 29, 27, 72, 102, 102, 102, 
    87, 91, 100, 104, 101, 86, 89, 101, 117, 116, 120, 90, 94, 97, 101, 
    0, 0, 74, 97, 97, 120, 114, 114, 106, 79, 20, 0, 0, 20, 95, 
    171, 174, 90, 42, 51, 0, 0, 0, 34, 90, 130, 155, 147, 118, 89, 
    0, 0, 0, 109, 93, 8, 19, 72, 101, 65, 17, 0, 13, 0, 1, 
    30, 128, 31, 40, 91, 197, 203, 60, 0, 0, 23, 65, 82, 118, 82, 
    121, 125, 169, 138, 78, 48, 27, 65, 78, 35, 41, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 54, 68, 
    60, 57, 107, 85, 58, 38, 143, 101, 62, 71, 109, 117, 74, 69, 115, 
    87, 36, 21, 44, 62, 62, 0, 110, 132, 101, 29, 44, 119, 119, 117, 
    104, 74, 63, 65, 71, 72, 58, 112, 75, 94, 168, 150, 111, 105, 100, 
    103, 119, 105, 96, 97, 95, 75, 98, 174, 182, 136, 109, 119, 116, 107, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 35, 63, 68, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41, 0, 47, 0, 0, 0, 0, 0, 0, 0, 
    82, 23, 0, 0, 0, 16, 0, 0, 0, 2, 59, 82, 85, 0, 0, 
    0, 0, 0, 42, 0, 141, 59, 40, 0, 13, 0, 0, 0, 0, 0, 
    94, 34, 0, 0, 22, 185, 0, 0, 0, 4, 68, 99, 53, 69, 0, 
    0, 0, 40, 0, 0, 0, 0, 37, 64, 58, 34, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 2, 69, 0, 14, 0, 44, 38, 63, 50, 
    0, 83, 61, 65, 52, 42, 54, 25, 10, 51, 32, 55, 0, 0, 0, 
    100, 22, 97, 100, 98, 93, 95, 87, 83, 91, 55, 13, 0, 0, 0, 
    58, 0, 16, 40, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71, 0, 24, 65, 24, 0, 0, 95, 79, 98, 114, 50, 0, 0, 0, 
    151, 1, 0, 12, 1, 0, 0, 8, 121, 11, 0, 0, 0, 0, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    9, 10, 10, 10, 10, 10, 10, 9, 13, 9, 5, 11, 11, 10, 9, 
    9, 10, 10, 10, 10, 10, 10, 12, 12, 5, 22, 11, 9, 10, 9, 
    11, 10, 11, 10, 8, 8, 11, 8, 18, 16, 15, 17, 11, 11, 9, 
    1, 3, 11, 11, 6, 9, 26, 15, 0, 0, 0, 0, 8, 10, 10, 
    41, 48, 31, 15, 11, 16, 10, 11, 0, 0, 0, 21, 34, 44, 13, 
    0, 0, 0, 29, 30, 31, 39, 34, 23, 6, 4, 0, 0, 0, 6, 
    27, 33, 29, 28, 0, 30, 29, 22, 0, 0, 11, 25, 34, 19, 30, 
    46, 14, 47, 42, 30, 5, 0, 0, 25, 27, 23, 24, 19, 9, 0, 
    34, 0, 0, 0, 0, 0, 9, 11, 0, 0, 0, 0, 3, 20, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 
    75, 61, 35, 41, 50, 36, 0, 0, 0, 0, 3, 4, 2, 13, 33, 
    116, 108, 76, 84, 103, 99, 28, 0, 0, 0, 0, 0, 12, 53, 59, 
    116, 123, 118, 123, 126, 122, 77, 30, 23, 37, 61, 95, 88, 71, 58, 
    115, 127, 124, 125, 128, 129, 98, 67, 93, 116, 113, 89, 92, 81, 56, 
    139, 142, 139, 135, 132, 130, 115, 113, 123, 109, 101, 106, 93, 75, 52, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 12, 13, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 14, 16, 17, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 7, 8, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 44, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 50, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 13, 0, 0, 24, 0, 0, 
    0, 0, 0, 0, 0, 211, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 0, 0, 0, 42, 41, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 16, 0, 0, 0, 
    16, 0, 1, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    64, 0, 45, 53, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74, 0, 0, 70, 31, 0, 0, 128, 103, 92, 79, 67, 0, 0, 0, 
    199, 1, 0, 19, 4, 0, 0, 121, 210, 112, 0, 0, 0, 0, 0, 
    203, 15, 0, 0, 0, 0, 0, 24, 3, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    176, 175, 175, 175, 174, 175, 175, 171, 164, 181, 190, 175, 174, 175, 175, 
    175, 174, 174, 174, 173, 173, 172, 170, 177, 207, 168, 167, 173, 174, 174, 
    170, 168, 171, 173, 171, 179, 178, 199, 204, 247, 191, 173, 175, 172, 177, 
    214, 210, 184, 168, 171, 191, 149, 211, 247, 281, 263, 207, 208, 198, 188, 
    157, 138, 175, 155, 171, 200, 171, 196, 213, 253, 262, 218, 172, 144, 199, 
    303, 278, 210, 127, 167, 169, 179, 183, 193, 259, 268, 270, 274, 199, 207, 
    180, 128, 174, 194, 272, 222, 182, 173, 177, 213, 203, 180, 179, 186, 159, 
    127, 229, 118, 75, 190, 266, 270, 237, 160, 171, 187, 193, 193, 230, 232, 
    101, 280, 259, 233, 243, 242, 243, 292, 297, 307, 325, 312, 267, 224, 208, 
    238, 257, 280, 291, 292, 303, 327, 294, 293, 292, 287, 276, 268, 236, 199, 
    68, 99, 124, 119, 105, 135, 229, 245, 255, 243, 241, 229, 222, 196, 142, 
    36, 27, 98, 69, 28, 25, 177, 248, 226, 215, 183, 180, 122, 86, 93, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 74, 123, 
    72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 52, 83, 141, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 50, 71, 108, 154, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 11, 9, 0, 0, 
    0, 1, 0, 6, 0, 18, 8, 4, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 35, 0, 0, 0, 0, 10, 15, 0, 2, 0, 
    0, 0, 14, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 5, 0, 0, 0, 0, 3, 6, 9, 1, 11, 10, 6, 0, 
    0, 3, 0, 1, 0, 0, 0, 0, 0, 8, 0, 0, 0, 2, 0, 
    7, 0, 0, 3, 2, 0, 0, 2, 2, 3, 0, 0, 0, 0, 0, 
    9, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    11, 13, 0, 0, 1, 0, 0, 0, 0, 3, 8, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 9, 0, 0, 0, 0, 
    13, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 
    25, 21, 0, 0, 0, 0, 10, 7, 11, 0, 0, 6, 6, 12, 0, 
    32, 48, 9, 24, 0, 27, 75, 54, 8, 0, 0, 0, 9, 4, 19, 
    137, 42, 34, 31, 5, 12, 16, 0, 5, 13, 21, 35, 38, 27, 10, 
    129, 5, 18, 5, 0, 0, 0, 1, 24, 23, 29, 18, 32, 29, 30, 
    69, 38, 37, 32, 32, 30, 28, 36, 36, 45, 51, 61, 69, 66, 59, 
    90, 106, 85, 94, 94, 98, 89, 86, 81, 85, 90, 93, 91, 59, 57, 
    117, 134, 104, 110, 126, 138, 156, 77, 95, 97, 95, 67, 62, 61, 54, 
    98, 129, 116, 117, 131, 134, 120, 49, 54, 51, 58, 73, 60, 58, 38, 
    68, 133, 133, 131, 134, 135, 122, 55, 67, 93, 83, 64, 52, 48, 31, 
    71, 120, 126, 128, 130, 132, 120, 98, 95, 81, 53, 51, 49, 41, 25, 
    
    -- channel=123
    548, 549, 549, 549, 550, 551, 551, 551, 550, 545, 550, 549, 549, 549, 552, 
    550, 551, 551, 550, 549, 549, 551, 550, 538, 451, 490, 548, 550, 550, 553, 
    546, 549, 554, 551, 556, 549, 547, 496, 422, 360, 415, 536, 553, 553, 557, 
    541, 545, 554, 558, 561, 501, 533, 474, 442, 414, 416, 530, 548, 552, 558, 
    285, 354, 538, 548, 552, 512, 543, 532, 541, 512, 436, 378, 353, 475, 556, 
    410, 461, 502, 452, 487, 365, 393, 428, 487, 484, 439, 432, 368, 502, 547, 
    220, 291, 387, 458, 412, 118, 158, 302, 484, 499, 444, 390, 395, 378, 443, 
    112, 306, 231, 397, 438, 409, 475, 396, 348, 313, 260, 264, 300, 357, 402, 
    349, 435, 429, 484, 512, 480, 475, 383, 381, 346, 370, 320, 299, 286, 284, 
    283, 272, 284, 294, 306, 309, 282, 255, 262, 203, 191, 151, 162, 182, 244, 
    0, 1, 0, 0, 0, 33, 68, 82, 84, 61, 55, 81, 145, 192, 245, 
    0, 0, 0, 0, 0, 0, 111, 57, 47, 71, 135, 200, 205, 216, 288, 
    0, 0, 0, 0, 0, 0, 203, 302, 283, 232, 167, 161, 200, 252, 352, 
    0, 0, 0, 0, 0, 0, 55, 259, 152, 118, 152, 207, 218, 277, 372, 
    0, 0, 0, 0, 0, 0, 0, 79, 97, 186, 207, 203, 247, 306, 392, 
    
    -- channel=124
    765, 766, 766, 766, 767, 769, 769, 767, 765, 764, 766, 770, 768, 766, 769, 
    767, 768, 768, 767, 765, 765, 767, 768, 755, 683, 714, 756, 765, 766, 769, 
    766, 765, 772, 769, 769, 767, 765, 727, 645, 569, 621, 767, 772, 772, 776, 
    750, 760, 778, 777, 774, 737, 749, 687, 626, 580, 562, 696, 780, 780, 785, 
    478, 553, 790, 766, 769, 741, 749, 752, 746, 728, 689, 635, 583, 701, 796, 
    577, 627, 715, 661, 728, 620, 675, 706, 751, 727, 623, 591, 516, 659, 779, 
    401, 457, 586, 658, 644, 217, 242, 364, 596, 731, 696, 640, 647, 624, 664, 
    191, 443, 366, 554, 636, 566, 630, 603, 540, 462, 371, 362, 403, 480, 556, 
    350, 645, 602, 664, 725, 729, 731, 633, 586, 564, 600, 548, 531, 506, 467, 
    464, 452, 456, 456, 458, 462, 425, 368, 385, 308, 315, 267, 270, 313, 379, 
    0, 66, 31, 48, 90, 133, 166, 186, 200, 151, 140, 156, 217, 279, 371, 
    0, 70, 98, 0, 0, 0, 152, 30, 30, 53, 131, 235, 315, 331, 423, 
    0, 0, 0, 0, 0, 0, 236, 344, 301, 274, 242, 232, 283, 395, 529, 
    18, 0, 0, 0, 0, 0, 28, 108, 35, 85, 187, 322, 381, 446, 577, 
    67, 0, 0, 0, 0, 0, 0, 50, 112, 283, 364, 380, 426, 494, 600, 
    
    -- channel=125
    483, 481, 481, 481, 481, 483, 482, 483, 480, 481, 476, 483, 483, 481, 482, 
    486, 483, 483, 483, 481, 482, 482, 485, 485, 475, 423, 460, 482, 482, 484, 
    483, 481, 484, 486, 482, 487, 477, 487, 435, 381, 353, 428, 487, 486, 487, 
    460, 474, 487, 489, 487, 499, 443, 461, 366, 344, 314, 382, 489, 488, 491, 
    327, 342, 442, 483, 485, 486, 449, 478, 449, 458, 445, 415, 393, 388, 487, 
    297, 310, 425, 444, 455, 449, 419, 431, 436, 457, 377, 338, 314, 320, 473, 
    260, 268, 359, 359, 427, 211, 113, 161, 300, 459, 452, 421, 402, 398, 382, 
    19, 183, 234, 297, 386, 323, 309, 394, 359, 316, 253, 216, 221, 260, 303, 
    0, 378, 322, 365, 417, 460, 457, 408, 315, 322, 320, 324, 303, 306, 290, 
    193, 269, 264, 267, 263, 270, 256, 208, 219, 178, 171, 149, 124, 151, 185, 
    22, 12, 27, 22, 45, 60, 73, 81, 92, 68, 52, 50, 64, 128, 185, 
    0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 78, 156, 183, 221, 
    3, 0, 0, 0, 0, 0, 27, 205, 171, 174, 174, 156, 169, 216, 284, 
    99, 0, 0, 0, 0, 0, 0, 111, 114, 83, 104, 176, 234, 254, 322, 
    126, 0, 0, 0, 0, 0, 0, 52, 59, 136, 229, 244, 253, 283, 337, 
    
    -- channel=126
    340, 337, 337, 337, 337, 338, 338, 341, 335, 336, 337, 338, 337, 337, 338, 
    341, 338, 338, 338, 336, 337, 336, 338, 334, 324, 271, 317, 338, 337, 339, 
    336, 336, 338, 339, 339, 341, 330, 332, 277, 256, 222, 284, 341, 338, 341, 
    322, 335, 339, 341, 344, 349, 289, 328, 272, 274, 252, 268, 340, 338, 342, 
    165, 173, 279, 332, 336, 342, 311, 338, 325, 333, 302, 253, 226, 220, 335, 
    256, 266, 312, 282, 289, 260, 232, 251, 273, 324, 283, 272, 267, 228, 327, 
    133, 128, 212, 239, 308, 147, 59, 113, 214, 322, 298, 262, 242, 246, 223, 
    0, 133, 143, 162, 260, 265, 261, 288, 218, 198, 168, 147, 152, 194, 214, 
    0, 293, 254, 279, 305, 319, 296, 281, 235, 230, 233, 230, 192, 179, 176, 
    119, 170, 172, 185, 188, 195, 202, 166, 167, 146, 127, 113, 91, 102, 122, 
    0, 0, 0, 0, 0, 0, 30, 44, 57, 47, 30, 33, 54, 100, 115, 
    0, 0, 2, 0, 0, 0, 0, 47, 15, 19, 44, 94, 119, 109, 119, 
    0, 0, 0, 0, 0, 0, 0, 191, 173, 145, 94, 55, 67, 103, 154, 
    13, 0, 0, 0, 0, 0, 0, 102, 39, 0, 12, 66, 100, 117, 177, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 36, 90, 93, 110, 142, 193, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    49, 76, 102, 103, 116, 125, 146, 138, 155, 155, 155, 167, 147, 154, 159, 
    71, 98, 134, 123, 147, 138, 149, 157, 158, 113, 160, 175, 151, 163, 165, 
    94, 110, 156, 144, 168, 149, 141, 155, 168, 62, 162, 183, 154, 175, 176, 
    108, 111, 153, 168, 173, 165, 151, 117, 71, 38, 46, 79, 184, 174, 189, 
    79, 76, 85, 116, 122, 129, 113, 77, 36, 28, 34, 58, 112, 98, 105, 
    35, 51, 35, 51, 50, 45, 42, 19, 37, 38, 76, 117, 55, 158, 38, 
    30, 24, 18, 44, 52, 27, 20, 12, 23, 42, 108, 141, 107, 109, 23, 
    16, 25, 34, 38, 50, 56, 57, 50, 74, 54, 115, 136, 114, 22, 52, 
    16, 34, 52, 56, 45, 53, 59, 62, 80, 60, 100, 103, 96, 87, 123, 
    0, 29, 43, 36, 43, 55, 69, 74, 94, 96, 91, 83, 81, 60, 64, 
    39, 25, 31, 33, 58, 80, 35, 13, 64, 93, 75, 52, 44, 37, 33, 
    57, 35, 4, 3, 14, 67, 46, 35, 46, 47, 41, 32, 16, 16, 9, 
    51, 40, 31, 26, 32, 35, 27, 34, 35, 31, 21, 30, 8, 9, 7, 
    9, 13, 16, 24, 30, 34, 27, 20, 40, 6, 17, 11, 7, 10, 11, 
    15, 18, 17, 19, 20, 21, 22, 18, 60, 0, 11, 6, 9, 15, 0, 
    
    -- channel=129
    91, 48, 79, 91, 104, 98, 104, 114, 95, 114, 109, 102, 101, 109, 100, 
    93, 54, 83, 96, 104, 102, 118, 117, 98, 132, 86, 108, 109, 121, 102, 
    100, 56, 81, 95, 100, 99, 122, 112, 101, 141, 66, 109, 117, 118, 104, 
    127, 81, 134, 138, 133, 114, 117, 103, 100, 111, 44, 80, 128, 138, 121, 
    124, 92, 109, 112, 134, 130, 116, 122, 81, 65, 51, 43, 39, 104, 85, 
    28, 23, 59, 25, 38, 34, 58, 73, 50, 42, 4, 39, 64, 100, 60, 
    47, 49, 65, 32, 56, 51, 46, 30, 10, 24, 32, 90, 125, 94, 100, 
    43, 41, 46, 42, 63, 63, 66, 76, 90, 106, 80, 92, 96, 66, 20, 
    89, 90, 69, 86, 97, 91, 68, 55, 52, 71, 38, 71, 84, 91, 104, 
    49, 43, 61, 79, 60, 48, 65, 90, 74, 77, 81, 110, 104, 103, 74, 
    59, 59, 74, 95, 93, 72, 84, 64, 21, 87, 99, 91, 67, 49, 64, 
    40, 61, 76, 47, 33, 53, 114, 69, 40, 57, 55, 38, 47, 39, 46, 
    57, 90, 102, 72, 59, 58, 58, 44, 49, 48, 39, 30, 55, 36, 29, 
    52, 52, 39, 33, 36, 35, 32, 34, 11, 34, 40, 40, 35, 27, 35, 
    34, 20, 13, 12, 14, 14, 20, 42, 17, 49, 40, 42, 29, 27, 55, 
    
    -- channel=130
    265, 265, 316, 318, 337, 332, 342, 337, 342, 350, 330, 351, 343, 354, 354, 
    262, 259, 313, 309, 328, 317, 326, 331, 337, 280, 269, 355, 341, 348, 354, 
    263, 247, 303, 307, 315, 306, 298, 269, 285, 216, 232, 302, 311, 319, 338, 
    249, 245, 286, 301, 300, 302, 280, 257, 160, 102, 127, 85, 177, 259, 267, 
    121, 128, 129, 146, 157, 168, 176, 156, 148, 146, 138, 177, 220, 217, 147, 
    143, 147, 154, 159, 206, 180, 196, 154, 147, 148, 205, 304, 234, 227, 149, 
    156, 132, 122, 172, 199, 213, 221, 219, 223, 218, 255, 267, 236, 185, 99, 
    199, 221, 257, 284, 278, 269, 256, 236, 223, 175, 178, 230, 245, 187, 220, 
    172, 158, 199, 245, 236, 206, 187, 191, 219, 225, 256, 250, 231, 209, 195, 
    175, 216, 236, 210, 204, 221, 225, 189, 173, 221, 239, 215, 156, 108, 101, 
    191, 205, 198, 167, 160, 185, 168, 107, 136, 165, 141, 106, 79, 66, 69, 
    168, 176, 153, 117, 144, 179, 139, 127, 124, 107, 73, 63, 64, 53, 39, 
    129, 120, 96, 99, 86, 77, 91, 93, 71, 66, 54, 66, 53, 49, 48, 
    45, 37, 41, 54, 57, 51, 56, 50, 85, 77, 55, 57, 44, 52, 54, 
    44, 48, 45, 51, 56, 61, 55, 42, 79, 43, 56, 54, 46, 54, 26, 
    
    -- channel=131
    122, 113, 189, 187, 206, 193, 210, 200, 210, 222, 194, 218, 201, 221, 212, 
    125, 111, 187, 175, 201, 179, 197, 202, 201, 162, 143, 221, 199, 219, 213, 
    122, 91, 172, 162, 189, 161, 166, 144, 160, 67, 127, 184, 176, 192, 204, 
    98, 78, 149, 151, 153, 152, 128, 108, 30, 0, 0, 0, 97, 139, 132, 
    0, 0, 0, 23, 27, 39, 35, 17, 0, 0, 0, 0, 38, 57, 6, 
    0, 0, 0, 0, 17, 0, 26, 0, 0, 0, 16, 110, 38, 72, 0, 
    0, 0, 0, 1, 45, 37, 49, 26, 36, 45, 103, 121, 53, 19, 0, 
    12, 22, 49, 90, 106, 109, 107, 92, 86, 37, 42, 78, 70, 0, 0, 
    27, 9, 54, 104, 100, 78, 64, 53, 68, 37, 74, 74, 64, 40, 38, 
    0, 44, 74, 65, 53, 74, 81, 56, 30, 75, 83, 59, 10, 0, 0, 
    40, 53, 54, 23, 34, 53, 32, 0, 0, 42, 4, 0, 0, 0, 0, 
    35, 31, 4, 0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=132
    148, 135, 161, 170, 175, 176, 186, 187, 184, 192, 187, 193, 192, 194, 187, 
    156, 142, 167, 177, 181, 178, 180, 179, 184, 190, 147, 187, 193, 192, 188, 
    158, 138, 168, 178, 186, 174, 178, 156, 165, 160, 130, 171, 190, 184, 181, 
    142, 126, 150, 148, 165, 161, 158, 163, 129, 72, 89, 96, 106, 158, 153, 
    75, 85, 85, 95, 99, 105, 104, 108, 84, 84, 75, 79, 112, 130, 103, 
    63, 82, 91, 69, 96, 99, 101, 88, 87, 89, 93, 140, 157, 104, 92, 
    78, 82, 62, 76, 95, 105, 104, 101, 115, 119, 138, 149, 121, 114, 76, 
    86, 95, 93, 115, 124, 134, 139, 140, 125, 128, 103, 122, 128, 102, 94, 
    92, 83, 88, 114, 125, 125, 127, 124, 125, 118, 126, 132, 126, 123, 110, 
    74, 90, 112, 113, 108, 127, 134, 130, 111, 126, 128, 125, 110, 87, 70, 
    89, 107, 110, 101, 97, 104, 125, 74, 84, 114, 104, 85, 78, 59, 59, 
    83, 100, 102, 68, 71, 101, 90, 78, 83, 80, 78, 63, 54, 46, 29, 
    72, 82, 66, 65, 70, 62, 57, 70, 66, 57, 54, 51, 39, 29, 28, 
    36, 30, 38, 42, 51, 53, 50, 53, 46, 66, 37, 35, 29, 30, 34, 
    28, 29, 37, 41, 43, 49, 51, 45, 43, 49, 30, 23, 28, 29, 29, 
    
    -- channel=133
    91, 29, 35, 59, 54, 57, 51, 74, 38, 54, 64, 48, 71, 59, 51, 
    86, 27, 23, 63, 42, 57, 46, 46, 43, 100, 0, 32, 73, 55, 41, 
    81, 26, 11, 58, 36, 53, 60, 23, 16, 151, 0, 6, 67, 38, 27, 
    66, 18, 11, 15, 36, 30, 61, 62, 62, 65, 0, 0, 0, 12, 2, 
    8, 3, 5, 0, 0, 0, 15, 61, 55, 39, 18, 11, 0, 31, 0, 
    0, 10, 47, 4, 28, 37, 31, 61, 32, 39, 0, 14, 98, 0, 97, 
    9, 30, 38, 0, 14, 61, 57, 68, 56, 46, 0, 13, 91, 21, 95, 
    45, 46, 43, 37, 46, 57, 63, 64, 40, 72, 0, 1, 41, 128, 31, 
    42, 29, 0, 30, 59, 51, 46, 53, 32, 82, 6, 30, 39, 51, 14, 
    69, 17, 31, 45, 42, 47, 46, 46, 19, 28, 33, 54, 43, 42, 2, 
    9, 47, 45, 55, 11, 3, 78, 61, 0, 7, 33, 42, 34, 23, 13, 
    0, 36, 75, 41, 26, 0, 62, 38, 6, 21, 31, 20, 23, 9, 15, 
    0, 20, 36, 15, 7, 7, 20, 13, 12, 8, 21, 0, 28, 2, 3, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 39, 4, 5, 7, 0, 0, 
    0, 0, 0, 0, 0, 2, 2, 8, 0, 61, 0, 2, 0, 0, 22, 
    
    -- channel=134
    109, 130, 144, 143, 149, 152, 159, 153, 166, 163, 158, 167, 163, 166, 170, 
    116, 134, 151, 144, 154, 151, 153, 155, 164, 131, 152, 174, 162, 163, 172, 
    118, 135, 155, 149, 156, 151, 142, 142, 149, 92, 141, 157, 151, 157, 169, 
    112, 127, 136, 143, 145, 148, 135, 123, 99, 68, 102, 93, 113, 134, 145, 
    76, 87, 91, 105, 101, 107, 105, 87, 75, 74, 80, 93, 134, 115, 106, 
    91, 93, 82, 101, 114, 106, 103, 76, 82, 82, 120, 147, 115, 123, 85, 
    88, 76, 70, 104, 109, 103, 106, 104, 114, 114, 140, 143, 107, 114, 50, 
    96, 103, 111, 127, 123, 122, 116, 106, 103, 82, 111, 127, 127, 94, 116, 
    76, 79, 105, 109, 102, 96, 98, 102, 116, 103, 139, 133, 122, 104, 110, 
    82, 100, 110, 101, 99, 107, 107, 93, 99, 115, 122, 103, 86, 69, 78, 
    91, 97, 91, 74, 82, 98, 84, 69, 99, 94, 82, 68, 59, 59, 56, 
    97, 87, 72, 70, 84, 102, 60, 66, 83, 73, 58, 61, 52, 51, 43, 
    77, 63, 46, 55, 61, 61, 59, 63, 58, 58, 48, 59, 44, 48, 50, 
    45, 40, 45, 51, 52, 55, 58, 52, 68, 57, 51, 50, 46, 52, 49, 
    48, 53, 54, 57, 57, 58, 55, 46, 74, 38, 51, 47, 48, 54, 35, 
    
    -- channel=135
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 7, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 71, 0, 0, 4, 0, 0, 
    14, 0, 0, 0, 0, 0, 4, 15, 25, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 18, 6, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 1, 0, 15, 0, 0, 0, 0, 49, 0, 76, 
    0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 18, 78, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 25, 0, 0, 0, 70, 0, 
    6, 0, 0, 0, 1, 0, 0, 0, 0, 16, 0, 0, 0, 19, 0, 
    5, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 12, 16, 20, 0, 
    0, 0, 0, 13, 0, 0, 20, 22, 0, 0, 4, 11, 19, 9, 9, 
    0, 0, 15, 2, 0, 0, 26, 11, 0, 0, 18, 0, 11, 3, 11, 
    0, 0, 9, 0, 0, 0, 2, 0, 4, 0, 10, 0, 17, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 3, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 44, 0, 0, 0, 0, 24, 
    
    -- channel=136
    471, 417, 519, 542, 565, 563, 592, 599, 585, 613, 595, 612, 606, 617, 601, 
    486, 429, 528, 549, 572, 555, 567, 582, 582, 562, 471, 602, 607, 614, 595, 
    493, 417, 521, 550, 574, 544, 549, 492, 520, 477, 391, 546, 581, 577, 577, 
    452, 382, 470, 488, 524, 511, 515, 476, 344, 241, 213, 216, 355, 492, 476, 
    235, 226, 253, 274, 304, 319, 331, 342, 264, 247, 220, 255, 318, 366, 275, 
    190, 233, 262, 217, 298, 294, 306, 279, 253, 260, 287, 441, 403, 372, 268, 
    227, 215, 194, 218, 303, 330, 333, 323, 339, 350, 390, 449, 432, 333, 192, 
    283, 306, 333, 376, 410, 430, 439, 417, 396, 360, 306, 383, 405, 307, 276, 
    283, 259, 284, 379, 401, 383, 373, 372, 380, 389, 380, 399, 387, 368, 352, 
    246, 296, 353, 344, 341, 387, 403, 377, 336, 391, 395, 384, 318, 243, 188, 
    289, 332, 335, 309, 290, 328, 348, 210, 216, 329, 298, 245, 198, 152, 131, 
    244, 302, 290, 196, 212, 286, 291, 224, 210, 218, 195, 153, 126, 92, 61, 
    206, 235, 210, 176, 166, 159, 162, 177, 158, 138, 125, 111, 93, 58, 55, 
    62, 59, 78, 93, 115, 114, 109, 113, 124, 148, 83, 70, 57, 57, 61, 
    49, 49, 66, 75, 91, 104, 105, 89, 94, 113, 58, 45, 50, 58, 40, 
    
    -- channel=137
    557, 525, 540, 503, 468, 411, 374, 352, 355, 354, 318, 319, 329, 335, 321, 
    476, 436, 432, 390, 361, 324, 320, 324, 324, 321, 303, 297, 297, 303, 295, 
    387, 354, 332, 283, 265, 267, 269, 275, 299, 295, 350, 315, 269, 245, 266, 
    289, 269, 223, 181, 151, 189, 203, 256, 301, 329, 343, 279, 269, 198, 152, 
    276, 258, 238, 213, 176, 194, 256, 333, 400, 421, 409, 313, 221, 155, 163, 
    373, 353, 346, 323, 348, 374, 460, 469, 417, 399, 372, 284, 173, 144, 204, 
    441, 381, 375, 423, 458, 482, 518, 499, 472, 438, 342, 222, 168, 144, 179, 
    496, 449, 480, 530, 543, 549, 558, 529, 486, 374, 259, 191, 206, 181, 179, 
    549, 489, 516, 567, 579, 561, 522, 452, 402, 335, 282, 259, 275, 257, 198, 
    518, 544, 549, 527, 531, 512, 472, 427, 389, 368, 335, 313, 290, 252, 230, 
    585, 573, 552, 505, 491, 487, 435, 360, 366, 371, 342, 317, 298, 276, 241, 
    527, 531, 503, 448, 445, 458, 413, 374, 350, 337, 336, 318, 292, 275, 226, 
    468, 467, 449, 426, 392, 358, 347, 354, 341, 323, 307, 301, 270, 264, 251, 
    315, 316, 319, 327, 318, 307, 317, 305, 319, 306, 274, 260, 262, 262, 250, 
    224, 233, 259, 267, 288, 298, 307, 259, 284, 284, 252, 247, 261, 260, 185, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 1, 0, 8, 
    0, 2, 0, 0, 0, 8, 9, 3, 10, 0, 48, 18, 10, 5, 19, 
    0, 27, 17, 16, 21, 26, 14, 38, 41, 0, 64, 34, 20, 29, 34, 
    18, 55, 53, 61, 56, 55, 35, 34, 40, 24, 35, 78, 92, 59, 86, 
    63, 76, 66, 87, 88, 91, 69, 24, 11, 0, 9, 26, 56, 44, 102, 
    16, 29, 7, 28, 4, 8, 0, 0, 1, 0, 15, 9, 22, 62, 49, 
    0, 18, 13, 16, 0, 0, 0, 0, 0, 0, 19, 45, 32, 77, 74, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 68, 50, 25, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 33, 29, 38, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 7, 14, 21, 42, 53, 71, 
    0, 0, 0, 0, 0, 0, 0, 12, 44, 29, 34, 33, 48, 51, 62, 
    0, 0, 0, 0, 0, 5, 1, 21, 31, 31, 40, 36, 43, 54, 62, 
    15, 8, 5, 20, 26, 34, 34, 31, 42, 39, 44, 52, 48, 57, 58, 
    52, 55, 49, 49, 48, 53, 48, 42, 50, 26, 52, 59, 57, 57, 58, 
    68, 68, 58, 56, 50, 47, 47, 53, 78, 34, 60, 62, 59, 58, 66, 
    
    -- channel=139
    205, 152, 211, 232, 245, 247, 265, 277, 258, 276, 280, 275, 270, 280, 262, 
    219, 164, 225, 245, 262, 255, 267, 273, 261, 300, 196, 267, 277, 289, 263, 
    234, 168, 228, 250, 272, 252, 272, 250, 240, 286, 144, 264, 280, 280, 264, 
    240, 159, 242, 249, 275, 249, 263, 236, 213, 136, 98, 118, 175, 266, 249, 
    149, 131, 148, 162, 186, 192, 184, 192, 115, 114, 94, 67, 142, 199, 144, 
    51, 67, 123, 70, 101, 97, 117, 121, 104, 99, 61, 158, 189, 183, 143, 
    89, 86, 87, 69, 107, 118, 111, 98, 93, 108, 131, 217, 224, 185, 129, 
    90, 95, 95, 122, 151, 164, 171, 178, 181, 201, 152, 178, 190, 141, 60, 
    119, 143, 104, 152, 180, 182, 168, 151, 143, 164, 137, 176, 175, 165, 201, 
    77, 73, 143, 156, 128, 138, 167, 188, 164, 173, 175, 190, 186, 153, 104, 
    108, 129, 137, 152, 153, 148, 175, 104, 55, 164, 175, 142, 105, 77, 83, 
    88, 125, 142, 74, 63, 104, 167, 113, 95, 100, 101, 81, 54, 46, 33, 
    89, 130, 131, 98, 96, 86, 70, 74, 88, 74, 49, 47, 58, 23, 20, 
    44, 36, 38, 37, 58, 60, 51, 49, 22, 73, 40, 33, 23, 18, 21, 
    23, 15, 18, 19, 22, 31, 41, 49, 31, 62, 28, 20, 17, 18, 44, 
    
    -- channel=140
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 
    8, 13, 7, 4, 0, 0, 0, 0, 0, 0, 0, 1, 6, 4, 6, 
    8, 4, 1, 0, 0, 0, 0, 4, 0, 0, 6, 6, 8, 5, 13, 
    
    -- channel=141
    227, 238, 272, 267, 271, 266, 272, 258, 272, 277, 273, 272, 258, 266, 265, 
    226, 236, 273, 254, 270, 252, 261, 270, 267, 242, 273, 277, 257, 270, 270, 
    221, 226, 265, 240, 255, 241, 237, 262, 280, 186, 272, 311, 262, 264, 270, 
    218, 209, 245, 252, 236, 235, 222, 204, 206, 162, 171, 197, 289, 266, 268, 
    200, 187, 190, 218, 219, 229, 228, 202, 163, 157, 164, 134, 182, 161, 174, 
    134, 137, 138, 141, 133, 138, 177, 169, 168, 152, 166, 174, 104, 181, 92, 
    161, 143, 133, 169, 188, 166, 163, 145, 136, 148, 198, 221, 160, 166, 107, 
    156, 142, 147, 181, 210, 222, 228, 223, 237, 196, 217, 199, 182, 77, 49, 
    192, 214, 222, 237, 240, 251, 239, 202, 194, 154, 168, 180, 187, 168, 201, 
    136, 167, 214, 215, 210, 203, 214, 222, 236, 215, 200, 191, 196, 165, 151, 
    227, 203, 207, 205, 234, 250, 182, 136, 167, 216, 210, 174, 142, 124, 108, 
    214, 203, 170, 141, 137, 198, 190, 162, 159, 151, 146, 137, 93, 95, 69, 
    197, 206, 192, 173, 171, 156, 129, 137, 146, 138, 103, 113, 90, 79, 69, 
    109, 111, 109, 115, 124, 128, 121, 107, 110, 91, 94, 79, 75, 74, 71, 
    71, 73, 78, 80, 86, 92, 103, 93, 134, 77, 76, 68, 74, 80, 51, 
    
    -- channel=142
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 0, 3, 0, 0, 
    15, 0, 0, 0, 0, 0, 3, 17, 27, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 14, 1, 0, 0, 0, 1, 0, 
    0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0, 0, 48, 0, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 90, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 75, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 23, 0, 
    0, 0, 0, 3, 0, 0, 22, 18, 0, 0, 5, 17, 16, 7, 0, 
    0, 0, 19, 0, 0, 0, 23, 12, 0, 0, 11, 1, 2, 0, 5, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 3, 0, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 15, 
    
    -- channel=143
    404, 388, 491, 475, 502, 483, 515, 508, 517, 528, 490, 535, 505, 532, 518, 
    406, 388, 489, 463, 506, 465, 488, 514, 504, 420, 435, 534, 496, 525, 514, 
    403, 356, 472, 460, 495, 458, 452, 411, 454, 315, 408, 482, 470, 496, 504, 
    357, 322, 395, 422, 430, 438, 417, 385, 232, 186, 195, 156, 380, 408, 393, 
    196, 186, 206, 232, 244, 261, 278, 265, 228, 213, 209, 255, 275, 298, 217, 
    222, 221, 217, 224, 301, 262, 286, 230, 231, 249, 314, 436, 277, 389, 152, 
    225, 189, 170, 249, 305, 315, 321, 312, 329, 332, 380, 379, 341, 204, 93, 
    272, 299, 346, 367, 387, 396, 396, 351, 352, 258, 289, 350, 339, 212, 297, 
    249, 225, 301, 374, 346, 331, 332, 339, 347, 334, 357, 338, 327, 298, 277, 
    232, 324, 333, 298, 336, 363, 357, 299, 294, 357, 344, 307, 235, 168, 155, 
    318, 309, 302, 257, 255, 331, 274, 159, 231, 292, 231, 187, 155, 125, 100, 
    289, 286, 240, 182, 225, 290, 221, 188, 194, 193, 154, 134, 110, 83, 51, 
    215, 196, 170, 155, 149, 149, 160, 162, 130, 128, 117, 108, 70, 66, 61, 
    64, 71, 88, 105, 111, 108, 111, 107, 164, 100, 84, 69, 63, 70, 68, 
    58, 67, 81, 91, 106, 110, 103, 73, 139, 63, 66, 55, 61, 76, 6, 
    
    -- channel=144
    649, 613, 735, 755, 781, 770, 794, 783, 782, 814, 788, 810, 797, 811, 803, 
    650, 610, 729, 738, 763, 739, 755, 771, 774, 718, 663, 802, 794, 804, 797, 
    646, 582, 702, 716, 736, 709, 699, 660, 701, 584, 571, 742, 750, 748, 770, 
    596, 537, 636, 662, 676, 671, 652, 598, 465, 343, 326, 331, 530, 638, 637, 
    351, 343, 355, 392, 422, 448, 467, 452, 371, 346, 327, 344, 420, 451, 373, 
    274, 314, 334, 309, 398, 385, 429, 391, 353, 345, 398, 566, 459, 473, 320, 
    334, 312, 282, 350, 449, 474, 477, 457, 454, 459, 528, 591, 533, 405, 244, 
    411, 425, 474, 538, 587, 606, 610, 578, 562, 475, 437, 512, 526, 371, 324, 
    435, 413, 462, 578, 591, 563, 534, 508, 513, 490, 490, 516, 511, 474, 450, 
    376, 445, 517, 509, 506, 533, 543, 507, 477, 527, 534, 507, 423, 321, 261, 
    459, 492, 490, 452, 440, 494, 464, 301, 325, 450, 412, 329, 255, 191, 166, 
    395, 455, 410, 303, 320, 417, 402, 314, 297, 293, 250, 201, 163, 124, 75, 
    327, 357, 317, 276, 259, 244, 237, 238, 215, 194, 159, 154, 122, 82, 71, 
    120, 116, 121, 137, 155, 153, 154, 147, 175, 171, 115, 100, 78, 76, 77, 
    60, 63, 79, 94, 112, 126, 129, 105, 156, 131, 86, 72, 68, 81, 34, 
    
    -- channel=145
    310, 233, 312, 334, 354, 350, 374, 392, 361, 391, 378, 386, 385, 394, 371, 
    316, 243, 315, 348, 362, 350, 364, 374, 361, 384, 257, 370, 388, 396, 367, 
    327, 236, 310, 350, 366, 348, 364, 303, 319, 358, 201, 337, 380, 370, 358, 
    311, 225, 305, 314, 345, 328, 343, 333, 218, 134, 72, 65, 190, 326, 290, 
    143, 125, 139, 146, 181, 192, 201, 232, 175, 162, 124, 147, 174, 236, 152, 
    90, 125, 178, 101, 170, 168, 188, 179, 152, 164, 140, 273, 280, 230, 187, 
    123, 123, 111, 95, 152, 193, 187, 182, 188, 198, 210, 270, 305, 210, 163, 
    164, 183, 209, 229, 252, 267, 279, 270, 252, 247, 161, 227, 258, 209, 151, 
    179, 154, 138, 225, 255, 240, 220, 217, 220, 265, 222, 245, 238, 245, 226, 
    130, 170, 215, 202, 194, 232, 259, 256, 206, 241, 242, 258, 216, 164, 104, 
    167, 195, 207, 208, 180, 189, 229, 112, 83, 208, 196, 158, 132, 95, 87, 
    112, 176, 186, 94, 103, 149, 217, 157, 115, 125, 130, 85, 72, 50, 32, 
    113, 156, 152, 117, 88, 76, 93, 108, 101, 74, 75, 58, 62, 26, 25, 
    16, 16, 35, 46, 70, 64, 50, 55, 58, 98, 42, 35, 27, 23, 31, 
    23, 15, 23, 27, 42, 56, 58, 52, 27, 82, 25, 19, 20, 22, 28, 
    
    -- channel=146
    86, 94, 78, 68, 56, 54, 50, 46, 52, 43, 45, 43, 43, 42, 38, 
    79, 86, 71, 60, 56, 49, 41, 41, 47, 44, 39, 34, 37, 37, 34, 
    72, 80, 67, 53, 59, 47, 48, 52, 53, 47, 80, 52, 39, 41, 38, 
    54, 62, 43, 25, 36, 40, 51, 66, 58, 42, 82, 58, 41, 44, 41, 
    54, 63, 53, 51, 32, 38, 40, 61, 88, 116, 114, 108, 111, 54, 55, 
    116, 127, 115, 106, 99, 108, 100, 104, 119, 124, 127, 105, 86, 68, 101, 
    122, 106, 98, 103, 89, 89, 101, 106, 120, 120, 108, 63, 44, 88, 64, 
    113, 107, 107, 114, 98, 98, 102, 101, 91, 87, 72, 53, 53, 58, 93, 
    99, 90, 82, 79, 86, 90, 96, 95, 101, 91, 103, 74, 66, 75, 79, 
    95, 117, 112, 91, 93, 112, 111, 103, 93, 83, 74, 71, 82, 77, 82, 
    106, 107, 104, 99, 102, 92, 90, 87, 112, 99, 85, 87, 109, 120, 118, 
    127, 105, 100, 102, 112, 120, 97, 113, 117, 110, 128, 125, 122, 129, 122, 
    128, 111, 111, 119, 119, 109, 108, 135, 131, 121, 131, 139, 122, 132, 134, 
    121, 120, 134, 142, 144, 138, 130, 133, 139, 146, 127, 127, 132, 139, 137, 
    135, 140, 146, 143, 147, 151, 151, 137, 138, 124, 129, 125, 139, 138, 130, 
    
    -- channel=147
    201, 116, 143, 158, 155, 143, 137, 162, 122, 137, 139, 124, 141, 144, 122, 
    185, 98, 118, 143, 133, 134, 137, 138, 122, 197, 58, 110, 141, 142, 112, 
    173, 87, 92, 125, 117, 123, 151, 115, 90, 257, 8, 91, 137, 120, 102, 
    165, 79, 110, 104, 123, 108, 142, 144, 165, 165, 92, 65, 24, 108, 73, 
    119, 92, 104, 76, 97, 94, 110, 170, 148, 146, 118, 72, 61, 131, 67, 
    87, 77, 146, 83, 114, 113, 137, 165, 124, 125, 43, 82, 159, 79, 163, 
    121, 118, 141, 86, 116, 154, 157, 153, 132, 123, 51, 96, 166, 106, 166, 
    143, 138, 139, 147, 156, 161, 163, 168, 150, 179, 68, 75, 117, 176, 82, 
    162, 162, 112, 152, 182, 172, 149, 134, 107, 159, 78, 112, 120, 120, 116, 
    170, 116, 154, 169, 143, 132, 140, 151, 109, 119, 123, 149, 140, 138, 90, 
    132, 161, 159, 172, 142, 115, 183, 150, 42, 111, 138, 140, 116, 103, 109, 
    89, 145, 193, 136, 118, 87, 180, 135, 99, 109, 115, 108, 108, 98, 99, 
    97, 144, 163, 131, 117, 107, 110, 101, 109, 105, 99, 82, 123, 90, 90, 
    101, 94, 91, 81, 90, 89, 90, 95, 59, 129, 96, 96, 93, 84, 86, 
    84, 73, 74, 73, 77, 81, 87, 96, 37, 140, 91, 95, 85, 79, 116, 
    
    -- channel=148
    5, 83, 57, 26, 15, 3, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 61, 40, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 
    0, 43, 26, 0, 0, 0, 0, 0, 9, 0, 121, 15, 0, 0, 0, 
    0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 70, 55, 54, 0, 0, 
    3, 25, 3, 32, 0, 2, 0, 0, 9, 38, 57, 42, 68, 0, 20, 
    81, 74, 17, 58, 46, 53, 71, 25, 49, 37, 96, 40, 0, 0, 0, 
    87, 47, 28, 111, 75, 36, 55, 42, 58, 51, 90, 3, 0, 6, 0, 
    69, 52, 72, 99, 74, 60, 48, 40, 37, 0, 33, 3, 0, 0, 3, 
    73, 51, 101, 75, 53, 45, 36, 15, 43, 0, 58, 14, 0, 0, 0, 
    38, 114, 90, 57, 49, 56, 46, 27, 33, 19, 18, 0, 0, 0, 15, 
    96, 71, 65, 34, 74, 63, 0, 0, 105, 45, 4, 0, 5, 14, 25, 
    141, 62, 12, 41, 65, 121, 0, 24, 58, 28, 25, 24, 27, 41, 16, 
    114, 58, 21, 57, 54, 39, 33, 54, 49, 35, 31, 63, 13, 47, 45, 
    57, 50, 52, 68, 59, 54, 54, 38, 72, 30, 40, 46, 41, 56, 50, 
    40, 57, 58, 60, 59, 61, 61, 32, 108, 0, 53, 44, 56, 59, 5, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 17, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 18, 26, 33, 
    10, 10, 16, 14, 8, 7, 9, 11, 16, 12, 20, 23, 30, 30, 31, 
    30, 30, 28, 26, 25, 23, 19, 18, 3, 21, 26, 29, 31, 30, 28, 
    
    -- channel=150
    23, 17, 21, 24, 22, 21, 21, 19, 18, 21, 27, 19, 18, 18, 18, 
    20, 16, 20, 21, 20, 19, 19, 20, 19, 27, 13, 18, 19, 20, 15, 
    20, 16, 18, 16, 17, 15, 17, 24, 20, 24, 15, 33, 22, 20, 17, 
    24, 9, 23, 21, 21, 13, 18, 13, 25, 5, 3, 10, 28, 28, 26, 
    19, 18, 9, 15, 16, 20, 16, 21, 11, 13, 15, 0, 8, 0, 1, 
    0, 0, 6, 0, 0, 0, 7, 14, 11, 3, 0, 1, 0, 7, 2, 
    8, 6, 0, 2, 3, 4, 0, 0, 0, 0, 4, 13, 8, 6, 7, 
    4, 0, 0, 5, 13, 16, 19, 22, 27, 26, 15, 6, 4, 0, 0, 
    19, 29, 6, 19, 27, 33, 24, 11, 6, 3, 0, 2, 7, 7, 16, 
    0, 2, 21, 20, 9, 10, 17, 28, 29, 13, 10, 16, 26, 15, 4, 
    17, 15, 17, 27, 30, 24, 19, 5, 0, 23, 26, 12, 10, 3, 8, 
    14, 16, 17, 3, 0, 9, 28, 18, 8, 5, 13, 7, 0, 0, 0, 
    17, 29, 28, 22, 19, 8, 0, 7, 12, 6, 0, 1, 2, 0, 0, 
    3, 2, 1, 1, 5, 7, 1, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 17, 26, 20, 28, 34, 37, 27, 31, 28, 
    0, 0, 0, 7, 23, 30, 41, 38, 29, 41, 22, 41, 40, 46, 40, 
    8, 2, 26, 45, 58, 51, 59, 46, 42, 47, 20, 43, 59, 68, 55, 
    50, 44, 84, 95, 101, 87, 73, 69, 27, 0, 0, 9, 59, 96, 98, 
    39, 38, 38, 56, 74, 72, 44, 21, 0, 0, 0, 11, 47, 86, 69, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 35, 76, 86, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 60, 76, 77, 79, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 40, 66, 60, 42, 40, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 26, 37, 32, 52, 65, 
    0, 0, 0, 0, 0, 0, 0, 3, 3, 7, 15, 35, 43, 46, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 22, 18, 28, 25, 47, 
    0, 0, 0, 0, 0, 0, 5, 9, 2, 5, 15, 8, 17, 25, 34, 
    0, 0, 0, 0, 0, 0, 0, 5, 13, 9, 17, 19, 26, 22, 23, 
    9, 8, 8, 9, 18, 19, 7, 11, 4, 13, 22, 26, 23, 23, 33, 
    38, 31, 22, 18, 13, 15, 14, 34, 22, 17, 28, 28, 24, 23, 53, 
    
    -- channel=152
    245, 193, 242, 268, 276, 280, 293, 306, 286, 305, 307, 303, 307, 309, 292, 
    263, 206, 253, 283, 287, 289, 297, 294, 289, 349, 240, 293, 315, 314, 295, 
    269, 207, 251, 283, 294, 283, 300, 273, 269, 335, 177, 271, 315, 302, 288, 
    258, 191, 249, 253, 284, 264, 279, 264, 271, 212, 175, 220, 196, 271, 257, 
    184, 172, 194, 195, 219, 221, 220, 232, 152, 137, 116, 90, 139, 235, 202, 
    79, 94, 140, 97, 130, 139, 146, 156, 132, 131, 83, 147, 236, 162, 175, 
    111, 131, 126, 104, 155, 168, 160, 145, 145, 152, 157, 237, 234, 202, 171, 
    117, 121, 100, 131, 170, 196, 207, 217, 205, 239, 179, 201, 215, 189, 100, 
    156, 167, 153, 186, 217, 221, 223, 208, 184, 185, 148, 199, 205, 195, 199, 
    137, 101, 155, 197, 183, 182, 195, 215, 185, 200, 204, 218, 209, 190, 142, 
    133, 169, 179, 180, 176, 177, 231, 169, 116, 188, 204, 186, 144, 107, 100, 
    114, 170, 196, 134, 113, 136, 182, 127, 128, 145, 138, 115, 96, 77, 60, 
    105, 152, 147, 116, 132, 135, 108, 103, 112, 109, 89, 74, 81, 46, 40, 
    83, 76, 71, 62, 77, 84, 87, 89, 46, 100, 64, 57, 47, 38, 43, 
    41, 35, 47, 50, 52, 55, 67, 71, 48, 101, 45, 40, 37, 35, 61, 
    
    -- channel=153
    150, 162, 206, 207, 230, 229, 241, 232, 242, 252, 233, 251, 239, 250, 259, 
    149, 166, 213, 206, 227, 219, 234, 240, 240, 167, 203, 266, 239, 252, 258, 
    162, 165, 215, 211, 222, 214, 206, 192, 208, 97, 193, 228, 213, 232, 254, 
    174, 186, 232, 247, 234, 232, 202, 175, 65, 31, 39, 18, 176, 206, 214, 
    83, 82, 82, 112, 124, 133, 125, 92, 83, 75, 76, 131, 156, 129, 103, 
    83, 95, 82, 93, 134, 108, 120, 78, 74, 73, 140, 234, 125, 205, 75, 
    87, 63, 57, 103, 118, 116, 120, 116, 115, 120, 181, 191, 182, 134, 31, 
    120, 138, 191, 194, 186, 165, 151, 131, 140, 85, 123, 183, 182, 98, 147, 
    106, 81, 117, 160, 142, 107, 79, 90, 136, 144, 188, 172, 158, 151, 142, 
    75, 155, 147, 109, 104, 125, 136, 110, 106, 142, 163, 147, 95, 52, 54, 
    108, 107, 108, 94, 92, 105, 67, 22, 71, 108, 73, 38, 27, 17, 31, 
    95, 85, 49, 34, 67, 117, 83, 67, 52, 41, 15, 0, 16, 7, 5, 
    77, 60, 42, 43, 14, 9, 41, 38, 17, 5, 6, 18, 9, 12, 14, 
    0, 0, 0, 11, 12, 2, 0, 0, 43, 12, 13, 19, 7, 15, 18, 
    10, 9, 0, 3, 9, 12, 2, 2, 40, 0, 25, 22, 10, 21, 0, 
    
    -- channel=154
    0, 27, 28, 0, 3, 0, 6, 0, 25, 6, 0, 11, 0, 0, 13, 
    0, 26, 39, 0, 10, 0, 6, 9, 18, 0, 66, 35, 0, 1, 18, 
    0, 21, 43, 0, 11, 0, 0, 30, 39, 0, 141, 56, 0, 9, 33, 
    0, 19, 34, 28, 3, 13, 0, 0, 0, 0, 44, 55, 139, 25, 46, 
    20, 28, 28, 71, 40, 50, 29, 0, 0, 0, 8, 5, 56, 0, 40, 
    35, 20, 0, 28, 17, 2, 8, 0, 0, 0, 50, 32, 0, 71, 0, 
    28, 0, 0, 64, 39, 0, 0, 0, 0, 0, 64, 27, 0, 6, 0, 
    0, 0, 11, 21, 11, 0, 0, 0, 0, 0, 57, 46, 0, 0, 0, 
    0, 6, 57, 29, 0, 0, 0, 0, 12, 0, 40, 8, 0, 0, 16, 
    0, 41, 20, 0, 0, 0, 0, 0, 14, 9, 7, 0, 0, 0, 6, 
    32, 0, 0, 0, 25, 35, 0, 0, 62, 30, 0, 0, 0, 0, 0, 
    90, 0, 0, 0, 8, 72, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    57, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    7, 7, 0, 12, 3, 3, 4, 0, 26, 0, 0, 0, 0, 1, 0, 
    0, 8, 4, 5, 2, 0, 0, 0, 73, 0, 6, 0, 1, 10, 0, 
    
    -- channel=155
    278, 243, 334, 353, 389, 394, 428, 436, 425, 449, 438, 455, 440, 456, 448, 
    297, 267, 361, 378, 414, 400, 418, 437, 427, 382, 333, 460, 447, 463, 449, 
    326, 272, 374, 402, 426, 404, 405, 359, 379, 316, 261, 414, 431, 442, 443, 
    334, 278, 377, 412, 430, 411, 398, 346, 195, 104, 67, 52, 262, 391, 390, 
    147, 136, 151, 183, 223, 236, 230, 212, 146, 124, 107, 160, 235, 267, 172, 
    89, 117, 150, 120, 184, 154, 170, 133, 125, 133, 174, 346, 275, 323, 167, 
    104, 92, 81, 105, 155, 176, 166, 163, 168, 186, 254, 334, 346, 234, 131, 
    145, 178, 222, 238, 255, 257, 254, 235, 241, 207, 206, 293, 310, 216, 196, 
    127, 130, 139, 220, 222, 203, 183, 193, 222, 264, 271, 286, 272, 259, 267, 
    90, 154, 205, 177, 171, 206, 236, 220, 207, 256, 267, 262, 205, 139, 102, 
    145, 158, 163, 160, 148, 184, 175, 71, 79, 195, 174, 122, 87, 59, 58, 
    103, 137, 119, 50, 76, 139, 169, 124, 95, 92, 70, 45, 26, 10, 0, 
    85, 107, 93, 70, 49, 37, 58, 66, 51, 36, 23, 22, 21, 0, 0, 
    0, 0, 0, 5, 23, 21, 10, 8, 41, 40, 11, 4, 0, 0, 0, 
    0, 0, 0, 0, 4, 15, 11, 10, 28, 15, 2, 0, 0, 0, 0, 
    
    -- channel=156
    423, 336, 410, 416, 424, 406, 414, 431, 398, 418, 404, 409, 414, 425, 401, 
    403, 317, 379, 394, 402, 379, 385, 405, 390, 402, 289, 391, 406, 414, 386, 
    386, 289, 346, 373, 375, 365, 376, 319, 331, 399, 223, 355, 389, 373, 366, 
    343, 250, 299, 311, 331, 324, 352, 338, 258, 222, 162, 99, 197, 313, 269, 
    186, 164, 178, 162, 188, 194, 230, 285, 263, 257, 228, 223, 214, 255, 149, 
    201, 207, 260, 205, 269, 254, 287, 290, 253, 263, 238, 335, 302, 258, 227, 
    233, 214, 213, 207, 264, 319, 323, 328, 320, 309, 267, 287, 334, 196, 197, 
    297, 308, 334, 356, 375, 383, 390, 365, 340, 307, 207, 242, 282, 286, 225, 
    284, 270, 254, 342, 362, 348, 328, 319, 296, 348, 278, 286, 286, 273, 249, 
    286, 293, 339, 317, 320, 338, 341, 312, 275, 309, 300, 298, 252, 204, 151, 
    307, 328, 319, 306, 264, 292, 317, 214, 158, 255, 248, 222, 189, 166, 141, 
    231, 293, 307, 220, 229, 230, 289, 241, 198, 200, 192, 176, 148, 127, 109, 
    204, 240, 241, 208, 180, 163, 178, 186, 172, 162, 152, 132, 144, 110, 111, 
    101, 101, 122, 128, 145, 140, 136, 140, 148, 178, 126, 113, 112, 108, 107, 
    99, 94, 107, 111, 128, 139, 139, 125, 97, 167, 105, 102, 103, 108, 94, 
    
    -- channel=157
    728, 707, 847, 843, 866, 840, 869, 848, 865, 887, 847, 880, 852, 882, 868, 
    716, 687, 829, 801, 842, 794, 818, 845, 846, 748, 724, 878, 840, 871, 858, 
    699, 641, 786, 764, 804, 758, 750, 722, 769, 580, 672, 832, 792, 809, 835, 
    636, 574, 690, 709, 716, 718, 693, 638, 483, 347, 370, 341, 614, 697, 687, 
    382, 365, 380, 433, 445, 482, 504, 494, 418, 410, 398, 393, 496, 467, 379, 
    354, 381, 390, 372, 469, 446, 516, 450, 423, 415, 491, 661, 451, 557, 317, 
    424, 354, 326, 437, 532, 540, 558, 527, 530, 539, 615, 645, 543, 429, 204, 
    494, 501, 574, 652, 693, 707, 707, 658, 648, 509, 493, 557, 559, 340, 356, 
    509, 488, 553, 678, 677, 648, 611, 573, 586, 536, 569, 570, 556, 502, 506, 
    428, 550, 632, 591, 584, 621, 631, 576, 549, 601, 594, 549, 460, 333, 284, 
    572, 584, 574, 521, 530, 589, 508, 316, 387, 527, 459, 357, 284, 226, 202, 
    522, 535, 464, 348, 385, 522, 454, 367, 357, 339, 294, 249, 193, 159, 93, 
    428, 432, 380, 340, 317, 288, 279, 295, 271, 240, 196, 204, 149, 119, 107, 
    156, 149, 165, 193, 211, 208, 205, 187, 241, 210, 155, 133, 112, 120, 116, 
    95, 105, 125, 140, 163, 181, 185, 142, 232, 139, 126, 102, 109, 128, 45, 
    
    -- channel=158
    61, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 
    64, 0, 0, 0, 0, 0, 0, 0, 0, 161, 0, 0, 0, 0, 0, 
    74, 0, 0, 0, 0, 0, 50, 0, 0, 372, 0, 0, 20, 0, 0, 
    84, 0, 0, 0, 7, 0, 58, 59, 114, 130, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 112, 40, 23, 0, 0, 0, 86, 0, 
    0, 0, 61, 0, 0, 0, 0, 49, 0, 0, 0, 0, 183, 0, 176, 
    0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 168, 5, 233, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 131, 0, 0, 0, 243, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 0, 0, 0, 16, 5, 
    22, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 47, 62, 100, 0, 
    0, 0, 0, 30, 0, 0, 123, 88, 0, 0, 38, 81, 51, 32, 42, 
    0, 0, 113, 0, 0, 0, 108, 29, 0, 0, 34, 27, 30, 11, 46, 
    0, 0, 59, 0, 0, 0, 0, 0, 0, 5, 12, 0, 76, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 77, 0, 1, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 25, 0, 144, 0, 0, 0, 0, 111, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 16, 19, 
    3, 3, 5, 5, 4, 3, 0, 0, 0, 0, 8, 12, 16, 19, 18, 
    23, 23, 17, 12, 8, 8, 7, 14, 7, 0, 18, 18, 21, 19, 33, 
    
    -- channel=160
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 9, 1, 9, 
    0, 0, 0, 0, 0, 7, 9, 4, 4, 16, 14, 14, 23, 15, 19, 
    0, 0, 0, 13, 12, 21, 22, 26, 15, 35, 0, 7, 28, 30, 24, 
    21, 19, 37, 57, 64, 47, 44, 13, 20, 24, 0, 26, 12, 42, 67, 
    28, 20, 34, 39, 63, 58, 39, 12, 0, 0, 0, 0, 0, 44, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 21, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 54, 62, 65, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 31, 38, 38, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 11, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 25, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=161
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=162
    0, 0, 18, 0, 6, 0, 4, 4, 10, 4, 0, 4, 0, 8, 0, 
    0, 0, 17, 0, 14, 0, 9, 16, 3, 0, 0, 10, 0, 10, 0, 
    0, 0, 11, 0, 17, 0, 11, 5, 0, 0, 22, 10, 0, 12, 1, 
    0, 0, 12, 4, 8, 2, 0, 4, 0, 0, 5, 0, 35, 17, 0, 
    0, 0, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 7, 16, 0, 
    14, 0, 2, 0, 18, 0, 7, 0, 0, 0, 0, 29, 0, 61, 0, 
    18, 0, 0, 17, 10, 0, 1, 0, 1, 5, 17, 6, 0, 0, 0, 
    0, 0, 10, 14, 10, 4, 0, 0, 3, 0, 10, 8, 0, 0, 10, 
    0, 1, 4, 11, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 7, 
    0, 15, 18, 1, 0, 1, 4, 0, 0, 8, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 10, 13, 0, 0, 0, 19, 0, 0, 0, 0, 4, 
    39, 0, 0, 0, 0, 27, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 2, 1, 0, 0, 1, 0, 15, 0, 3, 0, 0, 1, 0, 
    
    -- channel=163
    0, 0, 0, 3, 41, 53, 87, 97, 99, 106, 92, 119, 96, 115, 110, 
    0, 0, 50, 51, 95, 87, 112, 117, 106, 67, 78, 137, 109, 132, 123, 
    33, 17, 92, 103, 139, 113, 127, 98, 97, 29, 70, 97, 112, 149, 138, 
    72, 65, 141, 163, 178, 160, 138, 102, 0, 0, 0, 0, 100, 146, 150, 
    20, 10, 43, 70, 90, 87, 51, 11, 0, 0, 0, 38, 83, 139, 79, 
    0, 0, 0, 2, 31, 0, 0, 0, 0, 0, 16, 124, 99, 191, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 119, 130, 107, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 126, 113, 40, 138, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 38, 91, 89, 69, 72, 100, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 48, 52, 17, 11, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 13, 18, 27, 29, 
    11, 16, 15, 16, 14, 9, 3, 8, 7, 8, 18, 25, 28, 28, 32, 
    33, 30, 24, 21, 20, 18, 16, 24, 11, 15, 27, 32, 31, 26, 41, 
    
    -- channel=165
    260, 188, 264, 267, 276, 254, 262, 270, 249, 270, 255, 254, 250, 267, 245, 
    245, 172, 243, 241, 256, 230, 248, 264, 241, 257, 187, 248, 246, 268, 236, 
    231, 148, 211, 214, 228, 211, 233, 214, 216, 238, 143, 244, 240, 239, 226, 
    210, 123, 195, 201, 206, 191, 210, 178, 149, 143, 69, 71, 178, 214, 179, 
    128, 82, 111, 111, 133, 137, 150, 186, 131, 118, 100, 69, 71, 121, 60, 
    61, 56, 102, 58, 96, 92, 139, 153, 113, 106, 72, 130, 85, 142, 59, 
    105, 76, 92, 80, 144, 152, 160, 139, 118, 127, 112, 158, 179, 91, 49, 
    133, 125, 144, 169, 207, 218, 227, 212, 214, 180, 117, 127, 140, 71, 15, 
    173, 171, 161, 221, 238, 231, 204, 174, 149, 159, 103, 130, 144, 128, 143, 
    131, 139, 190, 194, 185, 179, 188, 187, 159, 174, 161, 169, 141, 105, 54, 
    182, 187, 188, 187, 179, 186, 176, 93, 48, 155, 148, 120, 70, 41, 25, 
    134, 168, 168, 95, 87, 127, 181, 102, 68, 83, 71, 50, 24, 3, 0, 
    113, 148, 155, 101, 83, 73, 62, 57, 56, 50, 24, 11, 18, 0, 0, 
    11, 13, 13, 14, 25, 23, 20, 19, 8, 27, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 3, 0, 23, 0, 0, 0, 0, 0, 
    
    -- channel=166
    352, 323, 431, 450, 483, 484, 518, 519, 519, 543, 527, 545, 522, 544, 532, 
    382, 344, 464, 465, 509, 486, 516, 530, 519, 486, 454, 553, 531, 557, 537, 
    404, 346, 470, 478, 518, 480, 493, 477, 488, 392, 381, 519, 517, 540, 533, 
    403, 335, 462, 491, 512, 485, 476, 394, 308, 242, 200, 258, 420, 489, 491, 
    262, 226, 276, 315, 348, 359, 343, 314, 193, 167, 153, 177, 274, 348, 277, 
    128, 144, 172, 160, 208, 194, 213, 190, 172, 166, 195, 332, 273, 380, 181, 
    160, 139, 145, 165, 250, 225, 227, 195, 197, 226, 307, 420, 381, 317, 134, 
    175, 189, 207, 246, 296, 315, 318, 303, 322, 291, 310, 370, 363, 193, 180, 
    204, 221, 256, 310, 315, 307, 297, 284, 295, 277, 291, 337, 333, 298, 349, 
    152, 185, 254, 273, 262, 272, 296, 299, 284, 330, 334, 329, 278, 222, 179, 
    216, 234, 244, 231, 253, 286, 258, 161, 172, 288, 266, 216, 142, 101, 91, 
    204, 225, 199, 131, 135, 233, 235, 148, 152, 170, 129, 97, 71, 42, 22, 
    166, 188, 173, 124, 134, 140, 115, 108, 101, 101, 61, 61, 45, 15, 1, 
    50, 47, 40, 47, 61, 66, 66, 61, 60, 60, 41, 26, 9, 8, 13, 
    8, 5, 11, 19, 26, 30, 38, 39, 76, 36, 19, 10, 2, 12, 4, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=168
    0, 0, 3, 6, 14, 19, 25, 27, 26, 30, 24, 31, 31, 32, 31, 
    0, 0, 8, 15, 21, 22, 23, 22, 27, 17, 0, 32, 33, 31, 34, 
    3, 0, 13, 22, 26, 25, 23, 3, 13, 0, 0, 12, 26, 23, 30, 
    4, 8, 18, 20, 25, 26, 19, 28, 0, 0, 0, 0, 0, 9, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 36, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 12, 8, 11, 0, 
    0, 0, 10, 17, 5, 1, 0, 0, 0, 0, 0, 2, 14, 2, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 24, 17, 2, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=169
    478, 438, 574, 579, 620, 608, 652, 651, 649, 676, 634, 680, 654, 682, 662, 
    487, 446, 582, 582, 631, 592, 623, 645, 640, 563, 499, 678, 651, 678, 660, 
    499, 421, 572, 585, 628, 584, 585, 513, 560, 428, 443, 602, 615, 630, 642, 
    461, 397, 520, 546, 571, 564, 542, 508, 286, 148, 153, 109, 381, 528, 505, 
    192, 189, 204, 248, 279, 305, 317, 303, 233, 220, 189, 257, 336, 367, 243, 
    183, 215, 240, 203, 317, 282, 314, 240, 229, 242, 309, 527, 390, 428, 203, 
    213, 177, 144, 224, 299, 328, 330, 318, 343, 351, 433, 475, 433, 296, 120, 
    280, 323, 388, 434, 454, 462, 459, 417, 401, 315, 299, 409, 424, 259, 306, 
    261, 228, 285, 405, 402, 368, 344, 347, 380, 393, 426, 423, 393, 368, 344, 
    205, 330, 378, 326, 334, 392, 412, 363, 322, 404, 410, 383, 284, 178, 135, 
    305, 323, 324, 282, 270, 332, 304, 123, 189, 321, 258, 177, 135, 85, 74, 
    252, 281, 239, 130, 181, 290, 251, 194, 176, 167, 130, 80, 58, 26, 0, 
    190, 194, 153, 133, 106, 85, 110, 133, 97, 72, 56, 58, 20, 0, 0, 
    0, 0, 7, 36, 59, 53, 44, 37, 98, 78, 20, 10, 0, 1, 6, 
    0, 0, 5, 17, 37, 53, 47, 15, 74, 15, 2, 0, 0, 6, 0, 
    
    -- channel=170
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=171
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 18, 0, 0, 78, 107, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 15, 134, 98, 77, 118, 120, 34, 37, 20, 
    70, 46, 113, 107, 76, 41, 30, 0, 226, 216, 140, 364, 328, 167, 191, 
    282, 226, 243, 292, 302, 301, 242, 179, 40, 4, 21, 0, 0, 28, 201, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 36, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 134, 127, 
    0, 0, 0, 0, 0, 0, 0, 0, 41, 99, 143, 59, 7, 0, 0, 
    56, 145, 72, 7, 44, 97, 68, 0, 0, 0, 0, 0, 1, 0, 123, 
    0, 0, 0, 40, 0, 0, 0, 81, 124, 3, 0, 53, 160, 191, 159, 
    0, 0, 0, 79, 173, 96, 37, 85, 31, 124, 190, 165, 106, 68, 88, 
    35, 25, 18, 23, 0, 23, 131, 42, 39, 66, 96, 70, 29, 46, 37, 
    102, 173, 186, 125, 147, 147, 55, 22, 103, 95, 27, 37, 54, 18, 0, 
    138, 137, 77, 50, 58, 81, 69, 44, 0, 0, 37, 29, 14, 0, 0, 
    10, 0, 0, 0, 0, 0, 1, 45, 62, 22, 21, 17, 3, 0, 57, 
    
    -- channel=172
    0, 0, 0, 0, 0, 20, 12, 26, 2, 16, 35, 17, 42, 20, 29, 
    10, 0, 0, 23, 0, 34, 15, 3, 14, 46, 0, 7, 52, 21, 32, 
    25, 19, 0, 39, 8, 36, 26, 1, 0, 89, 0, 0, 45, 15, 18, 
    39, 45, 21, 32, 40, 34, 41, 39, 28, 9, 0, 0, 0, 4, 22, 
    0, 2, 0, 0, 2, 0, 0, 0, 7, 0, 0, 14, 6, 36, 19, 
    0, 0, 11, 0, 0, 3, 0, 0, 0, 0, 0, 3, 111, 0, 97, 
    0, 3, 1, 0, 0, 0, 0, 3, 0, 0, 0, 18, 74, 58, 108, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 26, 0, 7, 42, 125, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 5, 26, 24, 45, 10, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 17, 25, 4, 
    0, 0, 0, 0, 0, 0, 5, 20, 0, 0, 0, 3, 1, 0, 2, 
    0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 2, 0, 0, 25, 
    
    -- channel=173
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=174
    0, 43, 43, 10, 13, 5, 11, 0, 28, 7, 0, 15, 0, 1, 14, 
    0, 36, 47, 0, 14, 0, 2, 6, 19, 0, 50, 31, 0, 0, 19, 
    0, 26, 47, 0, 10, 0, 0, 10, 28, 0, 124, 45, 0, 2, 29, 
    0, 20, 18, 14, 0, 8, 0, 0, 0, 0, 19, 0, 90, 2, 25, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 9, 19, 61, 0, 0, 
    40, 25, 0, 31, 22, 2, 13, 0, 0, 0, 77, 63, 0, 50, 0, 
    30, 0, 0, 65, 34, 0, 3, 0, 9, 12, 81, 19, 0, 0, 0, 
    11, 6, 35, 48, 29, 14, 0, 0, 1, 0, 38, 25, 0, 0, 6, 
    0, 0, 50, 30, 0, 0, 0, 0, 18, 0, 53, 5, 0, 0, 0, 
    0, 54, 34, 0, 4, 12, 4, 0, 8, 8, 4, 0, 0, 0, 0, 
    43, 5, 0, 0, 13, 34, 0, 0, 58, 14, 0, 0, 0, 0, 0, 
    91, 3, 0, 0, 10, 68, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 
    0, 6, 5, 6, 5, 4, 0, 0, 69, 0, 0, 0, 0, 7, 0, 
    
    -- channel=175
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    200, 219, 254, 238, 245, 235, 237, 222, 240, 239, 221, 238, 225, 234, 239, 
    192, 208, 244, 215, 232, 211, 217, 231, 231, 160, 239, 245, 217, 229, 237, 
    178, 189, 228, 202, 210, 200, 184, 194, 220, 100, 230, 236, 201, 214, 229, 
    153, 167, 175, 191, 173, 186, 171, 141, 100, 119, 126, 116, 219, 177, 183, 
    118, 107, 122, 134, 131, 134, 148, 127, 124, 113, 126, 147, 137, 115, 107, 
    138, 127, 98, 139, 149, 138, 152, 132, 130, 130, 187, 193, 72, 173, 46, 
    134, 108, 107, 156, 183, 168, 179, 172, 169, 167, 192, 173, 136, 88, 21, 
    161, 161, 181, 193, 207, 207, 206, 178, 186, 113, 162, 166, 150, 74, 122, 
    150, 144, 201, 215, 191, 184, 185, 181, 181, 150, 168, 153, 155, 129, 130, 
    153, 187, 183, 171, 196, 192, 177, 142, 161, 179, 168, 136, 106, 82, 91, 
    199, 181, 171, 142, 151, 195, 126, 99, 151, 145, 117, 102, 77, 72, 45, 
    185, 168, 126, 125, 140, 169, 112, 99, 109, 107, 76, 81, 61, 50, 37, 
    140, 118, 106, 97, 96, 103, 99, 90, 74, 81, 66, 68, 43, 49, 44, 
    56, 64, 65, 74, 68, 66, 73, 67, 102, 44, 58, 45, 46, 49, 43, 
    39, 45, 52, 57, 64, 63, 59, 44, 93, 34, 46, 42, 45, 55, 0, 
    
    -- channel=177
    37, 25, 49, 45, 62, 66, 85, 95, 88, 88, 83, 104, 95, 100, 97, 
    47, 42, 65, 69, 88, 79, 79, 94, 89, 43, 39, 98, 92, 98, 92, 
    68, 47, 83, 101, 112, 97, 91, 47, 60, 42, 32, 60, 85, 102, 96, 
    63, 52, 67, 86, 106, 106, 108, 95, 0, 0, 0, 0, 7, 68, 65, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 25, 19, 96, 82, 75, 3, 
    49, 63, 58, 54, 90, 57, 28, 6, 29, 58, 100, 185, 126, 150, 67, 
    17, 15, 5, 13, 10, 39, 37, 63, 86, 86, 95, 78, 126, 37, 28, 
    41, 77, 105, 76, 52, 43, 40, 20, 20, 8, 25, 80, 87, 108, 183, 
    0, 0, 0, 1, 0, 0, 0, 34, 60, 115, 121, 83, 65, 79, 58, 
    3, 53, 24, 0, 10, 50, 52, 15, 14, 56, 57, 47, 15, 0, 5, 
    0, 0, 0, 0, 0, 0, 6, 0, 10, 18, 0, 0, 19, 30, 30, 
    0, 0, 0, 0, 23, 11, 6, 29, 19, 18, 16, 15, 31, 26, 38, 
    0, 0, 0, 0, 0, 0, 19, 32, 6, 5, 36, 28, 27, 37, 47, 
    0, 0, 12, 24, 27, 19, 11, 24, 68, 42, 31, 34, 39, 47, 49, 
    51, 53, 50, 49, 55, 56, 40, 35, 33, 30, 38, 39, 42, 47, 39, 
    
    -- channel=178
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 88, 0, 0, 12, 0, 0, 
    41, 0, 0, 4, 0, 0, 14, 12, 0, 198, 0, 0, 28, 0, 0, 
    64, 0, 0, 0, 22, 0, 42, 15, 118, 128, 0, 60, 0, 10, 14, 
    65, 41, 46, 12, 48, 40, 42, 90, 43, 16, 0, 0, 0, 19, 18, 
    0, 0, 11, 0, 0, 0, 0, 34, 0, 0, 0, 0, 47, 0, 127, 
    0, 6, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 52, 182, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 93, 0, 0, 6, 115, 0, 
    4, 41, 0, 0, 9, 29, 23, 5, 0, 10, 0, 0, 0, 17, 30, 
    10, 0, 0, 10, 0, 0, 0, 32, 18, 0, 0, 33, 75, 102, 39, 
    0, 0, 0, 43, 14, 0, 67, 93, 0, 0, 69, 88, 58, 44, 35, 
    0, 0, 60, 30, 0, 0, 91, 35, 0, 20, 50, 41, 29, 23, 40, 
    0, 44, 83, 35, 38, 41, 20, 0, 32, 31, 25, 0, 58, 6, 2, 
    39, 37, 20, 0, 4, 13, 11, 20, 0, 37, 16, 13, 14, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 27, 0, 97, 0, 10, 0, 0, 69, 
    
    -- channel=179
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 4, 6, 4, 2, 39, 9, 7, 4, 7, 
    0, 19, 17, 23, 28, 26, 22, 32, 35, 20, 39, 24, 26, 32, 20, 
    24, 36, 31, 45, 52, 46, 46, 33, 35, 57, 39, 73, 76, 55, 71, 
    62, 63, 68, 70, 78, 73, 61, 40, 29, 17, 21, 49, 49, 65, 82, 
    36, 42, 29, 47, 16, 21, 0, 1, 24, 32, 35, 16, 41, 75, 57, 
    4, 30, 33, 12, 0, 0, 0, 0, 0, 0, 17, 41, 55, 67, 95, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 61, 62, 49, 54, 65, 
    0, 0, 0, 0, 0, 0, 0, 13, 13, 20, 25, 33, 35, 43, 64, 
    0, 0, 0, 0, 0, 0, 0, 8, 33, 23, 16, 25, 46, 69, 83, 
    0, 0, 0, 0, 0, 11, 4, 41, 52, 32, 42, 61, 73, 83, 75, 
    0, 0, 0, 19, 14, 3, 19, 37, 47, 58, 66, 74, 72, 77, 92, 
    16, 15, 27, 30, 48, 59, 56, 56, 60, 73, 79, 74, 75, 82, 82, 
    68, 77, 78, 74, 74, 80, 77, 79, 78, 57, 79, 77, 84, 82, 84, 
    94, 94, 90, 87, 83, 78, 78, 84, 87, 75, 76, 81, 83, 82, 93, 
    
    -- channel=180
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=181
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 192, 0, 0, 11, 0, 0, 
    38, 0, 0, 0, 0, 0, 27, 0, 37, 107, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 41, 27, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 0, 106, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 0, 208, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 2, 205, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 10, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 60, 1, 
    0, 0, 0, 0, 0, 0, 24, 66, 0, 0, 0, 45, 23, 20, 0, 
    0, 0, 16, 0, 0, 0, 36, 6, 0, 0, 0, 7, 2, 0, 32, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 1, 0, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 0, 0, 0, 0, 46, 
    
    -- channel=182
    388, 296, 341, 316, 299, 250, 232, 239, 210, 219, 186, 189, 202, 217, 184, 
    323, 227, 251, 235, 222, 186, 191, 203, 187, 225, 108, 167, 178, 191, 158, 
    256, 160, 171, 161, 153, 149, 173, 126, 134, 236, 116, 151, 158, 134, 132, 
    176, 93, 93, 63, 64, 79, 115, 164, 155, 165, 140, 41, 52, 87, 7, 
    102, 78, 79, 42, 31, 38, 95, 197, 233, 255, 222, 156, 78, 81, 10, 
    203, 180, 221, 157, 222, 222, 289, 297, 243, 244, 182, 185, 134, 64, 104, 
    254, 204, 205, 216, 255, 308, 334, 330, 316, 283, 170, 94, 114, 25, 76, 
    315, 297, 325, 358, 363, 364, 370, 342, 295, 232, 83, 60, 100, 131, 111, 
    331, 280, 269, 345, 367, 346, 312, 271, 225, 239, 159, 142, 149, 136, 82, 
    324, 339, 355, 321, 319, 322, 299, 256, 197, 213, 188, 184, 147, 113, 72, 
    353, 361, 343, 311, 269, 269, 285, 187, 138, 195, 175, 161, 147, 127, 106, 
    279, 312, 330, 245, 252, 240, 252, 214, 173, 168, 172, 157, 139, 121, 89, 
    238, 255, 251, 226, 187, 157, 169, 183, 167, 153, 146, 126, 130, 110, 110, 
    118, 117, 136, 141, 147, 136, 139, 139, 140, 173, 118, 109, 112, 111, 104, 
    84, 86, 106, 111, 131, 142, 146, 113, 85, 151, 102, 98, 108, 107, 70, 
    
    -- channel=183
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=184
    0, 9, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 14, 0, 4, 0, 3, 0, 0, 0, 2, 5, 0, 4, 0, 3, 
    0, 20, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 6, 0, 0, 
    0, 32, 4, 0, 0, 0, 0, 3, 17, 0, 7, 24, 0, 0, 4, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 20, 
    0, 5, 0, 0, 0, 0, 0, 0, 2, 0, 3, 0, 30, 0, 9, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 17, 34, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 13, 0, 0, 0, 13, 0, 
    7, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 1, 10, 6, 0, 0, 0, 7, 7, 7, 
    0, 0, 3, 5, 0, 0, 2, 4, 12, 0, 5, 0, 5, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 10, 7, 0, 4, 0, 0, 5, 0, 
    0, 6, 0, 9, 5, 0, 0, 3, 6, 0, 1, 8, 0, 0, 0, 
    2, 0, 0, 0, 3, 2, 0, 0, 0, 8, 0, 1, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 1, 5, 0, 10, 0, 0, 0, 0, 1, 
    
    -- channel=185
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=186
    2, 33, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 
    0, 29, 0, 0, 0, 0, 0, 0, 11, 35, 54, 29, 37, 0, 1, 
    47, 54, 36, 35, 24, 26, 29, 20, 58, 62, 77, 70, 55, 4, 31, 
    88, 77, 58, 84, 57, 52, 55, 51, 64, 64, 80, 36, 0, 38, 43, 
    73, 66, 70, 83, 51, 46, 44, 52, 47, 42, 36, 4, 4, 15, 58, 
    65, 60, 65, 52, 36, 26, 21, 17, 28, 9, 45, 23, 15, 35, 54, 
    46, 58, 57, 36, 20, 26, 27, 29, 30, 28, 40, 21, 21, 20, 27, 
    60, 66, 50, 33, 42, 32, 26, 22, 50, 29, 22, 12, 30, 41, 66, 
    71, 45, 37, 42, 49, 54, 17, 54, 72, 36, 37, 45, 63, 83, 81, 
    78, 51, 36, 69, 74, 53, 42, 73, 73, 60, 67, 86, 82, 97, 101, 
    81, 63, 67, 82, 77, 73, 78, 78, 83, 86, 89, 98, 94, 109, 112, 
    97, 101, 101, 103, 97, 98, 97, 90, 111, 78, 103, 103, 109, 112, 106, 
    112, 115, 111, 108, 106, 104, 101, 96, 116, 83, 108, 111, 113, 114, 98, 
    
    -- channel=187
    375, 384, 486, 494, 527, 523, 550, 533, 551, 572, 540, 573, 551, 568, 569, 
    389, 392, 500, 491, 529, 505, 526, 539, 544, 450, 480, 582, 551, 568, 575, 
    396, 378, 493, 489, 515, 489, 474, 452, 497, 308, 420, 528, 517, 531, 557, 
    370, 362, 446, 477, 475, 476, 437, 380, 241, 157, 164, 184, 384, 446, 459, 
    190, 181, 207, 252, 274, 292, 295, 243, 174, 148, 143, 202, 273, 291, 235, 
    133, 155, 146, 163, 224, 208, 231, 176, 163, 159, 252, 385, 256, 328, 124, 
    156, 130, 110, 187, 263, 254, 259, 237, 245, 257, 358, 407, 328, 254, 63, 
    208, 230, 273, 321, 354, 363, 360, 330, 329, 241, 281, 354, 347, 166, 200, 
    213, 195, 280, 347, 336, 309, 293, 285, 314, 277, 326, 337, 324, 286, 283, 
    169, 249, 288, 277, 285, 307, 316, 279, 270, 328, 338, 302, 222, 144, 122, 
    250, 260, 262, 218, 229, 286, 224, 109, 186, 256, 211, 147, 83, 42, 20, 
    218, 233, 172, 114, 141, 245, 179, 122, 129, 126, 72, 40, 15, 0, 0, 
    156, 152, 112, 89, 81, 83, 80, 76, 50, 40, 11, 17, 0, 0, 0, 
    0, 0, 0, 4, 12, 9, 14, 3, 49, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 
    
    -- channel=188
    566, 522, 679, 684, 729, 717, 768, 763, 765, 795, 764, 800, 761, 796, 771, 
    589, 543, 702, 694, 756, 707, 746, 776, 757, 700, 653, 800, 764, 803, 776, 
    607, 523, 700, 699, 756, 699, 706, 664, 708, 556, 586, 769, 753, 773, 769, 
    581, 491, 648, 683, 703, 683, 662, 599, 437, 298, 282, 303, 601, 697, 672, 
    352, 324, 356, 414, 451, 473, 471, 443, 319, 292, 275, 298, 409, 475, 369, 
    235, 260, 298, 262, 346, 316, 371, 319, 306, 306, 352, 547, 417, 536, 236, 
    277, 248, 217, 292, 382, 381, 371, 342, 357, 387, 500, 592, 519, 385, 204, 
    312, 338, 375, 434, 496, 524, 534, 504, 517, 440, 450, 520, 508, 287, 279, 
    341, 351, 391, 498, 500, 500, 487, 460, 461, 443, 463, 490, 484, 445, 468, 
    246, 348, 441, 426, 433, 465, 496, 479, 463, 513, 498, 479, 413, 311, 256, 
    404, 399, 410, 385, 404, 478, 415, 226, 280, 451, 403, 314, 243, 179, 155, 
    356, 381, 334, 214, 239, 378, 367, 280, 269, 270, 234, 190, 127, 99, 45, 
    295, 322, 286, 239, 234, 213, 193, 212, 197, 183, 134, 133, 89, 51, 38, 
    80, 80, 95, 114, 144, 148, 136, 126, 151, 128, 91, 63, 46, 47, 53, 
    42, 42, 60, 71, 89, 104, 112, 92, 156, 80, 53, 33, 39, 56, 7, 
    
    -- channel=189
    329, 259, 360, 392, 419, 425, 462, 480, 456, 488, 483, 490, 481, 493, 471, 
    363, 291, 392, 424, 453, 443, 465, 477, 462, 495, 380, 484, 492, 506, 472, 
    389, 298, 403, 443, 475, 447, 466, 425, 431, 446, 293, 453, 491, 493, 473, 
    384, 281, 398, 422, 465, 434, 447, 397, 325, 241, 165, 225, 343, 448, 426, 
    236, 206, 248, 270, 313, 320, 311, 317, 190, 158, 131, 134, 212, 326, 261, 
    88, 119, 174, 115, 179, 175, 188, 182, 153, 159, 128, 273, 305, 322, 212, 
    119, 129, 126, 107, 190, 201, 187, 165, 171, 198, 241, 366, 378, 285, 187, 
    135, 151, 155, 181, 236, 268, 284, 281, 286, 298, 256, 321, 331, 235, 150, 
    174, 183, 175, 246, 276, 279, 276, 268, 257, 273, 238, 298, 302, 287, 308, 
    118, 130, 201, 230, 220, 241, 271, 289, 261, 295, 294, 312, 281, 233, 168, 
    161, 195, 212, 218, 214, 237, 274, 163, 124, 266, 263, 222, 167, 115, 103, 
    130, 193, 205, 115, 107, 173, 237, 150, 137, 165, 154, 112, 82, 51, 32, 
    119, 173, 168, 115, 120, 126, 110, 107, 113, 101, 78, 55, 60, 13, 6, 
    37, 36, 41, 40, 65, 73, 67, 69, 44, 82, 40, 26, 14, 4, 11, 
    10, 2, 14, 19, 29, 36, 46, 51, 39, 76, 13, 3, 1, 4, 25, 
    
    -- channel=190
    279, 206, 289, 312, 329, 322, 338, 351, 325, 353, 341, 344, 346, 357, 339, 
    283, 209, 286, 312, 324, 313, 325, 333, 323, 340, 232, 336, 349, 357, 332, 
    283, 198, 272, 305, 315, 299, 315, 266, 270, 307, 153, 290, 333, 325, 315, 
    260, 180, 259, 271, 295, 276, 289, 252, 179, 124, 68, 74, 153, 268, 246, 
    105, 81, 108, 112, 145, 147, 155, 182, 117, 102, 77, 85, 118, 192, 99, 
    40, 59, 109, 57, 119, 110, 132, 134, 98, 98, 86, 204, 211, 173, 114, 
    81, 73, 70, 60, 134, 162, 165, 154, 149, 159, 166, 231, 247, 150, 77, 
    125, 137, 152, 181, 215, 227, 235, 226, 211, 203, 130, 179, 203, 158, 97, 
    142, 129, 125, 201, 226, 208, 193, 185, 177, 203, 161, 191, 193, 181, 172, 
    117, 121, 175, 184, 168, 189, 202, 192, 149, 193, 199, 205, 155, 107, 51, 
    127, 167, 171, 161, 137, 149, 190, 90, 43, 148, 141, 107, 59, 21, 16, 
    81, 142, 155, 72, 70, 109, 154, 83, 59, 72, 51, 23, 10, 0, 0, 
    58, 100, 93, 54, 44, 39, 36, 35, 25, 16, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    
    -- channel=191
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=192
    112, 90, 56, 84, 98, 91, 90, 96, 91, 94, 95, 95, 109, 119, 122, 
    100, 90, 78, 63, 107, 115, 112, 119, 118, 121, 120, 130, 114, 112, 117, 
    97, 86, 78, 93, 95, 102, 99, 117, 107, 104, 109, 120, 132, 114, 114, 
    85, 83, 62, 73, 85, 83, 81, 85, 79, 74, 94, 83, 114, 105, 107, 
    80, 81, 80, 64, 77, 79, 78, 82, 81, 79, 91, 112, 94, 101, 100, 
    105, 87, 89, 95, 79, 80, 85, 85, 79, 85, 93, 94, 97, 100, 102, 
    122, 49, 28, 90, 134, 110, 95, 95, 97, 93, 100, 98, 100, 101, 104, 
    132, 102, 100, 38, 33, 127, 151, 115, 100, 98, 102, 98, 97, 94, 94, 
    139, 125, 120, 114, 0, 69, 96, 134, 148, 124, 110, 94, 95, 98, 96, 
    144, 128, 122, 105, 0, 51, 69, 70, 70, 60, 100, 139, 151, 129, 104, 
    141, 116, 119, 78, 46, 0, 16, 90, 60, 19, 39, 21, 107, 95, 102, 
    143, 117, 121, 122, 123, 98, 99, 107, 80, 69, 79, 71, 66, 58, 70, 
    68, 48, 44, 54, 62, 57, 52, 58, 49, 55, 53, 57, 59, 51, 53, 
    54, 55, 51, 60, 62, 55, 53, 60, 62, 57, 60, 58, 57, 61, 87, 
    51, 51, 51, 58, 58, 55, 50, 65, 58, 56, 57, 66, 76, 86, 86, 
    
    -- channel=193
    73, 101, 92, 101, 98, 99, 95, 90, 86, 89, 94, 93, 88, 102, 100, 
    75, 87, 112, 186, 214, 217, 211, 208, 219, 212, 205, 168, 132, 120, 111, 
    75, 84, 132, 204, 183, 175, 187, 183, 168, 172, 167, 161, 131, 110, 111, 
    77, 88, 143, 198, 171, 162, 161, 175, 175, 196, 180, 172, 133, 112, 108, 
    87, 88, 97, 125, 107, 105, 98, 112, 118, 113, 103, 96, 118, 103, 104, 
    90, 107, 112, 106, 84, 87, 95, 106, 104, 90, 89, 96, 106, 103, 98, 
    87, 86, 66, 116, 149, 123, 113, 118, 114, 115, 114, 115, 111, 115, 114, 
    88, 103, 99, 66, 59, 122, 137, 123, 121, 121, 111, 111, 108, 107, 103, 
    92, 106, 107, 115, 119, 63, 71, 141, 166, 148, 121, 118, 114, 108, 107, 
    96, 113, 113, 144, 154, 64, 69, 70, 55, 89, 122, 170, 156, 129, 118, 
    97, 119, 113, 119, 56, 13, 0, 2, 27, 4, 0, 0, 13, 65, 105, 
    142, 177, 173, 174, 173, 178, 141, 135, 164, 154, 142, 147, 137, 159, 156, 
    71, 98, 94, 87, 79, 82, 88, 99, 121, 117, 120, 122, 129, 138, 125, 
    65, 83, 83, 62, 55, 56, 57, 51, 48, 38, 36, 38, 36, 17, 0, 
    44, 41, 43, 37, 35, 29, 32, 21, 21, 20, 26, 25, 0, 0, 2, 
    
    -- channel=194
    274, 312, 278, 275, 295, 298, 291, 289, 296, 296, 297, 293, 308, 330, 326, 
    273, 290, 293, 323, 329, 323, 311, 329, 330, 323, 329, 327, 341, 324, 331, 
    264, 282, 282, 348, 348, 369, 362, 385, 380, 375, 370, 372, 351, 322, 330, 
    273, 284, 291, 379, 345, 346, 335, 367, 355, 346, 350, 344, 360, 308, 316, 
    289, 288, 287, 291, 268, 260, 261, 284, 278, 265, 274, 296, 343, 311, 316, 
    294, 276, 240, 301, 317, 317, 332, 337, 331, 314, 316, 327, 310, 315, 321, 
    303, 293, 220, 150, 207, 306, 330, 334, 330, 321, 318, 314, 311, 310, 315, 
    310, 323, 305, 291, 172, 174, 264, 327, 324, 315, 315, 314, 316, 313, 314, 
    314, 327, 325, 316, 171, 131, 134, 134, 200, 271, 316, 332, 319, 307, 312, 
    314, 327, 327, 296, 115, 75, 108, 141, 132, 89, 86, 125, 203, 279, 324, 
    313, 332, 326, 305, 303, 271, 207, 271, 315, 237, 264, 226, 282, 322, 312, 
    198, 207, 184, 174, 170, 149, 184, 231, 213, 215, 231, 234, 255, 241, 241, 
    176, 200, 191, 174, 162, 154, 163, 172, 150, 138, 134, 131, 132, 131, 126, 
    84, 93, 86, 81, 70, 73, 78, 79, 73, 67, 67, 71, 74, 75, 102, 
    87, 86, 85, 84, 77, 106, 106, 103, 101, 96, 82, 70, 89, 94, 44, 
    
    -- channel=195
    120, 150, 105, 107, 122, 129, 122, 118, 122, 125, 130, 124, 139, 167, 160, 
    121, 153, 150, 102, 132, 133, 114, 131, 135, 136, 126, 125, 173, 170, 170, 
    115, 140, 163, 86, 103, 99, 90, 102, 109, 122, 114, 128, 161, 172, 175, 
    116, 138, 150, 93, 105, 105, 91, 122, 118, 116, 118, 129, 133, 163, 166, 
    126, 141, 137, 115, 95, 94, 94, 115, 109, 94, 101, 141, 154, 165, 161, 
    143, 135, 104, 137, 138, 138, 151, 154, 143, 138, 144, 159, 160, 159, 167, 
    157, 106, 47, 39, 92, 152, 171, 175, 169, 162, 162, 159, 160, 163, 164, 
    171, 172, 134, 46, 0, 60, 134, 171, 168, 156, 157, 156, 160, 156, 159, 
    179, 182, 179, 151, 0, 0, 0, 40, 86, 126, 155, 168, 161, 157, 159, 
    179, 178, 179, 162, 0, 0, 0, 0, 0, 0, 0, 39, 86, 134, 161, 
    175, 175, 176, 122, 46, 0, 0, 41, 62, 0, 8, 0, 92, 136, 149, 
    91, 89, 74, 66, 63, 17, 32, 85, 77, 62, 80, 74, 97, 98, 92, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=196
    120, 137, 140, 131, 117, 138, 139, 133, 139, 137, 140, 136, 139, 154, 159, 
    125, 142, 145, 107, 86, 75, 84, 85, 88, 90, 89, 95, 131, 150, 155, 
    121, 143, 152, 79, 83, 82, 82, 72, 92, 104, 100, 113, 121, 156, 157, 
    123, 136, 126, 74, 78, 83, 90, 82, 83, 82, 77, 93, 101, 149, 151, 
    132, 138, 140, 131, 118, 120, 119, 120, 121, 119, 123, 124, 143, 153, 150, 
    142, 148, 132, 127, 143, 142, 140, 140, 139, 143, 144, 151, 149, 152, 154, 
    149, 139, 140, 96, 87, 127, 144, 149, 151, 151, 147, 148, 150, 150, 148, 
    153, 158, 149, 149, 103, 78, 110, 145, 151, 146, 148, 148, 148, 148, 148, 
    156, 165, 167, 152, 123, 64, 80, 84, 99, 120, 127, 146, 148, 150, 147, 
    155, 163, 163, 170, 90, 36, 46, 56, 72, 68, 59, 87, 103, 126, 140, 
    147, 157, 160, 141, 110, 115, 70, 78, 128, 96, 102, 95, 107, 138, 139, 
    112, 116, 115, 111, 107, 91, 92, 101, 96, 97, 98, 96, 103, 94, 98, 
    80, 70, 71, 72, 75, 68, 63, 64, 66, 59, 58, 58, 57, 57, 49, 
    59, 51, 49, 52, 58, 49, 49, 53, 55, 55, 52, 52, 50, 51, 84, 
    54, 50, 48, 53, 53, 52, 57, 60, 63, 61, 60, 59, 58, 115, 119, 
    
    -- channel=197
    3, 43, 86, 38, 26, 48, 54, 44, 51, 46, 49, 49, 35, 42, 49, 
    9, 35, 77, 86, 0, 0, 17, 0, 10, 5, 11, 5, 28, 52, 51, 
    10, 42, 52, 40, 41, 16, 30, 0, 30, 34, 19, 9, 15, 56, 51, 
    23, 41, 94, 51, 43, 46, 58, 41, 49, 67, 37, 47, 5, 52, 50, 
    45, 41, 56, 75, 38, 38, 38, 34, 44, 49, 30, 15, 54, 52, 55, 
    43, 59, 45, 37, 65, 61, 55, 62, 70, 61, 54, 46, 54, 55, 53, 
    33, 104, 95, 0, 0, 20, 50, 59, 61, 65, 52, 58, 54, 53, 50, 
    20, 61, 89, 146, 49, 0, 0, 40, 61, 64, 54, 59, 56, 60, 55, 
    17, 51, 60, 78, 210, 0, 0, 0, 0, 13, 26, 59, 59, 56, 54, 
    17, 51, 56, 73, 196, 0, 0, 0, 0, 0, 0, 0, 0, 12, 43, 
    11, 51, 54, 112, 112, 142, 28, 0, 79, 97, 51, 60, 0, 26, 36, 
    0, 16, 15, 8, 1, 45, 10, 0, 29, 42, 20, 39, 24, 31, 29, 
    20, 23, 29, 21, 13, 17, 9, 0, 15, 0, 0, 0, 0, 1, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 4, 0, 7, 3, 3, 0, 0, 0, 17, 
    
    -- channel=198
    142, 144, 128, 130, 138, 143, 141, 143, 145, 145, 144, 143, 151, 156, 153, 
    139, 135, 127, 122, 123, 114, 111, 118, 116, 117, 117, 126, 146, 147, 150, 
    132, 131, 128, 124, 139, 158, 151, 162, 165, 161, 161, 163, 147, 145, 150, 
    132, 131, 120, 149, 145, 142, 146, 157, 145, 136, 142, 147, 161, 140, 145, 
    132, 132, 129, 128, 127, 127, 126, 134, 126, 126, 135, 145, 152, 141, 141, 
    137, 123, 112, 129, 140, 140, 145, 145, 140, 138, 143, 147, 140, 144, 146, 
    147, 131, 110, 97, 96, 132, 143, 143, 141, 137, 139, 137, 139, 139, 141, 
    153, 145, 132, 118, 105, 103, 123, 143, 142, 138, 141, 140, 139, 140, 141, 
    154, 150, 148, 141, 58, 87, 103, 88, 94, 115, 139, 143, 140, 137, 138, 
    154, 153, 149, 128, 35, 66, 78, 86, 95, 81, 78, 70, 96, 125, 140, 
    156, 150, 149, 131, 128, 123, 125, 153, 147, 125, 135, 132, 159, 160, 145, 
    106, 91, 87, 84, 85, 60, 83, 112, 96, 88, 104, 96, 115, 105, 103, 
    98, 91, 87, 85, 83, 75, 77, 84, 66, 62, 61, 61, 59, 56, 55, 
    72, 69, 64, 68, 67, 67, 66, 68, 66, 67, 68, 69, 70, 76, 103, 
    71, 72, 71, 75, 71, 82, 78, 84, 82, 79, 73, 68, 89, 95, 75, 
    
    -- channel=199
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 10, 0, 2, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 58, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 153, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 140, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 33, 62, 0, 0, 3, 35, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    2, 0, 4, 2, 1, 4, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 5, 
    
    -- channel=200
    411, 473, 450, 410, 411, 452, 450, 440, 448, 447, 455, 450, 466, 510, 519, 
    409, 468, 488, 372, 331, 334, 343, 339, 357, 364, 360, 370, 475, 510, 517, 
    402, 457, 480, 354, 379, 365, 355, 356, 401, 417, 411, 417, 451, 518, 520, 
    407, 450, 449, 342, 353, 364, 373, 360, 363, 364, 351, 387, 388, 496, 501, 
    438, 450, 469, 445, 394, 392, 394, 407, 411, 406, 405, 440, 488, 499, 498, 
    475, 470, 424, 454, 481, 475, 481, 489, 483, 481, 484, 484, 494, 499, 504, 
    490, 456, 370, 268, 328, 447, 491, 505, 507, 501, 492, 496, 495, 496, 495, 
    501, 522, 528, 454, 248, 253, 400, 496, 504, 494, 492, 493, 495, 493, 491, 
    511, 537, 541, 530, 344, 164, 183, 253, 347, 420, 455, 497, 495, 492, 489, 
    510, 531, 534, 524, 282, 96, 130, 164, 172, 148, 153, 272, 358, 438, 479, 
    492, 520, 527, 496, 412, 324, 204, 290, 412, 307, 307, 270, 341, 435, 459, 
    369, 380, 368, 354, 342, 333, 315, 330, 347, 344, 349, 357, 354, 343, 356, 
    249, 247, 246, 238, 234, 218, 207, 207, 207, 189, 184, 179, 183, 180, 157, 
    138, 125, 125, 125, 131, 112, 112, 119, 131, 120, 114, 118, 114, 122, 202, 
    130, 120, 119, 122, 121, 126, 139, 144, 151, 144, 135, 129, 145, 258, 236, 
    
    -- channel=201
    386, 451, 397, 310, 333, 340, 317, 317, 314, 317, 320, 316, 326, 334, 348, 
    441, 504, 441, 83, 76, 106, 89, 98, 90, 113, 127, 160, 347, 360, 363, 
    436, 505, 435, 83, 57, 40, 0, 11, 69, 79, 88, 123, 294, 385, 382, 
    436, 500, 328, 0, 96, 126, 82, 64, 105, 65, 61, 103, 189, 394, 412, 
    432, 489, 467, 378, 355, 357, 367, 351, 363, 344, 322, 369, 370, 420, 431, 
    406, 458, 443, 441, 427, 421, 414, 407, 408, 415, 399, 416, 420, 402, 420, 
    380, 397, 296, 283, 382, 422, 418, 420, 412, 407, 408, 413, 416, 411, 414, 
    387, 427, 370, 235, 210, 318, 367, 382, 384, 382, 385, 400, 413, 415, 438, 
    368, 380, 371, 331, 200, 155, 179, 261, 317, 355, 391, 400, 407, 414, 434, 
    334, 342, 361, 342, 179, 137, 133, 119, 133, 184, 270, 299, 333, 370, 406, 
    343, 359, 366, 304, 228, 181, 175, 202, 215, 191, 207, 179, 263, 304, 360, 
    330, 352, 339, 337, 338, 343, 348, 364, 397, 412, 410, 419, 427, 443, 436, 
    246, 287, 290, 272, 260, 265, 283, 307, 313, 314, 313, 322, 329, 316, 303, 
    133, 158, 163, 142, 115, 130, 140, 133, 127, 118, 121, 124, 124, 135, 225, 
    91, 128, 129, 119, 108, 124, 119, 105, 108, 114, 112, 104, 156, 280, 238, 
    
    -- channel=202
    18, 0, 0, 7, 17, 0, 2, 8, 3, 5, 4, 5, 6, 1, 2, 
    0, 0, 0, 36, 83, 77, 78, 81, 76, 77, 71, 74, 9, 0, 0, 
    0, 0, 0, 74, 53, 78, 80, 94, 66, 54, 64, 71, 26, 0, 0, 
    0, 0, 0, 88, 64, 48, 63, 64, 59, 55, 67, 45, 65, 0, 0, 
    0, 0, 0, 0, 5, 10, 3, 5, 3, 2, 13, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 66, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 53, 77, 42, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 82, 100, 98, 72, 27, 0, 0, 0, 0, 0, 
    11, 3, 0, 0, 14, 95, 94, 89, 89, 89, 106, 93, 66, 20, 0, 
    17, 0, 0, 0, 0, 0, 26, 44, 0, 4, 11, 16, 39, 7, 4, 
    65, 42, 53, 58, 61, 43, 43, 42, 19, 19, 11, 8, 0, 1, 5, 
    59, 31, 28, 37, 46, 46, 45, 45, 41, 50, 50, 54, 52, 50, 62, 
    100, 89, 86, 92, 96, 96, 92, 94, 92, 94, 96, 93, 93, 91, 71, 
    102, 88, 85, 92, 94, 85, 80, 89, 83, 84, 89, 97, 89, 52, 55, 
    
    -- channel=203
    168, 199, 194, 180, 182, 193, 196, 183, 188, 188, 194, 193, 186, 216, 227, 
    161, 201, 209, 225, 188, 222, 228, 214, 232, 231, 229, 217, 220, 231, 231, 
    163, 193, 215, 211, 214, 178, 195, 184, 198, 204, 201, 193, 232, 230, 232, 
    164, 187, 223, 168, 173, 178, 181, 177, 180, 197, 182, 197, 163, 223, 222, 
    184, 189, 197, 216, 180, 180, 172, 181, 191, 191, 185, 179, 215, 218, 219, 
    207, 212, 216, 195, 194, 189, 194, 205, 202, 200, 199, 207, 218, 217, 214, 
    211, 196, 154, 157, 188, 214, 216, 223, 223, 226, 221, 225, 224, 226, 224, 
    212, 228, 220, 184, 121, 142, 212, 234, 231, 225, 219, 220, 219, 217, 213, 
    221, 240, 244, 242, 192, 83, 113, 165, 215, 235, 213, 220, 221, 220, 217, 
    227, 240, 242, 257, 211, 63, 64, 82, 98, 112, 115, 194, 222, 227, 218, 
    219, 234, 237, 246, 114, 100, 30, 27, 131, 77, 65, 60, 69, 169, 197, 
    223, 246, 243, 238, 235, 222, 193, 197, 208, 181, 192, 183, 193, 185, 188, 
    115, 117, 115, 116, 115, 112, 107, 118, 133, 128, 131, 128, 136, 142, 133, 
    86, 86, 84, 76, 80, 66, 62, 66, 71, 64, 56, 60, 57, 50, 26, 
    66, 60, 57, 55, 57, 44, 56, 53, 60, 51, 57, 58, 43, 54, 141, 
    
    -- channel=204
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=205
    224, 232, 190, 177, 200, 201, 189, 191, 186, 190, 192, 192, 202, 218, 233, 
    232, 256, 230, 121, 148, 180, 170, 172, 173, 183, 183, 192, 237, 239, 238, 
    235, 248, 236, 126, 129, 120, 105, 121, 133, 129, 148, 163, 236, 246, 246, 
    221, 243, 192, 94, 128, 142, 128, 132, 139, 125, 130, 141, 170, 243, 245, 
    217, 237, 228, 197, 199, 199, 198, 197, 204, 200, 200, 224, 221, 237, 243, 
    233, 235, 252, 237, 203, 204, 209, 209, 204, 210, 213, 228, 240, 234, 237, 
    240, 181, 114, 197, 288, 266, 235, 234, 233, 229, 237, 239, 242, 244, 247, 
    252, 244, 205, 87, 91, 251, 298, 254, 232, 229, 232, 232, 234, 233, 238, 
    258, 252, 246, 221, 45, 114, 171, 249, 291, 272, 251, 225, 230, 237, 239, 
    254, 245, 245, 232, 80, 87, 104, 100, 115, 139, 224, 285, 305, 276, 242, 
    250, 239, 243, 184, 66, 0, 19, 83, 78, 33, 44, 27, 130, 179, 217, 
    281, 285, 287, 287, 292, 253, 243, 265, 249, 226, 241, 226, 235, 233, 242, 
    135, 135, 130, 134, 136, 134, 138, 164, 166, 174, 176, 184, 192, 186, 182, 
    101, 116, 111, 108, 97, 92, 94, 98, 94, 86, 85, 84, 82, 85, 114, 
    65, 78, 76, 79, 75, 71, 63, 72, 65, 61, 67, 78, 100, 128, 163, 
    
    -- channel=206
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 70, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 150, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 21, 61, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=207
    410, 430, 361, 355, 378, 400, 391, 390, 390, 393, 400, 390, 420, 448, 451, 
    408, 431, 420, 241, 297, 281, 268, 293, 286, 302, 302, 324, 439, 440, 449, 
    400, 423, 397, 255, 302, 319, 270, 312, 334, 343, 342, 346, 419, 450, 458, 
    393, 420, 356, 277, 311, 314, 304, 311, 314, 296, 321, 348, 370, 440, 441, 
    409, 418, 415, 353, 346, 338, 350, 356, 355, 342, 355, 416, 423, 437, 439, 
    444, 397, 344, 440, 423, 424, 430, 431, 422, 424, 428, 429, 435, 438, 448, 
    462, 386, 281, 196, 337, 426, 439, 444, 444, 430, 431, 430, 430, 429, 435, 
    479, 461, 455, 356, 137, 258, 403, 446, 432, 425, 431, 431, 435, 430, 434, 
    485, 474, 464, 446, 140, 160, 166, 227, 320, 377, 422, 433, 429, 428, 432, 
    484, 461, 463, 409, 87, 77, 135, 159, 149, 104, 144, 239, 335, 404, 432, 
    471, 450, 456, 406, 377, 239, 218, 357, 380, 243, 321, 241, 398, 397, 413, 
    321, 291, 278, 269, 262, 247, 256, 293, 278, 290, 291, 308, 296, 288, 305, 
    224, 222, 210, 202, 199, 189, 182, 183, 170, 162, 154, 155, 158, 147, 134, 
    101, 109, 109, 113, 107, 100, 105, 113, 118, 102, 106, 107, 104, 124, 244, 
    96, 105, 110, 113, 109, 137, 128, 142, 137, 133, 114, 114, 172, 267, 157, 
    
    -- channel=208
    581, 670, 611, 569, 596, 625, 612, 605, 610, 613, 623, 615, 640, 692, 705, 
    588, 673, 674, 534, 526, 554, 545, 555, 569, 577, 578, 587, 694, 708, 717, 
    580, 653, 663, 562, 539, 528, 503, 538, 571, 576, 573, 593, 669, 713, 723, 
    582, 646, 624, 515, 531, 541, 532, 535, 555, 541, 534, 565, 592, 693, 708, 
    612, 645, 659, 614, 563, 562, 563, 585, 591, 570, 568, 631, 684, 696, 703, 
    649, 646, 608, 652, 656, 653, 669, 679, 668, 657, 659, 681, 693, 694, 705, 
    667, 619, 473, 403, 542, 667, 703, 716, 713, 699, 694, 695, 693, 696, 703, 
    685, 720, 683, 529, 315, 423, 622, 707, 706, 690, 686, 688, 693, 689, 694, 
    694, 732, 734, 700, 378, 222, 281, 407, 540, 622, 673, 703, 696, 689, 694, 
    690, 721, 730, 690, 325, 133, 176, 218, 233, 227, 297, 438, 548, 642, 690, 
    676, 720, 723, 654, 510, 355, 254, 387, 492, 348, 368, 313, 462, 594, 652, 
    534, 565, 541, 525, 518, 475, 457, 517, 537, 527, 531, 540, 550, 555, 566, 
    341, 365, 350, 329, 314, 298, 300, 324, 325, 309, 304, 306, 317, 313, 291, 
    181, 190, 183, 169, 154, 140, 145, 148, 147, 125, 120, 125, 124, 132, 206, 
    139, 136, 135, 133, 127, 144, 153, 155, 156, 147, 134, 121, 155, 252, 231, 
    
    -- channel=209
    247, 286, 279, 243, 240, 267, 269, 256, 263, 258, 269, 265, 271, 314, 325, 
    238, 283, 307, 229, 201, 215, 223, 215, 232, 240, 235, 228, 300, 317, 320, 
    235, 280, 298, 240, 258, 242, 232, 230, 264, 279, 272, 270, 281, 326, 326, 
    241, 272, 284, 207, 214, 215, 236, 207, 211, 222, 207, 235, 210, 309, 309, 
    273, 272, 294, 290, 237, 234, 231, 242, 254, 250, 239, 257, 303, 309, 308, 
    300, 307, 275, 289, 304, 301, 302, 312, 312, 308, 305, 299, 305, 306, 308, 
    304, 281, 216, 130, 202, 280, 301, 313, 318, 320, 309, 316, 311, 310, 307, 
    306, 327, 354, 334, 139, 124, 247, 313, 316, 311, 307, 310, 311, 308, 303, 
    313, 339, 342, 344, 293, 83, 69, 134, 232, 285, 279, 308, 308, 307, 305, 
    316, 333, 338, 357, 250, 40, 67, 96, 82, 52, 44, 174, 246, 286, 301, 
    302, 320, 328, 323, 263, 216, 68, 116, 264, 173, 172, 125, 155, 244, 269, 
    252, 268, 261, 252, 239, 263, 240, 214, 226, 240, 226, 245, 219, 205, 217, 
    160, 157, 162, 160, 161, 156, 145, 132, 145, 131, 127, 119, 125, 127, 103, 
    75, 55, 63, 59, 69, 54, 54, 60, 77, 68, 61, 68, 61, 59, 99, 
    85, 65, 64, 64, 66, 61, 75, 72, 81, 76, 77, 77, 70, 157, 145, 
    
    -- channel=210
    70, 49, 53, 43, 37, 39, 40, 43, 43, 41, 39, 38, 40, 42, 47, 
    78, 67, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 36, 37, 
    82, 71, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 47, 41, 
    79, 67, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 43, 
    74, 67, 59, 38, 42, 41, 45, 33, 39, 40, 43, 44, 30, 50, 49, 
    73, 72, 68, 49, 67, 62, 56, 49, 53, 67, 63, 57, 47, 46, 48, 
    66, 46, 65, 67, 43, 39, 39, 38, 42, 46, 46, 47, 48, 45, 40, 
    65, 50, 61, 75, 96, 65, 41, 34, 33, 35, 44, 46, 48, 48, 49, 
    67, 47, 47, 45, 61, 97, 82, 53, 43, 39, 32, 34, 42, 49, 47, 
    60, 39, 39, 41, 39, 99, 92, 87, 90, 66, 55, 52, 52, 45, 37, 
    53, 32, 41, 30, 55, 94, 92, 89, 92, 100, 105, 100, 94, 62, 43, 
    65, 40, 45, 44, 44, 53, 76, 52, 26, 33, 46, 39, 37, 14, 21, 
    89, 68, 81, 93, 104, 104, 101, 92, 84, 89, 86, 86, 84, 78, 77, 
    89, 79, 85, 97, 103, 100, 104, 110, 117, 122, 124, 122, 119, 126, 166, 
    108, 114, 113, 117, 118, 113, 117, 121, 121, 124, 129, 135, 147, 189, 170, 
    
    -- channel=211
    108, 157, 177, 140, 130, 143, 145, 130, 138, 135, 139, 140, 121, 135, 138, 
    117, 149, 170, 204, 145, 159, 167, 150, 166, 160, 165, 139, 146, 151, 149, 
    116, 152, 166, 170, 166, 136, 155, 130, 146, 155, 139, 124, 146, 149, 151, 
    131, 153, 189, 152, 153, 154, 147, 150, 156, 177, 150, 162, 113, 153, 152, 
    153, 153, 158, 193, 147, 144, 140, 143, 157, 154, 136, 112, 165, 154, 158, 
    146, 169, 160, 151, 162, 156, 156, 168, 172, 160, 150, 151, 156, 153, 151, 
    131, 196, 163, 101, 99, 145, 160, 168, 166, 170, 159, 164, 160, 159, 156, 
    120, 161, 166, 198, 133, 57, 98, 153, 167, 166, 154, 161, 160, 162, 159, 
    116, 146, 151, 168, 269, 68, 52, 66, 102, 146, 146, 168, 165, 158, 161, 
    116, 144, 150, 178, 281, 76, 61, 75, 75, 97, 53, 85, 103, 132, 158, 
    117, 151, 149, 210, 145, 192, 85, 14, 135, 131, 96, 105, 24, 117, 136, 
    118, 156, 150, 144, 138, 171, 140, 127, 176, 166, 163, 170, 176, 180, 171, 
    111, 134, 137, 125, 111, 118, 120, 118, 141, 128, 133, 123, 128, 140, 130, 
    91, 86, 91, 70, 72, 73, 70, 65, 67, 65, 56, 62, 62, 50, 0, 
    82, 69, 71, 60, 62, 57, 69, 49, 66, 60, 62, 52, 28, 16, 85, 
    
    -- channel=212
    68, 30, 0, 4, 22, 1, 0, 3, 0, 1, 0, 0, 14, 9, 2, 
    78, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 2, 
    72, 51, 9, 0, 0, 0, 0, 0, 0, 0, 0, 6, 15, 2, 8, 
    65, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 8, 16, 
    37, 49, 15, 0, 15, 16, 15, 17, 9, 0, 14, 38, 15, 13, 18, 
    22, 25, 18, 13, 18, 21, 25, 12, 6, 15, 18, 36, 11, 8, 18, 
    26, 0, 0, 54, 56, 26, 15, 8, 3, 0, 11, 6, 11, 9, 14, 
    39, 6, 0, 0, 28, 105, 49, 3, 0, 0, 5, 4, 9, 7, 22, 
    36, 3, 0, 0, 0, 38, 77, 58, 26, 8, 21, 3, 5, 8, 17, 
    27, 0, 0, 0, 0, 26, 31, 16, 31, 25, 84, 36, 29, 17, 16, 
    37, 0, 0, 0, 0, 0, 32, 92, 0, 0, 21, 8, 117, 47, 28, 
    44, 3, 0, 1, 8, 0, 26, 67, 11, 11, 37, 20, 48, 33, 31, 
    27, 18, 16, 16, 21, 18, 35, 56, 18, 31, 28, 37, 32, 18, 25, 
    0, 13, 4, 11, 0, 13, 18, 18, 6, 8, 18, 17, 18, 18, 76, 
    0, 15, 15, 23, 9, 26, 14, 22, 7, 13, 14, 11, 39, 86, 18, 
    
    -- channel=213
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 13, 0, 0, 0, 11, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 5, 4, 5, 5, 
    2, 6, 5, 5, 7, 10, 7, 5, 6, 8, 6, 6, 6, 0, 0, 
    
    -- channel=214
    4, 18, 10, 5, 5, 9, 4, 3, 1, 2, 4, 4, 2, 11, 13, 
    10, 18, 17, 7, 4, 16, 16, 12, 15, 15, 18, 11, 12, 16, 17, 
    11, 17, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 16, 20, 16, 
    8, 15, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 17, 
    8, 14, 16, 14, 10, 12, 8, 6, 14, 10, 7, 6, 11, 17, 17, 
    11, 21, 33, 13, 8, 9, 9, 10, 11, 12, 10, 15, 15, 13, 13, 
    10, 3, 0, 14, 36, 24, 14, 16, 16, 16, 17, 18, 19, 20, 18, 
    12, 14, 10, 0, 0, 21, 36, 18, 14, 16, 14, 16, 16, 16, 15, 
    12, 16, 18, 13, 4, 0, 3, 25, 42, 32, 19, 15, 16, 18, 16, 
    9, 15, 15, 19, 17, 0, 0, 0, 0, 1, 18, 42, 42, 30, 17, 
    7, 16, 16, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    36, 46, 48, 47, 48, 41, 37, 35, 31, 31, 28, 27, 26, 24, 28, 
    0, 4, 5, 10, 11, 8, 11, 15, 21, 21, 24, 25, 26, 28, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    
    -- channel=215
    1, 0, 0, 20, 6, 2, 10, 6, 8, 6, 9, 8, 7, 17, 14, 
    0, 0, 0, 87, 128, 125, 124, 127, 129, 123, 115, 87, 22, 8, 8, 
    0, 0, 0, 97, 98, 107, 127, 115, 90, 95, 97, 94, 36, 3, 5, 
    0, 0, 5, 108, 77, 63, 75, 81, 70, 86, 85, 77, 46, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 10, 0, 2, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 4, 24, 29, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 4, 46, 34, 36, 32, 10, 0, 1, 0, 0, 0, 0, 0, 
    20, 13, 10, 16, 60, 68, 62, 59, 64, 42, 3, 0, 0, 0, 0, 
    31, 23, 14, 40, 68, 62, 77, 84, 68, 48, 36, 66, 63, 29, 0, 
    26, 10, 10, 12, 15, 26, 4, 9, 33, 7, 22, 7, 10, 8, 0, 
    59, 49, 57, 58, 55, 52, 50, 33, 7, 12, 3, 4, 0, 0, 0, 
    48, 27, 29, 40, 51, 49, 43, 33, 38, 39, 39, 37, 37, 41, 38, 
    73, 61, 64, 68, 78, 71, 68, 73, 76, 77, 76, 78, 74, 61, 29, 
    89, 70, 70, 75, 78, 70, 70, 75, 74, 73, 79, 84, 52, 36, 56, 
    
    -- channel=216
    185, 218, 238, 210, 206, 227, 234, 220, 227, 228, 233, 232, 218, 237, 248, 
    188, 230, 241, 222, 186, 199, 215, 192, 207, 211, 208, 191, 235, 255, 257, 
    189, 228, 245, 169, 163, 135, 138, 126, 143, 155, 151, 162, 208, 257, 256, 
    194, 219, 248, 167, 180, 176, 184, 170, 197, 208, 191, 201, 186, 255, 257, 
    213, 221, 228, 233, 203, 207, 205, 205, 214, 215, 206, 200, 226, 249, 249, 
    228, 241, 234, 202, 214, 206, 206, 215, 213, 215, 215, 228, 248, 250, 248, 
    236, 246, 241, 211, 181, 219, 242, 249, 249, 251, 243, 248, 250, 254, 253, 
    238, 255, 238, 204, 170, 151, 194, 247, 260, 254, 246, 247, 245, 247, 245, 
    242, 263, 272, 261, 249, 96, 148, 193, 202, 222, 221, 248, 251, 250, 247, 
    243, 266, 271, 294, 255, 79, 73, 85, 126, 173, 165, 203, 202, 217, 236, 
    235, 259, 266, 268, 148, 142, 80, 49, 140, 122, 88, 116, 94, 197, 231, 
    216, 241, 246, 242, 237, 215, 164, 179, 226, 193, 194, 184, 201, 214, 212, 
    129, 120, 118, 111, 109, 102, 94, 108, 132, 124, 128, 128, 133, 139, 135, 
    132, 119, 117, 106, 112, 97, 91, 91, 95, 87, 78, 77, 75, 73, 66, 
    91, 76, 73, 74, 76, 62, 75, 71, 83, 77, 77, 78, 62, 99, 170, 
    
    -- channel=217
    207, 226, 178, 203, 222, 215, 205, 210, 207, 208, 213, 209, 232, 253, 238, 
    193, 194, 212, 264, 329, 316, 290, 316, 319, 315, 302, 294, 276, 246, 242, 
    185, 178, 217, 338, 352, 382, 371, 403, 383, 379, 369, 354, 290, 235, 241, 
    190, 187, 229, 364, 321, 308, 308, 342, 320, 315, 326, 323, 304, 222, 223, 
    196, 189, 202, 209, 199, 190, 187, 216, 212, 192, 201, 241, 260, 222, 221, 
    205, 186, 162, 225, 225, 233, 250, 256, 247, 228, 232, 233, 220, 222, 224, 
    215, 168, 101, 100, 191, 229, 240, 244, 240, 231, 232, 227, 221, 223, 226, 
    224, 222, 226, 188, 94, 155, 229, 241, 236, 230, 229, 226, 226, 222, 220, 
    229, 232, 231, 231, 76, 96, 81, 118, 184, 217, 242, 243, 228, 216, 219, 
    237, 237, 238, 211, 32, 61, 95, 117, 79, 29, 66, 120, 179, 220, 238, 
    237, 244, 236, 204, 234, 150, 129, 237, 229, 139, 184, 125, 234, 230, 228, 
    169, 170, 147, 140, 138, 131, 163, 191, 167, 186, 184, 202, 193, 191, 192, 
    133, 160, 150, 136, 123, 120, 131, 134, 112, 106, 99, 97, 99, 99, 83, 
    38, 56, 51, 45, 32, 37, 45, 44, 38, 28, 33, 40, 40, 33, 34, 
    49, 53, 56, 52, 44, 67, 67, 64, 54, 53, 46, 32, 32, 30, 0, 
    
    -- channel=218
    68, 21, 0, 0, 39, 7, 0, 12, 0, 8, 6, 4, 24, 19, 8, 
    58, 27, 0, 0, 54, 41, 13, 37, 20, 30, 24, 44, 41, 11, 10, 
    56, 16, 0, 0, 14, 49, 10, 63, 32, 21, 24, 32, 58, 10, 10, 
    40, 19, 0, 21, 47, 34, 21, 53, 43, 18, 62, 40, 82, 11, 15, 
    10, 18, 0, 0, 11, 12, 8, 19, 10, 0, 18, 62, 4, 7, 7, 
    15, 0, 0, 10, 0, 0, 6, 0, 0, 0, 2, 14, 5, 2, 7, 
    31, 0, 0, 61, 97, 34, 12, 4, 0, 0, 6, 0, 4, 6, 13, 
    48, 0, 0, 0, 0, 131, 94, 15, 0, 0, 6, 0, 3, 0, 8, 
    49, 6, 0, 0, 0, 37, 83, 102, 71, 28, 34, 0, 0, 0, 5, 
    52, 10, 4, 0, 0, 29, 38, 21, 30, 31, 113, 81, 66, 36, 15, 
    61, 7, 6, 0, 0, 0, 11, 105, 0, 0, 0, 0, 122, 38, 32, 
    68, 19, 15, 20, 30, 0, 17, 68, 18, 1, 28, 10, 31, 31, 29, 
    10, 2, 0, 0, 0, 0, 5, 30, 0, 12, 9, 21, 19, 8, 21, 
    0, 19, 7, 12, 0, 8, 12, 12, 1, 0, 7, 3, 6, 14, 33, 
    0, 2, 4, 10, 0, 11, 0, 9, 0, 0, 0, 0, 28, 14, 0, 
    
    -- channel=219
    294, 333, 294, 295, 305, 325, 320, 314, 318, 316, 324, 319, 339, 382, 385, 
    279, 301, 334, 357, 364, 365, 361, 369, 384, 382, 376, 367, 381, 379, 383, 
    269, 290, 327, 391, 417, 422, 424, 434, 444, 447, 437, 428, 397, 376, 384, 
    271, 290, 333, 402, 367, 363, 375, 391, 368, 376, 375, 389, 354, 354, 353, 
    300, 292, 310, 320, 284, 275, 271, 295, 299, 291, 296, 324, 378, 348, 349, 
    336, 309, 279, 336, 337, 341, 355, 367, 360, 345, 350, 349, 346, 352, 353, 
    353, 303, 205, 139, 258, 343, 356, 366, 367, 361, 356, 356, 351, 351, 353, 
    361, 366, 383, 350, 138, 177, 330, 378, 367, 360, 357, 355, 353, 348, 341, 
    373, 391, 391, 395, 223, 121, 112, 167, 285, 341, 352, 363, 353, 345, 343, 
    384, 394, 392, 373, 187, 56, 105, 145, 117, 59, 66, 195, 294, 348, 359, 
    371, 386, 385, 373, 321, 233, 124, 225, 330, 204, 232, 164, 250, 322, 331, 
    282, 288, 272, 260, 252, 249, 252, 264, 244, 252, 253, 267, 255, 234, 248, 
    185, 190, 183, 179, 173, 165, 161, 157, 152, 136, 131, 125, 130, 133, 109, 
    79, 76, 73, 71, 73, 62, 65, 71, 76, 67, 64, 70, 67, 66, 92, 
    91, 76, 75, 76, 76, 87, 91, 96, 95, 85, 79, 75, 82, 105, 86, 
    
    -- channel=220
    309, 381, 369, 303, 307, 340, 334, 321, 329, 325, 332, 329, 334, 366, 374, 
    317, 376, 395, 264, 193, 217, 221, 209, 227, 235, 240, 238, 357, 374, 377, 
    314, 369, 372, 257, 284, 253, 239, 237, 290, 296, 290, 282, 326, 384, 384, 
    323, 368, 363, 230, 245, 257, 267, 242, 247, 253, 232, 275, 241, 370, 374, 
    355, 364, 383, 368, 311, 304, 307, 310, 320, 322, 305, 322, 375, 378, 381, 
    369, 370, 340, 384, 392, 387, 386, 394, 394, 390, 383, 370, 380, 379, 379, 
    362, 390, 289, 143, 241, 360, 378, 388, 390, 387, 376, 384, 379, 376, 374, 
    362, 399, 426, 411, 171, 146, 292, 376, 379, 376, 371, 378, 382, 382, 379, 
    361, 390, 394, 403, 336, 124, 88, 129, 241, 325, 353, 381, 378, 376, 377, 
    356, 376, 387, 378, 306, 83, 105, 133, 118, 85, 60, 166, 261, 338, 371, 
    342, 378, 380, 411, 355, 318, 175, 197, 346, 269, 270, 223, 220, 312, 329, 
    254, 286, 272, 259, 249, 286, 273, 261, 285, 300, 295, 317, 303, 289, 297, 
    203, 228, 231, 222, 210, 208, 203, 190, 200, 182, 180, 168, 174, 177, 153, 
    99, 97, 104, 98, 100, 92, 95, 97, 110, 103, 96, 104, 100, 110, 158, 
    109, 108, 110, 103, 106, 111, 121, 114, 125, 118, 112, 105, 129, 191, 184, 
    
    -- channel=221
    682, 758, 648, 613, 650, 679, 657, 653, 655, 660, 669, 660, 698, 759, 770, 
    697, 768, 738, 505, 540, 559, 534, 560, 567, 582, 581, 610, 758, 769, 781, 
    681, 748, 732, 522, 533, 534, 492, 539, 580, 590, 592, 620, 741, 780, 794, 
    676, 743, 646, 479, 534, 551, 522, 546, 552, 521, 532, 577, 630, 763, 776, 
    697, 738, 728, 658, 615, 612, 613, 635, 641, 613, 624, 704, 754, 767, 775, 
    740, 726, 677, 736, 730, 729, 747, 752, 737, 733, 737, 760, 761, 760, 778, 
    759, 659, 467, 438, 631, 753, 773, 783, 778, 762, 763, 763, 765, 764, 772, 
    786, 796, 740, 535, 324, 508, 722, 779, 763, 747, 751, 755, 762, 756, 768, 
    794, 809, 797, 753, 298, 259, 325, 460, 614, 697, 750, 764, 759, 756, 766, 
    786, 789, 793, 730, 237, 150, 209, 246, 257, 235, 336, 494, 634, 727, 764, 
    775, 781, 788, 684, 517, 342, 277, 461, 544, 354, 417, 328, 561, 665, 716, 
    627, 621, 594, 578, 572, 516, 534, 605, 588, 575, 602, 603, 623, 607, 621, 
    390, 406, 390, 375, 363, 347, 355, 386, 367, 356, 349, 354, 364, 352, 325, 
    183, 202, 191, 181, 163, 156, 162, 169, 166, 144, 144, 151, 148, 159, 281, 
    140, 157, 156, 158, 146, 174, 172, 182, 178, 168, 156, 145, 208, 338, 298, 
    
    -- channel=222
    0, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 160, 0, 0, 32, 0, 7, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 57, 72, 0, 45, 0, 2, 22, 0, 0, 0, 0, 0, 
    0, 0, 97, 19, 0, 0, 31, 0, 0, 72, 0, 23, 0, 0, 0, 
    0, 0, 0, 80, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 107, 129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 48, 246, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 498, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 176, 72, 244, 0, 0, 34, 82, 0, 14, 0, 0, 0, 
    0, 0, 3, 0, 0, 91, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 6, 0, 3, 0, 0, 22, 0, 0, 0, 0, 15, 0, 
    32, 0, 8, 0, 12, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 
    
    -- channel=223
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 4, 6, 7, 7, 12, 15, 13, 14, 13, 0, 
    1, 11, 13, 14, 14, 5, 7, 8, 3, 5, 12, 17, 6, 0, 0, 
    
    -- channel=224
    0, 0, 0, 8, 3, 0, 6, 5, 6, 7, 5, 8, 2, 0, 0, 
    0, 0, 0, 127, 129, 123, 132, 126, 130, 117, 114, 101, 5, 4, 4, 
    0, 0, 0, 137, 112, 119, 151, 137, 109, 105, 100, 90, 36, 0, 0, 
    0, 0, 3, 163, 116, 104, 106, 129, 118, 133, 130, 101, 86, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 4, 4, 7, 9, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 55, 20, 37, 44, 30, 13, 0, 0, 0, 0, 0, 
    0, 5, 0, 12, 86, 33, 30, 36, 35, 53, 42, 36, 18, 0, 0, 
    0, 3, 0, 18, 9, 2, 0, 0, 0, 12, 0, 0, 0, 0, 1, 
    17, 25, 29, 30, 32, 28, 0, 0, 18, 0, 0, 0, 0, 4, 0, 
    13, 8, 3, 1, 0, 0, 0, 2, 11, 8, 11, 11, 13, 18, 25, 
    53, 43, 39, 33, 36, 34, 27, 26, 23, 24, 20, 20, 20, 8, 0, 
    47, 25, 20, 20, 24, 18, 18, 17, 19, 15, 16, 16, 0, 0, 0, 
    
    -- channel=225
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=226
    22, 10, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    22, 9, 0, 0, 19, 3, 0, 4, 0, 1, 3, 0, 11, 0, 0, 
    21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 
    17, 10, 0, 0, 1, 0, 0, 0, 0, 0, 13, 16, 4, 4, 0, 
    14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 
    18, 2, 0, 9, 0, 0, 1, 0, 0, 0, 1, 6, 0, 0, 0, 
    20, 0, 0, 0, 17, 13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 2, 0, 0, 0, 24, 25, 4, 0, 0, 0, 0, 0, 0, 0, 
    29, 5, 0, 0, 0, 13, 14, 11, 10, 8, 5, 0, 0, 0, 0, 
    31, 4, 0, 0, 0, 0, 6, 4, 5, 0, 2, 9, 13, 8, 2, 
    28, 1, 0, 0, 0, 0, 4, 18, 9, 0, 13, 0, 41, 11, 7, 
    18, 0, 0, 0, 0, 0, 2, 19, 0, 0, 4, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 6, 
    
    -- channel=227
    60, 35, 16, 79, 77, 73, 79, 80, 80, 81, 84, 79, 92, 101, 88, 
    33, 0, 19, 169, 250, 207, 204, 217, 217, 208, 196, 171, 104, 79, 79, 
    28, 0, 30, 198, 235, 271, 275, 291, 247, 251, 251, 227, 130, 65, 70, 
    28, 0, 54, 276, 214, 198, 204, 237, 208, 221, 237, 215, 190, 57, 46, 
    37, 3, 7, 44, 52, 42, 40, 64, 53, 52, 74, 70, 82, 42, 37, 
    59, 14, 0, 42, 41, 44, 58, 63, 57, 46, 56, 50, 40, 51, 47, 
    76, 18, 30, 38, 35, 44, 53, 54, 55, 51, 53, 46, 43, 45, 45, 
    83, 48, 72, 95, 41, 61, 66, 72, 63, 60, 62, 53, 48, 43, 33, 
    97, 77, 73, 91, 16, 89, 72, 62, 64, 63, 59, 60, 52, 42, 34, 
    113, 93, 81, 85, 0, 59, 94, 108, 81, 37, 18, 42, 54, 56, 57, 
    108, 84, 79, 77, 125, 90, 97, 162, 140, 82, 116, 90, 142, 100, 79, 
    54, 29, 24, 23, 18, 12, 23, 31, 4, 0, 9, 8, 1, 0, 0, 
    60, 53, 48, 50, 53, 46, 40, 32, 18, 14, 8, 8, 4, 5, 3, 
    51, 57, 55, 61, 67, 62, 61, 66, 69, 65, 69, 69, 68, 58, 61, 
    76, 70, 73, 78, 76, 89, 86, 93, 87, 85, 78, 79, 57, 43, 0, 
    
    -- channel=228
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 18, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 6, 8, 12, 16, 18, 19, 18, 20, 22, 24, 23, 23, 13, 0, 
    23, 20, 22, 23, 24, 17, 19, 17, 15, 20, 26, 30, 1, 4, 0, 
    
    -- channel=229
    179, 236, 201, 168, 175, 194, 182, 175, 173, 176, 183, 181, 186, 213, 220, 
    194, 240, 250, 148, 145, 173, 166, 159, 174, 179, 178, 163, 230, 237, 232, 
    192, 232, 254, 138, 154, 119, 111, 113, 138, 151, 143, 137, 216, 240, 240, 
    191, 232, 234, 87, 132, 141, 122, 125, 136, 146, 136, 158, 131, 238, 238, 
    208, 226, 235, 219, 180, 176, 178, 184, 197, 190, 174, 202, 222, 238, 239, 
    225, 236, 227, 239, 215, 211, 218, 228, 223, 219, 214, 217, 238, 232, 232, 
    220, 206, 109, 117, 213, 243, 239, 247, 244, 240, 238, 242, 241, 242, 241, 
    226, 249, 242, 133, 30, 136, 228, 245, 241, 237, 229, 234, 237, 236, 236, 
    229, 244, 243, 245, 111, 10, 29, 137, 213, 235, 234, 238, 238, 236, 238, 
    226, 235, 242, 246, 138, 0, 1, 8, 2, 33, 84, 181, 220, 234, 237, 
    219, 238, 240, 235, 107, 17, 0, 13, 84, 23, 15, 0, 55, 145, 201, 
    210, 239, 230, 225, 221, 230, 188, 189, 230, 211, 215, 219, 214, 227, 228, 
    73, 100, 98, 89, 76, 77, 80, 95, 114, 107, 108, 108, 119, 121, 98, 
    0, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 40, 
    
    -- channel=230
    361, 406, 353, 364, 381, 396, 390, 386, 385, 392, 398, 395, 409, 444, 452, 
    359, 395, 402, 403, 433, 447, 443, 447, 459, 454, 458, 443, 451, 456, 461, 
    353, 382, 409, 402, 400, 391, 395, 413, 407, 414, 410, 415, 462, 452, 459, 
    348, 379, 395, 386, 394, 400, 378, 404, 407, 416, 420, 412, 429, 440, 444, 
    367, 379, 383, 377, 350, 348, 348, 370, 372, 363, 369, 402, 428, 430, 431, 
    407, 392, 370, 393, 377, 372, 392, 404, 391, 384, 393, 410, 427, 432, 435, 
    429, 360, 269, 317, 381, 423, 436, 444, 441, 431, 433, 430, 432, 438, 442, 
    448, 447, 418, 270, 189, 330, 429, 458, 449, 438, 433, 428, 427, 423, 422, 
    463, 473, 470, 461, 186, 159, 231, 345, 403, 420, 431, 438, 435, 428, 425, 
    469, 477, 473, 461, 199, 101, 135, 155, 172, 200, 262, 359, 401, 423, 434, 
    458, 469, 470, 424, 270, 134, 123, 225, 260, 169, 164, 152, 277, 370, 423, 
    394, 405, 395, 388, 385, 338, 298, 343, 367, 315, 343, 325, 345, 355, 364, 
    206, 215, 201, 192, 184, 171, 169, 200, 204, 197, 196, 202, 211, 209, 200, 
    138, 154, 143, 131, 125, 110, 107, 111, 109, 89, 86, 86, 86, 82, 102, 
    91, 89, 90, 92, 87, 92, 94, 101, 101, 91, 85, 85, 83, 119, 151, 
    
    -- channel=231
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 24, 18, 19, 12, 22, 20, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=232
    11, 5, 7, 0, 7, 8, 10, 8, 13, 10, 11, 10, 14, 23, 23, 
    2, 0, 3, 12, 19, 2, 2, 3, 3, 7, 2, 5, 24, 17, 20, 
    0, 0, 0, 11, 36, 55, 42, 52, 50, 49, 56, 52, 17, 21, 22, 
    5, 0, 0, 71, 42, 40, 49, 50, 46, 37, 38, 38, 42, 14, 12, 
    12, 0, 0, 8, 0, 0, 0, 0, 0, 0, 3, 4, 28, 7, 12, 
    13, 5, 0, 0, 22, 22, 25, 26, 26, 22, 22, 21, 8, 13, 14, 
    17, 6, 0, 0, 0, 0, 12, 14, 15, 16, 13, 13, 11, 9, 11, 
    17, 14, 20, 51, 2, 0, 0, 12, 16, 13, 16, 14, 13, 13, 12, 
    19, 19, 20, 18, 14, 0, 0, 0, 0, 0, 4, 14, 11, 9, 10, 
    23, 22, 22, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    20, 16, 17, 9, 42, 56, 7, 27, 60, 34, 41, 25, 27, 32, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    
    -- channel=233
    474, 524, 449, 432, 460, 487, 478, 469, 477, 476, 488, 477, 512, 571, 577, 
    464, 507, 512, 378, 400, 390, 384, 405, 413, 425, 425, 438, 558, 557, 571, 
    449, 495, 482, 416, 459, 481, 436, 482, 511, 520, 513, 521, 548, 570, 576, 
    451, 487, 459, 426, 429, 429, 437, 439, 432, 417, 432, 457, 479, 538, 548, 
    485, 489, 498, 464, 419, 408, 411, 437, 441, 421, 432, 496, 550, 542, 544, 
    527, 494, 424, 517, 533, 531, 546, 553, 542, 534, 539, 544, 535, 541, 551, 
    552, 462, 329, 205, 362, 513, 544, 556, 557, 545, 540, 541, 538, 536, 542, 
    570, 568, 567, 489, 190, 261, 467, 557, 548, 536, 539, 538, 542, 535, 536, 
    581, 592, 588, 566, 252, 150, 153, 225, 373, 471, 516, 547, 538, 530, 534, 
    584, 584, 587, 550, 152, 38, 111, 160, 144, 67, 89, 250, 392, 494, 540, 
    565, 571, 575, 510, 454, 332, 200, 363, 486, 292, 362, 260, 427, 494, 507, 
    390, 382, 359, 342, 329, 307, 333, 372, 340, 359, 366, 384, 377, 347, 368, 
    251, 254, 246, 235, 230, 214, 209, 207, 186, 166, 156, 151, 154, 145, 123, 
    71, 70, 66, 69, 69, 56, 62, 71, 81, 65, 64, 70, 68, 80, 196, 
    79, 75, 77, 82, 75, 101, 105, 114, 112, 105, 89, 87, 124, 244, 144, 
    
    -- channel=234
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=235
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 46, 141, 225, 216, 202, 210, 203, 202, 159, 0, 0, 0, 
    0, 0, 13, 90, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 2, 0, 1, 
    0, 0, 0, 0, 15, 35, 10, 6, 32, 18, 11, 0, 0, 0, 0, 
    0, 13, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 317, 327, 54, 0, 0, 0, 0, 0, 0, 0, 7, 13, 
    0, 0, 0, 0, 10, 332, 221, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 40, 231, 438, 367, 178, 40, 0, 0, 0, 0, 
    0, 0, 0, 45, 103, 112, 63, 11, 74, 284, 482, 500, 344, 127, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    322, 358, 390, 412, 433, 339, 220, 238, 290, 183, 189, 135, 160, 224, 218, 
    11, 1, 0, 1, 7, 15, 28, 107, 163, 195, 215, 243, 262, 269, 285, 
    139, 166, 151, 115, 96, 91, 77, 68, 45, 29, 25, 19, 19, 0, 0, 
    10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 
    
    -- channel=236
    0, 0, 52, 33, 15, 23, 32, 27, 36, 30, 29, 32, 21, 22, 22, 
    0, 0, 26, 168, 75, 87, 97, 87, 100, 83, 81, 74, 12, 28, 23, 
    0, 0, 24, 158, 131, 115, 156, 117, 122, 119, 103, 92, 17, 19, 21, 
    0, 0, 81, 165, 106, 102, 127, 118, 111, 135, 103, 93, 47, 11, 11, 
    0, 0, 10, 48, 17, 18, 15, 26, 22, 30, 15, 0, 30, 13, 10, 
    0, 3, 5, 0, 24, 27, 26, 33, 37, 23, 22, 14, 13, 18, 12, 
    0, 55, 73, 0, 0, 0, 17, 23, 26, 31, 19, 20, 15, 16, 12, 
    0, 14, 42, 127, 79, 0, 0, 13, 33, 30, 22, 22, 17, 20, 11, 
    0, 13, 26, 42, 205, 3, 0, 0, 0, 0, 4, 28, 22, 16, 12, 
    0, 22, 25, 45, 182, 14, 5, 25, 15, 0, 0, 0, 0, 0, 13, 
    0, 25, 22, 69, 113, 154, 48, 0, 75, 116, 54, 77, 0, 27, 10, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 11, 0, 8, 0, 2, 0, 
    23, 30, 33, 23, 17, 21, 17, 1, 11, 0, 0, 0, 0, 2, 0, 
    39, 12, 15, 12, 18, 15, 12, 11, 13, 18, 11, 13, 13, 3, 0, 
    57, 23, 18, 15, 21, 17, 30, 18, 28, 26, 25, 15, 0, 0, 0, 
    
    -- channel=237
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=238
    67, 18, 0, 0, 29, 0, 0, 4, 0, 2, 0, 0, 20, 17, 9, 
    62, 29, 0, 0, 13, 9, 0, 12, 0, 0, 0, 24, 31, 2, 5, 
    60, 23, 0, 0, 0, 12, 0, 26, 1, 0, 3, 14, 51, 4, 7, 
    46, 25, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 50, 5, 9, 
    21, 24, 0, 0, 0, 0, 0, 5, 0, 0, 5, 45, 2, 6, 6, 
    24, 0, 0, 18, 2, 5, 15, 3, 0, 1, 10, 20, 2, 0, 11, 
    35, 0, 0, 9, 61, 32, 10, 1, 0, 0, 4, 0, 1, 1, 6, 
    51, 4, 0, 0, 0, 90, 73, 13, 0, 0, 1, 0, 1, 0, 7, 
    55, 12, 0, 0, 0, 22, 52, 44, 34, 15, 28, 0, 0, 0, 4, 
    53, 8, 0, 0, 0, 0, 18, 10, 11, 0, 47, 22, 37, 29, 13, 
    58, 2, 2, 0, 0, 0, 19, 114, 0, 0, 23, 0, 129, 42, 23, 
    35, 0, 0, 0, 0, 0, 0, 44, 0, 0, 2, 0, 6, 0, 0, 
    5, 0, 0, 0, 0, 0, 2, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 53, 
    0, 0, 0, 1, 0, 11, 0, 10, 0, 0, 0, 0, 34, 40, 0, 
    
    -- channel=239
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=240
    208, 222, 177, 171, 193, 197, 185, 193, 187, 192, 191, 189, 209, 210, 211, 
    212, 229, 215, 107, 134, 138, 121, 137, 132, 138, 139, 161, 217, 217, 214, 
    212, 218, 210, 125, 144, 151, 126, 152, 163, 157, 162, 163, 207, 218, 221, 
    204, 221, 183, 129, 151, 160, 147, 158, 155, 141, 155, 163, 187, 214, 219, 
    201, 217, 218, 173, 179, 175, 184, 188, 181, 178, 181, 228, 207, 217, 218, 
    211, 191, 180, 230, 205, 207, 212, 211, 203, 204, 208, 208, 220, 219, 222, 
    219, 184, 114, 122, 203, 226, 223, 221, 218, 207, 213, 211, 212, 213, 218, 
    231, 224, 211, 110, 51, 171, 225, 223, 211, 207, 211, 210, 214, 213, 217, 
    232, 224, 217, 209, 1, 80, 98, 145, 179, 192, 223, 213, 210, 212, 215, 
    228, 216, 219, 175, 0, 49, 74, 74, 69, 67, 124, 149, 186, 209, 216, 
    227, 217, 218, 181, 166, 57, 108, 197, 142, 105, 128, 103, 203, 192, 207, 
    162, 154, 145, 143, 145, 131, 134, 163, 163, 157, 167, 169, 169, 179, 181, 
    103, 118, 107, 99, 91, 89, 93, 106, 95, 97, 94, 99, 103, 94, 90, 
    49, 68, 65, 64, 50, 52, 56, 58, 54, 44, 49, 46, 46, 59, 119, 
    30, 49, 51, 50, 46, 65, 53, 62, 53, 52, 41, 41, 82, 111, 49, 
    
    -- channel=241
    60, 48, 47, 63, 53, 63, 69, 70, 72, 67, 70, 65, 78, 87, 83, 
    41, 26, 49, 59, 65, 42, 45, 55, 52, 53, 53, 62, 61, 60, 66, 
    42, 27, 24, 86, 120, 133, 127, 131, 135, 137, 130, 107, 74, 63, 64, 
    44, 29, 42, 104, 85, 82, 97, 86, 69, 72, 86, 96, 68, 52, 42, 
    58, 32, 46, 40, 38, 30, 36, 37, 34, 37, 47, 55, 65, 51, 47, 
    77, 35, 3, 71, 85, 88, 85, 83, 86, 87, 86, 61, 49, 56, 58, 
    79, 65, 57, 0, 0, 36, 51, 54, 61, 59, 54, 52, 47, 42, 39, 
    76, 63, 126, 201, 25, 0, 19, 55, 50, 53, 58, 58, 56, 53, 45, 
    82, 74, 74, 97, 88, 64, 0, 0, 0, 25, 42, 55, 50, 49, 44, 
    89, 72, 69, 48, 32, 37, 65, 88, 45, 0, 0, 0, 0, 39, 49, 
    74, 63, 65, 97, 208, 199, 136, 182, 220, 166, 210, 152, 149, 91, 52, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 56, 59, 67, 74, 71, 58, 19, 7, 1, 0, 0, 0, 0, 0, 
    24, 13, 23, 41, 54, 46, 52, 61, 75, 77, 80, 82, 78, 90, 140, 
    87, 79, 82, 84, 90, 103, 106, 114, 113, 113, 103, 102, 120, 137, 47, 
    
    -- channel=242
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 108, 8, 66, 92, 47, 76, 65, 68, 34, 0, 0, 0, 
    0, 0, 4, 85, 9, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 1, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 48, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 248, 0, 0, 30, 32, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 329, 24, 0, 0, 0, 73, 39, 62, 21, 0, 0, 
    0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 84, 97, 98, 97, 132, 36, 0, 73, 43, 22, 22, 15, 41, 33, 
    0, 0, 3, 5, 0, 9, 1, 0, 58, 51, 61, 57, 66, 85, 80, 
    75, 44, 50, 29, 39, 28, 18, 13, 15, 16, 0, 0, 0, 0, 0, 
    46, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 
    
    -- channel=243
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 8, 23, 15, 11, 12, 12, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 5, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 14, 4, 3, 8, 0, 0, 1, 11, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 42, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 35, 43, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 85, 81, 70, 43, 3, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 58, 95, 98, 90, 88, 84, 75, 68, 43, 2, 0, 
    0, 0, 0, 0, 17, 9, 43, 42, 11, 41, 28, 42, 25, 0, 0, 
    33, 14, 30, 34, 35, 41, 23, 1, 0, 0, 0, 0, 0, 0, 0, 
    49, 22, 24, 39, 51, 51, 39, 29, 35, 40, 40, 42, 40, 37, 47, 
    105, 93, 95, 108, 118, 112, 107, 112, 117, 122, 121, 116, 115, 120, 127, 
    118, 107, 105, 112, 119, 108, 102, 114, 112, 113, 115, 129, 128, 107, 113, 
    
    -- channel=244
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 129, 0, 29, 63, 16, 47, 31, 39, 0, 0, 0, 0, 
    0, 0, 0, 126, 70, 11, 68, 8, 32, 21, 5, 0, 0, 0, 0, 
    0, 0, 50, 68, 24, 15, 53, 10, 23, 75, 20, 28, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 60, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 319, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 391, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 107, 96, 120, 0, 0, 0, 64, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 67, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 8, 0, 
    40, 7, 23, 6, 18, 7, 0, 0, 6, 9, 0, 0, 0, 0, 0, 
    54, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=246
    217, 294, 267, 175, 181, 209, 194, 182, 187, 184, 191, 188, 188, 209, 214, 
    251, 313, 290, 13, 0, 0, 0, 0, 0, 0, 0, 6, 206, 219, 220, 
    246, 311, 277, 3, 32, 13, 0, 0, 47, 59, 61, 62, 148, 238, 233, 
    256, 310, 213, 0, 17, 37, 32, 0, 17, 2, 0, 44, 49, 236, 248, 
    273, 301, 301, 262, 210, 205, 209, 201, 214, 207, 185, 201, 243, 260, 266, 
    256, 289, 254, 284, 293, 285, 277, 277, 280, 282, 266, 260, 263, 252, 257, 
    231, 278, 188, 60, 143, 244, 257, 264, 261, 260, 251, 260, 258, 251, 250, 
    230, 273, 270, 241, 80, 71, 160, 228, 238, 238, 237, 250, 261, 262, 272, 
    215, 233, 232, 224, 192, 26, 0, 24, 105, 185, 221, 252, 254, 254, 265, 
    193, 205, 223, 224, 151, 2, 6, 11, 6, 6, 3, 62, 127, 197, 245, 
    191, 220, 221, 232, 186, 195, 91, 79, 192, 136, 157, 113, 119, 176, 200, 
    134, 167, 152, 143, 136, 178, 185, 175, 208, 236, 230, 251, 248, 242, 239, 
    106, 150, 159, 143, 128, 130, 138, 134, 142, 127, 127, 119, 123, 120, 96, 
    0, 6, 17, 1, 0, 0, 7, 2, 11, 5, 2, 11, 10, 18, 93, 
    0, 17, 21, 9, 4, 15, 21, 4, 14, 15, 11, 0, 35, 148, 107, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=248
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 12, 6, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 41, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 24, 0, 0, 0, 3, 1, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 8, 9, 8, 8, 0, 5, 5, 0, 8, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 8, 
    
    -- channel=249
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=250
    39, 12, 0, 12, 22, 5, 2, 9, 6, 5, 2, 5, 9, 0, 0, 
    34, 11, 0, 0, 7, 18, 11, 18, 9, 11, 13, 28, 3, 0, 0, 
    34, 14, 0, 17, 15, 23, 22, 29, 21, 10, 15, 11, 23, 0, 0, 
    29, 17, 0, 1, 16, 14, 5, 12, 5, 0, 11, 4, 15, 0, 0, 
    17, 15, 6, 0, 19, 19, 21, 14, 14, 13, 17, 20, 1, 0, 0, 
    11, 0, 16, 24, 8, 12, 10, 5, 7, 9, 9, 4, 0, 0, 0, 
    8, 2, 0, 18, 51, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 5, 31, 55, 41, 1, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 75, 61, 37, 37, 24, 18, 0, 0, 0, 0, 
    2, 0, 0, 0, 5, 89, 89, 82, 68, 50, 56, 36, 42, 27, 6, 
    10, 0, 0, 0, 25, 33, 69, 73, 33, 46, 63, 52, 56, 16, 0, 
    33, 13, 17, 19, 23, 29, 51, 49, 23, 34, 34, 36, 32, 23, 23, 
    66, 61, 61, 67, 70, 74, 77, 72, 61, 68, 68, 68, 66, 62, 70, 
    70, 70, 72, 78, 75, 83, 82, 83, 81, 86, 90, 91, 93, 98, 93, 
    86, 90, 90, 90, 90, 94, 84, 89, 85, 86, 86, 90, 107, 70, 63, 
    
    -- channel=251
    396, 441, 376, 370, 401, 417, 404, 406, 407, 412, 416, 410, 443, 478, 482, 
    392, 436, 432, 353, 393, 397, 379, 404, 406, 409, 405, 417, 483, 483, 488, 
    382, 417, 433, 392, 395, 412, 385, 428, 432, 433, 437, 453, 468, 481, 494, 
    378, 415, 395, 406, 395, 400, 393, 414, 413, 398, 407, 413, 453, 462, 475, 
    396, 416, 422, 384, 362, 357, 361, 390, 380, 367, 376, 442, 464, 461, 464, 
    428, 406, 366, 431, 424, 425, 445, 452, 436, 426, 436, 453, 459, 463, 471, 
    454, 378, 260, 246, 359, 449, 473, 480, 475, 459, 462, 458, 458, 462, 470, 
    478, 481, 444, 295, 150, 293, 431, 483, 474, 457, 460, 456, 458, 454, 457, 
    488, 501, 495, 467, 122, 111, 171, 268, 358, 411, 457, 470, 460, 453, 457, 
    489, 497, 499, 454, 74, 25, 81, 110, 115, 103, 180, 275, 362, 429, 465, 
    482, 493, 493, 408, 328, 162, 140, 300, 311, 193, 219, 173, 347, 413, 445, 
    347, 349, 328, 319, 315, 262, 264, 329, 325, 308, 325, 324, 337, 342, 349, 
    188, 202, 185, 167, 157, 144, 145, 172, 155, 147, 140, 146, 154, 145, 130, 
    61, 74, 63, 58, 41, 35, 37, 42, 37, 18, 20, 21, 21, 26, 111, 
    28, 31, 30, 32, 24, 51, 45, 55, 47, 41, 25, 19, 51, 127, 51, 
    
    -- channel=252
    553, 602, 518, 506, 530, 562, 549, 539, 542, 546, 559, 551, 581, 643, 658, 
    552, 607, 602, 413, 458, 489, 482, 492, 505, 521, 518, 515, 641, 648, 659, 
    542, 590, 599, 430, 465, 452, 422, 453, 488, 504, 506, 529, 625, 662, 665, 
    529, 579, 540, 377, 426, 433, 427, 429, 435, 427, 441, 477, 494, 637, 641, 
    557, 574, 583, 530, 497, 492, 496, 510, 521, 506, 513, 577, 606, 634, 632, 
    616, 586, 554, 608, 574, 572, 586, 594, 580, 585, 593, 608, 626, 628, 635, 
    646, 523, 378, 353, 545, 631, 625, 634, 636, 624, 625, 628, 631, 635, 638, 
    673, 658, 632, 457, 214, 430, 634, 662, 633, 621, 622, 621, 625, 618, 618, 
    691, 692, 686, 653, 257, 220, 285, 429, 570, 614, 620, 623, 621, 623, 621, 
    692, 682, 684, 657, 239, 110, 182, 214, 224, 207, 294, 482, 593, 635, 627, 
    668, 664, 672, 586, 394, 215, 151, 315, 419, 227, 288, 206, 415, 524, 581, 
    567, 567, 560, 548, 540, 486, 465, 510, 492, 473, 486, 483, 483, 469, 494, 
    305, 301, 290, 290, 291, 272, 262, 285, 286, 276, 273, 277, 288, 280, 253, 
    161, 173, 167, 167, 163, 138, 140, 152, 159, 137, 133, 137, 133, 142, 240, 
    124, 130, 132, 139, 134, 141, 140, 159, 154, 144, 136, 145, 176, 299, 299, 
    
    -- channel=253
    297, 336, 323, 305, 303, 336, 341, 327, 331, 333, 343, 341, 341, 381, 392, 
    286, 332, 351, 300, 285, 302, 318, 302, 321, 327, 323, 307, 359, 389, 395, 
    282, 325, 355, 287, 294, 270, 274, 267, 294, 310, 302, 306, 344, 392, 393, 
    280, 315, 340, 259, 276, 272, 285, 271, 281, 300, 286, 310, 287, 379, 379, 
    308, 315, 333, 334, 293, 296, 291, 299, 311, 311, 306, 317, 352, 368, 367, 
    352, 350, 332, 323, 322, 316, 321, 334, 329, 329, 333, 339, 365, 369, 368, 
    370, 329, 273, 253, 293, 335, 357, 370, 372, 370, 363, 369, 370, 374, 374, 
    380, 388, 389, 302, 175, 223, 332, 380, 383, 376, 367, 367, 365, 363, 358, 
    391, 413, 415, 412, 285, 120, 168, 272, 332, 351, 342, 366, 369, 368, 361, 
    398, 414, 414, 430, 292, 81, 99, 121, 141, 169, 186, 299, 335, 351, 356, 
    384, 397, 407, 395, 243, 155, 74, 117, 232, 149, 133, 124, 175, 286, 339, 
    345, 355, 360, 353, 344, 329, 263, 267, 308, 278, 275, 273, 267, 275, 286, 
    183, 166, 163, 163, 164, 150, 133, 141, 165, 154, 155, 154, 162, 165, 149, 
    136, 120, 122, 113, 124, 100, 92, 98, 111, 97, 88, 92, 86, 86, 107, 
    107, 86, 84, 87, 90, 75, 87, 92, 102, 92, 93, 94, 86, 153, 207, 
    
    -- channel=254
    192, 268, 262, 228, 220, 253, 250, 237, 244, 244, 251, 248, 250, 285, 286, 
    199, 258, 294, 277, 220, 234, 236, 230, 251, 242, 245, 225, 272, 294, 296, 
    195, 249, 294, 243, 241, 207, 225, 203, 234, 250, 231, 239, 254, 298, 298, 
    205, 247, 302, 230, 219, 227, 227, 232, 233, 255, 226, 244, 211, 284, 285, 
    235, 247, 265, 269, 214, 213, 212, 228, 231, 229, 217, 231, 282, 287, 283, 
    255, 267, 237, 255, 268, 264, 271, 283, 279, 268, 269, 271, 284, 285, 286, 
    259, 273, 206, 125, 164, 256, 289, 301, 300, 296, 286, 288, 286, 288, 285, 
    264, 302, 303, 258, 103, 98, 209, 289, 300, 292, 283, 285, 286, 285, 279, 
    272, 306, 312, 312, 223, 29, 40, 107, 180, 239, 261, 295, 291, 284, 281, 
    271, 304, 308, 316, 199, 0, 5, 32, 33, 40, 38, 128, 181, 241, 278, 
    257, 304, 303, 312, 217, 161, 54, 80, 198, 129, 114, 96, 117, 224, 256, 
    182, 222, 208, 197, 188, 188, 157, 168, 206, 196, 196, 203, 206, 211, 212, 
    91, 115, 111, 98, 87, 79, 75, 82, 96, 79, 79, 74, 81, 88, 64, 
    16, 20, 19, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 4, 0, 0, 0, 0, 19, 54, 
    
    -- channel=255
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=256
    84, 55, 95, 88, 23, 105, 94, 110, 137, 148, 92, 161, 70, 116, 91, 
    102, 88, 99, 91, 21, 94, 87, 110, 117, 121, 97, 174, 90, 119, 101, 
    100, 118, 94, 76, 25, 102, 118, 105, 126, 65, 138, 183, 135, 130, 125, 
    64, 138, 84, 61, 68, 168, 147, 73, 129, 67, 159, 200, 166, 141, 72, 
    69, 187, 84, 73, 145, 158, 72, 119, 155, 167, 173, 214, 172, 138, 23, 
    54, 183, 158, 58, 157, 149, 106, 162, 156, 164, 148, 197, 167, 149, 22, 
    61, 143, 169, 145, 141, 155, 134, 136, 132, 145, 134, 149, 157, 162, 52, 
    89, 144, 138, 152, 145, 97, 160, 158, 151, 136, 125, 167, 109, 152, 38, 
    121, 139, 133, 148, 173, 103, 149, 149, 146, 155, 156, 149, 129, 128, 65, 
    125, 126, 96, 142, 138, 173, 140, 144, 154, 144, 140, 142, 92, 81, 141, 
    80, 149, 99, 141, 130, 108, 194, 157, 138, 136, 140, 140, 120, 117, 146, 
    132, 176, 141, 153, 126, 149, 173, 175, 148, 118, 147, 145, 144, 161, 158, 
    167, 256, 218, 192, 148, 173, 172, 137, 173, 143, 156, 121, 114, 147, 160, 
    84, 154, 273, 239, 198, 187, 186, 127, 141, 159, 153, 126, 72, 138, 164, 
    90, 82, 185, 286, 243, 206, 200, 193, 149, 155, 153, 130, 78, 113, 236, 
    
    -- channel=257
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 53, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 
    5, 0, 0, 0, 0, 1, 58, 0, 0, 0, 0, 0, 0, 0, 54, 
    0, 0, 0, 0, 43, 61, 50, 35, 65, 77, 63, 20, 9, 0, 29, 
    0, 0, 0, 3, 61, 43, 64, 85, 72, 45, 58, 80, 69, 0, 21, 
    0, 0, 0, 0, 39, 92, 69, 92, 74, 88, 90, 65, 125, 38, 0, 
    0, 0, 0, 0, 0, 68, 82, 82, 97, 102, 80, 88, 86, 0, 0, 
    15, 0, 0, 0, 0, 0, 46, 92, 103, 116, 95, 92, 64, 0, 0, 
    0, 0, 0, 0, 0, 0, 50, 111, 99, 101, 89, 102, 65, 0, 0, 
    8, 12, 0, 0, 0, 0, 48, 130, 93, 100, 105, 98, 88, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 102, 95, 106, 88, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 9, 97, 114, 61, 0, 0, 0, 
    
    -- channel=258
    65, 26, 41, 6, 0, 17, 22, 23, 16, 12, 6, 69, 25, 17, 43, 
    80, 47, 18, 26, 0, 0, 0, 34, 32, 37, 9, 94, 78, 92, 62, 
    17, 10, 29, 25, 0, 41, 39, 0, 19, 0, 26, 110, 127, 67, 67, 
    0, 77, 58, 48, 24, 37, 0, 0, 44, 46, 89, 67, 102, 102, 51, 
    12, 103, 81, 24, 79, 57, 12, 53, 50, 59, 41, 17, 97, 106, 9, 
    14, 83, 94, 82, 67, 106, 134, 156, 87, 81, 69, 95, 79, 86, 13, 
    48, 87, 86, 99, 131, 172, 185, 177, 150, 177, 203, 196, 99, 83, 29, 
    32, 71, 100, 97, 225, 146, 194, 206, 232, 241, 215, 227, 213, 97, 0, 
    86, 98, 60, 63, 142, 236, 224, 235, 245, 226, 201, 226, 164, 93, 27, 
    88, 50, 16, 49, 76, 127, 247, 268, 249, 256, 218, 202, 159, 74, 68, 
    37, 69, 35, 73, 69, 100, 214, 269, 258, 215, 222, 207, 166, 105, 94, 
    141, 222, 84, 55, 48, 102, 216, 249, 247, 218, 256, 218, 134, 110, 16, 
    53, 92, 125, 68, 45, 86, 164, 152, 166, 248, 247, 218, 149, 44, 0, 
    25, 0, 42, 112, 78, 35, 40, 91, 148, 230, 233, 189, 68, 20, 42, 
    0, 3, 0, 57, 128, 110, 43, 46, 58, 151, 148, 131, 92, 76, 108, 
    
    -- channel=259
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 25, 0, 7, 15, 3, 12, 11, 44, 8, 0, 0, 
    0, 0, 0, 0, 25, 7, 26, 25, 45, 43, 6, 36, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 31, 71, 53, 59, 16, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 69, 83, 69, 31, 24, 10, 0, 0, 0, 
    0, 51, 0, 0, 0, 0, 67, 78, 57, 18, 56, 21, 0, 0, 0, 
    0, 23, 7, 0, 0, 0, 30, 0, 5, 43, 60, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 53, 44, 0, 0, 0, 0, 
    0, 0, 0, 9, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    
    -- channel=260
    92, 69, 97, 103, 76, 61, 101, 90, 132, 120, 123, 107, 140, 71, 90, 
    111, 113, 113, 108, 71, 62, 68, 93, 117, 124, 116, 115, 135, 108, 132, 
    118, 100, 103, 93, 62, 66, 126, 133, 100, 108, 95, 130, 168, 150, 147, 
    90, 106, 124, 87, 57, 153, 176, 75, 102, 85, 124, 190, 168, 155, 136, 
    110, 129, 151, 92, 106, 158, 116, 92, 148, 164, 183, 161, 174, 153, 113, 
    93, 119, 155, 140, 161, 133, 83, 137, 169, 154, 133, 167, 184, 150, 112, 
    107, 119, 145, 172, 129, 106, 104, 117, 104, 101, 98, 137, 143, 169, 117, 
    117, 122, 156, 159, 130, 96, 106, 115, 111, 117, 120, 105, 147, 142, 108, 
    119, 155, 138, 141, 131, 125, 106, 108, 130, 124, 115, 133, 99, 111, 112, 
    152, 129, 130, 130, 131, 96, 119, 130, 122, 132, 119, 123, 99, 100, 107, 
    131, 118, 128, 112, 149, 143, 117, 143, 133, 118, 111, 112, 109, 102, 172, 
    128, 188, 192, 163, 145, 127, 146, 133, 120, 119, 118, 116, 122, 129, 174, 
    156, 156, 214, 222, 181, 145, 143, 115, 89, 114, 118, 110, 107, 101, 186, 
    122, 111, 158, 208, 227, 205, 179, 131, 134, 121, 122, 116, 79, 123, 136, 
    121, 93, 108, 183, 207, 236, 226, 204, 147, 100, 104, 90, 111, 114, 196, 
    
    -- channel=261
    9, 28, 0, 0, 65, 0, 0, 0, 0, 0, 43, 0, 116, 0, 0, 
    13, 29, 18, 0, 73, 0, 0, 0, 15, 0, 39, 0, 121, 0, 23, 
    3, 0, 5, 10, 57, 0, 0, 6, 0, 44, 0, 0, 76, 7, 24, 
    45, 0, 36, 22, 1, 0, 15, 43, 0, 49, 0, 0, 45, 19, 83, 
    45, 0, 95, 31, 0, 0, 87, 0, 0, 0, 3, 0, 26, 18, 140, 
    66, 0, 15, 109, 0, 0, 35, 0, 16, 0, 19, 0, 45, 7, 153, 
    70, 0, 0, 37, 27, 0, 16, 0, 2, 0, 6, 0, 38, 0, 132, 
    37, 0, 0, 15, 16, 42, 0, 3, 18, 15, 9, 0, 62, 3, 118, 
    5, 0, 14, 3, 0, 59, 0, 13, 7, 3, 27, 0, 36, 18, 75, 
    10, 18, 33, 0, 2, 0, 5, 8, 17, 27, 18, 24, 64, 19, 0, 
    75, 0, 46, 0, 0, 21, 0, 20, 35, 33, 5, 19, 34, 11, 0, 
    14, 7, 87, 0, 39, 0, 0, 1, 21, 51, 0, 20, 28, 0, 18, 
    0, 0, 51, 57, 39, 0, 0, 29, 0, 18, 9, 43, 45, 0, 6, 
    42, 0, 0, 13, 65, 24, 0, 43, 0, 0, 8, 42, 78, 0, 0, 
    59, 5, 0, 0, 19, 54, 45, 10, 21, 0, 0, 24, 63, 1, 0, 
    
    -- channel=262
    81, 65, 79, 70, 33, 77, 70, 79, 83, 84, 63, 116, 48, 83, 78, 
    96, 83, 77, 74, 32, 68, 62, 86, 78, 92, 62, 131, 70, 109, 88, 
    65, 63, 75, 65, 36, 88, 96, 71, 82, 55, 76, 145, 98, 103, 85, 
    54, 114, 82, 65, 70, 105, 70, 49, 95, 69, 117, 132, 100, 107, 60, 
    64, 125, 80, 68, 101, 105, 62, 94, 105, 112, 102, 119, 112, 107, 30, 
    53, 115, 103, 87, 118, 112, 82, 122, 104, 109, 91, 131, 105, 105, 27, 
    68, 114, 115, 103, 100, 120, 117, 126, 104, 113, 121, 135, 97, 112, 49, 
    71, 107, 114, 103, 131, 117, 133, 124, 134, 144, 134, 134, 116, 99, 45, 
    99, 114, 93, 98, 132, 108, 138, 134, 144, 140, 122, 139, 94, 88, 54, 
    100, 86, 71, 85, 97, 120, 133, 145, 140, 136, 131, 122, 92, 84, 103, 
    67, 94, 72, 104, 108, 102, 151, 147, 134, 123, 127, 122, 104, 98, 110, 
    121, 156, 107, 115, 83, 118, 143, 138, 136, 116, 140, 124, 100, 108, 92, 
    100, 126, 126, 117, 102, 105, 130, 99, 121, 129, 141, 120, 93, 98, 83, 
    64, 83, 119, 133, 118, 115, 111, 104, 141, 135, 130, 110, 60, 81, 108, 
    51, 61, 105, 134, 134, 135, 120, 123, 92, 105, 102, 101, 94, 110, 152, 
    
    -- channel=263
    0, 27, 0, 0, 54, 0, 1, 0, 0, 0, 29, 0, 82, 0, 0, 
    0, 31, 9, 0, 70, 0, 0, 0, 0, 0, 21, 0, 65, 0, 5, 
    12, 0, 0, 11, 60, 0, 0, 18, 0, 48, 0, 0, 27, 0, 0, 
    27, 0, 26, 14, 13, 0, 17, 40, 0, 32, 0, 0, 7, 0, 45, 
    40, 0, 47, 35, 0, 0, 58, 0, 0, 0, 0, 0, 1, 0, 94, 
    63, 0, 0, 63, 0, 0, 36, 0, 1, 0, 5, 0, 24, 0, 113, 
    57, 0, 0, 7, 15, 0, 5, 0, 0, 0, 0, 0, 22, 0, 95, 
    26, 0, 0, 0, 0, 50, 0, 0, 0, 0, 1, 0, 27, 0, 98, 
    0, 0, 9, 0, 0, 17, 0, 0, 0, 0, 13, 0, 19, 10, 53, 
    2, 7, 34, 0, 0, 0, 0, 0, 0, 0, 2, 7, 34, 8, 0, 
    47, 0, 34, 0, 0, 1, 0, 0, 4, 11, 0, 1, 21, 0, 0, 
    0, 0, 54, 0, 19, 0, 0, 0, 0, 24, 0, 7, 18, 0, 0, 
    0, 0, 8, 34, 23, 0, 0, 27, 0, 0, 0, 17, 34, 0, 3, 
    24, 0, 0, 0, 31, 13, 0, 21, 0, 0, 0, 34, 68, 0, 0, 
    47, 0, 0, 0, 0, 11, 20, 0, 32, 0, 0, 1, 41, 0, 0, 
    
    -- channel=264
    207, 132, 177, 189, 125, 89, 190, 168, 254, 240, 246, 223, 300, 120, 181, 
    256, 230, 230, 208, 117, 77, 126, 166, 256, 241, 239, 240, 348, 231, 279, 
    224, 190, 209, 182, 93, 115, 240, 242, 202, 186, 203, 288, 429, 321, 338, 
    177, 222, 258, 169, 106, 289, 314, 119, 175, 195, 278, 367, 434, 367, 312, 
    212, 298, 356, 192, 218, 342, 238, 173, 319, 336, 381, 340, 417, 372, 255, 
    185, 263, 392, 315, 311, 304, 255, 339, 368, 339, 310, 344, 420, 363, 256, 
    228, 257, 339, 418, 331, 292, 292, 300, 284, 291, 305, 344, 359, 378, 286, 
    240, 271, 338, 390, 375, 259, 299, 347, 346, 342, 324, 353, 383, 342, 216, 
    284, 337, 314, 329, 348, 361, 324, 353, 367, 362, 360, 352, 333, 275, 233, 
    338, 286, 250, 269, 294, 303, 355, 391, 393, 399, 351, 355, 282, 219, 256, 
    282, 256, 270, 271, 311, 303, 356, 434, 408, 368, 334, 337, 305, 269, 376, 
    347, 476, 421, 327, 335, 313, 383, 408, 389, 366, 362, 351, 320, 298, 374, 
    324, 409, 532, 474, 371, 349, 386, 320, 279, 370, 385, 339, 292, 214, 360, 
    247, 161, 354, 517, 501, 410, 377, 327, 310, 358, 371, 336, 202, 209, 303, 
    255, 148, 178, 405, 537, 535, 482, 417, 322, 293, 295, 271, 260, 259, 405, 
    
    -- channel=265
    143, 118, 167, 238, 178, 149, 145, 152, 129, 132, 148, 159, 62, 109, 140, 
    173, 135, 178, 240, 151, 126, 143, 146, 150, 160, 138, 157, 64, 159, 175, 
    171, 136, 197, 209, 132, 123, 156, 173, 192, 145, 143, 157, 125, 187, 194, 
    159, 166, 164, 143, 116, 140, 133, 94, 163, 122, 118, 145, 158, 196, 183, 
    181, 238, 194, 119, 124, 129, 74, 128, 128, 128, 111, 99, 134, 228, 167, 
    140, 230, 253, 158, 134, 44, 33, 122, 102, 64, 50, 107, 118, 250, 126, 
    142, 197, 230, 197, 10, 0, 0, 0, 0, 0, 0, 0, 80, 223, 143, 
    164, 201, 215, 198, 10, 0, 0, 0, 0, 0, 0, 30, 24, 173, 130, 
    179, 200, 210, 201, 102, 34, 0, 0, 0, 0, 0, 0, 30, 109, 147, 
    221, 174, 173, 193, 145, 86, 16, 21, 0, 0, 0, 0, 4, 131, 187, 
    169, 147, 150, 194, 186, 137, 71, 29, 30, 0, 0, 0, 0, 153, 246, 
    157, 91, 58, 184, 199, 163, 54, 0, 30, 18, 0, 0, 0, 118, 247, 
    168, 115, 50, 67, 121, 195, 72, 0, 35, 7, 0, 0, 0, 96, 239, 
    127, 89, 92, 64, 48, 88, 81, 75, 85, 0, 0, 0, 0, 167, 175, 
    126, 75, 77, 85, 74, 75, 85, 81, 49, 28, 17, 4, 65, 123, 123, 
    
    -- channel=266
    75, 86, 90, 72, 58, 116, 91, 104, 101, 115, 80, 118, 63, 119, 100, 
    65, 90, 77, 69, 70, 119, 101, 110, 85, 94, 77, 120, 52, 90, 67, 
    98, 114, 85, 75, 85, 105, 87, 87, 93, 87, 99, 115, 52, 73, 61, 
    68, 91, 70, 80, 106, 100, 100, 106, 115, 75, 87, 124, 65, 67, 41, 
    71, 87, 37, 85, 122, 82, 72, 118, 79, 103, 94, 131, 85, 63, 26, 
    83, 99, 54, 36, 90, 109, 109, 85, 88, 103, 99, 134, 89, 61, 35, 
    73, 83, 84, 57, 101, 136, 128, 111, 118, 127, 113, 109, 102, 76, 43, 
    81, 89, 79, 67, 88, 123, 130, 126, 115, 109, 113, 116, 77, 91, 65, 
    77, 70, 79, 75, 108, 83, 115, 110, 111, 120, 122, 119, 95, 103, 74, 
    73, 85, 94, 97, 94, 114, 102, 94, 102, 96, 112, 110, 94, 88, 85, 
    59, 109, 78, 72, 79, 85, 110, 84, 90, 99, 112, 112, 105, 82, 63, 
    59, 58, 76, 93, 65, 81, 98, 110, 98, 86, 98, 118, 126, 129, 62, 
    110, 134, 88, 97, 90, 95, 93, 127, 137, 97, 100, 103, 117, 137, 83, 
    73, 159, 158, 103, 86, 109, 112, 88, 101, 111, 111, 114, 114, 128, 73, 
    74, 104, 152, 158, 100, 77, 91, 100, 124, 125, 129, 117, 82, 59, 121, 
    
    -- channel=267
    80, 37, 53, 58, 70, 0, 79, 49, 115, 99, 115, 37, 187, 43, 45, 
    96, 64, 96, 68, 62, 28, 56, 27, 103, 79, 118, 43, 178, 45, 119, 
    114, 88, 71, 79, 45, 0, 53, 105, 80, 101, 64, 66, 205, 114, 129, 
    82, 37, 100, 75, 1, 87, 141, 70, 24, 70, 91, 106, 217, 142, 191, 
    83, 88, 155, 84, 46, 136, 129, 0, 124, 100, 162, 125, 189, 153, 176, 
    97, 91, 155, 107, 96, 124, 115, 139, 149, 147, 145, 84, 201, 146, 168, 
    83, 86, 129, 170, 167, 153, 130, 148, 141, 146, 141, 146, 171, 137, 148, 
    98, 91, 110, 165, 171, 130, 139, 159, 174, 145, 144, 172, 178, 150, 136, 
    90, 115, 145, 144, 163, 153, 159, 178, 179, 178, 176, 172, 198, 157, 101, 
    131, 143, 108, 103, 141, 156, 166, 178, 188, 212, 164, 183, 172, 80, 57, 
    156, 78, 114, 98, 99, 117, 139, 219, 207, 196, 177, 174, 156, 101, 141, 
    82, 162, 162, 107, 153, 108, 178, 212, 200, 185, 175, 184, 177, 123, 148, 
    162, 197, 228, 177, 149, 138, 194, 224, 149, 185, 205, 184, 168, 83, 138, 
    127, 87, 157, 207, 199, 155, 155, 131, 93, 191, 181, 188, 170, 41, 96, 
    141, 55, 65, 172, 230, 202, 179, 161, 154, 170, 196, 148, 76, 82, 112, 
    
    -- channel=268
    0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=269
    98, 57, 103, 129, 56, 115, 107, 133, 155, 170, 116, 182, 68, 127, 95, 
    125, 95, 123, 131, 48, 110, 110, 122, 132, 143, 114, 195, 70, 114, 129, 
    152, 156, 122, 120, 49, 92, 112, 131, 166, 94, 146, 198, 140, 158, 150, 
    87, 136, 100, 90, 62, 163, 161, 90, 135, 82, 141, 206, 200, 174, 123, 
    98, 221, 116, 85, 158, 164, 61, 97, 151, 162, 190, 222, 185, 187, 72, 
    87, 228, 210, 75, 142, 136, 85, 173, 153, 151, 124, 183, 179, 211, 42, 
    76, 171, 216, 189, 130, 124, 90, 109, 113, 127, 121, 132, 145, 201, 75, 
    123, 176, 181, 197, 131, 70, 136, 120, 117, 87, 98, 167, 106, 177, 80, 
    141, 164, 185, 197, 207, 110, 129, 134, 125, 136, 125, 146, 150, 172, 90, 
    174, 181, 137, 185, 172, 197, 152, 143, 144, 141, 130, 126, 88, 96, 152, 
    132, 158, 112, 170, 159, 143, 190, 168, 147, 141, 142, 117, 101, 134, 193, 
    133, 145, 104, 167, 165, 174, 187, 165, 159, 122, 135, 121, 121, 171, 212, 
    232, 305, 210, 159, 154, 199, 202, 156, 205, 142, 150, 108, 86, 163, 207, 
    109, 184, 303, 228, 159, 175, 184, 120, 140, 163, 149, 114, 83, 162, 189, 
    112, 77, 192, 306, 245, 180, 174, 180, 144, 177, 187, 141, 56, 104, 214, 
    
    -- channel=270
    0, 19, 0, 0, 53, 0, 5, 0, 0, 0, 39, 0, 106, 0, 0, 
    0, 18, 13, 0, 62, 0, 0, 0, 10, 0, 36, 0, 95, 0, 17, 
    13, 7, 2, 2, 54, 0, 0, 14, 0, 36, 0, 0, 51, 0, 7, 
    35, 0, 13, 24, 0, 0, 30, 44, 0, 40, 0, 0, 25, 0, 65, 
    34, 0, 66, 13, 0, 0, 69, 0, 0, 0, 9, 0, 8, 0, 115, 
    59, 0, 0, 74, 0, 0, 25, 0, 8, 0, 8, 0, 41, 0, 130, 
    54, 0, 0, 9, 5, 0, 2, 0, 0, 0, 0, 0, 23, 0, 103, 
    32, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 34, 0, 92, 
    0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 1, 0, 17, 24, 74, 
    0, 13, 31, 0, 0, 0, 0, 0, 0, 0, 0, 1, 47, 10, 0, 
    56, 0, 40, 0, 0, 15, 0, 0, 1, 0, 0, 0, 20, 0, 0, 
    0, 0, 64, 0, 22, 0, 0, 0, 0, 17, 0, 0, 28, 0, 13, 
    0, 0, 37, 39, 34, 0, 0, 27, 0, 0, 0, 19, 34, 0, 9, 
    35, 0, 0, 2, 47, 19, 0, 37, 0, 0, 0, 23, 84, 0, 0, 
    59, 24, 0, 0, 9, 33, 31, 0, 10, 0, 0, 24, 43, 0, 0, 
    
    -- channel=271
    194, 97, 191, 182, 51, 153, 164, 165, 208, 216, 181, 268, 157, 150, 179, 
    221, 173, 186, 199, 29, 102, 123, 182, 225, 216, 178, 300, 242, 250, 229, 
    158, 183, 195, 137, 27, 177, 241, 176, 211, 88, 251, 318, 338, 282, 291, 
    129, 296, 185, 138, 103, 302, 231, 55, 222, 163, 298, 356, 363, 319, 194, 
    141, 369, 275, 108, 261, 296, 128, 227, 282, 315, 312, 294, 345, 322, 104, 
    87, 326, 362, 224, 305, 255, 196, 332, 300, 279, 245, 347, 315, 333, 104, 
    158, 280, 319, 340, 236, 240, 253, 245, 231, 247, 265, 293, 288, 340, 154, 
    181, 284, 308, 332, 351, 127, 284, 291, 290, 292, 251, 334, 285, 311, 65, 
    270, 299, 240, 279, 276, 326, 262, 293, 301, 304, 286, 286, 228, 198, 173, 
    277, 213, 180, 269, 273, 248, 314, 346, 316, 321, 281, 276, 206, 194, 274, 
    171, 286, 198, 281, 251, 266, 371, 352, 338, 270, 278, 275, 232, 248, 339, 
    348, 447, 310, 292, 273, 282, 351, 347, 320, 271, 325, 269, 228, 282, 317, 
    252, 399, 445, 366, 288, 335, 303, 190, 269, 321, 306, 248, 202, 188, 293, 
    176, 117, 390, 466, 380, 330, 315, 285, 271, 305, 325, 220, 82, 241, 323, 
    159, 141, 177, 415, 474, 431, 380, 350, 226, 246, 219, 228, 205, 254, 425, 
    
    -- channel=272
    173, 82, 130, 144, 46, 56, 132, 137, 194, 203, 180, 229, 201, 93, 150, 
    240, 185, 170, 177, 41, 38, 89, 135, 204, 196, 169, 259, 273, 204, 237, 
    200, 172, 182, 161, 32, 73, 169, 167, 184, 129, 167, 306, 401, 289, 297, 
    112, 199, 214, 143, 72, 218, 198, 43, 152, 159, 241, 338, 422, 361, 272, 
    154, 320, 319, 139, 205, 289, 154, 137, 243, 277, 300, 297, 396, 381, 185, 
    145, 289, 397, 255, 259, 292, 267, 348, 333, 306, 279, 335, 375, 376, 172, 
    184, 256, 362, 412, 328, 319, 310, 323, 313, 338, 353, 376, 358, 370, 212, 
    207, 270, 347, 398, 421, 267, 346, 386, 389, 377, 363, 447, 409, 358, 155, 
    275, 321, 316, 329, 386, 418, 387, 422, 428, 430, 408, 414, 379, 286, 185, 
    332, 281, 217, 263, 305, 353, 432, 480, 470, 473, 412, 401, 306, 207, 239, 
    251, 254, 215, 256, 275, 302, 436, 518, 503, 431, 407, 389, 323, 276, 363, 
    348, 466, 331, 283, 312, 313, 448, 495, 482, 427, 432, 403, 312, 316, 328, 
    333, 453, 497, 382, 298, 358, 416, 358, 370, 456, 463, 389, 299, 205, 290, 
    192, 130, 370, 486, 405, 319, 317, 284, 316, 435, 454, 373, 188, 175, 265, 
    174, 62, 132, 401, 519, 460, 379, 336, 295, 337, 353, 300, 207, 205, 386, 
    
    -- channel=273
    134, 76, 105, 110, 103, 17, 132, 83, 159, 138, 181, 83, 262, 36, 103, 
    145, 137, 149, 123, 96, 19, 66, 70, 174, 140, 175, 83, 279, 120, 188, 
    153, 121, 129, 106, 71, 31, 138, 167, 106, 120, 116, 114, 314, 193, 234, 
    118, 95, 165, 114, 37, 160, 223, 72, 68, 133, 139, 197, 307, 232, 250, 
    143, 145, 264, 121, 119, 213, 171, 71, 197, 204, 256, 179, 278, 240, 227, 
    138, 122, 255, 219, 161, 171, 189, 216, 237, 203, 194, 183, 295, 222, 240, 
    160, 125, 179, 276, 221, 187, 185, 172, 174, 188, 192, 197, 238, 227, 240, 
    156, 142, 190, 254, 251, 143, 167, 227, 229, 203, 192, 217, 264, 220, 162, 
    168, 196, 193, 197, 196, 274, 186, 224, 223, 213, 233, 219, 236, 189, 184, 
    217, 177, 164, 164, 187, 156, 237, 244, 244, 268, 214, 235, 207, 131, 128, 
    198, 142, 191, 145, 177, 198, 180, 279, 270, 236, 212, 215, 207, 160, 237, 
    195, 296, 291, 186, 224, 165, 229, 261, 249, 245, 227, 232, 221, 191, 232, 
    194, 237, 364, 320, 250, 222, 242, 235, 155, 243, 239, 224, 215, 100, 236, 
    174, 59, 185, 338, 341, 263, 237, 225, 150, 224, 240, 232, 168, 117, 157, 
    206, 107, 46, 227, 362, 352, 315, 252, 214, 199, 203, 178, 166, 124, 197, 
    
    -- channel=274
    165, 173, 205, 209, 178, 203, 188, 192, 202, 185, 177, 190, 159, 172, 162, 
    170, 187, 201, 196, 168, 191, 165, 190, 190, 202, 182, 191, 141, 201, 192, 
    161, 160, 173, 174, 157, 199, 233, 219, 184, 170, 178, 196, 146, 195, 183, 
    183, 198, 178, 150, 170, 256, 238, 164, 195, 151, 219, 226, 150, 172, 149, 
    186, 202, 163, 169, 187, 206, 159, 196, 232, 226, 221, 210, 170, 161, 140, 
    158, 195, 178, 172, 226, 125, 110, 175, 186, 160, 152, 200, 174, 176, 144, 
    164, 194, 182, 167, 117, 84, 82, 102, 83, 75, 74, 105, 138, 201, 146, 
    164, 185, 172, 159, 67, 86, 62, 66, 67, 72, 74, 61, 79, 165, 142, 
    174, 195, 173, 171, 112, 45, 75, 51, 55, 40, 58, 72, 62, 140, 158, 
    177, 158, 165, 174, 143, 107, 51, 51, 48, 46, 51, 63, 68, 142, 186, 
    154, 170, 188, 193, 199, 136, 91, 55, 39, 48, 49, 53, 90, 159, 215, 
    158, 186, 209, 226, 175, 166, 91, 39, 46, 52, 52, 53, 100, 157, 229, 
    162, 143, 170, 226, 210, 184, 112, 59, 58, 42, 54, 46, 78, 174, 236, 
    163, 182, 164, 172, 222, 234, 203, 148, 148, 50, 47, 57, 86, 196, 204, 
    184, 187, 218, 190, 168, 213, 238, 213, 148, 81, 73, 77, 146, 205, 232, 
    
    -- channel=275
    49, 42, 2, 13, 104, 0, 28, 0, 0, 0, 60, 0, 152, 0, 8, 
    36, 11, 38, 22, 98, 0, 25, 0, 24, 0, 63, 0, 141, 0, 48, 
    38, 4, 26, 49, 79, 0, 0, 20, 0, 70, 0, 0, 104, 5, 38, 
    66, 0, 56, 63, 0, 0, 0, 53, 0, 57, 0, 0, 72, 27, 153, 
    55, 0, 103, 56, 0, 0, 107, 0, 0, 0, 0, 0, 33, 41, 202, 
    88, 0, 26, 86, 0, 0, 71, 4, 11, 8, 38, 0, 46, 21, 198, 
    67, 0, 0, 36, 58, 30, 41, 43, 49, 41, 49, 27, 54, 0, 151, 
    44, 0, 0, 28, 59, 68, 15, 42, 63, 48, 51, 40, 107, 27, 136, 
    9, 0, 34, 18, 1, 97, 44, 70, 59, 53, 60, 49, 108, 70, 75, 
    26, 41, 37, 0, 25, 13, 61, 63, 71, 97, 59, 76, 130, 45, 0, 
    106, 0, 50, 0, 0, 25, 0, 86, 96, 96, 68, 74, 82, 30, 6, 
    0, 3, 38, 0, 50, 0, 21, 66, 88, 104, 64, 75, 60, 0, 0, 
    0, 0, 10, 0, 4, 0, 29, 108, 14, 81, 81, 99, 97, 0, 0, 
    73, 0, 0, 0, 3, 0, 0, 38, 0, 62, 59, 97, 141, 0, 0, 
    83, 15, 0, 0, 0, 0, 0, 0, 16, 44, 67, 61, 52, 9, 0, 
    
    -- channel=276
    7, 0, 64, 47, 0, 111, 19, 53, 29, 22, 0, 113, 0, 70, 21, 
    7, 5, 10, 45, 0, 91, 15, 77, 0, 51, 0, 146, 0, 87, 2, 
    12, 4, 20, 23, 0, 76, 53, 28, 42, 0, 27, 133, 0, 22, 0, 
    0, 98, 0, 0, 18, 85, 0, 0, 117, 0, 68, 92, 0, 4, 0, 
    0, 132, 0, 0, 78, 11, 0, 86, 11, 39, 0, 34, 0, 7, 0, 
    0, 141, 0, 0, 81, 0, 0, 46, 0, 0, 0, 87, 0, 15, 0, 
    0, 98, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 
    0, 67, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    19, 48, 10, 1, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 0, 0, 50, 0, 32, 0, 0, 0, 0, 0, 0, 0, 2, 53, 
    0, 51, 0, 46, 50, 0, 57, 0, 0, 0, 0, 0, 0, 2, 51, 
    0, 12, 0, 61, 0, 43, 14, 0, 0, 0, 0, 0, 0, 32, 0, 
    42, 22, 0, 0, 0, 44, 0, 0, 7, 0, 0, 0, 0, 39, 23, 
    0, 93, 55, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 99, 5, 
    0, 0, 142, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 132, 
    
    -- channel=277
    4, 21, 10, 6, 29, 16, 5, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 28, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 23, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 2, 0, 11, 20, 0, 0, 12, 0, 19, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 1, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    
    -- channel=278
    0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    7, 8, 0, 1, 0, 0, 0, 0, 5, 3, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 10, 2, 10, 
    0, 2, 3, 0, 0, 0, 0, 0, 3, 0, 0, 13, 1, 3, 7, 
    2, 5, 8, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 14, 2, 
    0, 0, 11, 7, 1, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 8, 
    0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    1, 12, 3, 3, 17, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 14, 0, 2, 0, 0, 0, 0, 0, 0, 7, 10, 
    18, 26, 13, 0, 0, 11, 6, 13, 9, 0, 2, 0, 0, 0, 11, 
    3, 5, 23, 6, 0, 0, 2, 0, 0, 0, 0, 0, 7, 0, 0, 
    1, 0, 0, 21, 13, 0, 0, 0, 3, 2, 20, 0, 0, 0, 0, 
    
    -- channel=279
    77, 65, 70, 45, 63, 71, 88, 70, 98, 92, 94, 70, 129, 81, 75, 
    54, 68, 66, 49, 67, 83, 75, 70, 85, 79, 92, 71, 110, 66, 75, 
    92, 100, 66, 52, 71, 65, 69, 84, 64, 77, 90, 63, 104, 67, 85, 
    62, 59, 70, 85, 58, 87, 115, 85, 75, 81, 78, 93, 102, 75, 91, 
    65, 58, 72, 75, 101, 97, 96, 74, 83, 92, 120, 99, 103, 63, 81, 
    79, 65, 56, 61, 80, 123, 125, 112, 111, 123, 116, 107, 110, 58, 94, 
    72, 60, 51, 83, 142, 162, 154, 134, 139, 147, 136, 135, 108, 64, 84, 
    73, 59, 61, 78, 139, 112, 148, 158, 157, 140, 134, 122, 137, 85, 75, 
    62, 63, 61, 63, 96, 150, 125, 139, 146, 145, 146, 142, 128, 107, 88, 
    71, 74, 80, 88, 90, 87, 139, 128, 130, 144, 135, 144, 128, 78, 49, 
    79, 92, 83, 54, 64, 98, 100, 128, 129, 130, 144, 145, 133, 62, 64, 
    59, 106, 110, 69, 72, 65, 129, 152, 122, 125, 144, 155, 160, 109, 50, 
    101, 118, 143, 128, 102, 84, 117, 160, 128, 134, 131, 144, 157, 82, 78, 
    100, 108, 132, 139, 130, 114, 109, 99, 82, 143, 143, 149, 133, 101, 64, 
    101, 110, 98, 140, 140, 121, 117, 113, 128, 143, 148, 121, 84, 52, 95, 
    
    -- channel=280
    106, 76, 82, 106, 116, 18, 110, 79, 156, 147, 171, 74, 234, 72, 99, 
    130, 120, 138, 117, 110, 48, 91, 80, 139, 123, 162, 74, 221, 70, 158, 
    171, 130, 128, 122, 91, 26, 95, 149, 112, 166, 102, 96, 249, 171, 181, 
    131, 69, 156, 114, 48, 123, 213, 129, 82, 103, 118, 175, 247, 190, 240, 
    136, 111, 208, 130, 71, 176, 196, 42, 151, 149, 210, 183, 239, 205, 229, 
    150, 112, 200, 169, 146, 158, 127, 125, 199, 193, 193, 142, 259, 190, 218, 
    134, 115, 175, 222, 187, 152, 136, 172, 169, 146, 135, 179, 219, 198, 196, 
    160, 131, 177, 218, 152, 167, 145, 166, 154, 154, 175, 153, 215, 205, 204, 
    130, 169, 193, 191, 182, 166, 147, 168, 192, 201, 189, 184, 209, 180, 155, 
    184, 190, 179, 156, 174, 152, 164, 180, 194, 211, 182, 197, 185, 137, 110, 
    215, 118, 169, 118, 170, 166, 137, 219, 213, 210, 182, 183, 175, 131, 186, 
    125, 178, 234, 172, 192, 156, 180, 214, 208, 199, 170, 189, 193, 159, 218, 
    220, 218, 275, 261, 223, 160, 193, 229, 145, 181, 190, 192, 186, 135, 223, 
    176, 154, 197, 252, 281, 231, 220, 166, 128, 185, 187, 206, 189, 108, 147, 
    180, 89, 109, 210, 263, 280, 268, 240, 210, 165, 184, 163, 136, 125, 165, 
    
    -- channel=281
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 19, 0, 0, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 5, 6, 0, 
    0, 33, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 25, 0, 0, 0, 44, 107, 92, 0, 0, 0, 22, 0, 0, 0, 
    0, 11, 0, 14, 73, 139, 149, 115, 112, 157, 176, 124, 20, 0, 0, 
    0, 0, 0, 21, 184, 101, 168, 190, 195, 188, 159, 217, 131, 12, 0, 
    8, 0, 0, 0, 93, 191, 199, 209, 193, 186, 176, 169, 133, 23, 0, 
    0, 0, 0, 0, 5, 123, 197, 227, 216, 207, 179, 162, 102, 13, 0, 
    0, 15, 0, 0, 0, 15, 194, 206, 216, 179, 183, 174, 107, 28, 0, 
    60, 116, 0, 0, 0, 26, 161, 214, 202, 176, 215, 190, 94, 32, 0, 
    0, 41, 13, 0, 0, 30, 108, 119, 159, 211, 220, 172, 117, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 5, 89, 196, 206, 149, 17, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 130, 134, 82, 6, 0, 24, 
    
    -- channel=282
    0, 0, 16, 0, 0, 77, 0, 17, 0, 4, 0, 96, 0, 65, 0, 
    0, 0, 0, 0, 0, 61, 0, 38, 0, 0, 0, 135, 0, 51, 0, 
    0, 0, 0, 0, 0, 52, 0, 0, 18, 0, 32, 125, 0, 0, 0, 
    0, 88, 0, 0, 0, 47, 0, 0, 85, 0, 71, 58, 0, 0, 0, 
    0, 132, 0, 0, 50, 0, 0, 49, 0, 9, 0, 30, 0, 0, 0, 
    0, 141, 0, 0, 42, 0, 0, 30, 0, 0, 0, 64, 0, 0, 0, 
    0, 78, 46, 0, 0, 17, 0, 16, 0, 22, 10, 8, 0, 7, 0, 
    0, 52, 7, 0, 0, 0, 54, 14, 0, 2, 0, 68, 0, 2, 0, 
    0, 1, 0, 0, 63, 0, 54, 14, 14, 22, 0, 16, 0, 0, 0, 
    0, 0, 0, 27, 3, 103, 0, 26, 13, 0, 0, 0, 0, 0, 36, 
    0, 45, 0, 40, 0, 0, 132, 0, 0, 0, 9, 0, 0, 0, 1, 
    0, 3, 0, 5, 0, 39, 53, 25, 9, 0, 26, 0, 0, 22, 0, 
    28, 93, 0, 0, 0, 43, 21, 0, 82, 0, 32, 0, 0, 23, 0, 
    0, 74, 125, 0, 0, 0, 0, 0, 59, 38, 15, 0, 0, 42, 0, 
    0, 0, 137, 116, 0, 0, 0, 0, 0, 38, 31, 0, 0, 0, 132, 
    
    -- channel=283
    107, 36, 58, 28, 0, 5, 68, 53, 93, 90, 88, 100, 148, 31, 64, 
    121, 82, 74, 51, 0, 0, 27, 39, 114, 89, 92, 118, 210, 112, 127, 
    76, 78, 66, 42, 0, 29, 82, 66, 70, 25, 90, 147, 263, 136, 160, 
    35, 100, 100, 71, 12, 112, 85, 0, 41, 102, 135, 158, 259, 191, 146, 
    53, 152, 181, 61, 125, 163, 83, 58, 149, 152, 178, 146, 232, 191, 100, 
    57, 126, 202, 146, 125, 189, 208, 246, 195, 183, 171, 176, 222, 182, 110, 
    98, 117, 156, 224, 238, 270, 276, 236, 225, 265, 286, 262, 219, 169, 135, 
    86, 120, 153, 208, 345, 190, 278, 315, 346, 314, 267, 330, 301, 182, 56, 
    142, 154, 134, 153, 228, 341, 294, 339, 328, 320, 319, 305, 269, 182, 100, 
    158, 126, 81, 114, 172, 217, 336, 354, 350, 362, 307, 306, 242, 103, 104, 
    117, 133, 105, 130, 112, 176, 291, 375, 362, 317, 310, 307, 248, 153, 177, 
    207, 328, 218, 114, 157, 156, 313, 370, 343, 312, 341, 322, 264, 187, 125, 
    145, 265, 339, 235, 158, 192, 285, 274, 264, 346, 352, 311, 248, 91, 100, 
    99, 7, 202, 323, 256, 178, 175, 201, 188, 328, 341, 288, 156, 64, 124, 
    102, 53, 27, 234, 349, 286, 213, 189, 171, 254, 264, 231, 143, 106, 202, 
    
    -- channel=284
    166, 120, 129, 151, 148, 50, 144, 107, 145, 138, 182, 100, 243, 63, 124, 
    186, 151, 173, 162, 136, 41, 102, 86, 186, 146, 186, 95, 292, 139, 207, 
    140, 129, 153, 141, 114, 79, 151, 157, 144, 128, 139, 121, 308, 206, 231, 
    160, 135, 172, 148, 83, 153, 179, 106, 65, 183, 154, 150, 295, 238, 254, 
    169, 167, 295, 128, 124, 208, 191, 86, 207, 180, 213, 155, 251, 250, 255, 
    158, 133, 275, 269, 154, 152, 172, 220, 220, 183, 185, 144, 255, 244, 259, 
    187, 148, 191, 274, 191, 152, 164, 149, 145, 158, 184, 173, 221, 223, 265, 
    175, 162, 198, 244, 255, 120, 146, 178, 213, 189, 157, 204, 247, 212, 189, 
    196, 204, 197, 209, 166, 271, 164, 209, 195, 182, 195, 180, 205, 182, 210, 
    212, 190, 164, 157, 199, 134, 225, 230, 219, 242, 192, 202, 208, 150, 157, 
    217, 146, 193, 188, 170, 209, 166, 258, 253, 210, 192, 191, 189, 186, 243, 
    236, 293, 269, 170, 240, 172, 207, 221, 231, 231, 211, 191, 179, 166, 243, 
    154, 195, 323, 262, 221, 200, 219, 176, 137, 233, 217, 206, 176, 100, 211, 
    181, 11, 136, 292, 287, 218, 191, 230, 139, 194, 215, 187, 159, 93, 209, 
    201, 122, 11, 158, 311, 313, 268, 216, 151, 161, 161, 185, 188, 179, 150, 
    
    -- channel=285
    229, 99, 206, 216, 58, 136, 188, 198, 262, 264, 212, 324, 187, 163, 185, 
    297, 205, 236, 249, 32, 108, 138, 193, 264, 267, 207, 371, 270, 292, 298, 
    232, 211, 234, 205, 20, 141, 248, 228, 266, 137, 244, 422, 438, 358, 361, 
    139, 308, 252, 165, 85, 327, 258, 49, 231, 175, 342, 432, 491, 432, 296, 
    182, 467, 347, 158, 284, 372, 146, 195, 337, 352, 377, 383, 461, 452, 165, 
    138, 432, 484, 260, 354, 333, 264, 449, 380, 361, 306, 408, 422, 467, 138, 
    189, 367, 459, 471, 342, 330, 312, 341, 313, 354, 370, 401, 386, 453, 201, 
    227, 364, 415, 457, 461, 231, 373, 394, 402, 383, 357, 491, 403, 415, 124, 
    338, 402, 373, 394, 449, 408, 416, 436, 433, 431, 401, 437, 369, 324, 181, 
    398, 322, 241, 334, 361, 426, 448, 503, 481, 482, 410, 403, 291, 230, 316, 
    265, 328, 242, 360, 336, 333, 522, 544, 509, 432, 411, 387, 321, 325, 462, 
    407, 559, 352, 367, 372, 385, 512, 513, 497, 414, 457, 398, 306, 376, 408, 
    393, 554, 549, 428, 343, 452, 475, 345, 417, 466, 491, 367, 278, 251, 371, 
    215, 179, 479, 566, 443, 380, 371, 318, 374, 467, 464, 349, 144, 246, 356, 
    196, 94, 229, 523, 601, 517, 435, 409, 309, 373, 379, 301, 209, 278, 519, 
    
    -- channel=286
    8, 38, 0, 0, 209, 0, 0, 0, 0, 0, 115, 0, 395, 0, 0, 
    0, 0, 20, 0, 205, 0, 0, 0, 4, 0, 125, 0, 352, 0, 35, 
    5, 0, 0, 0, 151, 0, 0, 0, 0, 118, 0, 0, 187, 0, 7, 
    120, 0, 43, 58, 0, 0, 36, 137, 0, 91, 0, 0, 93, 0, 284, 
    76, 0, 199, 60, 0, 0, 271, 0, 0, 0, 0, 0, 16, 0, 461, 
    158, 0, 0, 193, 0, 0, 46, 0, 0, 0, 46, 0, 83, 0, 479, 
    112, 0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 55, 0, 357, 
    48, 0, 0, 0, 0, 57, 0, 0, 19, 0, 0, 0, 122, 0, 326, 
    0, 0, 0, 0, 0, 88, 0, 0, 0, 0, 18, 0, 103, 37, 169, 
    0, 11, 35, 0, 0, 0, 0, 0, 0, 48, 0, 41, 195, 0, 0, 
    198, 0, 81, 0, 0, 0, 0, 2, 30, 56, 0, 32, 84, 0, 0, 
    0, 0, 151, 0, 49, 0, 0, 0, 0, 85, 0, 30, 87, 0, 0, 
    0, 0, 39, 43, 36, 0, 0, 132, 0, 1, 0, 97, 138, 0, 0, 
    134, 0, 0, 0, 89, 0, 0, 66, 0, 0, 0, 105, 289, 0, 0, 
    195, 33, 0, 0, 0, 25, 19, 0, 1, 0, 0, 54, 88, 0, 0, 
    
    -- channel=287
    3, 20, 18, 6, 19, 44, 11, 22, 7, 2, 0, 6, 0, 32, 0, 
    0, 0, 0, 0, 19, 49, 22, 14, 0, 3, 0, 5, 0, 9, 0, 
    0, 2, 0, 5, 20, 34, 10, 7, 4, 6, 9, 0, 0, 0, 0, 
    11, 7, 0, 0, 22, 18, 0, 16, 10, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 13, 6, 0, 0, 14, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 22, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=288
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 17, 
    8, 0, 0, 0, 0, 19, 65, 0, 0, 0, 13, 0, 0, 0, 21, 
    0, 0, 0, 0, 54, 82, 89, 69, 79, 74, 73, 54, 22, 0, 13, 
    0, 0, 0, 0, 42, 108, 78, 93, 94, 89, 92, 64, 67, 0, 23, 
    0, 0, 0, 0, 32, 60, 82, 95, 91, 102, 103, 82, 99, 39, 0, 
    0, 0, 0, 0, 0, 51, 78, 67, 98, 90, 93, 89, 82, 0, 0, 
    0, 0, 0, 0, 0, 0, 31, 82, 77, 103, 93, 99, 78, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 96, 91, 88, 80, 103, 91, 0, 0, 
    0, 0, 0, 0, 0, 0, 32, 116, 81, 86, 93, 113, 89, 15, 0, 
    0, 1, 0, 0, 0, 0, 0, 9, 1, 86, 81, 113, 100, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 71, 84, 76, 20, 0, 0, 
    
    -- channel=289
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=290
    14, 0, 26, 4, 0, 23, 5, 0, 15, 2, 0, 10, 0, 26, 0, 
    0, 0, 0, 9, 0, 29, 6, 0, 8, 4, 0, 28, 0, 20, 7, 
    0, 0, 0, 0, 0, 18, 9, 0, 11, 0, 39, 16, 12, 1, 9, 
    0, 49, 0, 0, 0, 48, 4, 0, 29, 0, 57, 11, 19, 4, 11, 
    0, 70, 0, 0, 14, 13, 0, 2, 24, 8, 14, 0, 9, 4, 0, 
    0, 69, 8, 0, 43, 0, 0, 38, 2, 6, 2, 4, 0, 12, 0, 
    0, 44, 13, 0, 0, 2, 0, 8, 0, 1, 0, 4, 0, 10, 0, 
    0, 24, 0, 4, 22, 0, 19, 0, 0, 0, 0, 14, 0, 13, 0, 
    0, 7, 0, 0, 0, 0, 4, 0, 5, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 18, 10, 0, 10, 0, 7, 0, 0, 0, 0, 2, 
    0, 26, 0, 30, 0, 0, 40, 1, 1, 0, 0, 0, 0, 0, 31, 
    0, 44, 0, 0, 0, 2, 31, 13, 0, 0, 20, 0, 0, 8, 0, 
    10, 26, 0, 0, 0, 21, 3, 0, 2, 0, 10, 0, 0, 0, 2, 
    6, 5, 53, 9, 0, 0, 0, 0, 0, 18, 1, 0, 0, 18, 7, 
    0, 4, 36, 47, 8, 0, 0, 9, 0, 11, 9, 0, 0, 21, 66, 
    
    -- channel=291
    72, 28, 56, 0, 0, 57, 42, 31, 54, 37, 31, 63, 77, 60, 54, 
    40, 32, 14, 0, 0, 48, 26, 49, 47, 41, 38, 85, 104, 86, 43, 
    26, 33, 17, 0, 0, 74, 54, 18, 8, 0, 87, 77, 117, 38, 66, 
    0, 91, 45, 39, 25, 83, 25, 0, 84, 33, 120, 74, 94, 57, 39, 
    0, 84, 29, 42, 95, 66, 32, 87, 69, 82, 88, 39, 95, 45, 4, 
    0, 80, 37, 17, 95, 131, 152, 136, 89, 102, 107, 103, 81, 28, 18, 
    22, 70, 32, 56, 151, 215, 224, 194, 186, 201, 201, 191, 104, 41, 18, 
    13, 52, 44, 64, 210, 151, 232, 249, 242, 248, 219, 206, 187, 71, 0, 
    52, 53, 8, 28, 132, 198, 216, 227, 239, 237, 228, 204, 178, 78, 14, 
    42, 15, 5, 58, 54, 143, 209, 224, 230, 230, 209, 212, 159, 70, 61, 
    3, 91, 30, 54, 49, 59, 215, 219, 207, 209, 213, 226, 183, 67, 43, 
    96, 188, 97, 38, 18, 86, 193, 249, 203, 187, 251, 237, 200, 98, 0, 
    50, 121, 140, 98, 50, 71, 151, 183, 172, 219, 232, 218, 193, 53, 0, 
    50, 40, 126, 144, 112, 66, 85, 104, 132, 225, 220, 205, 101, 74, 24, 
    37, 67, 83, 132, 146, 110, 78, 86, 98, 186, 166, 144, 97, 73, 146, 
    
    -- channel=292
    9, 27, 20, 8, 31, 38, 20, 20, 10, 2, 8, 0, 11, 19, 17, 
    0, 14, 5, 5, 38, 40, 20, 20, 0, 6, 8, 0, 0, 7, 0, 
    12, 9, 4, 14, 39, 23, 5, 18, 0, 21, 8, 0, 0, 0, 0, 
    12, 0, 5, 11, 30, 0, 10, 20, 19, 2, 0, 0, 0, 0, 0, 
    14, 0, 0, 28, 8, 0, 4, 28, 0, 0, 0, 0, 0, 0, 4, 
    18, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 11, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 
    5, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 28, 0, 
    17, 29, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=293
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 35, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 54, 0, 5, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 3, 46, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 48, 89, 
    0, 21, 55, 0, 0, 9, 0, 0, 0, 0, 13, 0, 64, 67, 79, 
    0, 21, 89, 0, 0, 0, 10, 25, 10, 4, 14, 0, 53, 76, 51, 
    0, 0, 41, 81, 33, 3, 0, 0, 15, 22, 22, 5, 45, 36, 51, 
    0, 2, 12, 84, 56, 0, 12, 37, 33, 0, 2, 70, 51, 45, 9, 
    1, 10, 41, 53, 57, 59, 29, 60, 35, 47, 52, 30, 101, 44, 0, 
    36, 31, 0, 14, 30, 72, 55, 67, 79, 84, 42, 53, 39, 0, 0, 
    45, 0, 0, 16, 0, 0, 58, 103, 94, 87, 52, 47, 24, 7, 39, 
    15, 32, 0, 0, 51, 25, 62, 94, 93, 77, 60, 49, 21, 0, 43, 
    44, 98, 81, 3, 0, 43, 76, 73, 62, 78, 88, 49, 23, 0, 21, 
    8, 0, 45, 72, 22, 0, 0, 5, 0, 72, 68, 49, 12, 0, 0, 
    19, 0, 0, 40, 97, 35, 5, 0, 3, 59, 73, 30, 0, 0, 0, 
    
    -- channel=294
    109, 27, 65, 62, 5, 27, 77, 81, 150, 153, 119, 147, 157, 86, 85, 
    149, 86, 102, 89, 0, 34, 67, 77, 131, 119, 122, 171, 202, 110, 140, 
    140, 116, 101, 93, 0, 37, 80, 95, 119, 80, 139, 199, 295, 175, 200, 
    61, 121, 134, 76, 13, 142, 142, 36, 108, 69, 189, 214, 321, 235, 199, 
    68, 229, 171, 100, 121, 202, 115, 61, 171, 172, 228, 228, 297, 249, 131, 
    73, 226, 264, 105, 178, 234, 201, 237, 228, 241, 235, 207, 281, 247, 104, 
    76, 181, 252, 266, 273, 282, 252, 277, 273, 281, 274, 298, 275, 238, 130, 
    120, 180, 210, 278, 304, 223, 307, 332, 319, 303, 298, 347, 303, 249, 92, 
    163, 205, 214, 235, 325, 270, 322, 345, 349, 367, 348, 327, 343, 231, 75, 
    207, 202, 124, 185, 203, 330, 325, 358, 386, 379, 330, 332, 244, 127, 167, 
    168, 171, 128, 179, 187, 164, 366, 410, 375, 369, 335, 331, 268, 180, 217, 
    209, 310, 212, 174, 194, 241, 353, 420, 383, 331, 357, 344, 281, 222, 208, 
    268, 393, 364, 264, 192, 239, 339, 335, 328, 357, 390, 324, 257, 163, 184, 
    135, 148, 349, 364, 296, 216, 240, 190, 220, 371, 354, 322, 173, 111, 179, 
    125, 27, 164, 360, 392, 317, 261, 254, 231, 307, 318, 251, 120, 144, 287, 
    
    -- channel=295
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    
    -- channel=296
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 11, 10, 0, 3, 0, 0, 
    0, 0, 0, 7, 0, 0, 11, 22, 6, 0, 0, 11, 9, 0, 0, 
    0, 0, 0, 0, 5, 18, 26, 17, 2, 12, 25, 30, 0, 0, 0, 
    0, 0, 0, 0, 26, 14, 14, 29, 37, 42, 33, 17, 39, 0, 0, 
    0, 2, 0, 0, 1, 42, 25, 27, 37, 21, 20, 35, 2, 0, 0, 
    2, 0, 0, 0, 0, 0, 38, 38, 31, 37, 24, 22, 8, 0, 0, 
    0, 0, 0, 0, 2, 0, 8, 36, 31, 18, 22, 17, 15, 0, 6, 
    6, 55, 24, 2, 0, 0, 20, 24, 27, 20, 34, 28, 17, 10, 0, 
    0, 0, 25, 24, 6, 0, 10, 10, 0, 26, 24, 26, 16, 0, 0, 
    0, 0, 0, 16, 25, 10, 0, 9, 18, 20, 24, 21, 0, 0, 0, 
    0, 0, 0, 0, 23, 34, 14, 0, 0, 7, 0, 0, 12, 0, 13, 
    
    -- channel=297
    164, 45, 144, 114, 0, 59, 127, 107, 182, 170, 152, 205, 189, 67, 128, 
    198, 152, 147, 144, 0, 20, 46, 117, 198, 183, 149, 245, 275, 223, 224, 
    139, 127, 143, 93, 0, 90, 193, 151, 142, 52, 176, 283, 397, 267, 291, 
    65, 228, 178, 100, 26, 264, 203, 0, 151, 117, 267, 341, 394, 331, 219, 
    106, 328, 291, 85, 228, 285, 110, 158, 267, 304, 321, 258, 376, 336, 109, 
    68, 277, 362, 228, 278, 258, 236, 372, 326, 282, 244, 346, 360, 320, 116, 
    143, 243, 298, 364, 290, 302, 306, 291, 262, 306, 327, 353, 316, 341, 161, 
    151, 243, 304, 350, 425, 186, 330, 373, 385, 372, 327, 404, 384, 320, 43, 
    248, 302, 235, 264, 316, 419, 345, 383, 400, 379, 366, 379, 300, 227, 150, 
    292, 203, 153, 237, 264, 260, 409, 449, 416, 440, 360, 363, 264, 169, 223, 
    167, 243, 185, 239, 246, 274, 404, 471, 448, 362, 356, 347, 290, 236, 354, 
    331, 526, 352, 265, 260, 273, 422, 449, 416, 364, 417, 367, 290, 302, 281, 
    258, 396, 508, 411, 290, 331, 371, 287, 293, 411, 409, 339, 273, 150, 262, 
    155, 56, 347, 499, 437, 335, 307, 283, 292, 392, 411, 317, 114, 185, 248, 
    147, 89, 107, 403, 526, 492, 404, 344, 242, 298, 288, 251, 200, 202, 420, 
    
    -- channel=298
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=299
    0, 0, 0, 0, 0, 0, 0, 0, 9, 46, 0, 0, 0, 37, 0, 
    0, 0, 0, 0, 0, 39, 40, 0, 0, 0, 0, 0, 0, 0, 0, 
    112, 77, 0, 18, 0, 0, 0, 0, 19, 63, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 76, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 19, 
    13, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 0, 0, 0, 0, 32, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 12, 0, 0, 61, 
    0, 0, 56, 30, 112, 0, 0, 0, 0, 16, 5, 0, 134, 117, 0, 
    0, 80, 30, 28, 9, 197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 59, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 39, 23, 0, 0, 8, 19, 2, 0, 
    196, 219, 0, 0, 0, 0, 38, 221, 201, 0, 22, 0, 11, 81, 0, 
    0, 280, 227, 0, 0, 0, 0, 0, 0, 57, 0, 56, 142, 0, 0, 
    0, 0, 157, 156, 0, 0, 0, 0, 60, 142, 223, 49, 0, 0, 0, 
    
    -- channel=300
    0, 27, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 67, 0, 0, 
    0, 19, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 60, 0, 0, 
    0, 0, 0, 0, 56, 0, 0, 0, 0, 18, 0, 0, 9, 0, 0, 
    0, 0, 9, 15, 15, 0, 0, 19, 0, 38, 0, 0, 0, 0, 17, 
    16, 0, 26, 26, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 73, 
    55, 0, 0, 74, 0, 16, 70, 0, 0, 0, 0, 0, 0, 0, 101, 
    50, 0, 0, 0, 57, 55, 72, 46, 49, 46, 64, 38, 0, 0, 84, 
    8, 0, 0, 0, 45, 122, 23, 64, 81, 86, 85, 22, 89, 0, 84, 
    0, 0, 0, 0, 0, 101, 55, 71, 74, 62, 73, 61, 71, 5, 42, 
    0, 0, 0, 0, 0, 0, 73, 60, 75, 78, 76, 70, 78, 1, 0, 
    27, 0, 13, 0, 0, 19, 0, 67, 75, 75, 69, 69, 60, 0, 0, 
    0, 0, 33, 0, 0, 0, 2, 50, 65, 98, 54, 81, 65, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 75, 0, 72, 58, 107, 80, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 19, 6, 40, 58, 103, 95, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 29, 13, 25, 41, 59, 0, 0, 
    
    -- channel=301
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=302
    0, 0, 38, 11, 0, 98, 0, 38, 11, 20, 0, 127, 0, 67, 2, 
    0, 0, 0, 12, 0, 66, 1, 58, 0, 27, 0, 164, 0, 81, 0, 
    0, 0, 0, 0, 0, 79, 41, 0, 39, 0, 44, 155, 0, 10, 0, 
    0, 114, 0, 0, 2, 86, 0, 0, 101, 0, 96, 97, 0, 5, 0, 
    0, 156, 0, 0, 88, 13, 0, 84, 21, 48, 0, 55, 0, 0, 0, 
    0, 153, 7, 0, 74, 16, 0, 71, 0, 6, 0, 109, 0, 21, 0, 
    0, 98, 65, 0, 0, 8, 0, 12, 0, 10, 9, 25, 0, 39, 0, 
    0, 70, 35, 0, 1, 0, 40, 0, 0, 4, 0, 48, 0, 15, 0, 
    20, 33, 0, 3, 44, 0, 37, 0, 4, 1, 0, 14, 0, 0, 0, 
    3, 0, 0, 40, 7, 57, 0, 20, 0, 0, 0, 0, 0, 0, 57, 
    0, 63, 0, 61, 17, 0, 114, 0, 0, 0, 0, 0, 0, 12, 36, 
    25, 59, 0, 47, 0, 49, 55, 4, 0, 0, 20, 0, 0, 42, 0, 
    26, 85, 0, 0, 0, 57, 15, 0, 52, 0, 6, 0, 0, 34, 0, 
    0, 58, 123, 8, 0, 0, 2, 0, 69, 19, 1, 0, 0, 66, 45, 
    0, 0, 131, 126, 3, 0, 0, 0, 0, 10, 0, 0, 0, 30, 161, 
    
    -- channel=303
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=304
    62, 27, 57, 66, 0, 78, 40, 71, 58, 76, 32, 138, 0, 69, 62, 
    86, 51, 51, 71, 0, 40, 45, 79, 63, 72, 34, 155, 27, 97, 60, 
    42, 63, 67, 49, 0, 81, 76, 35, 91, 1, 99, 158, 79, 95, 90, 
    29, 129, 46, 35, 49, 94, 34, 3, 95, 52, 106, 126, 111, 110, 22, 
    32, 169, 64, 27, 104, 89, 0, 97, 84, 103, 81, 116, 100, 118, 0, 
    5, 156, 142, 52, 97, 94, 55, 112, 78, 79, 62, 129, 75, 132, 0, 
    33, 120, 139, 118, 64, 76, 75, 75, 76, 85, 99, 93, 75, 124, 14, 
    53, 120, 120, 125, 120, 36, 111, 99, 95, 97, 84, 141, 68, 100, 0, 
    105, 107, 90, 113, 134, 98, 104, 110, 100, 111, 99, 96, 88, 60, 29, 
    95, 76, 45, 101, 94, 136, 122, 129, 125, 105, 104, 86, 41, 60, 129, 
    33, 110, 42, 122, 94, 86, 180, 131, 118, 98, 103, 92, 60, 102, 107, 
    154, 138, 49, 98, 83, 131, 137, 128, 124, 94, 121, 84, 55, 86, 113, 
    95, 183, 123, 72, 67, 126, 124, 44, 138, 123, 117, 78, 32, 75, 83, 
    28, 45, 174, 150, 74, 76, 97, 89, 121, 116, 119, 61, 0, 85, 137, 
    18, 20, 85, 171, 153, 105, 82, 94, 58, 98, 78, 86, 53, 92, 157, 
    
    -- channel=305
    141, 128, 149, 112, 85, 127, 131, 118, 122, 112, 119, 133, 152, 94, 129, 
    133, 147, 125, 110, 86, 89, 88, 121, 151, 133, 130, 137, 204, 177, 143, 
    59, 100, 108, 76, 86, 163, 192, 121, 105, 63, 149, 145, 188, 147, 154, 
    114, 178, 118, 112, 129, 202, 142, 75, 117, 155, 191, 169, 160, 147, 88, 
    112, 145, 170, 93, 172, 174, 127, 181, 196, 200, 177, 137, 160, 122, 82, 
    84, 107, 146, 190, 184, 142, 163, 200, 181, 157, 155, 189, 153, 121, 125, 
    144, 127, 107, 149, 150, 159, 197, 148, 132, 143, 167, 160, 154, 141, 137, 
    108, 125, 121, 124, 215, 101, 151, 173, 202, 203, 145, 155, 166, 133, 62, 
    156, 144, 87, 104, 76, 202, 143, 160, 158, 139, 162, 136, 93, 88, 148, 
    113, 81, 87, 106, 123, 67, 158, 165, 148, 155, 144, 146, 140, 118, 143, 
    82, 154, 142, 146, 117, 142, 144, 150, 149, 114, 136, 155, 156, 145, 156, 
    210, 283, 244, 152, 136, 114, 147, 149, 128, 140, 167, 151, 160, 144, 137, 
    47, 110, 247, 236, 176, 151, 121, 73, 79, 161, 141, 148, 147, 98, 121, 
    117, 12, 113, 238, 247, 204, 170, 198, 138, 128, 156, 122, 84, 121, 175, 
    128, 163, 70, 138, 233, 254, 233, 187, 121, 99, 75, 129, 184, 184, 202, 
    
    -- channel=306
    0, 24, 0, 0, 106, 0, 0, 0, 0, 0, 49, 0, 161, 0, 0, 
    0, 0, 4, 0, 124, 0, 3, 0, 0, 0, 50, 0, 116, 0, 0, 
    30, 1, 0, 24, 108, 0, 0, 0, 0, 95, 0, 0, 38, 0, 0, 
    57, 0, 10, 24, 0, 0, 14, 126, 0, 42, 0, 0, 23, 0, 115, 
    46, 0, 49, 46, 0, 0, 137, 0, 0, 0, 0, 0, 1, 0, 220, 
    122, 0, 0, 53, 0, 0, 42, 0, 0, 0, 42, 0, 39, 0, 218, 
    52, 0, 0, 0, 38, 0, 0, 0, 13, 0, 0, 0, 52, 0, 170, 
    41, 0, 0, 0, 0, 80, 0, 0, 0, 0, 0, 0, 25, 0, 212, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 21, 0, 87, 66, 74, 
    0, 51, 45, 0, 0, 0, 0, 0, 0, 1, 0, 17, 82, 0, 0, 
    122, 0, 42, 0, 0, 0, 0, 0, 0, 42, 0, 13, 38, 0, 0, 
    0, 0, 33, 0, 25, 0, 0, 0, 11, 46, 0, 11, 56, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 107, 0, 0, 0, 49, 57, 0, 0, 
    49, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 72, 185, 0, 0, 
    90, 0, 0, 0, 0, 0, 0, 0, 38, 0, 37, 46, 8, 0, 0, 
    
    -- channel=307
    136, 152, 154, 155, 140, 173, 159, 169, 179, 193, 168, 172, 162, 172, 163, 
    136, 160, 160, 144, 147, 164, 165, 172, 168, 166, 170, 162, 163, 142, 143, 
    152, 181, 154, 137, 152, 179, 176, 165, 168, 150, 189, 155, 143, 156, 150, 
    157, 159, 136, 141, 167, 195, 217, 196, 172, 152, 165, 196, 153, 140, 114, 
    149, 149, 128, 142, 182, 176, 170, 183, 184, 192, 201, 223, 168, 128, 122, 
    147, 150, 147, 142, 169, 157, 137, 135, 172, 176, 178, 187, 181, 138, 130, 
    144, 140, 148, 137, 148, 147, 148, 130, 140, 128, 119, 135, 166, 154, 145, 
    159, 152, 141, 135, 109, 124, 137, 131, 126, 120, 116, 100, 111, 149, 147, 
    146, 143, 143, 154, 127, 102, 100, 107, 108, 118, 132, 112, 116, 151, 159, 
    131, 158, 161, 161, 144, 119, 107, 83, 100, 91, 115, 118, 117, 133, 171, 
    138, 168, 166, 151, 160, 138, 113, 88, 78, 103, 109, 120, 136, 141, 137, 
    143, 128, 194, 174, 147, 145, 110, 108, 92, 95, 99, 114, 165, 165, 185, 
    157, 194, 203, 221, 196, 146, 126, 124, 132, 97, 88, 113, 131, 197, 196, 
    151, 200, 236, 210, 224, 226, 206, 170, 127, 102, 106, 119, 146, 192, 205, 
    166, 190, 207, 238, 202, 209, 227, 217, 170, 133, 122, 155, 159, 161, 188, 
    
    -- channel=308
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=309
    0, 41, 0, 0, 100, 0, 0, 0, 0, 0, 36, 0, 175, 0, 0, 
    0, 0, 0, 0, 130, 0, 0, 0, 0, 0, 41, 0, 192, 0, 0, 
    0, 0, 0, 0, 126, 0, 0, 0, 0, 37, 0, 0, 56, 0, 0, 
    57, 0, 0, 37, 12, 0, 0, 123, 0, 111, 0, 0, 8, 0, 78, 
    30, 0, 95, 5, 0, 0, 146, 0, 0, 0, 0, 0, 0, 0, 228, 
    110, 0, 0, 137, 0, 0, 69, 0, 0, 0, 23, 0, 3, 0, 255, 
    87, 0, 0, 0, 30, 4, 48, 0, 17, 0, 14, 0, 34, 0, 218, 
    38, 0, 0, 0, 20, 63, 0, 0, 48, 10, 0, 0, 66, 0, 209, 
    0, 0, 0, 0, 0, 117, 0, 28, 0, 9, 54, 0, 78, 15, 136, 
    0, 5, 14, 0, 0, 0, 18, 0, 10, 28, 30, 34, 127, 0, 0, 
    98, 0, 32, 0, 0, 9, 0, 0, 33, 43, 27, 47, 61, 0, 0, 
    0, 0, 67, 0, 3, 0, 0, 0, 20, 83, 0, 31, 74, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 64, 0, 40, 0, 96, 80, 0, 0, 
    38, 0, 0, 0, 16, 0, 0, 56, 0, 0, 18, 78, 197, 0, 0, 
    74, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 100, 78, 0, 0, 
    
    -- channel=310
    64, 20, 58, 99, 94, 0, 49, 9, 21, 1, 68, 0, 77, 0, 23, 
    63, 29, 75, 104, 65, 0, 18, 0, 62, 38, 66, 0, 91, 38, 94, 
    45, 8, 67, 71, 35, 0, 47, 66, 45, 38, 30, 0, 108, 77, 107, 
    72, 41, 65, 48, 0, 33, 47, 0, 0, 47, 17, 0, 98, 88, 141, 
    78, 69, 155, 19, 0, 40, 37, 0, 53, 21, 37, 0, 53, 114, 148, 
    44, 44, 133, 121, 29, 0, 0, 43, 29, 0, 0, 0, 52, 114, 129, 
    66, 50, 58, 104, 0, 0, 0, 0, 0, 0, 0, 0, 6, 88, 119, 
    56, 54, 74, 85, 0, 0, 0, 0, 0, 0, 0, 0, 8, 56, 62, 
    64, 75, 65, 65, 0, 25, 0, 0, 0, 0, 0, 0, 0, 5, 84, 
    97, 46, 54, 51, 43, 0, 0, 0, 0, 0, 0, 0, 0, 37, 40, 
    85, 17, 59, 70, 50, 53, 0, 0, 0, 0, 0, 0, 0, 34, 133, 
    57, 65, 43, 40, 102, 24, 0, 0, 0, 0, 0, 0, 0, 0, 113, 
    9, 0, 26, 19, 38, 53, 0, 0, 0, 0, 0, 0, 0, 0, 103, 
    62, 0, 0, 9, 24, 9, 0, 32, 0, 0, 0, 0, 0, 15, 49, 
    73, 13, 0, 0, 20, 46, 39, 3, 0, 0, 0, 0, 21, 39, 0, 
    
    -- channel=311
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=312
    0, 7, 0, 0, 7, 0, 1, 7, 4, 5, 3, 10, 0, 0, 3, 
    0, 24, 0, 0, 20, 0, 0, 14, 0, 9, 0, 8, 0, 0, 0, 
    25, 12, 2, 6, 24, 0, 0, 13, 0, 22, 0, 7, 0, 5, 0, 
    0, 0, 7, 9, 13, 0, 18, 9, 3, 4, 0, 25, 0, 0, 0, 
    18, 0, 0, 11, 9, 0, 1, 6, 0, 10, 1, 15, 0, 0, 0, 
    28, 0, 0, 20, 0, 9, 0, 0, 13, 2, 0, 30, 0, 0, 0, 
    17, 0, 0, 13, 11, 4, 0, 0, 0, 0, 0, 9, 0, 7, 0, 
    18, 0, 19, 5, 0, 24, 0, 0, 0, 0, 9, 0, 10, 0, 24, 
    0, 7, 8, 0, 10, 13, 0, 0, 1, 0, 0, 10, 0, 1, 21, 
    15, 11, 24, 6, 0, 0, 11, 0, 0, 0, 2, 0, 0, 0, 0, 
    12, 0, 10, 0, 22, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 7, 0, 2, 0, 0, 0, 3, 0, 0, 1, 0, 1, 
    26, 0, 0, 14, 17, 0, 6, 6, 0, 0, 0, 0, 0, 1, 18, 
    1, 30, 0, 0, 8, 14, 6, 0, 21, 0, 0, 7, 0, 14, 0, 
    1, 5, 6, 0, 0, 10, 10, 1, 21, 0, 0, 0, 0, 0, 0, 
    
    -- channel=313
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=314
    78, 96, 92, 92, 79, 126, 84, 101, 64, 79, 55, 105, 15, 110, 86, 
    74, 71, 77, 84, 81, 118, 101, 97, 71, 77, 61, 102, 22, 90, 58, 
    51, 87, 81, 79, 95, 121, 85, 63, 101, 58, 90, 94, 5, 55, 39, 
    77, 101, 49, 81, 112, 74, 40, 98, 88, 88, 73, 55, 16, 44, 15, 
    71, 87, 34, 60, 103, 56, 50, 105, 66, 58, 34, 70, 23, 37, 20, 
    67, 87, 45, 48, 56, 51, 57, 71, 39, 49, 44, 66, 16, 50, 23, 
    66, 81, 60, 23, 33, 48, 51, 38, 39, 47, 54, 37, 34, 44, 35, 
    62, 78, 48, 27, 42, 35, 49, 27, 42, 33, 22, 48, 5, 45, 42, 
    72, 51, 50, 51, 31, 34, 39, 34, 19, 18, 20, 28, 13, 56, 66, 
    41, 55, 54, 61, 63, 43, 39, 22, 13, 11, 26, 19, 36, 64, 83, 
    38, 77, 57, 84, 45, 57, 45, 7, 11, 6, 30, 25, 33, 75, 42, 
    64, 26, 15, 57, 49, 53, 32, 8, 18, 14, 27, 17, 27, 66, 46, 
    31, 45, 6, 8, 34, 57, 27, 10, 62, 27, 17, 20, 26, 87, 38, 
    48, 73, 62, 20, 0, 30, 29, 53, 51, 25, 25, 10, 46, 79, 92, 
    45, 97, 85, 54, 14, 4, 11, 25, 28, 42, 38, 58, 56, 79, 42, 
    
    -- channel=315
    50, 0, 19, 7, 0, 0, 10, 28, 65, 74, 26, 145, 9, 12, 40, 
    99, 47, 25, 35, 0, 0, 0, 47, 61, 73, 17, 186, 83, 106, 82, 
    58, 42, 47, 16, 0, 5, 57, 25, 54, 0, 68, 216, 208, 137, 143, 
    0, 114, 68, 11, 0, 101, 41, 0, 85, 19, 133, 218, 233, 195, 73, 
    0, 214, 114, 13, 116, 140, 0, 66, 102, 155, 153, 165, 224, 211, 0, 
    0, 191, 221, 72, 137, 181, 142, 211, 168, 159, 127, 221, 196, 202, 0, 
    24, 145, 208, 227, 188, 220, 206, 214, 201, 230, 241, 257, 180, 206, 20, 
    54, 144, 200, 231, 286, 151, 261, 285, 272, 276, 263, 321, 254, 188, 0, 
    135, 176, 144, 166, 282, 275, 280, 300, 311, 316, 285, 297, 246, 135, 14, 
    173, 116, 57, 136, 146, 251, 318, 349, 345, 332, 289, 272, 150, 74, 136, 
    60, 139, 57, 128, 152, 153, 349, 375, 346, 298, 288, 267, 190, 142, 183, 
    222, 312, 145, 148, 123, 204, 328, 366, 342, 279, 325, 281, 189, 174, 143, 
    190, 322, 302, 202, 136, 208, 289, 219, 276, 324, 332, 261, 161, 90, 115, 
    32, 41, 267, 317, 216, 157, 179, 148, 228, 319, 323, 243, 31, 84, 130, 
    11, 0, 77, 295, 340, 269, 191, 187, 153, 238, 226, 175, 81, 81, 280, 
    
    -- channel=316
    240, 101, 216, 228, 81, 152, 224, 220, 333, 341, 282, 341, 291, 197, 209, 
    295, 221, 260, 257, 54, 130, 171, 215, 315, 300, 279, 377, 357, 275, 326, 
    290, 291, 257, 204, 41, 159, 271, 271, 301, 175, 324, 409, 509, 392, 414, 
    177, 319, 259, 189, 83, 391, 387, 118, 259, 202, 374, 497, 564, 459, 352, 
    204, 482, 388, 171, 328, 433, 222, 215, 394, 420, 489, 477, 531, 472, 225, 
    165, 449, 523, 281, 393, 385, 282, 469, 457, 435, 385, 474, 517, 490, 199, 
    205, 365, 467, 518, 401, 389, 354, 368, 359, 387, 387, 434, 449, 492, 253, 
    273, 378, 432, 511, 489, 230, 423, 438, 438, 395, 370, 489, 440, 462, 168, 
    345, 416, 392, 439, 465, 457, 400, 450, 461, 470, 446, 452, 416, 368, 245, 
    414, 371, 291, 398, 416, 408, 476, 502, 487, 508, 435, 442, 328, 249, 336, 
    314, 374, 291, 369, 363, 384, 512, 554, 518, 451, 442, 424, 359, 321, 482, 
    407, 575, 441, 394, 412, 403, 537, 552, 499, 432, 480, 436, 394, 414, 479, 
    471, 664, 689, 552, 432, 477, 513, 414, 449, 482, 487, 401, 343, 291, 466, 
    284, 266, 645, 697, 586, 497, 483, 376, 364, 490, 497, 393, 214, 321, 433, 
    276, 177, 298, 682, 726, 642, 574, 525, 383, 426, 432, 366, 235, 291, 568, 
    
    -- channel=317
    160, 87, 117, 136, 116, 31, 156, 119, 230, 224, 236, 144, 314, 102, 137, 
    190, 162, 192, 155, 105, 54, 121, 108, 220, 185, 228, 149, 334, 132, 225, 
    220, 187, 173, 146, 80, 47, 158, 205, 170, 183, 180, 187, 392, 254, 282, 
    161, 135, 206, 138, 53, 213, 304, 145, 118, 153, 208, 289, 414, 299, 315, 
    169, 216, 301, 164, 143, 288, 241, 85, 257, 257, 341, 310, 384, 313, 276, 
    170, 205, 329, 229, 232, 262, 218, 248, 308, 306, 297, 254, 397, 308, 268, 
    176, 187, 279, 352, 301, 268, 249, 262, 268, 262, 250, 282, 344, 305, 272, 
    209, 212, 260, 341, 308, 228, 268, 309, 295, 272, 270, 304, 325, 305, 231, 
    211, 253, 277, 292, 307, 291, 265, 308, 316, 335, 335, 301, 333, 266, 204, 
    272, 267, 232, 235, 272, 286, 290, 317, 341, 353, 307, 326, 276, 181, 184, 
    274, 209, 233, 207, 237, 243, 289, 372, 357, 342, 302, 312, 281, 205, 294, 
    234, 338, 357, 259, 300, 245, 321, 378, 346, 321, 305, 323, 312, 263, 326, 
    317, 410, 485, 416, 329, 296, 338, 350, 273, 321, 342, 308, 291, 195, 327, 
    238, 190, 372, 472, 445, 363, 352, 288, 212, 326, 330, 323, 247, 168, 244, 
    253, 121, 165, 399, 497, 455, 429, 378, 317, 290, 307, 270, 197, 184, 308, 
    
    -- channel=318
    13, 0, 0, 0, 0, 0, 0, 0, 10, 0, 35, 0, 110, 0, 0, 
    39, 2, 6, 0, 0, 0, 0, 0, 24, 0, 33, 0, 139, 0, 46, 
    26, 0, 0, 0, 0, 0, 0, 3, 0, 9, 0, 0, 176, 52, 87, 
    0, 0, 47, 2, 0, 0, 28, 0, 0, 16, 12, 24, 166, 102, 129, 
    12, 15, 125, 14, 0, 62, 56, 0, 37, 25, 71, 28, 130, 111, 117, 
    17, 0, 113, 88, 16, 81, 69, 75, 88, 84, 78, 19, 129, 99, 113, 
    30, 9, 63, 145, 124, 94, 91, 99, 95, 100, 108, 111, 111, 79, 108, 
    31, 17, 67, 127, 159, 78, 97, 136, 142, 131, 121, 138, 177, 80, 65, 
    40, 66, 71, 77, 113, 166, 123, 155, 158, 158, 153, 137, 159, 67, 37, 
    80, 62, 32, 27, 66, 96, 150, 177, 184, 194, 148, 154, 120, 22, 1, 
    91, 11, 41, 25, 42, 71, 115, 212, 203, 181, 145, 147, 113, 41, 84, 
    84, 158, 119, 27, 91, 63, 150, 199, 183, 179, 162, 158, 108, 40, 70, 
    74, 106, 191, 126, 77, 71, 150, 147, 88, 175, 184, 158, 117, 0, 55, 
    52, 0, 40, 164, 149, 73, 72, 76, 57, 161, 164, 154, 66, 0, 23, 
    52, 0, 0, 58, 185, 166, 118, 92, 85, 100, 114, 80, 44, 17, 48, 
    
    -- channel=319
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=320
    129, 156, 160, 163, 162, 160, 146, 141, 93, 88, 87, 75, 80, 100, 69, 
    177, 179, 169, 171, 180, 175, 161, 161, 115, 67, 95, 97, 108, 93, 91, 
    149, 188, 179, 190, 189, 189, 171, 180, 173, 92, 119, 89, 102, 108, 101, 
    142, 184, 184, 197, 193, 198, 178, 168, 180, 172, 145, 100, 94, 102, 106, 
    153, 175, 187, 191, 201, 189, 153, 150, 126, 174, 163, 97, 111, 108, 108, 
    179, 154, 187, 191, 189, 210, 125, 147, 130, 148, 117, 63, 103, 100, 109, 
    150, 202, 180, 169, 175, 190, 158, 100, 128, 130, 80, 43, 76, 99, 97, 
    89, 198, 166, 174, 199, 178, 171, 182, 163, 155, 78, 48, 89, 123, 61, 
    113, 180, 162, 130, 195, 184, 138, 174, 166, 145, 76, 43, 97, 159, 30, 
    104, 187, 159, 46, 203, 177, 110, 169, 82, 60, 45, 44, 100, 192, 28, 
    115, 168, 149, 41, 55, 93, 95, 139, 84, 48, 56, 77, 83, 197, 82, 
    125, 130, 151, 102, 84, 75, 90, 62, 26, 33, 25, 50, 96, 123, 152, 
    134, 136, 125, 182, 122, 114, 114, 75, 42, 30, 15, 38, 78, 69, 117, 
    112, 148, 121, 124, 111, 115, 139, 102, 97, 79, 81, 97, 83, 99, 96, 
    122, 129, 118, 129, 116, 129, 135, 129, 119, 105, 126, 138, 119, 107, 112, 
    
    -- channel=321
    94, 53, 124, 135, 131, 127, 133, 100, 110, 85, 105, 90, 86, 100, 115, 
    108, 118, 112, 121, 130, 130, 136, 135, 119, 70, 98, 123, 128, 125, 109, 
    113, 105, 110, 126, 125, 130, 138, 127, 132, 85, 85, 115, 139, 135, 118, 
    100, 98, 121, 121, 134, 147, 162, 137, 140, 147, 113, 120, 123, 114, 126, 
    101, 109, 119, 111, 132, 131, 131, 120, 127, 153, 134, 134, 106, 121, 125, 
    65, 98, 108, 120, 116, 69, 100, 146, 141, 114, 136, 118, 92, 105, 117, 
    45, 118, 126, 121, 76, 98, 124, 89, 58, 72, 119, 94, 66, 91, 116, 
    119, 92, 137, 110, 82, 121, 117, 122, 112, 108, 127, 99, 59, 80, 101, 
    166, 95, 127, 110, 128, 107, 177, 162, 163, 166, 173, 90, 41, 86, 123, 
    168, 98, 124, 157, 119, 121, 186, 140, 142, 100, 78, 90, 65, 72, 129, 
    181, 127, 137, 156, 31, 104, 152, 169, 183, 87, 86, 104, 75, 87, 151, 
    180, 153, 115, 101, 98, 98, 102, 120, 59, 50, 50, 44, 80, 103, 140, 
    164, 171, 122, 131, 125, 146, 153, 133, 77, 41, 33, 20, 52, 76, 102, 
    178, 162, 181, 115, 150, 125, 153, 178, 123, 114, 98, 86, 83, 89, 125, 
    166, 152, 178, 152, 132, 162, 166, 178, 154, 157, 148, 147, 146, 142, 114, 
    
    -- channel=322
    205, 225, 223, 244, 231, 223, 207, 202, 148, 127, 163, 158, 157, 187, 160, 
    227, 213, 229, 242, 249, 247, 239, 244, 194, 110, 147, 169, 210, 197, 173, 
    204, 212, 237, 245, 254, 248, 247, 231, 246, 211, 222, 204, 206, 194, 203, 
    190, 219, 233, 252, 251, 265, 257, 234, 237, 255, 237, 180, 176, 195, 202, 
    186, 230, 246, 247, 252, 257, 245, 272, 216, 243, 240, 151, 161, 179, 195, 
    167, 248, 256, 253, 219, 255, 242, 178, 177, 231, 211, 106, 133, 156, 185, 
    195, 242, 260, 246, 243, 253, 207, 249, 257, 250, 181, 116, 116, 153, 168, 
    206, 256, 257, 230, 280, 272, 284, 292, 262, 261, 199, 109, 119, 211, 155, 
    257, 295, 274, 199, 233, 240, 239, 200, 199, 157, 74, 63, 119, 230, 143, 
    262, 279, 270, 149, 133, 245, 202, 303, 229, 109, 117, 135, 140, 262, 172, 
    277, 269, 229, 115, 122, 61, 118, 203, 110, 87, 61, 110, 160, 235, 182, 
    259, 290, 222, 234, 200, 219, 232, 166, 47, 30, 33, 37, 117, 163, 199, 
    281, 290, 244, 209, 208, 229, 264, 226, 159, 117, 83, 80, 110, 125, 167, 
    256, 263, 250, 227, 177, 232, 273, 261, 223, 213, 202, 224, 204, 204, 178, 
    268, 303, 278, 286, 268, 285, 258, 244, 239, 234, 255, 265, 257, 226, 224, 
    
    -- channel=323
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 6, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 6, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 15, 0, 16, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 18, 40, 17, 0, 65, 0, 0, 18, 17, 0, 0, 0, 0, 0, 
    0, 44, 34, 3, 70, 56, 32, 67, 57, 47, 0, 0, 0, 0, 0, 
    0, 51, 47, 0, 76, 32, 21, 0, 8, 0, 0, 0, 0, 9, 0, 
    0, 48, 67, 0, 0, 39, 0, 42, 0, 0, 0, 0, 0, 39, 0, 
    0, 22, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 32, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=324
    75, 104, 70, 72, 71, 70, 57, 58, 53, 33, 31, 38, 31, 42, 35, 
    109, 106, 80, 81, 80, 78, 70, 62, 51, 35, 29, 28, 36, 43, 31, 
    111, 99, 95, 90, 91, 91, 80, 68, 69, 68, 52, 41, 32, 30, 43, 
    91, 102, 96, 94, 101, 87, 76, 73, 72, 70, 65, 60, 28, 33, 39, 
    85, 96, 101, 99, 100, 90, 80, 83, 80, 58, 73, 73, 39, 39, 41, 
    40, 97, 104, 108, 100, 106, 130, 86, 71, 61, 70, 35, 34, 38, 39, 
    72, 87, 118, 111, 100, 142, 100, 84, 94, 105, 74, 32, 33, 41, 35, 
    47, 72, 112, 96, 129, 127, 116, 111, 121, 117, 98, 42, 28, 56, 49, 
    43, 74, 111, 106, 127, 96, 112, 83, 83, 79, 38, 10, 30, 68, 70, 
    42, 74, 118, 105, 34, 108, 68, 62, 70, 19, 17, 23, 24, 73, 95, 
    58, 64, 107, 46, 43, 31, 22, 33, 17, 22, 18, 7, 33, 66, 94, 
    38, 64, 75, 87, 47, 29, 37, 28, 18, 9, 6, 17, 16, 52, 56, 
    54, 46, 81, 70, 92, 57, 31, 40, 29, 23, 21, 18, 35, 20, 53, 
    51, 42, 59, 65, 57, 47, 49, 44, 37, 43, 34, 46, 45, 51, 31, 
    34, 61, 45, 51, 58, 58, 51, 39, 47, 30, 42, 48, 52, 49, 42, 
    
    -- channel=325
    58, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 18, 
    0, 6, 0, 0, 0, 0, 0, 0, 25, 6, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 6, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 17, 0, 0, 64, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 52, 0, 18, 0, 11, 52, 0, 0, 0, 
    0, 0, 11, 13, 0, 0, 27, 56, 0, 0, 60, 39, 0, 0, 0, 
    5, 0, 21, 0, 0, 36, 14, 0, 12, 23, 87, 38, 0, 0, 37, 
    7, 0, 20, 36, 0, 0, 50, 0, 0, 0, 56, 4, 0, 0, 106, 
    18, 0, 16, 129, 0, 0, 68, 0, 52, 12, 3, 0, 0, 0, 148, 
    19, 0, 9, 130, 0, 0, 0, 0, 46, 4, 0, 0, 0, 0, 110, 
    8, 0, 0, 49, 32, 0, 0, 18, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 48, 1, 0, 36, 28, 6, 4, 0, 0, 0, 0, 
    0, 0, 23, 0, 28, 0, 0, 24, 0, 9, 0, 0, 4, 0, 2, 
    0, 0, 8, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 11, 0, 
    
    -- channel=326
    118, 137, 129, 135, 129, 130, 113, 120, 81, 87, 95, 94, 96, 106, 81, 
    133, 128, 138, 139, 141, 138, 132, 133, 100, 82, 95, 94, 107, 101, 97, 
    125, 136, 143, 144, 148, 145, 137, 141, 132, 105, 118, 103, 107, 103, 107, 
    117, 141, 140, 147, 146, 144, 139, 130, 140, 135, 134, 101, 100, 111, 109, 
    122, 136, 144, 150, 147, 146, 141, 148, 126, 137, 132, 84, 102, 102, 108, 
    133, 147, 152, 150, 140, 161, 136, 106, 98, 137, 117, 70, 95, 96, 107, 
    139, 145, 146, 139, 150, 155, 113, 121, 145, 144, 97, 71, 88, 97, 100, 
    104, 158, 136, 137, 164, 146, 150, 151, 139, 137, 92, 64, 91, 121, 90, 
    113, 161, 144, 116, 139, 149, 119, 116, 108, 93, 48, 53, 100, 137, 66, 
    122, 160, 144, 63, 113, 142, 95, 143, 110, 74, 76, 73, 100, 156, 71, 
    123, 145, 124, 51, 99, 77, 81, 119, 59, 66, 60, 73, 101, 153, 75, 
    122, 137, 125, 114, 101, 98, 109, 87, 59, 51, 47, 67, 91, 113, 102, 
    133, 136, 128, 124, 110, 117, 128, 99, 76, 73, 62, 67, 90, 90, 115, 
    120, 138, 112, 125, 91, 122, 137, 111, 109, 99, 96, 110, 101, 109, 92, 
    125, 140, 124, 133, 127, 134, 123, 119, 117, 112, 124, 132, 123, 111, 118, 
    
    -- channel=327
    47, 0, 4, 0, 0, 0, 11, 0, 34, 2, 0, 0, 0, 0, 25, 
    6, 7, 3, 0, 0, 0, 12, 0, 33, 31, 0, 0, 0, 3, 1, 
    34, 0, 0, 0, 0, 1, 10, 0, 6, 37, 0, 22, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 9, 9, 0, 0, 9, 46, 0, 0, 0, 
    2, 0, 0, 0, 0, 7, 2, 0, 26, 0, 0, 65, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 35, 13, 10, 0, 15, 53, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 19, 22, 0, 0, 52, 45, 0, 0, 0, 
    8, 0, 9, 0, 0, 13, 14, 0, 0, 0, 69, 48, 0, 0, 47, 
    14, 0, 2, 46, 0, 0, 53, 0, 0, 13, 57, 15, 0, 0, 90, 
    14, 0, 0, 114, 0, 0, 54, 0, 51, 29, 11, 4, 0, 0, 98, 
    20, 0, 0, 107, 0, 0, 0, 0, 58, 23, 0, 0, 0, 0, 61, 
    13, 0, 0, 30, 39, 1, 0, 21, 30, 6, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 59, 5, 0, 37, 29, 11, 14, 0, 0, 0, 0, 
    6, 0, 24, 0, 28, 0, 0, 23, 3, 14, 1, 0, 6, 0, 3, 
    0, 0, 8, 0, 4, 0, 0, 3, 0, 3, 0, 0, 7, 12, 0, 
    
    -- channel=328
    269, 272, 244, 249, 247, 227, 201, 183, 166, 105, 116, 117, 111, 142, 134, 
    325, 321, 258, 273, 275, 270, 241, 219, 179, 91, 100, 124, 154, 158, 132, 
    325, 304, 293, 294, 304, 297, 271, 240, 251, 208, 183, 157, 141, 145, 160, 
    289, 312, 301, 308, 321, 296, 281, 249, 253, 261, 231, 189, 124, 132, 158, 
    257, 301, 318, 308, 326, 306, 288, 293, 249, 227, 256, 222, 131, 149, 158, 
    142, 307, 335, 341, 311, 349, 378, 285, 237, 227, 231, 128, 110, 127, 145, 
    174, 298, 382, 347, 321, 391, 326, 294, 306, 315, 235, 104, 91, 125, 131, 
    171, 250, 366, 324, 392, 425, 364, 378, 392, 382, 298, 120, 91, 198, 155, 
    206, 271, 378, 298, 359, 323, 352, 266, 272, 243, 140, 29, 71, 233, 201, 
    204, 262, 397, 265, 183, 322, 271, 283, 228, 78, 72, 72, 80, 262, 291, 
    245, 241, 340, 188, 51, 72, 96, 141, 122, 48, 38, 60, 97, 229, 324, 
    216, 239, 274, 287, 177, 134, 149, 112, 19, 0, 0, 4, 58, 138, 242, 
    224, 239, 246, 281, 286, 204, 181, 174, 103, 59, 31, 29, 71, 67, 152, 
    216, 205, 249, 197, 214, 187, 216, 207, 171, 165, 143, 166, 161, 158, 155, 
    202, 240, 227, 228, 235, 244, 217, 203, 190, 164, 190, 217, 218, 197, 170, 
    
    -- channel=329
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 56, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=330
    156, 168, 194, 196, 196, 204, 202, 190, 154, 156, 147, 143, 142, 152, 137, 
    182, 182, 202, 191, 204, 205, 211, 211, 187, 159, 152, 156, 154, 152, 152, 
    161, 175, 198, 207, 205, 211, 211, 224, 209, 148, 153, 159, 163, 166, 157, 
    153, 167, 196, 206, 202, 224, 213, 216, 213, 198, 192, 176, 163, 166, 160, 
    166, 174, 189, 203, 206, 216, 176, 166, 174, 211, 199, 159, 163, 162, 159, 
    194, 160, 178, 193, 202, 185, 106, 147, 155, 171, 162, 143, 151, 161, 160, 
    162, 186, 153, 161, 170, 151, 146, 111, 106, 116, 123, 127, 133, 154, 156, 
    145, 179, 148, 162, 150, 132, 167, 142, 113, 110, 106, 124, 135, 138, 134, 
    168, 163, 136, 157, 144, 166, 155, 180, 171, 171, 143, 135, 148, 148, 105, 
    165, 178, 116, 114, 168, 160, 142, 152, 141, 150, 123, 120, 151, 154, 58, 
    164, 180, 127, 106, 138, 162, 166, 188, 175, 150, 137, 138, 149, 176, 73, 
    174, 165, 146, 117, 137, 134, 142, 141, 136, 127, 116, 132, 153, 177, 137, 
    186, 168, 159, 169, 164, 162, 162, 142, 119, 109, 101, 106, 139, 149, 152, 
    168, 182, 158, 177, 153, 154, 169, 162, 153, 134, 134, 136, 134, 151, 138, 
    163, 165, 166, 167, 153, 156, 185, 179, 173, 171, 174, 174, 166, 161, 168, 
    
    -- channel=331
    146, 124, 163, 152, 161, 152, 142, 118, 124, 77, 81, 77, 60, 84, 94, 
    174, 195, 149, 168, 172, 161, 161, 147, 137, 64, 70, 92, 106, 115, 86, 
    200, 162, 168, 177, 179, 186, 174, 149, 159, 111, 94, 110, 110, 109, 103, 
    159, 182, 179, 178, 192, 194, 188, 167, 162, 168, 145, 130, 101, 83, 106, 
    159, 160, 180, 182, 186, 198, 165, 148, 156, 151, 154, 168, 84, 111, 110, 
    33, 179, 165, 193, 195, 152, 202, 191, 170, 129, 155, 111, 74, 91, 99, 
    67, 158, 219, 199, 144, 207, 196, 145, 115, 140, 155, 77, 50, 79, 97, 
    128, 114, 213, 184, 182, 219, 198, 199, 211, 206, 174, 92, 48, 96, 107, 
    138, 135, 197, 179, 209, 169, 221, 199, 196, 201, 172, 47, 16, 114, 138, 
    155, 123, 204, 213, 122, 188, 199, 148, 175, 77, 31, 56, 42, 115, 189, 
    170, 141, 207, 174, 27, 78, 98, 131, 139, 57, 51, 57, 53, 116, 217, 
    161, 149, 162, 121, 126, 63, 87, 124, 25, 7, 14, 14, 34, 96, 161, 
    139, 165, 145, 175, 152, 159, 109, 112, 62, 28, 11, 1, 43, 47, 93, 
    160, 127, 179, 126, 155, 106, 139, 155, 99, 99, 79, 83, 86, 85, 131, 
    130, 145, 151, 136, 135, 159, 157, 154, 142, 116, 127, 139, 141, 138, 91, 
    
    -- channel=332
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 15, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=333
    17, 43, 47, 50, 39, 34, 22, 37, 22, 44, 40, 21, 21, 47, 27, 
    91, 81, 49, 51, 46, 34, 19, 25, 0, 6, 54, 44, 50, 32, 32, 
    74, 95, 63, 63, 62, 50, 24, 40, 32, 0, 20, 10, 38, 45, 37, 
    86, 101, 73, 76, 73, 55, 45, 41, 63, 48, 29, 3, 28, 30, 43, 
    101, 87, 78, 72, 68, 64, 64, 48, 34, 70, 67, 28, 58, 53, 50, 
    135, 64, 75, 80, 81, 110, 91, 130, 95, 78, 56, 22, 63, 45, 52, 
    105, 143, 113, 94, 88, 131, 111, 36, 57, 82, 42, 15, 47, 39, 45, 
    24, 137, 107, 113, 144, 112, 79, 132, 141, 125, 38, 35, 72, 55, 10, 
    18, 124, 105, 87, 177, 138, 77, 140, 143, 141, 83, 28, 72, 111, 2, 
    16, 119, 141, 21, 197, 159, 63, 74, 4, 26, 8, 3, 68, 139, 10, 
    32, 111, 139, 0, 30, 90, 75, 100, 51, 34, 57, 52, 41, 161, 68, 
    47, 59, 106, 20, 0, 0, 5, 11, 4, 21, 25, 57, 71, 94, 119, 
    42, 55, 63, 131, 48, 59, 33, 0, 0, 0, 0, 7, 44, 33, 83, 
    40, 84, 51, 67, 52, 33, 60, 13, 18, 11, 4, 13, 2, 23, 43, 
    30, 41, 31, 37, 35, 39, 44, 54, 38, 25, 35, 44, 29, 21, 31, 
    
    -- channel=334
    43, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 18, 
    0, 9, 0, 0, 0, 0, 2, 0, 33, 12, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 3, 0, 1, 34, 0, 3, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 7, 0, 0, 70, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 22, 0, 27, 0, 5, 54, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 15, 30, 0, 0, 44, 35, 0, 0, 0, 
    1, 0, 5, 0, 0, 0, 0, 0, 0, 0, 65, 40, 0, 0, 26, 
    0, 0, 0, 30, 0, 0, 35, 0, 0, 6, 68, 18, 0, 0, 95, 
    10, 0, 0, 126, 0, 0, 52, 0, 39, 23, 0, 0, 0, 0, 116, 
    8, 0, 0, 115, 0, 0, 0, 0, 60, 21, 0, 0, 0, 0, 86, 
    0, 0, 0, 21, 14, 0, 0, 25, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 44, 5, 0, 23, 20, 2, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 20, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    
    -- channel=335
    174, 225, 169, 193, 181, 160, 142, 143, 98, 74, 100, 93, 101, 126, 88, 
    249, 229, 187, 205, 210, 199, 157, 168, 116, 39, 98, 96, 137, 114, 104, 
    207, 262, 215, 222, 231, 210, 190, 167, 192, 153, 167, 95, 102, 115, 129, 
    194, 238, 224, 242, 231, 212, 188, 170, 187, 199, 157, 104, 93, 115, 126, 
    187, 252, 242, 232, 246, 220, 215, 246, 142, 186, 194, 107, 118, 112, 130, 
    219, 221, 284, 252, 207, 339, 255, 186, 162, 203, 148, 40, 100, 99, 123, 
    193, 280, 281, 264, 272, 304, 239, 255, 289, 260, 126, 48, 84, 109, 99, 
    108, 282, 272, 244, 356, 323, 261, 332, 309, 312, 178, 50, 97, 210, 61, 
    150, 286, 298, 170, 337, 274, 206, 191, 216, 142, 33, 13, 107, 254, 78, 
    136, 282, 327, 82, 222, 258, 146, 304, 91, 34, 58, 55, 102, 317, 146, 
    164, 223, 263, 48, 60, 40, 70, 117, 37, 9, 23, 73, 95, 263, 213, 
    144, 197, 240, 223, 94, 131, 121, 45, 0, 1, 0, 7, 92, 100, 247, 
    177, 190, 179, 238, 171, 133, 169, 113, 74, 53, 26, 58, 70, 57, 132, 
    148, 180, 159, 148, 150, 164, 186, 138, 143, 124, 123, 161, 131, 132, 118, 
    176, 202, 168, 184, 183, 184, 153, 142, 134, 118, 156, 180, 158, 134, 149, 
    
    -- channel=336
    252, 268, 259, 271, 254, 233, 208, 202, 163, 116, 142, 133, 130, 183, 157, 
    351, 322, 269, 289, 291, 277, 239, 236, 172, 78, 127, 158, 202, 191, 160, 
    332, 317, 306, 314, 323, 307, 274, 247, 258, 201, 208, 180, 182, 185, 198, 
    305, 330, 320, 335, 339, 324, 302, 264, 277, 291, 251, 186, 150, 167, 199, 
    296, 335, 339, 328, 342, 329, 316, 325, 258, 274, 294, 203, 151, 180, 198, 
    212, 339, 363, 362, 321, 387, 411, 331, 260, 273, 264, 117, 125, 145, 180, 
    223, 373, 425, 384, 358, 436, 379, 331, 342, 353, 253, 110, 101, 135, 157, 
    202, 343, 421, 374, 461, 473, 408, 459, 466, 451, 310, 121, 113, 231, 154, 
    256, 371, 440, 329, 425, 409, 393, 322, 345, 304, 156, 26, 98, 299, 190, 
    261, 364, 480, 252, 259, 396, 305, 358, 241, 97, 74, 71, 115, 350, 273, 
    306, 340, 415, 172, 68, 106, 142, 216, 143, 43, 42, 77, 123, 330, 341, 
    287, 319, 345, 295, 181, 166, 185, 125, 0, 0, 0, 0, 87, 191, 309, 
    298, 318, 305, 353, 290, 240, 246, 197, 107, 52, 8, 15, 79, 88, 186, 
    281, 298, 307, 260, 256, 229, 294, 264, 212, 198, 167, 193, 175, 181, 187, 
    272, 323, 298, 298, 293, 304, 278, 261, 242, 219, 245, 275, 267, 228, 214, 
    
    -- channel=337
    187, 168, 166, 165, 168, 147, 141, 110, 129, 65, 66, 67, 52, 77, 101, 
    220, 227, 164, 175, 180, 180, 169, 144, 138, 57, 45, 76, 97, 107, 79, 
    228, 190, 188, 189, 198, 193, 187, 149, 178, 158, 108, 112, 87, 93, 102, 
    193, 191, 196, 197, 213, 200, 194, 175, 161, 173, 143, 143, 76, 68, 95, 
    156, 188, 206, 194, 211, 216, 189, 188, 163, 137, 170, 196, 78, 96, 97, 
    19, 181, 199, 225, 200, 217, 263, 202, 185, 133, 154, 102, 53, 78, 83, 
    53, 175, 255, 235, 188, 247, 221, 211, 175, 190, 173, 77, 35, 70, 78, 
    114, 106, 252, 203, 238, 285, 245, 248, 258, 254, 239, 105, 31, 114, 111, 
    150, 137, 250, 208, 233, 174, 261, 177, 192, 177, 133, 21, 0, 120, 184, 
    139, 118, 263, 247, 74, 207, 213, 187, 172, 50, 35, 54, 17, 125, 259, 
    178, 126, 228, 178, 0, 6, 49, 59, 118, 39, 19, 32, 42, 90, 275, 
    145, 148, 167, 202, 127, 89, 96, 87, 1, 0, 0, 0, 0, 55, 163, 
    143, 150, 148, 172, 229, 154, 105, 129, 81, 32, 7, 0, 17, 17, 63, 
    152, 105, 183, 113, 155, 106, 122, 153, 110, 114, 94, 105, 108, 98, 112, 
    121, 148, 153, 145, 155, 155, 148, 140, 126, 105, 120, 135, 145, 137, 102, 
    
    -- channel=338
    37, 85, 17, 9, 12, 15, 14, 36, 54, 66, 44, 50, 52, 49, 44, 
    31, 32, 15, 18, 7, 8, 6, 3, 24, 74, 51, 37, 28, 29, 40, 
    37, 35, 19, 8, 7, 2, 0, 9, 7, 52, 58, 35, 19, 20, 29, 
    36, 48, 15, 12, 9, 0, 0, 2, 0, 0, 14, 26, 24, 26, 22, 
    40, 27, 18, 13, 5, 2, 0, 4, 15, 0, 4, 37, 45, 36, 25, 
    40, 20, 19, 15, 18, 39, 49, 43, 21, 20, 13, 40, 66, 46, 31, 
    95, 11, 22, 16, 33, 50, 26, 35, 69, 61, 34, 57, 82, 55, 39, 
    30, 35, 13, 32, 41, 27, 18, 28, 42, 37, 41, 73, 86, 56, 58, 
    0, 32, 17, 41, 34, 2, 0, 14, 10, 23, 23, 68, 91, 48, 47, 
    0, 24, 24, 24, 65, 32, 0, 10, 18, 43, 64, 79, 82, 54, 53, 
    0, 8, 29, 21, 86, 47, 1, 0, 0, 73, 85, 62, 70, 49, 42, 
    0, 0, 31, 38, 61, 50, 49, 38, 80, 102, 111, 112, 60, 48, 26, 
    0, 0, 17, 24, 33, 10, 0, 22, 76, 103, 115, 122, 98, 47, 50, 
    0, 0, 0, 13, 11, 10, 0, 0, 22, 41, 53, 64, 63, 61, 45, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 23, 
    
    -- channel=339
    83, 0, 43, 33, 44, 35, 50, 31, 93, 49, 61, 68, 51, 44, 97, 
    25, 44, 22, 33, 32, 28, 44, 34, 88, 62, 37, 62, 62, 83, 64, 
    81, 10, 19, 21, 24, 28, 45, 7, 46, 86, 33, 80, 69, 66, 65, 
    60, 24, 27, 12, 29, 28, 52, 40, 24, 48, 47, 86, 70, 44, 62, 
    40, 18, 24, 18, 15, 41, 55, 52, 67, 20, 38, 126, 34, 62, 62, 
    0, 57, 9, 34, 30, 0, 106, 79, 85, 30, 85, 123, 30, 51, 49, 
    0, 0, 66, 62, 6, 42, 73, 109, 39, 51, 128, 109, 34, 41, 60, 
    97, 0, 80, 47, 7, 71, 57, 61, 79, 87, 149, 112, 20, 34, 106, 
    97, 0, 74, 80, 35, 15, 116, 60, 66, 89, 158, 85, 0, 4, 172, 
    115, 0, 79, 210, 0, 34, 145, 46, 149, 91, 67, 91, 0, 0, 225, 
    115, 20, 91, 214, 19, 35, 59, 38, 127, 78, 59, 56, 28, 0, 198, 
    99, 72, 60, 83, 109, 71, 64, 129, 74, 55, 70, 23, 4, 13, 74, 
    58, 90, 65, 32, 76, 92, 65, 117, 102, 78, 77, 41, 19, 41, 26, 
    102, 36, 117, 45, 103, 57, 52, 121, 75, 93, 74, 56, 71, 45, 104, 
    82, 63, 97, 71, 77, 84, 74, 84, 80, 77, 60, 60, 83, 92, 45, 
    
    -- channel=340
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    121, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 18, 0, 
    0, 39, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 48, 55, 0, 
    0, 0, 0, 0, 61, 6, 0, 0, 0, 0, 2, 0, 19, 84, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 52, 26, 34, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 50, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=341
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 16, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 10, 5, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 27, 32, 35, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 32, 40, 37, 3, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=342
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=343
    209, 220, 245, 254, 259, 260, 257, 224, 192, 159, 162, 161, 152, 163, 162, 
    234, 250, 249, 251, 266, 270, 278, 273, 238, 156, 158, 174, 187, 186, 168, 
    216, 228, 252, 263, 264, 276, 281, 270, 271, 210, 189, 193, 192, 192, 185, 
    191, 217, 252, 261, 272, 291, 282, 272, 261, 262, 233, 213, 185, 181, 184, 
    190, 222, 251, 257, 272, 265, 221, 216, 221, 249, 241, 214, 181, 184, 184, 
    162, 205, 227, 248, 248, 203, 164, 178, 208, 194, 197, 159, 153, 178, 181, 
    153, 210, 214, 219, 196, 200, 194, 166, 136, 150, 161, 132, 128, 169, 174, 
    184, 179, 209, 191, 189, 200, 229, 192, 162, 163, 169, 139, 125, 163, 155, 
    218, 182, 188, 189, 204, 178, 224, 222, 213, 195, 172, 129, 122, 161, 158, 
    215, 174, 164, 190, 142, 196, 210, 218, 202, 142, 121, 143, 141, 155, 145, 
    225, 191, 173, 161, 118, 122, 167, 194, 189, 143, 122, 140, 153, 157, 158, 
    216, 209, 168, 184, 184, 177, 182, 169, 112, 97, 91, 97, 135, 167, 175, 
    231, 215, 193, 187, 216, 214, 199, 190, 147, 111, 97, 96, 124, 138, 153, 
    215, 201, 218, 200, 193, 192, 206, 224, 186, 178, 175, 179, 176, 182, 172, 
    207, 215, 219, 213, 202, 219, 230, 223, 217, 206, 218, 219, 214, 210, 192, 
    
    -- channel=344
    132, 101, 121, 110, 122, 116, 105, 92, 116, 60, 55, 67, 54, 61, 77, 
    162, 172, 122, 131, 129, 124, 117, 99, 114, 72, 46, 59, 61, 86, 64, 
    194, 144, 142, 144, 146, 147, 139, 114, 110, 95, 53, 74, 70, 70, 73, 
    165, 152, 153, 144, 161, 149, 144, 131, 120, 124, 121, 123, 69, 60, 78, 
    137, 142, 154, 158, 157, 158, 140, 128, 143, 105, 127, 161, 56, 76, 77, 
    23, 165, 156, 171, 176, 136, 197, 169, 139, 93, 138, 121, 48, 67, 68, 
    48, 128, 198, 185, 139, 205, 188, 136, 105, 137, 153, 83, 44, 60, 71, 
    104, 77, 195, 166, 166, 201, 174, 172, 195, 188, 182, 91, 29, 59, 104, 
    96, 87, 184, 187, 193, 173, 219, 176, 173, 190, 168, 55, 10, 83, 158, 
    118, 95, 195, 236, 64, 158, 175, 72, 155, 79, 28, 33, 13, 70, 204, 
    130, 106, 202, 172, 52, 109, 85, 105, 122, 57, 51, 21, 32, 73, 213, 
    110, 114, 141, 120, 83, 21, 40, 93, 55, 23, 18, 23, 15, 84, 121, 
    97, 112, 145, 135, 140, 102, 62, 82, 48, 25, 19, 3, 30, 42, 95, 
    126, 84, 140, 112, 136, 81, 88, 115, 69, 66, 46, 42, 57, 57, 80, 
    87, 98, 107, 90, 99, 107, 116, 99, 101, 81, 78, 89, 102, 104, 61, 
    
    -- channel=345
    192, 223, 248, 279, 254, 250, 239, 215, 144, 143, 180, 161, 165, 206, 170, 
    232, 219, 244, 262, 278, 278, 270, 281, 199, 112, 170, 203, 239, 211, 193, 
    191, 223, 250, 270, 277, 273, 274, 273, 272, 196, 239, 222, 237, 228, 224, 
    168, 220, 248, 275, 272, 297, 297, 267, 278, 285, 243, 190, 203, 222, 227, 
    191, 243, 257, 252, 278, 274, 265, 281, 227, 295, 265, 149, 187, 204, 220, 
    211, 227, 267, 262, 225, 251, 203, 199, 185, 255, 220, 102, 159, 175, 211, 
    215, 262, 249, 236, 236, 224, 194, 216, 238, 218, 160, 111, 126, 165, 191, 
    204, 289, 250, 226, 261, 263, 276, 276, 232, 230, 170, 102, 130, 221, 151, 
    291, 308, 266, 176, 219, 231, 245, 209, 214, 168, 81, 63, 136, 233, 115, 
    283, 299, 254, 102, 204, 243, 219, 353, 208, 115, 130, 141, 168, 268, 112, 
    306, 288, 211, 93, 93, 76, 164, 238, 154, 87, 75, 144, 178, 260, 143, 
    301, 304, 227, 219, 199, 243, 251, 158, 41, 35, 31, 40, 144, 185, 213, 
    325, 317, 235, 245, 222, 246, 304, 237, 148, 98, 59, 68, 118, 134, 170, 
    290, 312, 277, 230, 206, 249, 314, 287, 247, 227, 213, 233, 205, 214, 198, 
    306, 335, 318, 318, 284, 313, 294, 290, 268, 272, 295, 301, 282, 247, 254, 
    
    -- channel=346
    0, 37, 23, 37, 13, 26, 6, 32, 0, 25, 30, 8, 25, 57, 0, 
    10, 0, 16, 27, 34, 22, 5, 32, 0, 0, 58, 38, 45, 10, 21, 
    0, 41, 24, 34, 33, 19, 4, 48, 7, 0, 47, 0, 44, 35, 26, 
    0, 42, 24, 44, 20, 28, 18, 17, 51, 23, 9, 0, 26, 54, 38, 
    24, 42, 23, 29, 30, 29, 19, 25, 0, 81, 30, 0, 48, 36, 38, 
    165, 7, 54, 23, 14, 67, 0, 29, 0, 74, 6, 0, 65, 29, 51, 
    177, 82, 5, 0, 32, 36, 0, 0, 47, 22, 0, 0, 43, 35, 41, 
    0, 176, 0, 28, 63, 0, 0, 43, 6, 0, 0, 0, 54, 59, 0, 
    7, 139, 9, 0, 72, 56, 0, 41, 38, 20, 0, 0, 102, 110, 0, 
    0, 158, 15, 0, 202, 62, 0, 88, 0, 0, 0, 0, 98, 160, 0, 
    0, 109, 11, 0, 62, 73, 43, 125, 0, 0, 28, 42, 61, 190, 0, 
    15, 52, 44, 0, 0, 6, 31, 0, 0, 10, 5, 57, 88, 95, 40, 
    47, 42, 23, 75, 0, 3, 52, 0, 0, 0, 0, 18, 73, 26, 92, 
    26, 92, 0, 38, 0, 38, 85, 0, 13, 0, 0, 27, 0, 32, 12, 
    37, 66, 13, 42, 7, 36, 40, 30, 26, 25, 49, 52, 16, 0, 42, 
    
    -- channel=347
    330, 312, 342, 364, 357, 338, 318, 275, 214, 158, 193, 177, 167, 209, 198, 
    366, 374, 352, 368, 386, 383, 370, 361, 283, 126, 169, 210, 257, 244, 209, 
    341, 351, 370, 391, 400, 401, 390, 358, 385, 282, 263, 251, 248, 251, 250, 
    305, 349, 376, 398, 407, 422, 408, 367, 370, 386, 329, 261, 223, 224, 249, 
    297, 349, 390, 386, 413, 408, 371, 376, 313, 355, 355, 269, 210, 235, 249, 
    212, 352, 381, 405, 371, 390, 354, 295, 304, 312, 293, 163, 165, 202, 230, 
    191, 368, 407, 386, 352, 380, 343, 329, 307, 312, 254, 135, 120, 186, 207, 
    244, 319, 398, 353, 404, 435, 416, 412, 380, 381, 292, 140, 130, 263, 188, 
    332, 354, 400, 301, 367, 344, 380, 324, 324, 271, 177, 66, 101, 282, 205, 
    335, 329, 393, 250, 229, 361, 339, 414, 289, 128, 113, 131, 140, 318, 261, 
    367, 330, 341, 217, 57, 66, 173, 240, 213, 96, 62, 137, 161, 287, 312, 
    353, 345, 319, 322, 255, 237, 247, 191, 27, 2, 1, 4, 121, 188, 308, 
    363, 373, 297, 335, 334, 319, 320, 276, 160, 88, 37, 36, 92, 125, 177, 
    328, 332, 352, 275, 279, 279, 335, 339, 271, 250, 231, 251, 235, 231, 241, 
    338, 359, 362, 353, 339, 362, 341, 340, 311, 289, 323, 345, 331, 300, 271, 
    
    -- channel=348
    145, 91, 80, 79, 81, 55, 57, 45, 85, 46, 60, 61, 49, 54, 91, 
    126, 132, 75, 87, 83, 78, 65, 53, 72, 31, 37, 53, 74, 80, 61, 
    148, 114, 91, 87, 95, 82, 81, 38, 86, 119, 73, 72, 52, 62, 74, 
    141, 119, 99, 93, 98, 80, 81, 68, 65, 86, 72, 76, 53, 38, 64, 
    109, 111, 113, 92, 97, 101, 123, 130, 87, 49, 83, 130, 49, 64, 70, 
    1, 128, 113, 123, 101, 144, 221, 131, 141, 90, 99, 87, 42, 51, 55, 
    6, 111, 178, 163, 128, 162, 167, 206, 167, 163, 150, 85, 45, 49, 53, 
    85, 60, 182, 141, 177, 221, 159, 188, 217, 225, 202, 99, 50, 107, 88, 
    95, 100, 194, 134, 168, 122, 164, 94, 118, 100, 109, 40, 5, 97, 167, 
    98, 66, 223, 191, 50, 142, 164, 151, 119, 51, 60, 65, 19, 103, 262, 
    115, 72, 179, 181, 0, 0, 32, 0, 78, 35, 26, 51, 33, 54, 268, 
    96, 94, 138, 176, 104, 85, 72, 81, 21, 15, 34, 0, 9, 9, 149, 
    76, 105, 90, 118, 146, 108, 80, 106, 91, 70, 53, 42, 19, 28, 29, 
    91, 59, 125, 61, 118, 78, 72, 106, 86, 99, 89, 90, 97, 65, 104, 
    88, 90, 105, 94, 117, 103, 73, 85, 73, 62, 70, 83, 94, 94, 64, 
    
    -- channel=349
    192, 257, 211, 229, 202, 182, 149, 167, 110, 96, 124, 104, 105, 173, 117, 
    314, 279, 218, 243, 244, 218, 172, 183, 98, 35, 122, 137, 187, 154, 131, 
    286, 303, 260, 265, 275, 247, 202, 185, 212, 147, 196, 132, 150, 154, 169, 
    255, 320, 277, 294, 291, 256, 235, 196, 237, 241, 188, 114, 113, 137, 170, 
    276, 310, 299, 280, 288, 275, 273, 291, 192, 236, 244, 135, 141, 157, 175, 
    239, 296, 331, 324, 264, 402, 393, 322, 220, 266, 218, 53, 131, 122, 163, 
    267, 372, 401, 350, 333, 449, 337, 304, 359, 357, 199, 66, 98, 119, 136, 
    156, 383, 390, 355, 480, 452, 368, 474, 471, 454, 254, 85, 124, 246, 104, 
    202, 399, 421, 275, 460, 383, 323, 303, 329, 275, 96, 0, 120, 332, 109, 
    192, 387, 481, 149, 343, 408, 232, 380, 169, 47, 49, 60, 135, 416, 206, 
    245, 338, 406, 81, 59, 81, 102, 195, 66, 12, 34, 82, 117, 397, 300, 
    227, 287, 338, 250, 147, 145, 161, 79, 0, 0, 0, 2, 99, 186, 321, 
    244, 280, 261, 347, 227, 206, 212, 142, 74, 39, 1, 25, 93, 55, 190, 
    222, 272, 248, 218, 207, 200, 274, 191, 176, 170, 139, 189, 146, 165, 174, 
    228, 287, 235, 259, 247, 267, 220, 214, 193, 160, 205, 241, 217, 175, 186, 
    
    -- channel=350
    176, 0, 38, 0, 55, 29, 64, 0, 144, 0, 0, 30, 0, 0, 95, 
    0, 76, 7, 19, 21, 28, 73, 20, 168, 55, 0, 0, 0, 58, 8, 
    139, 0, 0, 3, 7, 38, 85, 0, 54, 142, 0, 65, 4, 10, 5, 
    82, 0, 13, 0, 20, 25, 69, 46, 0, 36, 46, 148, 42, 0, 0, 
    0, 0, 2, 0, 4, 41, 45, 14, 94, 0, 0, 264, 0, 7, 0, 
    0, 53, 0, 16, 45, 0, 133, 33, 124, 0, 80, 218, 0, 0, 0, 
    0, 0, 51, 64, 0, 0, 82, 136, 0, 0, 202, 141, 0, 0, 0, 
    88, 0, 74, 0, 0, 63, 29, 0, 12, 46, 255, 146, 0, 0, 142, 
    77, 0, 29, 92, 0, 0, 179, 6, 5, 67, 293, 92, 0, 0, 337, 
    134, 0, 8, 455, 0, 0, 255, 0, 239, 97, 26, 61, 0, 0, 466, 
    118, 0, 47, 475, 0, 0, 15, 0, 222, 70, 1, 0, 0, 0, 376, 
    83, 0, 0, 113, 141, 0, 0, 177, 83, 5, 32, 0, 0, 0, 9, 
    0, 32, 0, 0, 120, 92, 0, 146, 105, 47, 48, 0, 0, 0, 0, 
    78, 0, 132, 0, 135, 0, 0, 146, 24, 57, 33, 0, 39, 0, 96, 
    27, 0, 72, 0, 33, 34, 32, 56, 49, 33, 0, 0, 51, 99, 0, 
    
    -- channel=351
    0, 8, 8, 10, 8, 15, 15, 13, 8, 28, 25, 19, 19, 18, 10, 
    0, 0, 2, 4, 5, 6, 13, 16, 10, 25, 32, 24, 17, 13, 17, 
    0, 0, 0, 0, 0, 2, 3, 17, 6, 0, 18, 14, 23, 19, 12, 
    0, 1, 0, 0, 0, 0, 0, 6, 11, 0, 2, 4, 24, 21, 14, 
    1, 0, 0, 0, 0, 0, 0, 0, 2, 12, 0, 0, 26, 22, 16, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 9, 39, 26, 20, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 35, 26, 24, 
    4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 35, 11, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 31, 40, 0, 0, 
    0, 0, 0, 0, 38, 0, 0, 0, 0, 20, 26, 35, 42, 0, 0, 
    0, 0, 0, 0, 30, 30, 25, 23, 17, 34, 41, 42, 32, 9, 0, 
    0, 0, 0, 0, 13, 14, 18, 25, 36, 47, 51, 57, 41, 25, 0, 
    0, 0, 0, 0, 0, 10, 5, 4, 14, 28, 36, 40, 46, 29, 18, 
    0, 2, 0, 0, 0, 3, 4, 0, 3, 7, 13, 13, 11, 17, 19, 
    0, 0, 0, 0, 0, 0, 2, 8, 7, 6, 11, 4, 0, 6, 7, 
    
    -- channel=352
    192, 122, 201, 202, 212, 213, 212, 179, 153, 116, 129, 125, 122, 122, 134, 
    164, 182, 208, 204, 216, 221, 237, 223, 207, 127, 117, 144, 146, 153, 145, 
    166, 156, 196, 214, 214, 232, 236, 233, 230, 157, 129, 166, 169, 168, 150, 
    166, 153, 198, 204, 217, 246, 249, 229, 217, 225, 212, 190, 162, 156, 160, 
    144, 157, 192, 210, 218, 227, 194, 181, 196, 215, 205, 174, 133, 151, 152, 
    105, 179, 174, 200, 207, 150, 113, 137, 159, 155, 177, 161, 103, 139, 145, 
    63, 160, 168, 167, 155, 134, 156, 119, 81, 105, 147, 117, 81, 124, 140, 
    163, 119, 166, 161, 119, 151, 184, 142, 118, 115, 129, 105, 76, 103, 140, 
    205, 128, 151, 161, 104, 163, 193, 185, 160, 162, 165, 103, 62, 104, 132, 
    222, 140, 118, 161, 86, 134, 203, 142, 196, 137, 94, 94, 78, 95, 112, 
    216, 169, 129, 176, 68, 113, 150, 189, 198, 116, 82, 100, 102, 108, 118, 
    228, 186, 138, 137, 159, 125, 135, 155, 91, 57, 42, 47, 96, 132, 130, 
    209, 217, 170, 149, 168, 181, 190, 179, 107, 67, 51, 33, 63, 118, 122, 
    204, 197, 207, 169, 159, 162, 182, 217, 163, 139, 131, 117, 125, 125, 139, 
    208, 183, 217, 196, 179, 197, 212, 215, 200, 201, 193, 195, 196, 185, 161, 
    
    -- channel=353
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=354
    0, 10, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 7, 0, 8, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 1, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 1, 0, 6, 0, 0, 2, 0, 1, 
    8, 0, 9, 0, 0, 5, 0, 0, 0, 11, 0, 0, 13, 0, 3, 
    46, 1, 0, 0, 0, 14, 0, 0, 22, 0, 0, 0, 0, 3, 1, 
    0, 41, 0, 0, 13, 0, 0, 16, 0, 2, 0, 0, 0, 25, 0, 
    0, 34, 0, 0, 57, 0, 0, 4, 8, 0, 0, 0, 7, 34, 0, 
    0, 32, 0, 0, 58, 8, 0, 49, 0, 0, 0, 7, 14, 51, 0, 
    0, 10, 5, 0, 11, 0, 0, 27, 0, 0, 0, 8, 4, 45, 0, 
    0, 9, 5, 0, 0, 0, 1, 0, 0, 0, 0, 3, 9, 0, 27, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 5, 16, 0, 21, 
    0, 0, 0, 0, 0, 4, 14, 0, 0, 0, 0, 12, 0, 1, 9, 
    0, 12, 0, 0, 0, 8, 0, 0, 0, 0, 2, 3, 0, 0, 0, 
    
    -- channel=355
    320, 342, 372, 403, 403, 400, 382, 335, 257, 207, 244, 233, 238, 257, 222, 
    343, 362, 382, 402, 425, 431, 429, 423, 352, 199, 236, 260, 293, 280, 257, 
    306, 361, 388, 414, 421, 433, 438, 429, 425, 304, 318, 290, 306, 296, 285, 
    270, 340, 385, 412, 419, 450, 443, 408, 407, 416, 370, 306, 281, 297, 293, 
    262, 351, 392, 404, 434, 417, 361, 381, 337, 404, 372, 267, 265, 274, 285, 
    269, 336, 399, 393, 374, 357, 247, 251, 269, 327, 302, 194, 226, 254, 280, 
    269, 336, 342, 338, 329, 317, 272, 269, 289, 274, 222, 160, 181, 254, 260, 
    280, 337, 326, 303, 323, 329, 362, 333, 267, 268, 232, 149, 168, 284, 216, 
    363, 342, 322, 252, 310, 294, 328, 316, 288, 234, 160, 137, 181, 293, 180, 
    359, 347, 276, 199, 240, 288, 289, 397, 304, 174, 174, 200, 205, 316, 180, 
    371, 335, 259, 183, 165, 149, 221, 327, 230, 154, 130, 195, 227, 292, 210, 
    353, 364, 276, 301, 272, 284, 301, 241, 114, 95, 79, 100, 201, 237, 278, 
    384, 381, 309, 296, 299, 313, 361, 309, 202, 149, 119, 125, 175, 191, 261, 
    353, 353, 342, 294, 267, 329, 367, 359, 308, 273, 274, 296, 274, 284, 254, 
    372, 382, 373, 373, 336, 385, 374, 360, 342, 337, 367, 375, 352, 331, 312, 
    
    -- channel=356
    19, 24, 28, 29, 29, 34, 42, 35, 43, 44, 38, 36, 39, 35, 40, 
    11, 12, 24, 20, 23, 30, 39, 33, 43, 52, 40, 44, 33, 33, 39, 
    5, 8, 18, 18, 15, 22, 29, 39, 33, 30, 35, 42, 39, 38, 33, 
    8, 4, 14, 15, 16, 23, 29, 34, 29, 24, 23, 40, 36, 39, 33, 
    6, 9, 11, 11, 17, 18, 7, 6, 25, 28, 26, 37, 41, 36, 30, 
    17, 0, 5, 6, 12, 0, 0, 21, 18, 13, 21, 42, 41, 41, 34, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 40, 40, 42, 38, 
    29, 3, 0, 0, 0, 0, 0, 0, 0, 0, 12, 45, 34, 17, 41, 
    36, 0, 0, 14, 0, 0, 10, 12, 7, 15, 31, 54, 41, 5, 30, 
    19, 1, 0, 23, 20, 0, 15, 7, 30, 44, 50, 53, 41, 0, 4, 
    22, 9, 0, 25, 35, 39, 34, 30, 48, 53, 53, 46, 42, 2, 0, 
    20, 15, 0, 14, 34, 44, 46, 40, 57, 64, 61, 56, 43, 35, 0, 
    25, 10, 13, 4, 36, 24, 24, 41, 45, 45, 53, 50, 48, 39, 34, 
    25, 19, 23, 20, 20, 25, 19, 26, 34, 36, 39, 35, 37, 41, 28, 
    19, 17, 21, 24, 16, 18, 29, 28, 28, 34, 30, 23, 26, 30, 35, 
    
    -- channel=357
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 43, 52, 11, 0, 0, 0, 0, 0, 0, 
    0, 4, 38, 13, 0, 28, 37, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 43, 16, 24, 62, 0, 57, 76, 70, 26, 0, 0, 0, 0, 
    0, 0, 48, 0, 67, 17, 41, 31, 44, 41, 35, 0, 0, 0, 0, 
    0, 0, 83, 21, 46, 29, 47, 16, 0, 0, 0, 0, 0, 0, 56, 
    0, 0, 72, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 103, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=358
    270, 259, 308, 318, 319, 304, 275, 250, 196, 136, 168, 149, 153, 193, 159, 
    344, 350, 315, 340, 350, 338, 312, 303, 232, 103, 163, 192, 225, 212, 184, 
    332, 351, 340, 365, 369, 370, 342, 329, 323, 192, 216, 193, 227, 225, 211, 
    305, 356, 358, 373, 387, 387, 375, 323, 342, 352, 296, 218, 193, 205, 229, 
    291, 344, 369, 371, 394, 370, 333, 331, 288, 340, 327, 227, 189, 213, 225, 
    236, 346, 383, 385, 368, 369, 332, 335, 275, 289, 283, 160, 163, 179, 214, 
    226, 376, 413, 373, 336, 407, 357, 260, 282, 302, 233, 105, 113, 170, 193, 
    225, 348, 396, 368, 402, 422, 382, 419, 400, 382, 255, 110, 118, 223, 160, 
    285, 350, 396, 303, 413, 393, 382, 378, 362, 330, 210, 64, 108, 295, 155, 
    296, 361, 403, 226, 323, 367, 323, 347, 267, 120, 77, 86, 129, 338, 211, 
    325, 350, 380, 191, 75, 169, 194, 313, 202, 69, 75, 115, 132, 336, 298, 
    322, 328, 329, 256, 192, 154, 189, 167, 22, 3, 0, 25, 129, 219, 324, 
    314, 352, 306, 361, 263, 260, 275, 208, 94, 37, 3, 12, 94, 109, 240, 
    308, 330, 329, 264, 262, 260, 322, 291, 222, 190, 170, 189, 169, 185, 211, 
    310, 321, 319, 312, 281, 334, 317, 307, 279, 256, 280, 308, 288, 258, 223, 
    
    -- channel=359
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=360
    42, 56, 44, 53, 48, 46, 38, 32, 15, 3, 7, 10, 4, 16, 12, 
    50, 47, 47, 49, 53, 57, 60, 52, 38, 9, 0, 8, 21, 22, 12, 
    41, 34, 54, 52, 60, 54, 58, 53, 59, 44, 33, 34, 24, 18, 25, 
    29, 36, 47, 55, 56, 60, 59, 57, 49, 48, 49, 37, 13, 20, 21, 
    15, 39, 51, 55, 54, 70, 52, 62, 43, 42, 51, 32, 11, 16, 18, 
    0, 42, 53, 61, 49, 60, 44, 16, 21, 37, 35, 0, 0, 11, 15, 
    21, 32, 50, 47, 48, 49, 16, 46, 45, 48, 22, 0, 0, 9, 11, 
    26, 27, 45, 34, 54, 50, 68, 52, 37, 35, 37, 2, 0, 25, 21, 
    45, 47, 51, 40, 27, 18, 45, 19, 14, 5, 0, 0, 0, 23, 23, 
    41, 37, 41, 27, 0, 44, 20, 50, 45, 0, 0, 5, 0, 31, 28, 
    51, 36, 23, 0, 0, 0, 0, 6, 0, 0, 0, 0, 12, 16, 14, 
    33, 51, 17, 45, 31, 29, 36, 15, 0, 0, 0, 0, 0, 6, 0, 
    50, 44, 40, 11, 58, 40, 36, 38, 17, 0, 0, 0, 0, 0, 7, 
    42, 27, 37, 33, 6, 27, 36, 41, 31, 28, 22, 34, 32, 33, 8, 
    30, 54, 42, 50, 47, 45, 44, 35, 33, 31, 41, 44, 45, 35, 35, 
    
    -- channel=361
    263, 321, 277, 307, 289, 262, 232, 212, 150, 92, 126, 118, 110, 168, 130, 
    365, 348, 292, 315, 329, 321, 283, 275, 198, 53, 107, 134, 197, 179, 139, 
    325, 346, 333, 343, 358, 340, 318, 279, 310, 232, 230, 175, 170, 171, 192, 
    277, 338, 339, 366, 365, 358, 329, 297, 302, 316, 259, 187, 134, 160, 185, 
    261, 347, 365, 353, 376, 370, 330, 363, 253, 288, 309, 204, 150, 167, 185, 
    190, 328, 390, 389, 330, 437, 391, 284, 251, 284, 246, 69, 111, 135, 168, 
    228, 368, 420, 389, 364, 434, 328, 341, 366, 357, 210, 62, 72, 133, 140, 
    182, 344, 405, 349, 472, 462, 418, 461, 430, 425, 289, 81, 79, 255, 123, 
    261, 381, 427, 290, 431, 350, 360, 287, 304, 230, 60, 0, 72, 306, 155, 
    245, 360, 448, 208, 213, 381, 253, 413, 223, 38, 45, 69, 94, 372, 247, 
    298, 317, 365, 100, 36, 2, 71, 174, 81, 10, 0, 53, 114, 310, 307, 
    253, 317, 311, 310, 171, 179, 200, 105, 0, 0, 0, 0, 59, 141, 289, 
    298, 303, 280, 313, 306, 245, 248, 199, 100, 37, 0, 0, 58, 46, 161, 
    266, 268, 282, 233, 214, 230, 284, 253, 209, 192, 170, 219, 188, 194, 166, 
    258, 327, 283, 301, 290, 303, 273, 245, 232, 198, 252, 282, 266, 227, 217, 
    
    -- channel=362
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=363
    0, 0, 17, 0, 0, 16, 23, 13, 27, 47, 20, 0, 0, 8, 7, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 15, 54, 63, 16, 12, 14, 
    25, 0, 0, 14, 0, 9, 0, 28, 0, 0, 0, 0, 54, 60, 0, 
    21, 16, 22, 10, 27, 38, 50, 31, 62, 17, 0, 0, 41, 13, 33, 
    83, 0, 0, 7, 3, 25, 0, 0, 11, 95, 44, 45, 46, 62, 39, 
    85, 0, 0, 0, 58, 0, 0, 195, 87, 6, 63, 99, 59, 46, 45, 
    3, 85, 16, 0, 0, 24, 72, 0, 0, 0, 8, 20, 6, 6, 55, 
    0, 48, 24, 57, 0, 0, 0, 0, 0, 0, 0, 42, 21, 0, 0, 
    0, 0, 0, 70, 105, 99, 95, 251, 227, 317, 316, 99, 13, 0, 0, 
    19, 32, 0, 70, 300, 100, 112, 0, 1, 105, 0, 0, 26, 0, 0, 
    24, 97, 107, 71, 0, 310, 231, 268, 247, 87, 136, 64, 0, 123, 0, 
    86, 16, 52, 0, 0, 0, 0, 42, 56, 56, 41, 95, 80, 174, 93, 
    13, 39, 32, 138, 0, 37, 0, 0, 0, 0, 0, 0, 14, 35, 118, 
    71, 110, 75, 65, 91, 0, 33, 14, 0, 0, 0, 0, 0, 0, 33, 
    6, 0, 12, 0, 0, 0, 64, 94, 51, 35, 0, 0, 0, 0, 0, 
    
    -- channel=364
    173, 109, 151, 137, 149, 147, 149, 119, 126, 89, 89, 101, 92, 84, 122, 
    124, 133, 152, 144, 144, 161, 180, 155, 160, 115, 64, 99, 100, 122, 109, 
    137, 81, 145, 143, 145, 162, 176, 158, 154, 166, 104, 157, 119, 112, 116, 
    141, 94, 135, 133, 151, 171, 176, 167, 136, 153, 165, 166, 116, 105, 112, 
    97, 102, 133, 141, 148, 155, 148, 133, 169, 124, 140, 158, 80, 101, 104, 
    0, 141, 109, 139, 143, 64, 128, 80, 124, 92, 133, 136, 50, 94, 94, 
    3, 70, 121, 123, 111, 72, 122, 133, 67, 93, 151, 117, 55, 81, 96, 
    142, 11, 126, 104, 67, 131, 162, 77, 89, 91, 157, 112, 46, 61, 146, 
    162, 50, 119, 147, 11, 95, 170, 81, 76, 86, 114, 72, 20, 27, 178, 
    175, 35, 88, 197, 0, 76, 183, 74, 191, 106, 92, 83, 36, 0, 174, 
    177, 77, 80, 181, 45, 26, 82, 65, 140, 93, 46, 49, 77, 0, 124, 
    174, 129, 74, 155, 162, 127, 131, 126, 78, 35, 31, 13, 30, 66, 37, 
    162, 147, 128, 69, 179, 150, 132, 164, 126, 84, 67, 35, 32, 92, 36, 
    155, 113, 163, 127, 120, 115, 118, 181, 131, 133, 125, 103, 130, 109, 97, 
    141, 143, 175, 149, 160, 151, 154, 149, 148, 158, 140, 137, 160, 152, 123, 
    
    -- channel=365
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=366
    0, 38, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 28, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 15, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 1, 0, 0, 34, 0, 0, 0, 0, 
    0, 13, 0, 9, 0, 0, 0, 0, 4, 0, 0, 0, 0, 14, 0, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 16, 0, 0, 
    133, 0, 17, 0, 0, 48, 0, 0, 0, 34, 0, 0, 28, 0, 13, 
    155, 49, 0, 0, 14, 14, 0, 0, 38, 13, 0, 0, 17, 6, 0, 
    0, 140, 0, 0, 52, 0, 0, 26, 0, 0, 0, 0, 35, 42, 0, 
    0, 116, 0, 0, 44, 21, 0, 0, 0, 0, 0, 0, 84, 86, 0, 
    0, 120, 0, 0, 132, 32, 0, 65, 0, 0, 0, 0, 76, 139, 0, 
    0, 69, 0, 0, 48, 3, 0, 47, 0, 0, 0, 5, 40, 151, 0, 
    0, 16, 9, 0, 0, 6, 20, 0, 0, 0, 0, 24, 54, 49, 4, 
    3, 0, 0, 26, 0, 0, 9, 0, 0, 0, 0, 20, 48, 0, 46, 
    0, 38, 0, 9, 0, 7, 39, 0, 0, 0, 0, 26, 0, 19, 0, 
    0, 28, 0, 6, 0, 0, 0, 0, 0, 0, 7, 11, 0, 0, 14, 
    
    -- channel=367
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=368
    25, 44, 30, 40, 28, 20, 9, 24, 0, 20, 33, 18, 36, 44, 15, 
    60, 42, 38, 44, 39, 35, 9, 21, 0, 0, 43, 32, 45, 21, 33, 
    28, 78, 46, 48, 50, 35, 19, 32, 26, 3, 45, 8, 28, 35, 34, 
    57, 69, 50, 58, 47, 35, 28, 18, 42, 41, 27, 0, 22, 39, 40, 
    55, 75, 58, 51, 56, 34, 60, 67, 17, 57, 46, 0, 42, 31, 41, 
    143, 56, 86, 57, 41, 115, 59, 58, 39, 73, 27, 0, 43, 26, 44, 
    93, 116, 79, 65, 93, 81, 72, 62, 103, 89, 14, 0, 39, 32, 29, 
    16, 136, 74, 81, 128, 99, 61, 111, 108, 103, 14, 0, 57, 75, 0, 
    29, 125, 96, 27, 113, 121, 29, 58, 68, 34, 0, 0, 70, 111, 0, 
    23, 127, 119, 0, 142, 92, 27, 105, 0, 1, 25, 0, 58, 149, 0, 
    29, 94, 85, 0, 20, 34, 40, 58, 0, 0, 13, 39, 37, 136, 29, 
    45, 57, 87, 55, 0, 31, 28, 0, 0, 2, 0, 19, 64, 45, 95, 
    50, 63, 45, 98, 22, 25, 67, 5, 0, 5, 0, 24, 29, 32, 59, 
    31, 85, 32, 41, 27, 55, 69, 18, 39, 21, 27, 40, 23, 29, 25, 
    62, 59, 47, 55, 51, 52, 33, 41, 28, 35, 45, 54, 36, 20, 46, 
    
    -- channel=369
    236, 249, 204, 215, 222, 210, 211, 185, 158, 122, 135, 140, 141, 138, 138, 
    206, 217, 215, 223, 234, 241, 234, 229, 217, 122, 119, 130, 156, 151, 143, 
    181, 210, 219, 224, 230, 235, 239, 216, 248, 239, 213, 171, 137, 147, 157, 
    165, 195, 211, 227, 220, 233, 216, 215, 198, 220, 203, 174, 144, 146, 144, 
    152, 201, 220, 219, 236, 222, 193, 220, 170, 177, 190, 161, 139, 139, 145, 
    133, 194, 224, 217, 198, 239, 174, 101, 151, 170, 141, 101, 119, 137, 137, 
    127, 172, 191, 196, 212, 171, 168, 227, 222, 183, 136, 108, 114, 145, 126, 
    149, 160, 183, 168, 206, 218, 218, 191, 167, 183, 167, 103, 115, 199, 127, 
    184, 183, 189, 136, 148, 139, 148, 103, 112, 60, 44, 79, 108, 163, 135, 
    167, 162, 164, 114, 78, 135, 143, 252, 150, 90, 123, 138, 119, 184, 164, 
    172, 141, 124, 130, 80, 0, 62, 59, 86, 84, 59, 116, 133, 124, 166, 
    157, 162, 158, 235, 195, 212, 190, 124, 71, 71, 72, 47, 99, 74, 161, 
    181, 175, 141, 153, 194, 160, 177, 194, 171, 147, 126, 134, 105, 105, 80, 
    144, 134, 160, 133, 148, 170, 163, 178, 181, 180, 197, 213, 206, 180, 156, 
    181, 186, 179, 189, 197, 187, 166, 159, 160, 156, 183, 189, 184, 178, 176, 
    
    -- channel=370
    83, 0, 17, 0, 12, 7, 33, 0, 82, 12, 0, 5, 0, 0, 52, 
    0, 26, 6, 0, 0, 0, 23, 0, 73, 46, 0, 7, 0, 22, 11, 
    65, 0, 0, 0, 0, 14, 23, 0, 12, 38, 0, 30, 0, 12, 0, 
    70, 0, 4, 0, 7, 14, 34, 25, 0, 14, 28, 73, 18, 0, 0, 
    28, 0, 0, 0, 0, 9, 0, 0, 43, 0, 3, 129, 0, 8, 0, 
    0, 19, 0, 0, 35, 0, 36, 49, 66, 0, 37, 142, 0, 1, 0, 
    0, 0, 17, 14, 0, 0, 81, 10, 0, 0, 104, 85, 0, 0, 0, 
    43, 0, 32, 18, 0, 16, 6, 0, 6, 6, 100, 89, 0, 0, 76, 
    27, 0, 0, 81, 0, 0, 95, 47, 40, 103, 222, 73, 0, 0, 155, 
    59, 0, 0, 223, 0, 0, 156, 0, 114, 91, 4, 1, 0, 0, 176, 
    46, 0, 35, 261, 0, 46, 48, 0, 167, 58, 27, 0, 0, 0, 158, 
    66, 0, 5, 7, 69, 0, 0, 82, 64, 18, 19, 0, 0, 0, 3, 
    0, 14, 6, 1, 52, 32, 0, 53, 34, 3, 7, 0, 0, 4, 0, 
    29, 0, 76, 0, 83, 0, 0, 63, 0, 11, 0, 0, 0, 0, 46, 
    5, 0, 32, 0, 2, 0, 19, 35, 28, 24, 0, 0, 16, 35, 0, 
    
    -- channel=371
    177, 153, 161, 160, 173, 173, 174, 163, 152, 136, 127, 128, 131, 116, 122, 
    163, 177, 179, 167, 172, 177, 179, 170, 172, 144, 131, 125, 118, 121, 129, 
    149, 175, 173, 177, 175, 183, 180, 186, 185, 147, 126, 122, 120, 131, 123, 
    167, 158, 173, 175, 175, 183, 171, 176, 169, 167, 163, 152, 131, 129, 124, 
    147, 155, 170, 180, 183, 174, 145, 140, 143, 156, 161, 154, 141, 131, 125, 
    173, 145, 160, 167, 185, 174, 97, 119, 152, 132, 128, 149, 134, 139, 128, 
    113, 160, 138, 146, 160, 134, 149, 110, 102, 108, 116, 121, 127, 141, 125, 
    117, 129, 129, 145, 133, 128, 138, 118, 106, 107, 107, 121, 132, 124, 116, 
    120, 113, 116, 138, 131, 145, 120, 155, 139, 135, 145, 144, 133, 126, 112, 
    116, 122, 98, 116, 142, 125, 128, 108, 112, 135, 122, 111, 123, 127, 92, 
    107, 122, 110, 135, 117, 139, 134, 126, 152, 140, 130, 131, 119, 124, 108, 
    119, 105, 127, 132, 121, 109, 103, 118, 140, 137, 126, 133, 140, 125, 138, 
    118, 114, 121, 139, 144, 120, 114, 119, 116, 117, 118, 125, 119, 135, 127, 
    104, 118, 116, 129, 128, 125, 105, 116, 122, 106, 122, 115, 123, 122, 116, 
    119, 93, 112, 111, 115, 106, 125, 126, 124, 122, 123, 125, 120, 127, 126, 
    
    -- channel=372
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=373
    207, 0, 86, 61, 101, 77, 116, 47, 132, 40, 44, 60, 41, 0, 115, 
    57, 101, 91, 75, 77, 92, 118, 87, 168, 73, 0, 43, 32, 79, 65, 
    112, 25, 63, 75, 73, 101, 128, 71, 113, 155, 0, 92, 41, 69, 55, 
    143, 13, 74, 52, 77, 104, 119, 109, 56, 104, 111, 145, 81, 24, 48, 
    63, 22, 64, 65, 80, 82, 95, 60, 106, 30, 75, 195, 15, 47, 49, 
    0, 88, 12, 61, 95, 0, 79, 20, 149, 0, 82, 194, 0, 45, 22, 
    0, 0, 63, 84, 34, 0, 141, 137, 0, 0, 161, 136, 0, 19, 32, 
    91, 0, 89, 51, 0, 90, 71, 0, 29, 57, 172, 120, 0, 0, 109, 
    110, 0, 58, 99, 0, 39, 138, 36, 47, 66, 239, 114, 0, 0, 237, 
    152, 0, 34, 277, 0, 0, 243, 0, 151, 131, 73, 40, 0, 0, 276, 
    125, 0, 46, 358, 0, 0, 90, 0, 231, 85, 22, 39, 0, 0, 243, 
    149, 18, 47, 140, 123, 58, 15, 121, 94, 28, 28, 0, 0, 0, 62, 
    69, 90, 34, 28, 139, 101, 65, 146, 106, 56, 44, 0, 0, 61, 0, 
    88, 16, 141, 35, 149, 42, 0, 163, 83, 78, 81, 9, 71, 0, 90, 
    103, 10, 133, 56, 97, 61, 77, 108, 91, 104, 55, 54, 95, 115, 37, 
    
    -- channel=374
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=375
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=376
    0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 4, 0, 4, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 4, 9, 1, 0, 7, 
    0, 0, 0, 25, 0, 0, 10, 0, 0, 6, 0, 0, 6, 0, 14, 
    0, 0, 0, 21, 0, 13, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 10, 2, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 9, 0, 16, 0, 
    1, 0, 8, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=377
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=378
    43, 47, 44, 42, 41, 43, 52, 65, 57, 88, 84, 79, 83, 76, 73, 
    25, 23, 43, 35, 35, 34, 39, 50, 54, 81, 89, 78, 76, 65, 78, 
    14, 34, 31, 31, 28, 27, 29, 40, 48, 61, 71, 67, 67, 73, 71, 
    34, 31, 29, 30, 20, 27, 25, 40, 41, 40, 45, 44, 75, 74, 67, 
    51, 32, 25, 27, 19, 27, 34, 34, 27, 48, 42, 34, 82, 73, 70, 
    108, 28, 17, 18, 21, 47, 8, 24, 50, 61, 37, 62, 88, 79, 74, 
    76, 51, 8, 17, 39, 5, 25, 47, 43, 33, 35, 78, 92, 80, 74, 
    58, 68, 10, 31, 28, 2, 14, 24, 14, 20, 13, 74, 107, 77, 55, 
    48, 65, 11, 19, 20, 34, 0, 29, 34, 29, 51, 101, 111, 69, 32, 
    43, 58, 12, 0, 91, 35, 22, 63, 24, 88, 97, 92, 109, 78, 8, 
    31, 56, 16, 36, 94, 72, 76, 54, 59, 96, 98, 107, 94, 79, 11, 
    49, 41, 50, 32, 66, 89, 77, 71, 98, 114, 119, 112, 110, 70, 63, 
    46, 45, 33, 49, 27, 58, 64, 57, 88, 105, 107, 119, 97, 100, 58, 
    36, 59, 31, 58, 48, 59, 52, 42, 68, 70, 82, 80, 76, 72, 76, 
    54, 42, 43, 50, 52, 37, 41, 50, 54, 59, 58, 54, 48, 51, 72, 
    
    -- channel=379
    178, 219, 220, 243, 223, 208, 172, 167, 85, 62, 94, 76, 87, 136, 82, 
    283, 255, 238, 254, 259, 253, 217, 216, 115, 21, 91, 112, 156, 131, 112, 
    231, 271, 267, 278, 289, 273, 244, 240, 230, 128, 168, 126, 147, 142, 146, 
    226, 269, 273, 297, 298, 294, 272, 229, 254, 257, 213, 125, 106, 140, 157, 
    209, 281, 292, 289, 308, 285, 267, 280, 203, 262, 253, 104, 120, 130, 151, 
    225, 267, 323, 307, 265, 338, 276, 236, 178, 236, 194, 33, 84, 99, 143, 
    211, 328, 334, 298, 300, 342, 269, 221, 267, 276, 142, 19, 50, 95, 113, 
    138, 323, 320, 291, 382, 363, 328, 369, 346, 326, 175, 23, 63, 180, 73, 
    208, 333, 344, 223, 341, 342, 287, 260, 262, 203, 36, 0, 76, 258, 59, 
    206, 335, 364, 88, 224, 319, 203, 307, 152, 21, 18, 7, 82, 319, 99, 
    245, 300, 298, 24, 29, 52, 95, 208, 62, 0, 0, 30, 86, 301, 171, 
    235, 273, 254, 216, 101, 114, 141, 48, 0, 0, 0, 0, 68, 152, 225, 
    263, 273, 241, 276, 210, 182, 224, 128, 28, 0, 0, 0, 33, 47, 162, 
    226, 275, 231, 207, 155, 197, 262, 201, 161, 127, 108, 142, 113, 136, 105, 
    236, 281, 248, 257, 234, 260, 235, 219, 195, 185, 214, 240, 217, 170, 178, 
    
    -- channel=380
    270, 318, 300, 324, 312, 285, 249, 233, 175, 120, 145, 125, 119, 178, 137, 
    418, 411, 318, 345, 353, 334, 285, 282, 188, 57, 144, 156, 210, 186, 149, 
    377, 421, 368, 383, 391, 373, 331, 301, 316, 199, 209, 151, 177, 190, 194, 
    344, 411, 390, 408, 414, 390, 352, 316, 338, 341, 264, 181, 148, 162, 197, 
    338, 400, 414, 399, 422, 388, 352, 357, 267, 325, 336, 231, 185, 193, 207, 
    292, 363, 427, 429, 392, 473, 424, 375, 325, 309, 270, 107, 155, 162, 194, 
    268, 457, 484, 445, 401, 510, 421, 325, 348, 366, 230, 72, 107, 156, 163, 
    183, 408, 466, 416, 535, 518, 434, 511, 502, 487, 295, 101, 129, 261, 113, 
    236, 412, 467, 337, 562, 450, 407, 407, 420, 354, 182, 26, 117, 353, 151, 
    232, 397, 515, 237, 374, 464, 309, 413, 204, 72, 43, 54, 130, 420, 247, 
    285, 359, 460, 140, 56, 123, 163, 249, 144, 36, 52, 95, 118, 393, 365, 
    264, 313, 376, 294, 143, 129, 154, 104, 0, 0, 0, 7, 115, 203, 382, 
    287, 306, 302, 404, 304, 257, 234, 153, 63, 12, 0, 4, 83, 75, 220, 
    265, 300, 299, 262, 266, 235, 290, 237, 190, 167, 146, 186, 156, 175, 189, 
    256, 302, 272, 279, 273, 296, 276, 262, 239, 192, 244, 279, 252, 223, 202, 
    
    -- channel=381
    261, 217, 257, 253, 263, 246, 227, 187, 185, 103, 109, 107, 94, 119, 127, 
    319, 335, 264, 279, 289, 279, 259, 234, 209, 95, 95, 123, 139, 154, 124, 
    337, 307, 294, 308, 314, 316, 296, 259, 267, 180, 139, 141, 140, 150, 146, 
    287, 306, 314, 314, 335, 322, 310, 272, 273, 276, 235, 208, 135, 124, 153, 
    260, 292, 319, 318, 339, 327, 286, 270, 253, 247, 263, 259, 128, 152, 156, 
    119, 296, 321, 343, 334, 318, 335, 302, 257, 212, 239, 167, 104, 129, 141, 
    110, 290, 371, 345, 287, 369, 333, 249, 220, 247, 233, 106, 70, 117, 132, 
    164, 210, 360, 317, 340, 391, 333, 344, 352, 343, 281, 119, 63, 155, 146, 
    202, 213, 347, 295, 362, 318, 370, 311, 311, 301, 234, 56, 32, 193, 205, 
    216, 221, 360, 306, 206, 300, 304, 239, 231, 104, 46, 49, 48, 204, 282, 
    247, 222, 338, 246, 24, 130, 147, 183, 201, 61, 54, 63, 63, 195, 336, 
    229, 220, 267, 235, 153, 79, 96, 129, 35, 2, 0, 1, 50, 137, 258, 
    212, 237, 233, 290, 266, 203, 164, 154, 67, 16, 0, 0, 45, 62, 151, 
    228, 200, 261, 188, 243, 170, 199, 216, 149, 130, 103, 111, 115, 117, 160, 
    200, 207, 224, 203, 203, 227, 227, 221, 197, 165, 179, 206, 206, 197, 144, 
    
    -- channel=382
    106, 72, 91, 93, 94, 79, 66, 41, 45, 0, 10, 9, 2, 21, 32, 
    127, 131, 89, 106, 108, 104, 91, 78, 55, 0, 0, 22, 44, 50, 22, 
    142, 110, 109, 115, 120, 120, 113, 77, 92, 67, 44, 45, 41, 38, 43, 
    113, 121, 120, 118, 137, 127, 127, 89, 94, 112, 81, 63, 25, 20, 45, 
    90, 115, 130, 117, 137, 119, 121, 120, 103, 83, 92, 90, 10, 33, 44, 
    0, 132, 134, 142, 121, 104, 184, 124, 98, 71, 95, 30, 0, 11, 30, 
    0, 105, 181, 158, 109, 170, 154, 130, 110, 121, 107, 8, 0, 4, 23, 
    62, 60, 181, 133, 156, 214, 168, 171, 190, 186, 152, 16, 0, 47, 44, 
    97, 84, 184, 122, 157, 132, 196, 113, 122, 107, 65, 0, 0, 61, 95, 
    106, 72, 195, 153, 22, 131, 159, 122, 117, 0, 0, 0, 0, 60, 172, 
    133, 82, 165, 115, 0, 0, 17, 41, 45, 0, 0, 0, 0, 42, 189, 
    113, 109, 108, 131, 64, 29, 37, 26, 0, 0, 0, 0, 0, 9, 100, 
    103, 121, 100, 109, 116, 85, 76, 72, 5, 0, 0, 0, 0, 0, 19, 
    107, 83, 134, 60, 97, 69, 94, 114, 55, 58, 35, 39, 39, 29, 51, 
    98, 112, 121, 103, 103, 126, 97, 96, 81, 68, 75, 91, 97, 83, 42, 
    
    -- channel=383
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=384
    247, 248, 271, 269, 251, 223, 223, 195, 179, 146, 138, 121, 45, 72, 88, 
    241, 217, 202, 186, 172, 154, 157, 147, 136, 123, 126, 71, 22, 71, 92, 
    168, 147, 140, 128, 130, 120, 123, 130, 128, 130, 108, 43, 54, 106, 102, 
    109, 109, 111, 110, 120, 121, 125, 131, 136, 132, 30, 52, 96, 113, 105, 
    102, 107, 109, 110, 121, 134, 142, 136, 128, 67, 0, 51, 90, 99, 102, 
    107, 106, 108, 110, 119, 123, 137, 139, 159, 135, 101, 0, 87, 66, 86, 
    110, 106, 102, 110, 114, 97, 54, 12, 36, 100, 158, 0, 0, 62, 63, 
    109, 105, 114, 77, 46, 70, 35, 25, 65, 126, 118, 19, 0, 30, 63, 
    102, 109, 47, 64, 19, 53, 101, 179, 147, 137, 78, 0, 41, 49, 104, 
    112, 148, 0, 29, 0, 44, 126, 127, 106, 96, 164, 47, 71, 74, 64, 
    137, 130, 0, 0, 0, 37, 107, 106, 43, 0, 47, 177, 64, 55, 5, 
    91, 17, 48, 0, 22, 65, 131, 102, 0, 19, 3, 95, 80, 0, 17, 
    63, 39, 59, 0, 54, 40, 109, 90, 0, 54, 0, 11, 106, 0, 36, 
    51, 49, 54, 23, 72, 84, 91, 84, 11, 61, 10, 0, 36, 0, 20, 
    55, 15, 0, 0, 0, 0, 0, 0, 1, 55, 20, 0, 10, 14, 28, 
    
    -- channel=385
    258, 270, 284, 283, 286, 272, 264, 253, 238, 220, 197, 176, 125, 112, 170, 
    284, 272, 284, 294, 285, 263, 253, 237, 223, 206, 166, 143, 87, 95, 191, 
    255, 272, 268, 263, 240, 236, 235, 216, 208, 194, 143, 100, 84, 137, 195, 
    224, 232, 231, 231, 230, 237, 231, 209, 196, 174, 116, 58, 163, 194, 206, 
    226, 242, 244, 244, 239, 227, 193, 191, 128, 119, 55, 45, 171, 197, 193, 
    240, 246, 241, 238, 209, 137, 107, 130, 156, 164, 52, 53, 72, 163, 187, 
    243, 249, 247, 209, 172, 131, 131, 106, 99, 0, 63, 136, 12, 107, 149, 
    247, 246, 180, 143, 105, 72, 57, 0, 0, 0, 78, 200, 109, 16, 34, 
    253, 194, 102, 89, 82, 27, 0, 50, 103, 118, 140, 153, 83, 10, 64, 
    203, 99, 88, 45, 66, 30, 0, 86, 92, 160, 155, 94, 42, 76, 124, 
    176, 150, 130, 59, 44, 0, 0, 76, 162, 114, 49, 101, 124, 130, 139, 
    172, 49, 77, 60, 1, 10, 3, 76, 160, 37, 48, 5, 96, 122, 60, 
    139, 61, 57, 24, 0, 0, 6, 75, 136, 21, 50, 31, 82, 108, 55, 
    124, 92, 90, 82, 77, 136, 149, 161, 169, 40, 85, 57, 45, 55, 33, 
    125, 65, 7, 8, 0, 2, 9, 21, 25, 36, 94, 52, 19, 16, 10, 
    
    -- channel=386
    394, 364, 362, 346, 335, 316, 311, 288, 283, 224, 224, 214, 122, 92, 199, 
    358, 344, 334, 333, 319, 296, 293, 271, 261, 248, 247, 180, 77, 149, 232, 
    276, 277, 283, 291, 279, 282, 286, 268, 266, 269, 223, 101, 138, 214, 237, 
    252, 276, 282, 281, 289, 301, 314, 305, 286, 271, 92, 59, 203, 228, 230, 
    275, 293, 294, 294, 303, 303, 272, 308, 336, 313, 138, 119, 211, 228, 224, 
    294, 301, 293, 285, 298, 320, 308, 276, 229, 178, 298, 119, 61, 203, 213, 
    300, 303, 291, 280, 269, 180, 101, 9, 43, 166, 323, 207, 58, 70, 148, 
    301, 302, 287, 267, 152, 143, 129, 201, 308, 381, 331, 147, 101, 86, 202, 
    303, 308, 171, 103, 59, 43, 134, 352, 323, 318, 292, 110, 233, 269, 278, 
    324, 402, 148, 94, 20, 48, 186, 288, 279, 195, 205, 316, 317, 253, 184, 
    318, 169, 96, 67, 9, 107, 223, 270, 180, 20, 45, 156, 214, 143, 20, 
    247, 112, 139, 46, 63, 136, 246, 286, 104, 81, 52, 108, 187, 68, 42, 
    190, 124, 145, 80, 176, 249, 291, 263, 104, 125, 120, 66, 110, 3, 48, 
    175, 129, 71, 19, 33, 23, 22, 22, 0, 111, 75, 18, 9, 0, 33, 
    175, 125, 72, 70, 46, 54, 51, 45, 30, 52, 54, 4, 13, 16, 31, 
    
    -- channel=387
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 41, 35, 52, 0, 82, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 211, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 191, 189, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 216, 195, 185, 164, 0, 0, 0, 88, 
    0, 87, 0, 0, 0, 0, 6, 166, 147, 104, 84, 50, 87, 79, 37, 
    0, 16, 0, 0, 0, 0, 53, 137, 86, 0, 0, 80, 71, 19, 0, 
    0, 0, 0, 0, 0, 0, 97, 144, 0, 0, 0, 0, 35, 0, 0, 
    0, 0, 0, 0, 0, 34, 148, 126, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=388
    19, 17, 21, 18, 12, 3, 4, 0, 0, 0, 1, 0, 9, 8, 0, 
    1, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 27, 22, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 20, 20, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 5, 25, 60, 45, 40, 7, 0, 0, 
    0, 0, 0, 0, 0, 3, 78, 111, 117, 78, 125, 102, 6, 21, 0, 
    0, 0, 0, 0, 14, 49, 56, 31, 15, 24, 148, 124, 46, 3, 0, 
    0, 0, 0, 27, 36, 41, 42, 50, 91, 187, 175, 132, 37, 1, 47, 
    0, 0, 33, 31, 52, 33, 36, 163, 185, 169, 180, 51, 0, 68, 105, 
    0, 59, 94, 34, 25, 13, 63, 149, 155, 161, 97, 119, 132, 128, 126, 
    0, 65, 74, 46, 6, 17, 93, 148, 165, 30, 59, 59, 131, 117, 43, 
    0, 37, 64, 37, 12, 63, 102, 160, 109, 31, 24, 43, 82, 77, 8, 
    0, 26, 63, 44, 55, 101, 145, 151, 108, 31, 53, 39, 55, 30, 4, 
    0, 16, 53, 37, 53, 54, 61, 61, 20, 40, 33, 22, 12, 0, 1, 
    0, 10, 23, 41, 22, 24, 27, 17, 12, 15, 30, 6, 4, 6, 12, 
    
    -- channel=389
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 88, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 30, 40, 172, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 26, 0, 0, 0, 269, 35, 0, 0, 
    0, 0, 0, 0, 24, 0, 36, 11, 0, 0, 52, 195, 74, 0, 0, 
    0, 0, 11, 0, 50, 0, 0, 0, 42, 56, 112, 201, 0, 0, 0, 
    0, 0, 194, 0, 60, 0, 0, 1, 48, 71, 0, 128, 37, 48, 55, 
    0, 0, 129, 21, 19, 0, 0, 32, 107, 90, 0, 0, 82, 59, 96, 
    0, 8, 6, 82, 0, 0, 0, 56, 236, 0, 22, 0, 0, 142, 0, 
    0, 0, 0, 96, 0, 24, 0, 57, 236, 0, 64, 0, 0, 123, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 82, 0, 44, 43, 0, 9, 0, 
    0, 13, 17, 35, 5, 3, 4, 2, 0, 0, 9, 27, 0, 0, 0, 
    
    -- channel=390
    169, 171, 179, 177, 168, 160, 159, 145, 143, 113, 112, 100, 77, 83, 94, 
    180, 168, 162, 155, 147, 138, 138, 129, 125, 114, 128, 97, 48, 90, 103, 
    141, 131, 129, 130, 127, 125, 126, 124, 120, 125, 109, 74, 89, 107, 106, 
    116, 119, 122, 119, 126, 126, 134, 135, 135, 128, 60, 68, 87, 104, 104, 
    118, 121, 122, 120, 128, 129, 135, 146, 173, 150, 75, 91, 115, 111, 108, 
    120, 123, 122, 120, 132, 156, 155, 142, 124, 91, 130, 61, 78, 103, 104, 
    125, 123, 114, 123, 127, 114, 65, 35, 41, 128, 175, 51, 64, 67, 90, 
    124, 120, 131, 130, 93, 89, 78, 122, 177, 204, 160, 41, 31, 70, 120, 
    121, 133, 107, 78, 48, 68, 116, 177, 159, 149, 126, 31, 110, 136, 144, 
    134, 189, 66, 70, 27, 56, 138, 149, 134, 90, 99, 119, 159, 127, 88, 
    140, 107, 25, 50, 27, 90, 160, 135, 73, 19, 70, 107, 92, 68, 21, 
    109, 67, 73, 36, 63, 102, 148, 137, 25, 62, 46, 109, 90, 31, 39, 
    95, 73, 87, 52, 123, 134, 168, 130, 23, 90, 64, 61, 82, 3, 55, 
    87, 65, 50, 24, 53, 39, 37, 34, 0, 81, 49, 29, 49, 17, 51, 
    88, 72, 67, 57, 55, 58, 55, 49, 44, 69, 36, 24, 42, 44, 54, 
    
    -- channel=391
    0, 6, 0, 1, 7, 6, 0, 16, 0, 0, 4, 5, 29, 0, 0, 
    0, 11, 8, 7, 3, 5, 0, 6, 0, 2, 0, 37, 29, 0, 0, 
    3, 6, 3, 5, 0, 0, 0, 0, 0, 0, 0, 35, 4, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 55, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 55, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 8, 0, 150, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 4, 30, 0, 0, 0, 161, 53, 0, 0, 
    0, 1, 0, 7, 1, 0, 10, 0, 0, 0, 0, 144, 57, 0, 0, 
    0, 0, 26, 0, 37, 0, 0, 0, 0, 0, 25, 147, 0, 0, 0, 
    0, 0, 139, 0, 61, 0, 0, 0, 0, 52, 0, 42, 0, 0, 28, 
    0, 0, 65, 15, 31, 0, 0, 0, 55, 64, 0, 0, 27, 26, 76, 
    0, 10, 0, 64, 0, 0, 0, 0, 148, 0, 19, 0, 0, 101, 11, 
    0, 0, 0, 63, 0, 0, 0, 0, 160, 0, 32, 8, 0, 106, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 65, 0, 23, 52, 0, 25, 0, 
    0, 4, 0, 17, 0, 0, 0, 1, 2, 0, 15, 32, 0, 0, 0, 
    
    -- channel=392
    189, 185, 195, 185, 168, 139, 138, 119, 92, 89, 74, 60, 51, 37, 36, 
    167, 169, 137, 95, 84, 74, 76, 71, 61, 58, 74, 74, 14, 30, 40, 
    111, 75, 58, 47, 46, 50, 52, 64, 64, 68, 135, 117, 70, 88, 66, 
    30, 31, 40, 42, 49, 57, 81, 103, 115, 111, 79, 25, 67, 56, 41, 
    32, 32, 37, 42, 53, 100, 145, 149, 201, 246, 153, 104, 98, 52, 40, 
    33, 36, 43, 44, 55, 159, 336, 385, 371, 335, 430, 208, 52, 113, 34, 
    41, 43, 40, 42, 135, 159, 156, 52, 26, 100, 494, 399, 50, 52, 41, 
    44, 43, 82, 155, 144, 130, 144, 171, 317, 500, 553, 423, 100, 6, 172, 
    38, 53, 109, 123, 128, 55, 140, 512, 570, 559, 530, 197, 94, 225, 366, 
    29, 302, 260, 79, 41, 9, 172, 478, 494, 458, 403, 446, 410, 400, 345, 
    59, 260, 238, 86, 0, 43, 233, 466, 427, 92, 64, 244, 408, 326, 120, 
    18, 89, 220, 88, 17, 149, 313, 502, 342, 61, 56, 71, 287, 207, 8, 
    1, 95, 212, 119, 163, 313, 409, 468, 319, 108, 145, 40, 157, 80, 0, 
    18, 69, 133, 69, 86, 124, 146, 150, 97, 83, 109, 23, 0, 0, 0, 
    56, 48, 63, 77, 29, 38, 34, 14, 0, 21, 66, 0, 0, 0, 0, 
    
    -- channel=393
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 41, 119, 209, 320, 94, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 161, 164, 117, 238, 404, 224, 123, 43, 0, 
    0, 0, 0, 0, 13, 68, 132, 172, 185, 350, 431, 308, 126, 100, 74, 
    0, 0, 0, 161, 187, 166, 236, 378, 380, 394, 338, 83, 34, 184, 251, 
    0, 0, 183, 243, 158, 189, 338, 427, 444, 402, 376, 284, 310, 344, 279, 
    0, 220, 332, 225, 135, 213, 386, 440, 396, 237, 245, 410, 421, 361, 161, 
    0, 214, 345, 194, 178, 324, 433, 446, 282, 195, 177, 261, 389, 253, 83, 
    0, 213, 357, 242, 305, 371, 420, 434, 288, 240, 211, 183, 316, 195, 44, 
    0, 143, 306, 291, 337, 349, 353, 349, 259, 249, 221, 153, 166, 140, 95, 
    0, 74, 218, 225, 223, 223, 203, 179, 142, 186, 206, 126, 115, 113, 119, 
    
    -- channel=394
    362, 386, 398, 412, 399, 375, 363, 347, 327, 255, 264, 245, 164, 152, 209, 
    389, 361, 353, 355, 335, 312, 303, 297, 278, 260, 246, 196, 120, 144, 222, 
    308, 299, 298, 290, 280, 267, 267, 266, 260, 257, 195, 106, 133, 184, 225, 
    253, 258, 257, 257, 262, 262, 256, 252, 252, 248, 125, 118, 187, 236, 241, 
    241, 258, 260, 259, 261, 255, 230, 227, 196, 135, 63, 106, 192, 228, 237, 
    256, 257, 257, 256, 253, 190, 122, 103, 110, 70, 0, 30, 143, 147, 217, 
    260, 256, 253, 245, 205, 138, 88, 89, 107, 104, 0, 0, 85, 118, 164, 
    257, 256, 228, 164, 93, 111, 66, 24, 6, 11, 0, 0, 58, 106, 69, 
    254, 239, 152, 95, 56, 103, 96, 13, 1, 0, 0, 29, 83, 55, 19, 
    254, 138, 5, 67, 71, 110, 98, 0, 0, 15, 43, 0, 0, 0, 30, 
    254, 89, 0, 52, 94, 74, 59, 0, 0, 51, 102, 87, 0, 14, 57, 
    218, 86, 4, 37, 87, 53, 37, 0, 0, 74, 66, 113, 20, 2, 104, 
    184, 78, 12, 26, 39, 0, 0, 0, 0, 63, 27, 92, 72, 45, 120, 
    158, 106, 57, 77, 87, 86, 90, 87, 55, 80, 49, 77, 98, 100, 108, 
    143, 98, 50, 44, 61, 57, 62, 70, 82, 100, 80, 89, 100, 101, 102, 
    
    -- channel=395
    203, 216, 221, 218, 209, 183, 177, 165, 144, 143, 117, 102, 86, 33, 77, 
    195, 181, 186, 162, 152, 136, 133, 125, 111, 106, 90, 82, 34, 21, 89, 
    158, 147, 125, 119, 110, 106, 109, 106, 106, 102, 105, 79, 40, 78, 107, 
    89, 93, 99, 99, 101, 108, 111, 115, 114, 116, 104, 4, 83, 108, 98, 
    90, 98, 101, 105, 105, 118, 133, 128, 99, 100, 43, 35, 97, 89, 87, 
    99, 101, 103, 105, 98, 78, 122, 192, 236, 233, 147, 121, 30, 96, 75, 
    101, 105, 111, 92, 91, 143, 136, 75, 51, 0, 194, 202, 13, 63, 58, 
    103, 107, 81, 96, 89, 52, 86, 0, 0, 107, 234, 295, 76, 0, 19, 
    104, 88, 79, 59, 108, 32, 0, 185, 274, 259, 285, 134, 27, 1, 154, 
    83, 69, 147, 27, 45, 0, 5, 216, 209, 273, 234, 177, 139, 173, 190, 
    56, 216, 144, 53, 2, 0, 0, 202, 264, 105, 50, 114, 222, 188, 160, 
    77, 20, 104, 65, 0, 34, 63, 214, 253, 18, 21, 16, 130, 168, 0, 
    40, 45, 97, 36, 0, 63, 126, 193, 198, 20, 55, 11, 97, 94, 8, 
    39, 53, 109, 70, 93, 147, 163, 168, 137, 36, 79, 27, 29, 0, 0, 
    56, 39, 0, 0, 0, 0, 0, 0, 0, 14, 67, 13, 0, 0, 0, 
    
    -- channel=396
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 16, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 18, 
    0, 0, 13, 23, 28, 33, 28, 26, 36, 1, 0, 8, 31, 36, 22, 
    0, 0, 0, 0, 0, 0, 0, 5, 12, 16, 16, 19, 24, 22, 15, 
    
    -- channel=397
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 44, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 58, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 63, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 78, 159, 235, 248, 172, 0, 90, 6, 0, 
    0, 0, 0, 0, 17, 128, 132, 94, 81, 147, 260, 12, 0, 81, 10, 
    0, 0, 0, 6, 62, 81, 67, 18, 6, 152, 251, 145, 37, 32, 44, 
    0, 0, 17, 111, 86, 100, 141, 263, 289, 282, 213, 0, 16, 45, 162, 
    0, 72, 15, 94, 33, 84, 216, 266, 252, 263, 326, 130, 138, 183, 171, 
    25, 245, 116, 65, 27, 61, 182, 245, 201, 114, 137, 316, 226, 197, 109, 
    5, 74, 138, 32, 43, 136, 248, 242, 79, 63, 35, 174, 209, 75, 29, 
    4, 90, 156, 28, 90, 103, 208, 227, 46, 102, 29, 57, 209, 49, 42, 
    0, 77, 159, 133, 209, 253, 269, 265, 136, 135, 77, 17, 89, 32, 32, 
    13, 27, 38, 12, 36, 38, 33, 28, 22, 99, 95, 32, 21, 24, 38, 
    
    -- channel=398
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 35, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 52, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 125, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 22, 0, 0, 0, 192, 14, 0, 0, 
    0, 0, 0, 0, 14, 0, 17, 0, 0, 0, 0, 133, 73, 0, 0, 
    0, 0, 16, 0, 34, 0, 0, 0, 0, 0, 32, 135, 0, 0, 0, 
    0, 0, 141, 0, 50, 0, 0, 0, 0, 23, 0, 66, 0, 0, 19, 
    0, 0, 104, 8, 26, 0, 0, 0, 58, 82, 0, 0, 29, 25, 86, 
    0, 3, 0, 55, 0, 0, 0, 0, 169, 0, 8, 0, 0, 99, 1, 
    0, 0, 0, 56, 0, 0, 0, 0, 172, 0, 30, 0, 0, 109, 0, 
    0, 0, 0, 22, 0, 0, 0, 0, 86, 0, 18, 36, 0, 21, 0, 
    0, 10, 0, 6, 0, 0, 0, 0, 0, 0, 13, 37, 0, 0, 0, 
    
    -- channel=399
    105, 73, 87, 65, 52, 37, 49, 24, 23, 24, 26, 28, 1, 31, 2, 
    68, 68, 21, 5, 5, 2, 12, 7, 8, 15, 56, 16, 0, 45, 2, 
    27, 0, 0, 0, 0, 5, 5, 20, 23, 34, 133, 56, 43, 73, 18, 
    0, 0, 0, 0, 9, 17, 47, 64, 69, 69, 11, 39, 48, 13, 0, 
    0, 0, 0, 0, 19, 65, 104, 115, 200, 197, 118, 71, 41, 11, 3, 
    0, 0, 0, 2, 43, 188, 324, 287, 259, 254, 475, 0, 64, 56, 0, 
    1, 0, 0, 28, 130, 104, 111, 0, 44, 240, 517, 221, 0, 53, 3, 
    1, 2, 86, 109, 98, 134, 126, 264, 401, 524, 481, 185, 50, 38, 239, 
    0, 60, 55, 129, 55, 73, 212, 560, 473, 488, 404, 20, 158, 278, 345, 
    42, 406, 73, 96, 0, 51, 290, 452, 439, 287, 377, 383, 369, 335, 238, 
    99, 190, 174, 53, 0, 147, 329, 429, 270, 6, 56, 367, 312, 225, 0, 
    40, 104, 253, 1, 72, 209, 413, 434, 114, 93, 44, 121, 321, 45, 20, 
    21, 124, 251, 63, 263, 344, 430, 414, 116, 165, 102, 21, 222, 0, 4, 
    26, 94, 113, 35, 79, 91, 105, 95, 28, 153, 80, 0, 0, 0, 0, 
    53, 54, 89, 79, 48, 61, 47, 27, 7, 51, 50, 0, 0, 0, 28, 
    
    -- channel=400
    202, 178, 182, 163, 149, 127, 131, 105, 105, 106, 76, 81, 57, 38, 48, 
    168, 166, 139, 113, 106, 94, 97, 82, 77, 72, 94, 75, 4, 53, 61, 
    131, 107, 93, 80, 77, 84, 87, 83, 86, 95, 186, 114, 60, 109, 86, 
    63, 73, 83, 81, 87, 103, 126, 135, 135, 145, 72, 44, 109, 86, 60, 
    77, 82, 88, 92, 108, 147, 179, 203, 258, 271, 149, 109, 105, 64, 56, 
    86, 91, 91, 88, 122, 231, 403, 452, 471, 452, 535, 174, 71, 118, 54, 
    93, 99, 91, 98, 201, 243, 239, 94, 72, 230, 675, 423, 36, 78, 48, 
    101, 103, 144, 201, 162, 176, 179, 210, 362, 634, 738, 492, 122, 35, 208, 
    100, 135, 145, 182, 142, 85, 227, 684, 757, 763, 695, 236, 180, 306, 482, 
    124, 420, 255, 135, 35, 37, 326, 657, 679, 608, 596, 564, 525, 525, 444, 
    184, 396, 296, 104, 0, 75, 373, 638, 539, 154, 136, 458, 563, 429, 149, 
    106, 157, 289, 77, 25, 221, 492, 673, 356, 94, 54, 172, 433, 227, 12, 
    58, 164, 297, 134, 229, 404, 571, 640, 331, 168, 156, 64, 262, 81, 0, 
    57, 140, 200, 120, 176, 248, 280, 285, 152, 162, 158, 12, 0, 0, 0, 
    94, 83, 73, 60, 20, 31, 24, 7, 0, 46, 103, 0, 0, 0, 0, 
    
    -- channel=401
    145, 149, 142, 139, 132, 108, 100, 99, 66, 59, 54, 54, 60, 0, 23, 
    120, 129, 103, 77, 67, 59, 53, 57, 45, 45, 40, 62, 16, 0, 29, 
    86, 56, 44, 38, 32, 35, 34, 44, 47, 42, 121, 84, 30, 44, 60, 
    15, 18, 27, 30, 31, 39, 53, 68, 76, 82, 79, 0, 34, 41, 34, 
    17, 21, 26, 32, 33, 79, 99, 84, 92, 152, 112, 41, 63, 36, 29, 
    23, 26, 32, 33, 26, 74, 235, 300, 289, 259, 302, 170, 4, 78, 21, 
    28, 31, 40, 21, 100, 85, 89, 9, 0, 0, 264, 359, 9, 22, 14, 
    29, 34, 50, 109, 91, 70, 93, 48, 121, 272, 341, 366, 114, 0, 76, 
    29, 24, 60, 58, 97, 0, 6, 311, 369, 352, 355, 151, 17, 104, 216, 
    2, 175, 225, 19, 36, 0, 26, 279, 307, 330, 279, 344, 251, 247, 243, 
    17, 158, 220, 54, 0, 0, 40, 281, 327, 64, 0, 91, 286, 235, 106, 
    3, 43, 146, 69, 0, 51, 127, 317, 308, 20, 31, 0, 179, 175, 0, 
    0, 46, 116, 72, 38, 155, 192, 279, 290, 29, 101, 2, 72, 95, 0, 
    0, 43, 92, 63, 33, 68, 88, 94, 116, 17, 64, 18, 0, 0, 0, 
    32, 23, 5, 41, 0, 5, 2, 0, 0, 0, 64, 2, 0, 0, 0, 
    
    -- channel=402
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 74, 56, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 61, 66, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 95, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 103, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 42, 59, 54, 49, 95, 101, 81, 0, 0, 
    0, 0, 0, 0, 0, 25, 40, 63, 67, 98, 96, 32, 132, 69, 7, 
    0, 0, 0, 0, 56, 81, 100, 104, 131, 145, 72, 65, 64, 116, 81, 
    0, 0, 35, 66, 110, 114, 114, 114, 65, 38, 31, 4, 37, 101, 98, 
    0, 4, 89, 113, 110, 135, 125, 78, 61, 74, 52, 45, 95, 83, 73, 
    0, 69, 69, 121, 115, 134, 145, 82, 70, 50, 105, 69, 64, 81, 67, 
    0, 89, 117, 122, 133, 145, 111, 85, 74, 111, 120, 134, 72, 91, 97, 
    2, 97, 121, 111, 140, 124, 119, 67, 72, 120, 111, 124, 113, 87, 107, 
    26, 91, 129, 116, 128, 84, 72, 61, 59, 112, 85, 118, 133, 113, 126, 
    32, 81, 124, 142, 151, 147, 146, 136, 137, 137, 103, 118, 143, 144, 144, 
    
    -- channel=403
    0, 3, 0, 0, 11, 16, 7, 33, 31, 68, 56, 60, 114, 26, 65, 
    6, 26, 39, 46, 53, 56, 46, 53, 52, 58, 40, 102, 108, 8, 72, 
    49, 70, 58, 71, 59, 66, 63, 53, 55, 47, 78, 107, 63, 29, 83, 
    62, 65, 68, 71, 61, 67, 63, 58, 49, 55, 167, 10, 49, 63, 73, 
    69, 73, 74, 78, 63, 62, 52, 62, 40, 118, 142, 31, 65, 70, 63, 
    73, 79, 76, 76, 59, 42, 53, 96, 106, 156, 116, 219, 6, 92, 71, 
    74, 82, 93, 67, 59, 98, 142, 120, 87, 0, 74, 328, 90, 62, 63, 
    77, 87, 57, 94, 122, 49, 128, 44, 12, 14, 146, 319, 167, 52, 23, 
    87, 70, 103, 76, 153, 39, 0, 39, 142, 152, 225, 257, 88, 37, 99, 
    66, 10, 265, 70, 134, 27, 0, 123, 138, 191, 113, 190, 122, 140, 159, 
    14, 138, 226, 118, 86, 15, 0, 134, 243, 180, 42, 0, 196, 171, 210, 
    87, 81, 132, 163, 42, 35, 0, 146, 348, 72, 103, 0, 111, 251, 60, 
    80, 90, 108, 145, 11, 94, 51, 139, 315, 45, 147, 64, 50, 201, 42, 
    80, 92, 113, 108, 63, 99, 105, 119, 202, 36, 145, 119, 63, 78, 49, 
    86, 113, 83, 97, 73, 73, 77, 81, 75, 32, 117, 99, 56, 52, 37, 
    
    -- channel=404
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 4, 20, 0, 0, 0, 34, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 167, 127, 0, 32, 10, 0, 
    0, 0, 0, 0, 0, 26, 0, 22, 85, 188, 23, 0, 0, 49, 47, 
    0, 0, 0, 24, 0, 61, 128, 149, 23, 0, 0, 0, 14, 103, 55, 
    0, 81, 0, 76, 0, 100, 229, 64, 19, 0, 0, 0, 67, 19, 0, 
    47, 49, 0, 23, 0, 109, 255, 38, 0, 0, 115, 163, 0, 0, 0, 
    0, 44, 29, 0, 67, 157, 190, 26, 0, 47, 8, 209, 38, 0, 0, 
    9, 57, 67, 0, 141, 75, 156, 14, 0, 90, 0, 74, 124, 0, 40, 
    1, 55, 59, 24, 120, 63, 48, 28, 0, 116, 0, 0, 73, 0, 49, 
    0, 5, 31, 34, 58, 57, 49, 39, 30, 115, 13, 0, 42, 44, 57, 
    
    -- channel=405
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 17, 29, 1, 3, 
    0, 0, 0, 0, 0, 0, 4, 47, 14, 0, 0, 0, 42, 31, 23, 
    0, 0, 0, 0, 1, 8, 0, 0, 0, 0, 0, 0, 2, 9, 0, 
    0, 0, 14, 10, 30, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 22, 44, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 25, 46, 0, 0, 0, 0, 30, 31, 0, 0, 0, 39, 
    0, 7, 0, 34, 23, 0, 0, 0, 0, 12, 28, 23, 0, 23, 28, 
    11, 0, 0, 7, 0, 0, 0, 0, 0, 7, 5, 36, 12, 46, 42, 
    5, 22, 36, 49, 48, 48, 45, 44, 45, 4, 16, 46, 50, 48, 43, 
    
    -- channel=406
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 30, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 7, 2, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 43, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 10, 31, 25, 27, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 17, 15, 49, 49, 0, 0, 7, 15, 
    0, 40, 12, 0, 0, 0, 0, 17, 35, 9, 0, 31, 31, 22, 27, 
    0, 0, 1, 0, 0, 0, 0, 19, 24, 0, 0, 0, 8, 19, 0, 
    0, 0, 4, 0, 0, 0, 0, 11, 9, 0, 0, 0, 14, 9, 0, 
    0, 0, 22, 19, 30, 43, 49, 49, 33, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    
    -- channel=407
    504, 514, 531, 537, 516, 477, 460, 436, 390, 318, 324, 265, 159, 155, 253, 
    491, 464, 454, 443, 414, 383, 376, 361, 336, 323, 274, 210, 127, 167, 272, 
    376, 362, 358, 353, 339, 329, 330, 329, 321, 306, 197, 109, 151, 231, 282, 
    305, 314, 316, 317, 326, 327, 324, 321, 315, 280, 129, 101, 245, 287, 294, 
    299, 318, 320, 321, 320, 314, 285, 272, 221, 168, 68, 98, 228, 279, 281, 
    316, 318, 317, 316, 285, 197, 139, 139, 134, 82, 43, 64, 95, 204, 255, 
    320, 318, 316, 280, 216, 126, 71, 50, 77, 0, 0, 56, 46, 93, 180, 
    317, 313, 237, 175, 98, 93, 60, 6, 0, 4, 0, 50, 103, 54, 73, 
    314, 254, 124, 52, 57, 48, 0, 30, 22, 6, 31, 60, 64, 33, 32, 
    265, 142, 44, 26, 55, 55, 0, 0, 0, 32, 34, 34, 4, 4, 55, 
    225, 58, 38, 43, 61, 18, 0, 0, 40, 27, 33, 4, 4, 32, 67, 
    204, 44, 14, 35, 38, 8, 0, 0, 32, 47, 46, 19, 10, 34, 85, 
    163, 43, 0, 1, 0, 0, 0, 0, 28, 20, 35, 49, 39, 51, 94, 
    158, 81, 43, 47, 35, 38, 43, 44, 59, 44, 30, 54, 54, 67, 74, 
    147, 73, 5, 22, 20, 21, 31, 41, 53, 46, 71, 69, 69, 68, 65, 
    
    -- channel=408
    60, 84, 87, 95, 94, 77, 69, 69, 54, 83, 50, 35, 69, 8, 11, 
    78, 77, 69, 50, 41, 36, 32, 36, 27, 23, 19, 63, 27, 0, 12, 
    64, 56, 30, 20, 15, 13, 14, 20, 19, 13, 67, 61, 18, 8, 31, 
    8, 1, 6, 8, 5, 10, 13, 31, 31, 43, 112, 14, 27, 40, 20, 
    0, 0, 5, 9, 4, 25, 53, 53, 61, 116, 80, 27, 39, 19, 13, 
    0, 2, 9, 11, 5, 25, 76, 119, 173, 171, 125, 189, 18, 42, 14, 
    4, 6, 16, 0, 38, 115, 178, 144, 85, 0, 194, 254, 60, 38, 13, 
    6, 12, 0, 53, 96, 46, 86, 17, 22, 127, 266, 313, 77, 0, 10, 
    7, 0, 96, 73, 117, 57, 7, 154, 285, 290, 334, 215, 4, 19, 130, 
    0, 26, 194, 45, 76, 3, 6, 235, 252, 304, 196, 166, 137, 192, 226, 
    0, 177, 187, 78, 27, 0, 34, 232, 324, 169, 123, 108, 251, 233, 185, 
    12, 65, 108, 93, 0, 44, 84, 244, 297, 37, 48, 29, 148, 207, 14, 
    0, 51, 101, 85, 5, 94, 163, 250, 266, 16, 85, 47, 93, 132, 2, 
    1, 41, 108, 87, 107, 171, 194, 205, 155, 38, 103, 60, 42, 24, 0, 
    14, 44, 36, 35, 9, 12, 19, 18, 15, 17, 69, 34, 0, 0, 0, 
    
    -- channel=409
    539, 518, 531, 517, 497, 472, 464, 427, 410, 321, 306, 290, 146, 154, 268, 
    526, 499, 492, 498, 476, 440, 430, 396, 377, 349, 332, 213, 75, 202, 319, 
    413, 410, 432, 429, 407, 406, 404, 379, 370, 367, 274, 113, 153, 283, 320, 
    369, 399, 404, 400, 409, 420, 429, 403, 380, 339, 76, 80, 270, 314, 324, 
    393, 419, 421, 417, 428, 413, 364, 379, 371, 291, 103, 140, 283, 318, 321, 
    417, 427, 415, 404, 402, 368, 351, 301, 239, 176, 224, 8, 110, 247, 302, 
    426, 428, 405, 384, 343, 176, 59, 0, 28, 136, 257, 98, 16, 113, 213, 
    427, 418, 380, 295, 128, 144, 85, 122, 225, 286, 215, 87, 72, 69, 203, 
    427, 394, 171, 101, 21, 17, 116, 300, 226, 219, 175, 50, 229, 236, 231, 
    423, 426, 55, 64, 0, 42, 161, 194, 186, 130, 193, 244, 240, 171, 121, 
    394, 156, 35, 24, 0, 68, 162, 173, 80, 0, 0, 170, 127, 75, 0, 
    291, 76, 97, 0, 39, 95, 187, 185, 0, 53, 26, 76, 135, 0, 48, 
    230, 100, 97, 12, 118, 152, 192, 159, 6, 101, 62, 30, 90, 0, 58, 
    206, 130, 41, 0, 1, 0, 0, 0, 0, 81, 41, 0, 0, 0, 30, 
    208, 98, 23, 23, 10, 15, 11, 12, 5, 42, 45, 0, 0, 3, 18, 
    
    -- channel=410
    87, 74, 99, 86, 73, 75, 89, 54, 84, 59, 36, 60, 8, 49, 29, 
    98, 70, 73, 84, 83, 73, 82, 62, 66, 47, 82, 0, 0, 81, 45, 
    78, 66, 78, 69, 74, 67, 69, 60, 59, 71, 82, 0, 0, 72, 34, 
    68, 72, 71, 63, 72, 74, 75, 65, 56, 61, 0, 46, 42, 54, 41, 
    73, 74, 73, 68, 86, 80, 80, 78, 83, 0, 0, 44, 48, 44, 55, 
    75, 72, 69, 66, 102, 109, 91, 28, 47, 0, 0, 0, 94, 1, 49, 
    75, 70, 58, 89, 101, 59, 0, 0, 20, 183, 155, 0, 0, 77, 38, 
    73, 67, 102, 44, 0, 43, 0, 9, 66, 119, 6, 0, 0, 42, 76, 
    70, 99, 26, 42, 0, 51, 127, 158, 19, 0, 0, 0, 81, 64, 70, 
    114, 170, 0, 41, 0, 68, 208, 69, 3, 0, 60, 0, 22, 0, 0, 
    170, 101, 0, 0, 0, 78, 202, 25, 0, 0, 78, 239, 0, 0, 0, 
    102, 0, 20, 0, 32, 114, 170, 0, 0, 17, 0, 179, 36, 0, 0, 
    72, 41, 60, 0, 100, 23, 123, 0, 0, 76, 0, 10, 137, 0, 44, 
    49, 53, 30, 0, 83, 64, 54, 35, 0, 97, 0, 0, 57, 0, 29, 
    43, 2, 0, 0, 0, 0, 0, 0, 0, 98, 0, 0, 5, 9, 26, 
    
    -- channel=411
    591, 587, 606, 595, 569, 518, 504, 466, 417, 329, 322, 276, 139, 123, 237, 
    575, 544, 518, 492, 463, 421, 410, 384, 355, 330, 311, 210, 64, 131, 276, 
    423, 397, 392, 387, 365, 359, 360, 352, 343, 341, 265, 151, 147, 247, 301, 
    313, 334, 344, 344, 357, 371, 390, 384, 376, 336, 115, 33, 234, 286, 295, 
    323, 348, 354, 356, 369, 385, 374, 387, 386, 326, 125, 111, 271, 291, 282, 
    347, 357, 354, 350, 347, 346, 387, 406, 365, 322, 366, 85, 74, 251, 254, 
    360, 361, 348, 328, 307, 210, 104, 0, 13, 68, 348, 286, 0, 78, 178, 
    360, 358, 332, 286, 161, 143, 126, 125, 227, 352, 376, 272, 107, 17, 177, 
    355, 335, 156, 101, 67, 5, 84, 405, 414, 403, 367, 123, 164, 200, 298, 
    346, 414, 166, 30, 0, 0, 121, 321, 322, 279, 331, 385, 316, 272, 223, 
    302, 231, 142, 21, 0, 20, 114, 302, 239, 10, 0, 175, 261, 180, 57, 
    232, 51, 137, 14, 0, 71, 201, 328, 186, 28, 8, 15, 196, 88, 12, 
    164, 77, 125, 29, 88, 188, 246, 286, 159, 74, 77, 0, 97, 12, 8, 
    149, 93, 61, 4, 2, 28, 45, 49, 46, 53, 53, 0, 0, 0, 0, 
    168, 75, 0, 2, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 0, 
    
    -- channel=412
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 46, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 125, 45, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 17, 60, 132, 164, 66, 18, 0, 0, 
    0, 0, 0, 0, 0, 51, 201, 262, 241, 291, 397, 198, 22, 66, 0, 
    0, 0, 0, 0, 29, 86, 121, 55, 44, 50, 327, 454, 54, 54, 7, 
    0, 0, 0, 78, 125, 96, 164, 192, 240, 313, 408, 392, 175, 44, 144, 
    0, 0, 47, 110, 154, 57, 85, 348, 402, 410, 407, 217, 104, 172, 277, 
    0, 164, 288, 95, 100, 28, 101, 350, 374, 326, 323, 434, 325, 318, 260, 
    0, 178, 305, 122, 55, 85, 120, 360, 345, 153, 13, 145, 353, 271, 165, 
    0, 99, 242, 151, 69, 127, 213, 387, 388, 96, 100, 7, 262, 247, 48, 
    0, 114, 218, 183, 156, 285, 273, 355, 365, 122, 184, 49, 121, 167, 11, 
    5, 77, 138, 112, 71, 95, 109, 115, 182, 87, 149, 79, 13, 40, 22, 
    43, 85, 114, 129, 93, 100, 88, 74, 56, 22, 113, 69, 30, 31, 38, 
    
    -- channel=413
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 34, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 162, 99, 39, 64, 0, 
    0, 0, 0, 0, 0, 0, 14, 21, 34, 57, 44, 52, 38, 0, 0, 
    0, 0, 0, 0, 0, 46, 110, 123, 189, 204, 130, 105, 37, 0, 0, 
    0, 0, 0, 0, 25, 191, 434, 505, 537, 519, 643, 66, 88, 68, 0, 
    0, 0, 0, 1, 166, 257, 232, 54, 64, 316, 839, 333, 13, 93, 1, 
    0, 0, 75, 162, 155, 197, 201, 249, 444, 779, 829, 463, 81, 51, 251, 
    0, 46, 104, 212, 153, 117, 307, 863, 853, 839, 723, 93, 199, 361, 577, 
    22, 481, 202, 180, 5, 85, 461, 777, 754, 650, 697, 581, 614, 590, 462, 
    148, 490, 280, 121, 0, 149, 514, 735, 557, 94, 163, 612, 608, 454, 103, 
    75, 160, 378, 57, 66, 336, 636, 761, 297, 124, 63, 273, 512, 191, 0, 
    38, 207, 401, 111, 335, 497, 703, 704, 252, 246, 159, 74, 381, 16, 0, 
    38, 175, 267, 139, 255, 302, 326, 319, 123, 241, 164, 0, 40, 0, 0, 
    79, 81, 98, 83, 58, 71, 57, 29, 0, 114, 124, 0, 0, 0, 9, 
    
    -- channel=414
    36, 96, 65, 93, 131, 110, 72, 132, 54, 115, 90, 53, 135, 0, 60, 
    83, 111, 129, 115, 106, 100, 71, 97, 71, 74, 7, 127, 122, 0, 66, 
    83, 120, 85, 101, 66, 68, 66, 61, 58, 27, 0, 138, 35, 0, 104, 
    53, 47, 55, 68, 45, 56, 43, 54, 43, 23, 260, 0, 0, 62, 89, 
    39, 53, 57, 69, 29, 29, 18, 24, 0, 125, 169, 0, 60, 76, 55, 
    48, 61, 68, 70, 0, 0, 0, 0, 0, 88, 0, 435, 0, 103, 58, 
    55, 67, 97, 20, 0, 0, 108, 124, 24, 0, 0, 667, 59, 0, 34, 
    55, 80, 0, 24, 107, 0, 98, 0, 0, 0, 0, 547, 245, 0, 0, 
    69, 0, 53, 0, 184, 0, 0, 0, 0, 0, 206, 504, 0, 0, 0, 
    0, 0, 479, 0, 185, 0, 0, 0, 0, 108, 0, 170, 0, 0, 102, 
    0, 0, 341, 75, 70, 0, 0, 0, 283, 269, 0, 0, 117, 121, 368, 
    0, 0, 13, 238, 0, 0, 0, 0, 695, 0, 63, 0, 0, 434, 4, 
    0, 0, 0, 173, 0, 0, 0, 0, 622, 0, 146, 0, 0, 372, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 317, 0, 130, 143, 0, 59, 0, 
    4, 52, 0, 44, 0, 0, 0, 10, 20, 0, 66, 117, 0, 0, 0, 
    
    -- channel=415
    61, 61, 71, 67, 64, 65, 68, 62, 59, 51, 52, 47, 40, 57, 58, 
    62, 53, 66, 66, 66, 64, 68, 62, 62, 59, 48, 35, 33, 57, 56, 
    59, 58, 63, 65, 64, 59, 62, 59, 58, 55, 15, 28, 40, 53, 52, 
    60, 61, 59, 59, 60, 56, 49, 46, 46, 38, 18, 39, 42, 51, 57, 
    61, 60, 57, 56, 56, 47, 40, 29, 0, 0, 0, 42, 51, 59, 58, 
    57, 57, 57, 58, 49, 9, 0, 0, 0, 0, 0, 0, 48, 39, 56, 
    57, 55, 54, 53, 21, 9, 0, 2, 16, 0, 0, 0, 30, 48, 61, 
    55, 53, 38, 14, 4, 11, 0, 0, 0, 0, 0, 0, 0, 37, 4, 
    54, 40, 9, 3, 12, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 12, 22, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 14, 35, 18, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    37, 0, 0, 14, 30, 2, 0, 0, 0, 15, 20, 20, 0, 0, 34, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 23, 0, 0, 57, 
    39, 13, 6, 8, 13, 0, 0, 0, 0, 10, 0, 31, 50, 38, 56, 
    35, 15, 10, 14, 32, 28, 30, 33, 42, 42, 20, 38, 55, 55, 50, 
    
    -- channel=416
    466, 498, 512, 528, 515, 480, 458, 442, 403, 335, 321, 271, 152, 122, 237, 
    510, 477, 476, 475, 448, 411, 392, 377, 349, 320, 277, 218, 102, 102, 271, 
    386, 399, 391, 388, 364, 348, 348, 335, 321, 314, 170, 96, 122, 177, 275, 
    321, 333, 335, 337, 340, 346, 339, 328, 315, 283, 136, 48, 197, 279, 299, 
    312, 342, 346, 345, 342, 319, 274, 291, 251, 198, 60, 42, 223, 285, 282, 
    336, 347, 342, 339, 313, 226, 96, 77, 74, 61, 0, 69, 67, 179, 260, 
    348, 348, 341, 307, 208, 132, 72, 65, 57, 0, 0, 32, 24, 58, 173, 
    346, 345, 270, 189, 109, 55, 41, 0, 0, 0, 0, 45, 47, 28, 2, 
    344, 298, 149, 48, 23, 6, 0, 0, 0, 0, 8, 131, 78, 0, 0, 
    323, 108, 62, 0, 33, 2, 0, 0, 0, 3, 4, 0, 0, 0, 18, 
    259, 69, 0, 0, 26, 0, 0, 0, 0, 63, 7, 0, 0, 0, 76, 
    235, 22, 0, 17, 0, 0, 0, 0, 41, 0, 12, 0, 0, 29, 39, 
    186, 14, 0, 0, 0, 0, 0, 0, 29, 0, 3, 10, 0, 47, 42, 
    153, 47, 0, 0, 0, 10, 16, 27, 46, 0, 21, 24, 14, 23, 22, 
    135, 67, 0, 0, 0, 0, 0, 0, 7, 7, 11, 31, 10, 8, 4, 
    
    -- channel=417
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=418
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 20, 0, 6, 0, 42, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 1, 0, 0, 5, 2, 85, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 22, 57, 5, 0, 0, 0, 32, 
    0, 0, 0, 0, 0, 2, 0, 96, 12, 0, 8, 0, 22, 3, 37, 
    0, 58, 0, 3, 0, 3, 21, 45, 0, 0, 4, 0, 14, 0, 0, 
    0, 30, 0, 0, 0, 21, 29, 20, 8, 0, 6, 68, 0, 0, 0, 
    18, 0, 53, 0, 0, 52, 35, 1, 0, 7, 0, 19, 23, 0, 0, 
    0, 8, 55, 0, 29, 23, 52, 0, 0, 20, 0, 0, 71, 0, 6, 
    0, 15, 25, 0, 20, 9, 3, 0, 0, 40, 0, 0, 23, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 20, 1, 0, 0, 0, 2, 
    
    -- channel=419
    827, 826, 862, 855, 822, 761, 743, 689, 628, 505, 499, 428, 210, 209, 392, 
    817, 766, 744, 731, 690, 633, 623, 587, 549, 515, 469, 324, 138, 252, 443, 
    595, 586, 595, 591, 567, 551, 557, 545, 528, 514, 332, 127, 224, 376, 447, 
    504, 528, 532, 533, 549, 558, 567, 558, 538, 471, 145, 103, 362, 451, 469, 
    506, 541, 543, 543, 551, 543, 481, 491, 468, 383, 111, 134, 383, 451, 451, 
    536, 544, 539, 535, 505, 436, 324, 233, 165, 82, 124, 14, 127, 324, 410, 
    548, 544, 531, 489, 397, 176, 64, 0, 64, 61, 121, 37, 16, 126, 277, 
    541, 535, 454, 332, 167, 137, 75, 100, 185, 145, 51, 0, 55, 63, 191, 
    535, 475, 207, 81, 13, 24, 45, 157, 67, 61, 57, 28, 204, 157, 126, 
    499, 414, 11, 22, 0, 37, 22, 58, 20, 0, 32, 89, 103, 48, 52, 
    435, 76, 0, 9, 9, 51, 33, 23, 0, 0, 0, 39, 0, 0, 0, 
    358, 29, 42, 0, 36, 34, 37, 18, 0, 36, 32, 21, 27, 0, 68, 
    280, 58, 26, 0, 48, 44, 54, 8, 0, 48, 39, 17, 51, 0, 96, 
    254, 105, 0, 0, 0, 0, 0, 0, 0, 45, 7, 6, 23, 9, 62, 
    238, 101, 13, 17, 0, 6, 14, 21, 33, 51, 17, 11, 43, 44, 53, 
    
    -- channel=420
    93, 96, 98, 104, 103, 101, 97, 98, 90, 72, 80, 79, 55, 56, 81, 
    90, 94, 96, 101, 97, 94, 92, 92, 88, 86, 68, 66, 64, 58, 79, 
    85, 84, 90, 91, 90, 87, 88, 86, 85, 81, 51, 36, 49, 65, 79, 
    85, 88, 86, 88, 87, 84, 71, 71, 74, 72, 43, 41, 67, 75, 84, 
    84, 87, 86, 86, 82, 79, 56, 39, 4, 9, 22, 37, 55, 77, 83, 
    86, 86, 86, 85, 68, 27, 10, 7, 0, 0, 0, 20, 50, 49, 77, 
    85, 85, 86, 74, 57, 7, 0, 20, 27, 0, 0, 0, 45, 42, 62, 
    84, 83, 60, 39, 21, 24, 0, 0, 0, 0, 0, 0, 35, 38, 5, 
    85, 60, 35, 20, 18, 24, 2, 0, 0, 0, 0, 0, 3, 0, 0, 
    66, 0, 0, 18, 44, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 0, 0, 26, 56, 16, 0, 0, 0, 0, 12, 0, 0, 0, 8, 
    63, 19, 0, 30, 39, 0, 0, 0, 0, 22, 41, 11, 0, 0, 55, 
    66, 18, 0, 9, 0, 0, 0, 0, 0, 6, 14, 40, 0, 32, 58, 
    62, 35, 13, 33, 12, 0, 0, 0, 18, 5, 6, 51, 41, 60, 59, 
    52, 29, 17, 33, 38, 33, 37, 42, 51, 44, 34, 55, 63, 61, 55, 
    
    -- channel=421
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 32, 99, 146, 206, 164, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 67, 8, 0, 0, 219, 159, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 10, 0, 0, 64, 245, 263, 8, 0, 0, 
    0, 0, 0, 23, 36, 0, 0, 191, 256, 277, 254, 67, 0, 0, 125, 
    0, 0, 63, 0, 0, 0, 0, 234, 236, 251, 271, 168, 111, 159, 146, 
    0, 166, 150, 0, 0, 0, 0, 221, 236, 65, 0, 168, 225, 177, 81, 
    0, 0, 121, 0, 0, 11, 95, 229, 210, 0, 0, 0, 158, 109, 0, 
    0, 2, 107, 0, 0, 69, 122, 209, 160, 0, 4, 0, 87, 34, 0, 
    0, 0, 74, 26, 51, 123, 142, 150, 125, 0, 39, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    
    -- channel=422
    457, 456, 494, 482, 461, 412, 409, 360, 329, 317, 258, 212, 101, 101, 171, 
    458, 424, 408, 382, 357, 319, 319, 289, 266, 242, 228, 156, 36, 99, 196, 
    337, 326, 301, 287, 272, 263, 270, 261, 253, 249, 213, 99, 92, 189, 216, 
    234, 243, 249, 248, 260, 274, 284, 287, 280, 256, 110, 50, 194, 230, 219, 
    234, 251, 257, 260, 273, 292, 293, 312, 304, 262, 71, 68, 201, 212, 201, 
    250, 257, 256, 256, 257, 281, 311, 328, 370, 355, 298, 58, 95, 181, 183, 
    260, 263, 256, 239, 247, 244, 215, 95, 86, 125, 468, 187, 0, 104, 129, 
    264, 262, 238, 212, 167, 127, 112, 67, 170, 320, 462, 329, 40, 4, 124, 
    260, 245, 146, 146, 94, 54, 127, 437, 495, 508, 452, 151, 149, 137, 317, 
    248, 333, 108, 65, 0, 10, 151, 442, 417, 409, 429, 282, 285, 317, 296, 
    258, 355, 146, 38, 0, 1, 177, 396, 352, 100, 103, 351, 339, 283, 130, 
    198, 56, 181, 17, 0, 114, 277, 403, 223, 26, 15, 118, 269, 133, 0, 
    128, 95, 186, 6, 79, 187, 334, 384, 163, 84, 56, 5, 214, 20, 7, 
    107, 104, 141, 46, 130, 215, 238, 244, 116, 93, 95, 0, 28, 0, 0, 
    124, 53, 7, 0, 0, 0, 0, 0, 0, 54, 49, 0, 0, 0, 0, 
    
    -- channel=423
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 26, 78, 13, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=424
    125, 127, 121, 122, 113, 102, 95, 90, 78, 31, 45, 45, 21, 0, 23, 
    122, 113, 101, 96, 87, 76, 71, 68, 58, 53, 57, 41, 0, 0, 41, 
    70, 58, 63, 67, 59, 58, 58, 57, 57, 55, 62, 0, 3, 24, 42, 
    41, 51, 54, 56, 58, 61, 74, 71, 68, 68, 0, 0, 4, 36, 41, 
    46, 56, 58, 59, 60, 74, 61, 67, 81, 89, 17, 0, 44, 42, 41, 
    56, 59, 58, 58, 59, 71, 84, 74, 34, 0, 37, 18, 0, 29, 31, 
    60, 59, 59, 50, 68, 0, 0, 0, 0, 0, 16, 24, 0, 0, 3, 
    58, 60, 66, 69, 8, 0, 0, 5, 57, 87, 22, 0, 0, 0, 16, 
    57, 60, 31, 0, 0, 0, 0, 50, 31, 10, 9, 0, 8, 51, 23, 
    57, 112, 22, 0, 0, 0, 0, 2, 3, 0, 0, 55, 53, 11, 0, 
    69, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=425
    345, 317, 332, 310, 288, 247, 246, 208, 184, 123, 122, 119, 45, 0, 66, 
    298, 292, 240, 210, 191, 166, 167, 150, 135, 124, 148, 90, 0, 35, 88, 
    194, 144, 139, 132, 128, 131, 134, 139, 141, 149, 234, 66, 47, 133, 123, 
    93, 108, 120, 121, 135, 151, 181, 201, 200, 202, 25, 0, 98, 104, 90, 
    107, 118, 123, 130, 150, 212, 232, 243, 308, 320, 121, 77, 127, 100, 88, 
    120, 127, 129, 126, 159, 281, 467, 477, 433, 344, 553, 67, 15, 131, 72, 
    132, 131, 129, 135, 247, 161, 95, 0, 0, 138, 589, 338, 0, 16, 32, 
    132, 138, 189, 229, 124, 136, 116, 202, 405, 653, 602, 308, 55, 0, 229, 
    129, 170, 107, 96, 41, 0, 139, 679, 628, 603, 531, 33, 146, 311, 428, 
    156, 531, 165, 44, 0, 0, 248, 529, 523, 415, 436, 521, 487, 414, 317, 
    214, 248, 176, 19, 0, 57, 298, 499, 375, 0, 0, 297, 391, 273, 0, 
    110, 67, 226, 0, 0, 170, 402, 534, 188, 31, 0, 61, 315, 64, 0, 
    47, 94, 219, 25, 205, 352, 476, 478, 178, 111, 96, 0, 171, 0, 0, 
    44, 79, 88, 0, 23, 33, 54, 48, 0, 95, 31, 0, 0, 0, 0, 
    81, 36, 5, 25, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    
    -- channel=426
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=427
    13, 101, 151, 181, 186, 175, 171, 151, 167, 211, 128, 82, 112, 107, 54, 
    151, 108, 161, 183, 176, 152, 144, 126, 109, 83, 15, 49, 36, 0, 43, 
    212, 231, 172, 146, 123, 93, 91, 71, 61, 41, 42, 33, 0, 0, 56, 
    111, 91, 81, 74, 69, 67, 22, 0, 1, 33, 137, 78, 49, 100, 95, 
    72, 85, 91, 90, 80, 53, 45, 6, 0, 0, 0, 0, 18, 72, 77, 
    80, 82, 82, 90, 60, 0, 0, 0, 233, 284, 0, 0, 142, 0, 70, 
    80, 87, 99, 65, 28, 251, 298, 322, 216, 0, 0, 0, 0, 157, 77, 
    93, 87, 0, 0, 22, 0, 0, 0, 0, 0, 0, 178, 0, 0, 0, 
    101, 25, 59, 128, 111, 112, 0, 0, 30, 38, 21, 42, 0, 0, 0, 
    34, 0, 0, 36, 67, 77, 0, 19, 0, 302, 307, 0, 0, 0, 111, 
    124, 428, 34, 19, 38, 0, 0, 0, 185, 289, 290, 377, 113, 185, 323, 
    157, 9, 0, 0, 0, 0, 0, 0, 43, 0, 0, 186, 64, 111, 13, 
    106, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 234, 140, 58, 
    36, 90, 220, 241, 393, 581, 624, 639, 372, 63, 87, 38, 197, 83, 15, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 124, 139, 48, 0, 0, 0, 
    
    -- channel=428
    336, 351, 333, 345, 336, 317, 292, 298, 255, 209, 205, 180, 107, 78, 176, 
    334, 327, 332, 323, 299, 280, 263, 257, 238, 224, 188, 152, 86, 94, 203, 
    254, 267, 271, 269, 249, 249, 246, 232, 228, 222, 89, 99, 111, 142, 207, 
    225, 240, 244, 247, 245, 251, 245, 239, 226, 198, 88, 33, 161, 202, 210, 
    232, 251, 254, 251, 246, 219, 188, 202, 190, 180, 105, 89, 176, 203, 201, 
    250, 256, 254, 245, 215, 142, 79, 82, 33, 6, 0, 239, 15, 164, 191, 
    253, 259, 250, 215, 122, 54, 14, 43, 2, 0, 0, 221, 87, 13, 134, 
    256, 256, 180, 155, 78, 42, 45, 26, 17, 0, 4, 126, 123, 26, 25, 
    257, 200, 108, 0, 37, 0, 0, 0, 1, 3, 57, 239, 58, 39, 3, 
    223, 32, 189, 0, 80, 0, 0, 0, 0, 25, 0, 125, 31, 22, 46, 
    124, 0, 64, 27, 52, 0, 0, 0, 35, 85, 0, 0, 25, 20, 92, 
    105, 39, 0, 84, 0, 0, 0, 0, 155, 3, 33, 0, 0, 106, 53, 
    91, 0, 0, 93, 0, 0, 0, 0, 173, 0, 72, 31, 0, 122, 23, 
    100, 5, 0, 6, 0, 0, 0, 0, 38, 0, 30, 59, 0, 33, 15, 
    98, 58, 11, 29, 6, 3, 12, 19, 21, 0, 15, 53, 12, 11, 0, 
    
    -- channel=429
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=430
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 56, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 35, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 4, 24, 0, 0, 19, 0, 0, 0, 
    0, 0, 0, 0, 19, 53, 56, 5, 9, 0, 34, 0, 40, 0, 0, 
    0, 0, 0, 7, 34, 7, 0, 0, 0, 182, 148, 0, 0, 15, 0, 
    0, 0, 25, 0, 0, 22, 0, 47, 113, 174, 18, 0, 0, 34, 74, 
    0, 23, 0, 2, 0, 28, 125, 179, 19, 0, 0, 0, 56, 84, 70, 
    34, 150, 0, 29, 0, 56, 219, 62, 3, 0, 27, 0, 38, 0, 0, 
    106, 35, 0, 0, 0, 91, 224, 27, 0, 0, 40, 190, 0, 0, 0, 
    38, 0, 13, 0, 33, 115, 189, 7, 0, 12, 0, 162, 30, 0, 0, 
    20, 28, 50, 0, 122, 57, 138, 0, 0, 75, 0, 1, 108, 0, 18, 
    11, 31, 8, 0, 53, 7, 0, 0, 0, 92, 0, 0, 27, 0, 13, 
    2, 0, 0, 0, 0, 2, 0, 0, 0, 71, 0, 0, 0, 1, 21, 
    
    -- channel=431
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    
    -- channel=432
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 10, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 25, 69, 35, 27, 42, 4, 0, 0, 
    0, 0, 0, 0, 0, 82, 126, 106, 103, 129, 203, 0, 72, 13, 0, 
    0, 0, 0, 0, 33, 51, 53, 20, 36, 197, 265, 20, 0, 53, 10, 
    0, 0, 29, 25, 46, 71, 50, 142, 197, 216, 231, 34, 4, 36, 128, 
    0, 11, 2, 90, 15, 58, 173, 259, 213, 238, 153, 0, 102, 136, 168, 
    7, 178, 0, 72, 0, 48, 205, 229, 222, 120, 223, 159, 163, 162, 95, 
    48, 111, 62, 23, 0, 100, 216, 214, 79, 34, 54, 256, 145, 103, 0, 
    0, 61, 126, 0, 52, 121, 257, 209, 0, 53, 26, 117, 178, 0, 23, 
    7, 72, 140, 35, 158, 174, 222, 207, 0, 112, 37, 17, 137, 0, 17, 
    7, 46, 63, 32, 72, 88, 91, 87, 25, 99, 49, 0, 23, 2, 12, 
    20, 21, 64, 31, 35, 41, 30, 22, 11, 61, 23, 0, 1, 4, 24, 
    
    -- channel=433
    377, 346, 341, 330, 312, 283, 277, 265, 224, 168, 201, 186, 84, 89, 173, 
    306, 298, 267, 247, 234, 221, 221, 218, 207, 213, 204, 143, 100, 134, 186, 
    195, 176, 195, 199, 203, 203, 207, 219, 219, 220, 151, 94, 150, 193, 192, 
    179, 194, 198, 203, 210, 214, 229, 241, 239, 207, 63, 61, 170, 178, 187, 
    188, 196, 195, 199, 204, 218, 202, 209, 246, 216, 140, 118, 158, 180, 179, 
    197, 197, 197, 197, 194, 216, 225, 160, 57, 41, 221, 70, 58, 145, 159, 
    200, 195, 191, 189, 161, 23, 0, 0, 4, 66, 89, 164, 51, 45, 107, 
    192, 194, 201, 153, 74, 101, 99, 206, 286, 217, 73, 20, 91, 86, 184, 
    185, 194, 69, 35, 31, 26, 74, 162, 57, 52, 43, 33, 138, 183, 125, 
    204, 254, 78, 31, 32, 42, 53, 42, 41, 0, 13, 189, 142, 70, 20, 
    138, 0, 45, 35, 52, 112, 64, 51, 0, 0, 0, 0, 5, 0, 0, 
    114, 43, 76, 45, 93, 55, 64, 64, 33, 68, 65, 0, 37, 1, 81, 
    99, 53, 54, 72, 132, 143, 77, 43, 56, 83, 92, 25, 0, 6, 65, 
    111, 62, 0, 0, 0, 0, 0, 0, 0, 36, 26, 44, 0, 43, 67, 
    117, 79, 75, 99, 76, 80, 76, 69, 71, 16, 25, 53, 77, 79, 86, 
    
    -- channel=434
    3, 46, 23, 51, 67, 58, 34, 67, 35, 90, 53, 29, 65, 0, 27, 
    31, 39, 61, 56, 49, 48, 28, 45, 32, 32, 0, 57, 76, 0, 22, 
    49, 77, 47, 49, 32, 28, 26, 22, 20, 5, 0, 72, 6, 0, 42, 
    25, 22, 25, 30, 14, 18, 0, 0, 0, 0, 152, 0, 6, 43, 45, 
    12, 24, 28, 32, 7, 0, 0, 0, 0, 0, 36, 0, 0, 23, 23, 
    21, 27, 29, 30, 0, 0, 0, 0, 2, 104, 0, 221, 0, 0, 24, 
    24, 31, 42, 0, 0, 42, 113, 165, 56, 0, 0, 242, 50, 0, 5, 
    27, 36, 0, 0, 35, 0, 40, 0, 0, 0, 0, 315, 119, 0, 0, 
    33, 0, 30, 0, 113, 0, 0, 0, 0, 0, 89, 329, 0, 0, 0, 
    0, 0, 218, 0, 136, 0, 0, 0, 0, 133, 31, 0, 0, 0, 68, 
    0, 75, 166, 36, 68, 0, 0, 0, 147, 258, 3, 0, 92, 100, 287, 
    0, 0, 0, 135, 0, 0, 0, 0, 352, 0, 31, 0, 0, 250, 23, 
    0, 0, 0, 90, 0, 0, 0, 0, 308, 0, 30, 0, 0, 255, 0, 
    0, 0, 34, 101, 24, 112, 134, 161, 260, 0, 94, 97, 13, 67, 0, 
    0, 19, 0, 0, 0, 0, 0, 0, 4, 0, 55, 87, 0, 0, 0, 
    
    -- channel=435
    236, 254, 269, 280, 271, 250, 244, 236, 210, 185, 196, 170, 119, 136, 151, 
    251, 233, 219, 209, 199, 188, 186, 190, 179, 175, 165, 144, 130, 112, 145, 
    186, 180, 173, 167, 168, 156, 158, 172, 167, 165, 115, 115, 129, 127, 145, 
    153, 147, 146, 149, 153, 149, 150, 158, 165, 158, 121, 122, 132, 155, 162, 
    134, 140, 141, 143, 143, 149, 146, 143, 133, 98, 86, 89, 133, 153, 154, 
    137, 137, 140, 146, 137, 121, 66, 53, 57, 67, 27, 55, 130, 114, 140, 
    140, 134, 139, 138, 110, 87, 84, 105, 116, 92, 0, 16, 84, 98, 125, 
    136, 136, 132, 92, 101, 99, 83, 75, 44, 0, 0, 2, 82, 105, 69, 
    129, 129, 97, 95, 78, 112, 102, 0, 0, 0, 0, 68, 59, 39, 6, 
    129, 65, 37, 70, 98, 109, 61, 0, 0, 0, 39, 0, 0, 1, 28, 
    121, 45, 52, 70, 120, 97, 31, 0, 0, 98, 86, 54, 0, 30, 92, 
    119, 78, 38, 77, 107, 49, 27, 0, 25, 84, 94, 80, 31, 42, 122, 
    118, 70, 34, 68, 56, 5, 0, 0, 29, 71, 57, 87, 67, 91, 120, 
    109, 78, 63, 88, 77, 76, 78, 78, 96, 74, 68, 99, 114, 128, 117, 
    101, 90, 88, 77, 90, 89, 92, 96, 110, 100, 80, 126, 125, 126, 125, 
    
    -- channel=436
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 6, 19, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 13, 10, 5, 
    
    -- channel=437
    186, 233, 213, 240, 255, 233, 201, 235, 162, 182, 163, 125, 86, 46, 125, 
    233, 232, 237, 235, 219, 205, 177, 192, 164, 162, 109, 113, 123, 0, 132, 
    176, 216, 201, 200, 172, 169, 166, 158, 149, 136, 0, 146, 73, 21, 149, 
    153, 156, 159, 168, 152, 160, 148, 146, 134, 98, 153, 0, 86, 137, 161, 
    138, 159, 163, 169, 145, 119, 94, 120, 87, 92, 120, 0, 97, 140, 132, 
    155, 166, 168, 164, 118, 28, 0, 0, 0, 71, 0, 246, 0, 109, 126, 
    162, 169, 173, 133, 0, 0, 62, 117, 44, 0, 0, 441, 20, 0, 86, 
    163, 176, 93, 34, 71, 0, 66, 0, 0, 0, 0, 276, 212, 0, 0, 
    168, 120, 34, 0, 83, 0, 0, 0, 0, 0, 68, 436, 0, 0, 0, 
    137, 0, 270, 0, 144, 0, 0, 0, 0, 0, 0, 148, 0, 0, 12, 
    0, 0, 238, 14, 93, 0, 0, 0, 51, 273, 0, 0, 44, 31, 261, 
    16, 9, 0, 143, 0, 0, 0, 0, 383, 0, 39, 0, 0, 232, 73, 
    23, 0, 0, 152, 0, 0, 0, 0, 377, 0, 69, 0, 0, 291, 0, 
    28, 0, 0, 41, 0, 0, 0, 0, 263, 0, 92, 98, 0, 92, 0, 
    36, 47, 8, 0, 0, 0, 0, 0, 12, 0, 33, 119, 0, 0, 0, 
    
    -- channel=438
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 37, 45, 114, 267, 77, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 230, 306, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 53, 97, 122, 220, 279, 270, 75, 0, 22, 
    0, 0, 0, 28, 93, 9, 9, 234, 239, 242, 250, 39, 0, 77, 146, 
    0, 0, 182, 76, 50, 7, 64, 256, 270, 232, 178, 268, 225, 220, 158, 
    0, 53, 252, 104, 13, 64, 113, 271, 285, 81, 11, 101, 271, 209, 62, 
    0, 52, 224, 108, 42, 137, 174, 286, 285, 63, 65, 0, 210, 185, 0, 
    0, 67, 205, 142, 142, 246, 222, 260, 279, 84, 136, 26, 103, 104, 0, 
    0, 4, 127, 103, 84, 84, 88, 87, 125, 66, 97, 45, 0, 7, 0, 
    0, 0, 93, 128, 96, 100, 78, 56, 28, 2, 78, 20, 0, 0, 0, 
    
    -- channel=439
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=440
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 11, 0, 0, 73, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 15, 35, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 32, 0, 0, 0, 
    0, 0, 26, 0, 21, 1, 13, 0, 0, 25, 0, 8, 0, 0, 19, 
    0, 0, 1, 11, 14, 0, 8, 0, 15, 24, 26, 0, 7, 17, 13, 
    0, 16, 0, 12, 0, 0, 0, 0, 0, 0, 0, 12, 0, 10, 12, 
    0, 0, 0, 18, 0, 0, 0, 0, 17, 0, 3, 31, 0, 27, 3, 
    0, 0, 0, 24, 11, 6, 10, 12, 0, 0, 0, 10, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 0, 0, 0, 
    
    -- channel=441
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=442
    29, 25, 20, 23, 27, 38, 40, 46, 57, 58, 70, 83, 83, 103, 86, 
    31, 31, 35, 47, 53, 60, 61, 65, 70, 76, 87, 70, 111, 106, 81, 
    54, 56, 62, 67, 72, 73, 71, 72, 74, 82, 75, 88, 94, 82, 75, 
    79, 79, 77, 76, 75, 73, 70, 63, 64, 70, 77, 111, 81, 74, 78, 
    81, 78, 76, 75, 76, 65, 64, 64, 62, 23, 73, 93, 65, 77, 83, 
    79, 76, 74, 74, 87, 81, 45, 35, 33, 54, 57, 11, 114, 66, 83, 
    75, 74, 72, 91, 70, 72, 51, 66, 92, 144, 16, 0, 88, 100, 89, 
    75, 74, 94, 64, 67, 92, 90, 112, 77, 28, 0, 0, 85, 136, 93, 
    74, 97, 66, 89, 73, 111, 129, 31, 0, 0, 0, 11, 108, 85, 46, 
    107, 67, 21, 104, 92, 130, 139, 8, 0, 0, 49, 29, 33, 20, 2, 
    105, 55, 43, 84, 120, 146, 105, 11, 0, 69, 77, 95, 7, 8, 55, 
    104, 100, 71, 78, 137, 103, 88, 1, 0, 110, 98, 123, 61, 23, 115, 
    114, 106, 81, 86, 120, 65, 35, 1, 0, 120, 72, 101, 92, 70, 121, 
    106, 106, 81, 99, 96, 71, 63, 57, 73, 117, 81, 94, 118, 121, 131, 
    99, 108, 110, 98, 123, 120, 115, 117, 118, 119, 97, 117, 132, 131, 131, 
    
    -- channel=443
    319, 300, 322, 302, 275, 244, 246, 199, 190, 145, 116, 100, 0, 25, 61, 
    303, 278, 249, 229, 211, 182, 184, 154, 142, 119, 138, 47, 0, 51, 90, 
    201, 178, 174, 158, 151, 150, 152, 144, 139, 145, 152, 23, 22, 116, 103, 
    121, 135, 142, 137, 153, 166, 189, 188, 182, 168, 0, 0, 99, 111, 96, 
    133, 145, 150, 150, 173, 196, 206, 228, 277, 232, 31, 42, 119, 99, 94, 
    147, 153, 150, 145, 171, 254, 339, 331, 324, 264, 354, 0, 34, 106, 79, 
    157, 158, 140, 145, 203, 157, 96, 0, 0, 187, 501, 138, 0, 16, 45, 
    161, 155, 178, 176, 90, 100, 47, 120, 282, 470, 501, 188, 0, 0, 159, 
    156, 171, 80, 88, 0, 0, 161, 517, 513, 521, 421, 35, 130, 224, 329, 
    171, 419, 37, 29, 0, 0, 245, 449, 448, 345, 392, 348, 349, 326, 248, 
    235, 235, 74, 0, 0, 11, 287, 412, 269, 0, 33, 336, 311, 219, 0, 
    106, 45, 133, 0, 0, 114, 372, 432, 61, 0, 0, 108, 263, 0, 0, 
    50, 55, 147, 0, 138, 245, 399, 408, 50, 73, 17, 0, 152, 0, 0, 
    37, 43, 49, 0, 44, 90, 110, 110, 0, 72, 6, 0, 0, 0, 0, 
    57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=444
    260, 247, 288, 267, 240, 195, 205, 156, 134, 138, 103, 67, 32, 60, 32, 
    230, 215, 174, 131, 116, 96, 108, 89, 77, 71, 87, 38, 0, 44, 30, 
    165, 109, 78, 56, 60, 58, 62, 77, 76, 79, 183, 104, 35, 106, 70, 
    38, 34, 44, 42, 56, 68, 93, 116, 126, 128, 53, 39, 97, 73, 42, 
    33, 32, 40, 47, 68, 131, 198, 185, 214, 191, 70, 74, 90, 50, 38, 
    34, 36, 45, 49, 76, 192, 392, 474, 537, 502, 573, 19, 91, 114, 25, 
    42, 43, 42, 56, 176, 243, 230, 54, 69, 190, 680, 308, 0, 89, 35, 
    47, 46, 95, 139, 147, 158, 143, 151, 266, 577, 692, 421, 85, 0, 196, 
    40, 70, 76, 170, 122, 89, 193, 732, 749, 743, 649, 72, 86, 212, 453, 
    40, 409, 133, 94, 0, 27, 321, 653, 636, 577, 645, 490, 447, 474, 417, 
    125, 412, 273, 66, 0, 58, 324, 608, 516, 93, 119, 520, 516, 414, 118, 
    54, 92, 304, 4, 0, 217, 491, 625, 276, 66, 12, 159, 434, 150, 0, 
    6, 127, 304, 25, 185, 327, 525, 581, 223, 145, 85, 8, 324, 10, 0, 
    10, 105, 212, 106, 208, 287, 326, 322, 149, 177, 105, 0, 8, 0, 0, 
    53, 24, 16, 1, 0, 0, 0, 0, 0, 46, 94, 0, 0, 0, 0, 
    
    -- channel=445
    268, 301, 328, 333, 318, 272, 261, 240, 194, 189, 154, 115, 87, 46, 67, 
    297, 280, 253, 217, 195, 170, 165, 158, 134, 119, 108, 109, 22, 0, 74, 
    211, 183, 150, 131, 119, 110, 112, 123, 117, 109, 146, 104, 43, 75, 109, 
    90, 84, 91, 93, 98, 107, 120, 139, 148, 141, 125, 2, 79, 110, 100, 
    72, 80, 89, 95, 99, 139, 171, 169, 169, 194, 91, 34, 112, 98, 86, 
    80, 85, 93, 98, 91, 124, 233, 292, 334, 328, 266, 143, 51, 105, 70, 
    90, 92, 98, 80, 130, 172, 197, 104, 64, 0, 344, 319, 0, 66, 52, 
    92, 94, 90, 122, 127, 80, 103, 18, 77, 238, 402, 419, 70, 0, 55, 
    88, 76, 108, 107, 122, 39, 33, 327, 447, 451, 453, 204, 17, 46, 230, 
    54, 168, 196, 23, 33, 0, 33, 362, 373, 416, 364, 285, 228, 278, 294, 
    51, 275, 220, 46, 0, 0, 47, 344, 399, 134, 68, 217, 336, 291, 180, 
    50, 36, 154, 56, 0, 50, 152, 363, 343, 12, 20, 4, 218, 206, 0, 
    14, 47, 137, 43, 8, 129, 235, 349, 292, 22, 68, 0, 137, 101, 0, 
    10, 44, 119, 69, 95, 185, 218, 228, 173, 29, 97, 13, 0, 0, 0, 
    40, 18, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 
    
    -- channel=446
    102, 91, 98, 86, 82, 61, 57, 46, 26, 32, 13, 0, 0, 0, 0, 
    80, 83, 77, 54, 44, 32, 32, 20, 13, 5, 0, 0, 0, 0, 1, 
    45, 43, 30, 23, 13, 19, 20, 15, 15, 10, 1, 17, 0, 9, 18, 
    5, 8, 14, 15, 19, 29, 39, 41, 37, 19, 0, 0, 20, 9, 4, 
    13, 16, 20, 22, 26, 38, 52, 66, 75, 110, 29, 0, 27, 7, 0, 
    17, 21, 22, 19, 10, 36, 122, 165, 169, 171, 203, 107, 0, 49, 0, 
    20, 28, 24, 4, 20, 46, 63, 0, 0, 0, 238, 286, 0, 0, 0, 
    27, 26, 3, 44, 36, 3, 25, 9, 76, 189, 308, 304, 38, 0, 21, 
    27, 1, 0, 3, 31, 0, 0, 227, 316, 325, 344, 161, 10, 39, 170, 
    0, 89, 147, 0, 0, 0, 0, 251, 270, 273, 210, 251, 188, 207, 188, 
    0, 116, 139, 0, 0, 0, 0, 247, 277, 42, 0, 60, 240, 181, 71, 
    0, 0, 84, 10, 0, 0, 78, 271, 259, 0, 0, 0, 127, 134, 0, 
    0, 0, 67, 15, 0, 117, 167, 252, 226, 0, 38, 0, 14, 32, 0, 
    0, 0, 22, 0, 0, 29, 46, 59, 55, 0, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=447
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=448
    80, 75, 86, 81, 116, 134, 96, 78, 65, 68, 58, 47, 42, 42, 32, 
    78, 72, 85, 84, 134, 176, 163, 134, 81, 71, 67, 63, 64, 62, 56, 
    78, 77, 69, 104, 147, 178, 198, 203, 155, 104, 103, 100, 88, 77, 70, 
    80, 80, 40, 93, 168, 179, 191, 216, 205, 177, 152, 121, 85, 73, 80, 
    95, 109, 82, 84, 164, 198, 192, 192, 223, 219, 218, 182, 121, 102, 107, 
    132, 134, 85, 67, 140, 194, 189, 195, 209, 217, 223, 218, 165, 128, 109, 
    125, 120, 112, 23, 121, 194, 193, 210, 204, 188, 208, 226, 176, 133, 87, 
    125, 127, 126, 133, 61, 120, 156, 212, 218, 189, 204, 212, 188, 130, 88, 
    142, 147, 135, 112, 163, 107, 164, 185, 216, 196, 202, 207, 203, 146, 97, 
    159, 176, 176, 142, 198, 152, 182, 184, 214, 205, 208, 207, 197, 111, 77, 
    176, 159, 77, 155, 187, 194, 189, 189, 214, 209, 200, 198, 176, 122, 77, 
    155, 125, 94, 117, 107, 178, 179, 96, 178, 199, 187, 183, 151, 148, 85, 
    104, 105, 98, 106, 103, 113, 169, 138, 171, 209, 182, 190, 156, 132, 132, 
    96, 106, 118, 110, 107, 112, 117, 145, 158, 176, 189, 182, 168, 128, 128, 
    98, 98, 102, 94, 109, 125, 119, 113, 112, 117, 134, 142, 125, 114, 103, 
    
    -- channel=449
    21, 22, 29, 44, 12, 0, 12, 24, 23, 25, 26, 27, 23, 21, 19, 
    20, 23, 29, 11, 0, 0, 0, 0, 11, 18, 9, 9, 10, 23, 34, 
    20, 24, 45, 7, 0, 0, 0, 0, 0, 4, 22, 35, 49, 66, 67, 
    14, 10, 24, 0, 0, 0, 0, 0, 0, 0, 0, 24, 56, 55, 50, 
    0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 63, 60, 
    43, 56, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 83, 86, 
    64, 68, 63, 31, 4, 0, 0, 0, 0, 0, 0, 0, 0, 69, 86, 
    35, 43, 63, 64, 17, 0, 0, 0, 0, 0, 0, 0, 0, 4, 51, 
    31, 28, 25, 4, 45, 48, 26, 0, 0, 0, 0, 0, 0, 1, 96, 
    34, 70, 119, 122, 25, 80, 0, 0, 0, 0, 0, 0, 0, 26, 93, 
    106, 135, 91, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 80, 
    142, 122, 87, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 82, 
    66, 51, 51, 47, 47, 0, 0, 0, 0, 0, 0, 0, 0, 52, 78, 
    37, 40, 54, 77, 72, 60, 0, 3, 0, 0, 0, 0, 0, 65, 74, 
    69, 81, 74, 73, 71, 69, 48, 68, 59, 40, 14, 31, 51, 78, 94, 
    
    -- channel=450
    92, 83, 106, 102, 72, 66, 73, 75, 72, 64, 55, 44, 39, 53, 55, 
    89, 83, 93, 61, 39, 11, 20, 34, 56, 74, 82, 96, 106, 124, 116, 
    74, 75, 57, 39, 0, 0, 0, 0, 64, 125, 123, 127, 121, 116, 97, 
    73, 88, 97, 22, 0, 0, 0, 0, 11, 41, 72, 85, 125, 115, 109, 
    174, 207, 167, 23, 0, 10, 31, 0, 0, 0, 0, 35, 131, 159, 156, 
    220, 209, 145, 39, 19, 36, 0, 0, 0, 0, 0, 0, 99, 176, 164, 
    181, 184, 179, 126, 37, 15, 0, 0, 12, 0, 0, 0, 50, 128, 115, 
    177, 206, 197, 167, 163, 103, 57, 16, 19, 0, 0, 0, 0, 70, 118, 
    216, 268, 308, 230, 211, 174, 126, 37, 0, 0, 0, 0, 0, 46, 102, 
    362, 381, 297, 203, 128, 129, 93, 22, 0, 0, 0, 0, 0, 42, 117, 
    358, 318, 131, 42, 8, 0, 0, 2, 1, 0, 0, 0, 0, 109, 130, 
    180, 133, 123, 108, 9, 0, 30, 39, 0, 0, 24, 13, 32, 124, 134, 
    95, 106, 119, 130, 107, 72, 45, 24, 0, 10, 47, 0, 44, 113, 132, 
    104, 118, 97, 80, 92, 114, 79, 37, 12, 2, 0, 0, 5, 96, 124, 
    91, 79, 86, 99, 125, 133, 96, 94, 98, 75, 51, 46, 60, 106, 123, 
    
    -- channel=451
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 25, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 36, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 87, 106, 36, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    179, 216, 172, 60, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    228, 197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    93, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=452
    88, 86, 81, 83, 102, 112, 98, 75, 71, 69, 58, 50, 42, 36, 34, 
    87, 85, 83, 75, 114, 123, 124, 111, 70, 63, 64, 61, 61, 59, 57, 
    83, 80, 75, 78, 112, 128, 138, 137, 103, 95, 94, 89, 75, 66, 57, 
    80, 80, 67, 80, 124, 134, 137, 141, 140, 113, 116, 101, 66, 65, 59, 
    101, 120, 136, 91, 123, 129, 154, 157, 152, 153, 144, 128, 86, 73, 73, 
    137, 141, 125, 89, 111, 139, 160, 160, 151, 155, 157, 144, 105, 78, 74, 
    129, 125, 117, 110, 89, 122, 156, 154, 149, 154, 153, 150, 125, 78, 66, 
    127, 129, 140, 105, 113, 101, 137, 147, 162, 166, 158, 157, 130, 91, 67, 
    140, 145, 157, 181, 163, 147, 118, 153, 163, 167, 165, 162, 141, 111, 58, 
    184, 203, 196, 188, 160, 144, 127, 159, 166, 170, 170, 170, 148, 84, 24, 
    204, 203, 161, 133, 154, 140, 147, 124, 159, 163, 154, 157, 130, 71, 41, 
    171, 130, 114, 116, 123, 129, 119, 109, 122, 143, 146, 154, 108, 66, 60, 
    104, 100, 90, 96, 91, 104, 109, 112, 128, 150, 165, 160, 122, 70, 56, 
    84, 92, 97, 76, 52, 63, 84, 104, 107, 123, 128, 150, 125, 60, 53, 
    77, 57, 47, 41, 39, 60, 81, 58, 49, 60, 75, 79, 65, 41, 32, 
    
    -- channel=453
    7, 10, 0, 7, 0, 0, 10, 2, 7, 0, 0, 2, 0, 0, 0, 
    7, 13, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 6, 
    2, 4, 7, 0, 0, 0, 0, 0, 0, 0, 5, 2, 4, 6, 4, 
    0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 6, 0, 
    3, 10, 68, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    10, 21, 100, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    16, 22, 40, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    10, 13, 28, 41, 95, 0, 3, 0, 0, 8, 0, 0, 0, 0, 1, 
    8, 11, 54, 77, 38, 61, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    35, 38, 59, 122, 0, 70, 0, 20, 0, 0, 0, 0, 0, 6, 0, 
    57, 83, 144, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    53, 47, 66, 32, 35, 0, 0, 19, 0, 0, 0, 0, 0, 0, 24, 
    19, 5, 6, 2, 30, 2, 0, 10, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=454
    81, 78, 88, 81, 85, 90, 81, 72, 71, 69, 63, 56, 55, 61, 59, 
    81, 76, 83, 78, 79, 88, 81, 84, 71, 75, 80, 81, 83, 86, 80, 
    76, 75, 64, 71, 74, 84, 88, 91, 98, 96, 97, 94, 87, 82, 74, 
    77, 84, 76, 76, 76, 91, 97, 103, 104, 94, 93, 90, 88, 81, 81, 
    118, 128, 95, 66, 77, 101, 108, 99, 101, 100, 97, 95, 105, 98, 100, 
    132, 126, 84, 72, 89, 117, 99, 87, 103, 103, 100, 105, 112, 110, 103, 
    116, 114, 107, 77, 80, 94, 83, 96, 107, 99, 96, 104, 104, 103, 85, 
    118, 126, 117, 103, 99, 116, 101, 107, 110, 95, 93, 97, 94, 99, 87, 
    137, 158, 165, 143, 128, 107, 108, 105, 107, 96, 96, 93, 100, 92, 77, 
    185, 188, 152, 96, 126, 94, 117, 93, 105, 100, 101, 90, 94, 80, 79, 
    175, 150, 87, 83, 87, 77, 87, 91, 101, 98, 95, 90, 92, 95, 89, 
    105, 91, 74, 91, 75, 82, 103, 85, 89, 99, 105, 101, 91, 106, 86, 
    77, 87, 91, 93, 77, 85, 96, 78, 89, 111, 108, 97, 94, 102, 96, 
    88, 91, 84, 75, 79, 86, 95, 83, 80, 90, 82, 85, 90, 93, 98, 
    76, 72, 76, 80, 96, 97, 87, 85, 86, 82, 84, 80, 76, 90, 88, 
    
    -- channel=455
    0, 1, 0, 1, 0, 0, 14, 1, 4, 0, 4, 7, 3, 0, 2, 
    0, 2, 0, 4, 0, 0, 2, 6, 11, 0, 0, 0, 0, 0, 3, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 6, 
    0, 0, 13, 3, 0, 0, 0, 0, 0, 0, 0, 9, 0, 5, 2, 
    0, 0, 29, 44, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 40, 57, 0, 0, 4, 9, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 75, 0, 0, 8, 0, 0, 6, 4, 0, 0, 0, 16, 
    0, 0, 1, 18, 51, 0, 1, 0, 0, 12, 8, 0, 0, 0, 4, 
    0, 0, 0, 47, 0, 34, 0, 16, 0, 2, 5, 8, 0, 10, 14, 
    0, 0, 22, 58, 0, 33, 0, 29, 0, 0, 0, 17, 0, 22, 4, 
    0, 17, 103, 0, 2, 4, 0, 0, 0, 0, 0, 7, 5, 0, 21, 
    22, 11, 46, 9, 25, 0, 0, 25, 0, 0, 0, 1, 22, 0, 27, 
    11, 0, 0, 0, 23, 8, 0, 14, 0, 0, 0, 7, 24, 0, 0, 
    0, 0, 1, 8, 0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 0, 
    5, 1, 0, 5, 0, 0, 3, 7, 1, 0, 0, 0, 2, 0, 0, 
    
    -- channel=456
    212, 202, 198, 209, 228, 244, 213, 177, 161, 148, 121, 97, 74, 63, 61, 
    207, 199, 193, 169, 232, 236, 249, 212, 151, 145, 140, 141, 146, 150, 144, 
    190, 188, 161, 146, 202, 214, 227, 234, 218, 238, 235, 225, 195, 175, 143, 
    180, 186, 163, 130, 193, 217, 231, 254, 244, 238, 261, 234, 179, 169, 150, 
    277, 338, 354, 171, 194, 251, 308, 286, 270, 260, 263, 264, 220, 208, 204, 
    388, 401, 371, 177, 204, 266, 308, 293, 280, 278, 269, 259, 242, 234, 221, 
    363, 358, 356, 249, 176, 239, 297, 281, 292, 292, 274, 258, 255, 212, 183, 
    349, 370, 387, 343, 293, 217, 283, 281, 325, 325, 285, 259, 246, 194, 175, 
    395, 435, 501, 461, 453, 363, 309, 305, 313, 326, 305, 281, 254, 221, 143, 
    576, 625, 594, 541, 421, 400, 305, 319, 312, 327, 327, 301, 249, 163, 79, 
    644, 625, 402, 316, 305, 287, 269, 251, 304, 312, 295, 280, 228, 178, 117, 
    479, 379, 324, 300, 232, 203, 239, 196, 208, 261, 296, 300, 207, 175, 163, 
    268, 251, 241, 253, 251, 218, 216, 226, 232, 288, 348, 319, 245, 158, 173, 
    211, 227, 227, 175, 131, 173, 174, 205, 190, 209, 254, 277, 239, 142, 135, 
    181, 133, 114, 105, 104, 164, 181, 140, 112, 125, 137, 156, 138, 102, 94, 
    
    -- channel=457
    188, 178, 169, 165, 91, 46, 95, 137, 146, 137, 137, 137, 127, 118, 110, 
    188, 175, 154, 110, 22, 0, 0, 0, 79, 98, 72, 72, 76, 83, 80, 
    178, 169, 128, 70, 0, 0, 0, 0, 0, 75, 62, 46, 55, 67, 45, 
    152, 148, 94, 7, 0, 0, 0, 0, 0, 0, 14, 0, 45, 50, 0, 
    151, 167, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    177, 185, 147, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    192, 182, 169, 53, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    175, 162, 143, 84, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    153, 150, 152, 96, 58, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    221, 239, 237, 157, 64, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    286, 268, 117, 67, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    268, 229, 166, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    177, 162, 132, 92, 45, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    98, 78, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=458
    72, 75, 83, 78, 100, 117, 101, 88, 83, 88, 90, 89, 92, 94, 90, 
    73, 72, 85, 99, 120, 155, 143, 135, 109, 91, 96, 93, 91, 88, 88, 
    79, 78, 90, 123, 143, 172, 185, 192, 157, 94, 97, 100, 105, 100, 106, 
    85, 81, 67, 127, 164, 172, 185, 200, 202, 164, 127, 122, 108, 98, 113, 
    61, 52, 43, 121, 166, 159, 150, 175, 205, 205, 196, 166, 126, 120, 130, 
    60, 61, 31, 111, 135, 150, 149, 167, 183, 197, 210, 196, 165, 143, 134, 
    65, 64, 51, 61, 134, 163, 159, 175, 167, 165, 189, 204, 176, 148, 121, 
    65, 63, 65, 82, 62, 119, 136, 183, 166, 147, 178, 200, 173, 144, 116, 
    66, 55, 24, 58, 72, 85, 122, 163, 168, 146, 167, 183, 178, 156, 149, 
    19, 20, 41, 38, 99, 89, 134, 161, 167, 150, 159, 176, 183, 155, 158, 
    11, 14, 59, 105, 152, 155, 174, 175, 171, 166, 167, 176, 179, 151, 150, 
    57, 60, 75, 81, 110, 176, 154, 125, 166, 171, 153, 151, 176, 172, 145, 
    85, 85, 83, 93, 95, 116, 155, 141, 151, 160, 123, 146, 170, 180, 162, 
    94, 101, 117, 137, 150, 138, 144, 150, 170, 174, 153, 152, 171, 182, 180, 
    119, 140, 154, 161, 173, 154, 153, 166, 177, 168, 169, 171, 171, 187, 180, 
    
    -- channel=459
    92, 88, 85, 102, 107, 109, 99, 90, 75, 68, 61, 51, 37, 26, 21, 
    90, 87, 89, 70, 112, 113, 122, 103, 80, 63, 51, 44, 46, 53, 59, 
    85, 86, 92, 69, 94, 92, 106, 100, 85, 99, 100, 106, 98, 97, 87, 
    77, 75, 63, 44, 79, 78, 81, 106, 117, 120, 126, 129, 91, 85, 79, 
    74, 100, 169, 79, 76, 90, 118, 120, 118, 116, 125, 129, 108, 104, 102, 
    166, 183, 206, 69, 68, 85, 134, 127, 114, 115, 120, 111, 117, 132, 125, 
    174, 171, 164, 112, 75, 112, 142, 121, 120, 120, 122, 102, 128, 126, 117, 
    149, 154, 181, 161, 142, 46, 118, 113, 133, 140, 124, 109, 114, 96, 82, 
    162, 166, 171, 160, 202, 176, 136, 137, 129, 137, 123, 118, 104, 107, 121, 
    197, 255, 303, 301, 216, 234, 143, 153, 123, 132, 133, 130, 107, 94, 63, 
    294, 312, 248, 178, 152, 171, 139, 119, 130, 138, 142, 119, 95, 90, 80, 
    306, 240, 153, 155, 109, 79, 80, 97, 82, 97, 113, 128, 105, 98, 103, 
    138, 136, 118, 116, 126, 95, 111, 103, 91, 98, 140, 140, 124, 96, 105, 
    95, 104, 132, 130, 94, 93, 82, 104, 95, 101, 131, 123, 120, 95, 93, 
    118, 108, 84, 73, 67, 101, 101, 96, 79, 76, 80, 98, 93, 76, 82, 
    
    -- channel=460
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=461
    123, 117, 124, 125, 138, 123, 102, 107, 92, 92, 84, 73, 62, 56, 39, 
    122, 111, 117, 111, 124, 145, 131, 102, 84, 82, 59, 50, 49, 54, 53, 
    119, 115, 100, 120, 114, 110, 118, 107, 95, 98, 98, 94, 89, 91, 78, 
    107, 104, 45, 66, 111, 97, 91, 103, 109, 135, 138, 104, 82, 72, 60, 
    94, 112, 97, 71, 102, 142, 121, 101, 108, 113, 134, 118, 91, 61, 59, 
    173, 186, 126, 55, 85, 131, 139, 126, 114, 103, 103, 125, 104, 83, 74, 
    189, 179, 153, 26, 93, 173, 141, 127, 127, 111, 105, 125, 111, 108, 87, 
    167, 162, 162, 145, 38, 64, 89, 119, 150, 131, 112, 110, 115, 92, 62, 
    173, 171, 140, 107, 161, 90, 126, 106, 156, 145, 120, 109, 124, 97, 68, 
    184, 231, 271, 215, 220, 146, 157, 116, 147, 151, 136, 117, 117, 53, 17, 
    277, 264, 162, 185, 183, 179, 152, 138, 148, 150, 136, 109, 84, 50, 12, 
    302, 249, 147, 135, 88, 114, 114, 70, 125, 132, 129, 110, 60, 80, 22, 
    160, 158, 135, 120, 96, 81, 129, 97, 122, 152, 148, 139, 73, 53, 66, 
    112, 113, 122, 106, 79, 68, 70, 85, 94, 132, 171, 135, 91, 48, 58, 
    104, 88, 56, 30, 45, 73, 68, 44, 30, 43, 71, 79, 47, 28, 29, 
    
    -- channel=462
    0, 0, 0, 0, 0, 0, 6, 1, 1, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 15, 7, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 17, 0, 5, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 34, 47, 0, 0, 0, 21, 6, 2, 0, 5, 0, 0, 0, 
    0, 0, 61, 39, 1, 0, 11, 27, 1, 7, 11, 0, 0, 0, 0, 
    0, 0, 2, 84, 0, 0, 27, 3, 0, 17, 17, 0, 0, 0, 13, 
    0, 0, 0, 10, 67, 0, 9, 0, 0, 26, 23, 8, 0, 0, 0, 
    0, 0, 0, 23, 11, 42, 0, 24, 0, 18, 20, 22, 0, 0, 7, 
    0, 0, 0, 94, 0, 54, 0, 48, 0, 4, 12, 32, 1, 14, 0, 
    0, 14, 110, 8, 6, 24, 9, 4, 0, 4, 13, 25, 0, 0, 2, 
    29, 26, 45, 18, 39, 0, 0, 29, 0, 0, 0, 14, 9, 0, 29, 
    6, 0, 0, 0, 24, 9, 0, 26, 0, 0, 6, 15, 27, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 1, 0, 0, 15, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=463
    186, 169, 186, 173, 190, 215, 168, 156, 136, 127, 103, 79, 66, 70, 63, 
    182, 170, 176, 129, 185, 193, 206, 170, 126, 133, 130, 139, 143, 144, 128, 
    165, 166, 110, 134, 154, 172, 178, 196, 210, 217, 200, 192, 158, 137, 106, 
    163, 176, 136, 91, 161, 185, 192, 199, 191, 211, 224, 173, 159, 135, 124, 
    282, 328, 263, 88, 153, 249, 261, 195, 210, 203, 219, 222, 193, 173, 167, 
    343, 340, 269, 81, 188, 261, 227, 219, 230, 205, 205, 222, 205, 193, 168, 
    305, 300, 303, 143, 139, 212, 226, 228, 254, 216, 201, 215, 197, 180, 124, 
    313, 332, 314, 280, 201, 202, 212, 232, 284, 244, 206, 199, 212, 162, 150, 
    357, 412, 469, 324, 398, 265, 284, 208, 268, 256, 234, 209, 219, 162, 80, 
    531, 544, 438, 394, 328, 295, 247, 221, 266, 267, 259, 215, 196, 99, 59, 
    543, 488, 187, 242, 232, 205, 211, 192, 253, 247, 224, 212, 173, 158, 62, 
    333, 273, 251, 230, 138, 161, 238, 114, 187, 229, 253, 228, 133, 158, 104, 
    215, 207, 206, 216, 195, 157, 181, 181, 197, 270, 292, 232, 172, 119, 156, 
    186, 196, 169, 112, 103, 158, 135, 157, 148, 167, 219, 216, 162, 96, 107, 
    124, 84, 88, 73, 88, 148, 134, 89, 78, 100, 110, 117, 95, 67, 67, 
    
    -- channel=464
    230, 213, 229, 239, 219, 213, 195, 181, 161, 142, 115, 87, 59, 55, 46, 
    223, 207, 210, 166, 178, 161, 170, 144, 133, 138, 125, 128, 136, 153, 147, 
    200, 197, 154, 130, 104, 82, 84, 97, 161, 231, 233, 228, 208, 195, 154, 
    182, 193, 149, 69, 58, 66, 78, 104, 124, 186, 232, 206, 200, 182, 149, 
    304, 375, 346, 99, 62, 149, 191, 131, 105, 107, 141, 180, 215, 221, 207, 
    466, 483, 388, 123, 108, 178, 190, 145, 129, 111, 98, 129, 209, 256, 239, 
    444, 439, 418, 228, 131, 179, 179, 141, 173, 153, 107, 112, 177, 220, 197, 
    414, 444, 447, 384, 260, 176, 187, 162, 212, 194, 119, 93, 134, 154, 175, 
    468, 535, 590, 480, 476, 352, 288, 191, 195, 199, 149, 104, 122, 155, 140, 
    703, 778, 745, 603, 436, 382, 273, 205, 187, 203, 188, 126, 106, 94, 75, 
    831, 787, 452, 306, 253, 203, 170, 162, 186, 192, 176, 122, 100, 144, 98, 
    618, 489, 378, 297, 138, 64, 154, 121, 106, 142, 191, 172, 111, 164, 141, 
    317, 297, 283, 282, 238, 160, 161, 141, 122, 187, 258, 200, 143, 127, 168, 
    229, 244, 230, 177, 140, 166, 131, 133, 103, 134, 186, 161, 126, 101, 127, 
    187, 136, 106, 87, 102, 165, 150, 105, 79, 80, 85, 107, 89, 76, 83, 
    
    -- channel=465
    130, 124, 114, 129, 136, 155, 139, 115, 101, 90, 75, 59, 42, 26, 27, 
    126, 125, 115, 87, 151, 147, 175, 141, 99, 80, 74, 77, 84, 89, 90, 
    114, 115, 107, 83, 123, 132, 136, 146, 145, 156, 150, 147, 127, 115, 92, 
    107, 104, 98, 53, 111, 125, 133, 154, 152, 152, 170, 156, 113, 103, 93, 
    151, 201, 268, 113, 119, 150, 199, 184, 174, 166, 168, 183, 137, 131, 132, 
    241, 253, 277, 105, 120, 134, 193, 196, 178, 173, 177, 157, 148, 153, 148, 
    226, 223, 230, 184, 93, 141, 206, 178, 184, 187, 179, 156, 174, 139, 125, 
    210, 224, 255, 236, 216, 91, 178, 170, 210, 220, 187, 166, 162, 112, 107, 
    235, 246, 298, 292, 318, 268, 200, 196, 195, 212, 199, 186, 157, 148, 104, 
    353, 401, 399, 425, 260, 308, 173, 221, 195, 206, 212, 205, 158, 111, 50, 
    410, 424, 278, 189, 196, 195, 182, 157, 194, 205, 192, 182, 144, 121, 77, 
    337, 244, 234, 205, 149, 111, 143, 121, 101, 149, 187, 193, 136, 101, 124, 
    173, 156, 141, 157, 186, 151, 126, 159, 137, 165, 230, 209, 179, 95, 114, 
    122, 140, 152, 118, 72, 111, 96, 126, 119, 120, 157, 178, 161, 92, 77, 
    122, 83, 65, 65, 51, 100, 120, 91, 67, 76, 71, 92, 92, 60, 61, 
    
    -- channel=466
    136, 136, 123, 123, 150, 153, 147, 137, 135, 139, 137, 138, 139, 133, 132, 
    136, 136, 130, 139, 173, 189, 184, 178, 142, 134, 131, 132, 134, 126, 121, 
    139, 136, 131, 149, 194, 212, 218, 203, 165, 145, 130, 120, 107, 99, 98, 
    140, 136, 115, 177, 226, 217, 211, 204, 188, 163, 159, 129, 92, 102, 104, 
    132, 136, 132, 162, 223, 206, 207, 211, 211, 213, 208, 170, 107, 86, 89, 
    104, 96, 96, 148, 188, 214, 213, 214, 206, 209, 213, 203, 118, 63, 66, 
    91, 85, 93, 101, 154, 179, 202, 217, 206, 204, 212, 222, 147, 82, 75, 
    107, 98, 99, 101, 120, 160, 170, 198, 213, 213, 222, 224, 186, 131, 97, 
    101, 80, 78, 121, 109, 107, 124, 191, 219, 217, 224, 233, 216, 148, 71, 
    84, 71, 66, 76, 139, 107, 158, 183, 225, 223, 220, 237, 217, 112, 55, 
    40, 41, 63, 124, 167, 180, 186, 162, 211, 211, 196, 215, 185, 97, 73, 
    58, 50, 74, 129, 172, 211, 177, 157, 192, 205, 196, 195, 142, 90, 66, 
    101, 110, 101, 110, 124, 158, 167, 166, 222, 219, 203, 207, 144, 88, 75, 
    113, 119, 119, 93, 77, 95, 135, 149, 169, 175, 183, 200, 159, 77, 74, 
    106, 84, 77, 77, 73, 86, 105, 81, 86, 109, 132, 119, 97, 67, 58, 
    
    -- channel=467
    62, 63, 50, 70, 21, 9, 46, 59, 65, 58, 63, 67, 61, 54, 63, 
    62, 67, 53, 31, 3, 0, 0, 0, 47, 49, 45, 45, 47, 57, 69, 
    56, 61, 74, 4, 0, 0, 0, 0, 0, 37, 43, 53, 63, 77, 76, 
    49, 48, 87, 0, 0, 0, 0, 0, 0, 0, 0, 40, 66, 69, 55, 
    35, 42, 125, 29, 0, 0, 0, 0, 0, 0, 0, 0, 32, 55, 47, 
    67, 78, 166, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 67, 
    79, 85, 98, 132, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 84, 
    58, 62, 83, 74, 126, 0, 0, 0, 0, 0, 0, 0, 0, 5, 51, 
    51, 52, 79, 67, 64, 95, 5, 0, 0, 0, 0, 0, 0, 0, 73, 
    70, 97, 129, 171, 20, 113, 0, 0, 0, 0, 0, 0, 0, 27, 57, 
    127, 161, 176, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 65, 
    149, 132, 101, 76, 28, 0, 0, 24, 0, 0, 0, 0, 0, 0, 74, 
    74, 69, 64, 52, 74, 23, 0, 0, 0, 0, 0, 0, 0, 8, 30, 
    48, 43, 48, 58, 40, 36, 6, 0, 0, 0, 0, 0, 0, 18, 18, 
    62, 58, 39, 38, 15, 30, 23, 33, 24, 13, 0, 0, 20, 18, 42, 
    
    -- channel=468
    17, 13, 31, 8, 0, 0, 0, 1, 8, 13, 12, 10, 16, 28, 15, 
    17, 7, 24, 5, 0, 0, 0, 0, 0, 4, 4, 7, 13, 18, 6, 
    18, 10, 1, 13, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    16, 18, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 27, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 1, 21, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=469
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 15, 23, 25, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 14, 15, 11, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=470
    0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 6, 1, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 36, 36, 13, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 26, 19, 3, 14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 27, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=471
    62, 65, 68, 72, 101, 119, 99, 82, 74, 79, 78, 74, 75, 73, 71, 
    62, 66, 76, 77, 133, 156, 161, 140, 98, 83, 88, 88, 88, 89, 91, 
    66, 69, 87, 111, 145, 177, 193, 202, 156, 106, 107, 115, 108, 105, 109, 
    72, 69, 77, 106, 156, 175, 191, 217, 213, 162, 137, 135, 112, 104, 123, 
    58, 62, 104, 126, 158, 164, 171, 198, 227, 223, 206, 181, 144, 144, 154, 
    74, 74, 84, 101, 140, 140, 157, 188, 203, 220, 233, 197, 177, 169, 155, 
    70, 72, 71, 103, 124, 160, 187, 192, 178, 184, 215, 204, 189, 156, 127, 
    70, 73, 93, 101, 118, 106, 168, 194, 179, 174, 200, 210, 182, 140, 127, 
    77, 65, 56, 86, 135, 148, 158, 184, 170, 164, 188, 201, 178, 167, 175, 
    52, 66, 78, 128, 115, 155, 143, 192, 172, 163, 183, 199, 186, 173, 169, 
    48, 68, 84, 109, 152, 169, 180, 180, 187, 183, 189, 195, 188, 177, 167, 
    80, 63, 90, 106, 129, 163, 153, 136, 150, 162, 163, 180, 194, 184, 182, 
    79, 80, 80, 101, 126, 146, 158, 157, 148, 150, 147, 165, 205, 196, 181, 
    91, 109, 134, 153, 153, 154, 148, 170, 180, 168, 153, 165, 191, 205, 191, 
    134, 152, 165, 174, 176, 172, 177, 193, 195, 184, 178, 188, 196, 201, 195, 
    
    -- channel=472
    119, 118, 106, 122, 135, 138, 131, 105, 98, 92, 81, 71, 55, 40, 40, 
    118, 117, 110, 105, 139, 143, 147, 129, 98, 83, 74, 63, 56, 56, 64, 
    115, 111, 116, 92, 136, 134, 149, 143, 99, 103, 109, 112, 106, 103, 96, 
    104, 102, 97, 86, 129, 134, 134, 142, 155, 142, 143, 145, 99, 95, 80, 
    99, 117, 184, 117, 123, 115, 154, 169, 160, 159, 160, 149, 105, 102, 96, 
    181, 207, 230, 119, 110, 124, 194, 182, 158, 163, 169, 153, 123, 121, 122, 
    200, 200, 187, 167, 114, 136, 186, 166, 160, 170, 167, 148, 151, 120, 124, 
    179, 179, 206, 153, 151, 89, 161, 153, 173, 191, 175, 162, 148, 113, 91, 
    185, 191, 204, 232, 210, 207, 146, 182, 181, 194, 179, 173, 142, 127, 111, 
    216, 262, 317, 323, 238, 242, 160, 201, 180, 188, 186, 189, 155, 120, 49, 
    324, 345, 333, 250, 215, 210, 181, 158, 177, 186, 186, 182, 140, 84, 65, 
    335, 291, 200, 169, 177, 141, 115, 143, 142, 154, 158, 174, 132, 82, 100, 
    182, 164, 148, 135, 125, 112, 127, 139, 129, 138, 186, 188, 141, 91, 85, 
    122, 120, 142, 136, 101, 94, 101, 126, 127, 146, 171, 178, 155, 83, 81, 
    122, 111, 88, 70, 49, 87, 110, 91, 74, 81, 94, 114, 104, 62, 62, 
    
    -- channel=473
    35, 28, 58, 56, 14, 4, 11, 27, 26, 20, 14, 7, 7, 24, 22, 
    31, 27, 46, 9, 0, 0, 0, 0, 12, 32, 38, 56, 71, 91, 84, 
    20, 26, 17, 0, 0, 0, 0, 0, 17, 74, 79, 87, 90, 89, 73, 
    22, 34, 36, 0, 0, 0, 0, 0, 0, 0, 18, 32, 95, 86, 88, 
    109, 139, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 139, 140, 
    150, 135, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 165, 152, 
    117, 118, 116, 38, 10, 0, 0, 0, 0, 0, 0, 0, 8, 114, 96, 
    105, 137, 130, 134, 73, 50, 0, 0, 0, 0, 0, 0, 0, 28, 96, 
    143, 185, 215, 122, 141, 97, 90, 0, 0, 0, 0, 0, 0, 16, 96, 
    275, 289, 217, 113, 57, 64, 37, 0, 0, 0, 0, 0, 0, 13, 135, 
    255, 221, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98, 134, 
    96, 54, 83, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 128, 123, 
    46, 50, 65, 89, 75, 25, 0, 0, 0, 0, 0, 0, 7, 108, 142, 
    59, 80, 62, 58, 80, 103, 38, 7, 0, 0, 0, 0, 0, 102, 131, 
    68, 66, 85, 107, 141, 130, 79, 94, 100, 67, 32, 32, 56, 127, 143, 
    
    -- channel=474
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 10, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    13, 11, 0, 0, 0, 27, 0, 0, 0, 0, 2, 0, 7, 0, 1, 
    15, 3, 0, 0, 0, 50, 0, 0, 0, 0, 0, 11, 28, 14, 0, 
    6, 0, 0, 0, 28, 36, 0, 0, 0, 0, 0, 11, 0, 30, 0, 
    6, 9, 0, 0, 0, 31, 0, 1, 0, 0, 0, 0, 0, 8, 0, 
    18, 30, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 4, 0, 0, 
    25, 21, 0, 0, 12, 0, 27, 0, 0, 0, 0, 0, 0, 0, 9, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 0, 21, 4, 0, 0, 0, 52, 0, 
    0, 0, 0, 0, 0, 0, 29, 0, 0, 27, 0, 0, 0, 24, 27, 
    0, 4, 0, 0, 8, 9, 0, 0, 0, 19, 4, 0, 0, 2, 40, 
    0, 0, 5, 5, 44, 34, 0, 0, 6, 5, 19, 8, 0, 25, 23, 
    
    -- channel=475
    114, 105, 122, 129, 128, 149, 120, 102, 85, 76, 58, 39, 26, 27, 25, 
    110, 104, 114, 81, 128, 127, 151, 121, 86, 86, 87, 95, 107, 121, 116, 
    94, 99, 82, 80, 85, 96, 104, 127, 158, 171, 175, 177, 157, 146, 121, 
    93, 103, 98, 38, 58, 83, 107, 151, 157, 156, 172, 166, 154, 137, 139, 
    186, 239, 247, 83, 63, 140, 176, 150, 158, 150, 151, 181, 199, 208, 211, 
    285, 284, 255, 74, 104, 131, 137, 137, 153, 154, 150, 146, 206, 254, 230, 
    252, 252, 255, 157, 80, 140, 158, 141, 161, 151, 149, 132, 185, 208, 168, 
    237, 266, 278, 281, 232, 120, 170, 165, 183, 163, 138, 123, 143, 142, 156, 
    287, 331, 381, 292, 359, 270, 247, 181, 154, 152, 144, 127, 127, 151, 167, 
    442, 490, 441, 403, 277, 307, 206, 190, 147, 148, 162, 134, 113, 124, 145, 
    481, 459, 234, 155, 150, 154, 139, 150, 164, 159, 161, 128, 122, 189, 166, 
    326, 236, 215, 202, 87, 61, 138, 93, 76, 116, 160, 166, 149, 202, 199, 
    156, 158, 158, 181, 192, 143, 143, 135, 101, 142, 186, 161, 192, 183, 215, 
    139, 164, 169, 152, 139, 173, 132, 135, 111, 99, 124, 123, 149, 182, 181, 
    146, 131, 134, 143, 162, 193, 170, 168, 154, 135, 113, 128, 142, 164, 173, 
    
    -- channel=476
    166, 158, 146, 159, 139, 143, 137, 139, 136, 122, 109, 100, 86, 76, 81, 
    164, 161, 142, 112, 128, 90, 129, 107, 107, 117, 107, 112, 118, 124, 124, 
    147, 151, 123, 92, 88, 67, 55, 56, 100, 162, 158, 149, 134, 130, 108, 
    139, 144, 152, 51, 64, 64, 57, 55, 52, 90, 138, 132, 124, 122, 102, 
    198, 238, 272, 112, 60, 103, 139, 98, 65, 57, 67, 113, 121, 122, 114, 
    256, 262, 309, 109, 107, 91, 125, 116, 92, 73, 61, 66, 85, 121, 123, 
    241, 241, 260, 212, 64, 92, 134, 98, 112, 112, 83, 51, 93, 104, 119, 
    231, 242, 250, 244, 247, 87, 131, 86, 131, 150, 99, 62, 90, 87, 108, 
    252, 277, 344, 270, 303, 234, 173, 119, 117, 148, 118, 93, 80, 88, 74, 
    375, 404, 370, 405, 224, 274, 131, 142, 116, 138, 133, 111, 72, 69, 35, 
    420, 416, 276, 164, 124, 126, 96, 94, 114, 120, 116, 99, 66, 91, 55, 
    318, 258, 239, 216, 132, 54, 100, 102, 56, 84, 128, 130, 64, 55, 96, 
    179, 173, 164, 161, 184, 132, 85, 122, 92, 109, 181, 139, 105, 37, 79, 
    139, 140, 129, 92, 57, 95, 76, 80, 63, 54, 107, 120, 84, 38, 28, 
    109, 68, 46, 38, 21, 71, 78, 51, 26, 37, 29, 41, 45, 11, 22, 
    
    -- channel=477
    273, 250, 276, 274, 250, 249, 222, 214, 191, 173, 142, 108, 81, 80, 62, 
    267, 243, 255, 182, 208, 205, 202, 175, 157, 164, 146, 149, 163, 182, 167, 
    240, 236, 176, 156, 123, 111, 113, 123, 203, 273, 266, 255, 227, 210, 158, 
    220, 234, 150, 77, 87, 97, 101, 129, 145, 227, 267, 220, 215, 187, 151, 
    358, 439, 374, 77, 96, 219, 237, 139, 126, 132, 174, 212, 242, 216, 204, 
    527, 534, 400, 96, 139, 247, 222, 162, 162, 126, 116, 171, 233, 251, 228, 
    491, 479, 453, 174, 151, 237, 205, 175, 220, 169, 125, 151, 196, 236, 190, 
    463, 491, 482, 413, 249, 202, 197, 191, 272, 223, 137, 120, 173, 181, 179, 
    526, 594, 639, 473, 522, 347, 318, 194, 252, 236, 175, 131, 174, 178, 120, 
    783, 863, 797, 606, 492, 400, 312, 198, 240, 250, 225, 148, 146, 79, 44, 
    897, 829, 380, 318, 278, 222, 199, 182, 231, 235, 202, 137, 122, 146, 69, 
    655, 501, 368, 330, 126, 94, 214, 110, 138, 184, 233, 198, 103, 177, 97, 
    336, 332, 306, 305, 255, 176, 202, 155, 166, 257, 313, 228, 138, 116, 165, 
    254, 272, 248, 172, 126, 165, 134, 148, 116, 167, 231, 185, 133, 81, 114, 
    196, 125, 84, 57, 91, 169, 138, 77, 52, 69, 92, 107, 63, 45, 55, 
    
    -- channel=478
    0, 0, 0, 0, 0, 0, 16, 0, 8, 0, 8, 21, 9, 0, 8, 
    0, 5, 0, 0, 0, 0, 4, 0, 8, 0, 0, 0, 0, 0, 4, 
    0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 39, 
    0, 0, 95, 0, 0, 0, 0, 0, 0, 0, 0, 39, 2, 24, 15, 
    0, 0, 165, 87, 0, 0, 0, 5, 0, 0, 0, 0, 0, 7, 1, 
    0, 0, 270, 71, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 37, 252, 0, 0, 21, 0, 0, 0, 3, 0, 0, 0, 73, 
    0, 0, 4, 32, 243, 0, 16, 0, 0, 20, 4, 0, 0, 0, 5, 
    0, 0, 0, 27, 43, 147, 0, 12, 0, 0, 0, 0, 0, 0, 86, 
    0, 0, 11, 293, 0, 235, 0, 66, 0, 0, 0, 22, 0, 75, 34, 
    0, 80, 336, 51, 0, 44, 0, 0, 0, 0, 0, 7, 0, 14, 67, 
    108, 108, 92, 73, 111, 0, 0, 71, 0, 0, 0, 11, 30, 0, 126, 
    10, 0, 0, 0, 74, 13, 0, 44, 0, 0, 0, 0, 65, 0, 0, 
    0, 0, 5, 50, 0, 0, 0, 0, 0, 0, 0, 0, 27, 18, 0, 
    26, 40, 17, 24, 0, 0, 10, 45, 14, 0, 0, 0, 43, 0, 18, 
    
    -- channel=479
    0, 0, 0, 0, 3, 0, 0, 0, 4, 11, 13, 21, 26, 29, 28, 
    0, 0, 0, 7, 17, 23, 14, 13, 8, 13, 11, 11, 11, 10, 10, 
    0, 0, 10, 25, 32, 39, 43, 33, 7, 0, 0, 0, 0, 2, 11, 
    0, 0, 0, 43, 44, 38, 38, 43, 29, 9, 2, 0, 0, 5, 16, 
    0, 0, 0, 25, 41, 28, 15, 32, 39, 36, 28, 9, 0, 0, 5, 
    0, 0, 0, 15, 25, 24, 10, 21, 28, 39, 37, 27, 6, 0, 0, 
    0, 0, 0, 0, 27, 27, 15, 25, 16, 23, 37, 34, 11, 4, 3, 
    0, 0, 0, 0, 0, 12, 11, 27, 9, 10, 33, 35, 22, 12, 4, 
    0, 0, 0, 0, 0, 0, 0, 17, 10, 8, 22, 32, 28, 14, 21, 
    0, 0, 0, 0, 0, 0, 7, 6, 11, 8, 14, 26, 27, 18, 33, 
    0, 0, 0, 0, 0, 12, 13, 22, 16, 10, 18, 22, 24, 17, 31, 
    0, 0, 0, 0, 10, 40, 11, 16, 35, 20, 11, 14, 24, 25, 12, 
    0, 0, 0, 0, 0, 15, 30, 11, 34, 16, 0, 13, 17, 29, 21, 
    0, 0, 1, 11, 16, 13, 22, 26, 29, 23, 14, 14, 24, 33, 31, 
    10, 20, 25, 32, 36, 23, 18, 29, 37, 35, 36, 29, 29, 41, 38, 
    
    -- channel=480
    0, 0, 3, 8, 9, 16, 20, 10, 4, 5, 11, 9, 10, 11, 15, 
    0, 0, 1, 20, 10, 22, 23, 28, 27, 14, 22, 19, 17, 20, 28, 
    0, 0, 19, 6, 18, 20, 29, 43, 37, 11, 23, 37, 46, 49, 58, 
    0, 0, 22, 17, 0, 10, 26, 49, 67, 48, 25, 57, 56, 50, 60, 
    0, 0, 4, 36, 4, 0, 4, 36, 52, 51, 43, 47, 67, 85, 87, 
    6, 13, 26, 37, 5, 0, 13, 15, 29, 46, 51, 38, 79, 112, 106, 
    17, 24, 22, 42, 26, 12, 16, 18, 15, 26, 45, 32, 65, 92, 87, 
    6, 14, 23, 45, 45, 16, 35, 34, 8, 7, 28, 31, 33, 60, 67, 
    8, 15, 8, 29, 20, 49, 39, 51, 6, 0, 11, 21, 18, 53, 114, 
    0, 1, 37, 34, 31, 59, 43, 52, 1, 0, 5, 17, 21, 84, 127, 
    18, 30, 86, 41, 18, 45, 27, 47, 16, 13, 30, 26, 43, 85, 128, 
    39, 52, 31, 16, 20, 10, 12, 37, 13, 10, 8, 26, 84, 105, 126, 
    21, 17, 30, 31, 38, 23, 32, 35, 0, 0, 0, 14, 77, 122, 115, 
    29, 30, 49, 84, 102, 78, 64, 51, 45, 26, 12, 6, 58, 133, 129, 
    59, 92, 107, 115, 122, 101, 88, 123, 127, 97, 77, 82, 106, 138, 147, 
    
    -- channel=481
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=482
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 1, 5, 0, 0, 4, 0, 2, 0, 0, 0, 
    0, 2, 0, 0, 0, 6, 2, 5, 1, 3, 0, 0, 0, 0, 0, 
    5, 10, 12, 0, 0, 26, 10, 0, 2, 0, 4, 0, 0, 0, 0, 
    9, 3, 0, 0, 5, 26, 0, 0, 8, 0, 5, 5, 0, 0, 0, 
    0, 0, 0, 0, 10, 17, 0, 3, 13, 0, 0, 0, 0, 5, 0, 
    1, 1, 2, 0, 0, 0, 0, 6, 14, 0, 0, 0, 11, 0, 0, 
    8, 9, 5, 0, 17, 0, 21, 0, 8, 0, 0, 0, 8, 0, 0, 
    13, 16, 0, 0, 3, 10, 3, 0, 8, 1, 1, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 11, 1, 2, 0, 0, 3, 0, 
    0, 0, 0, 3, 0, 0, 15, 0, 14, 2, 5, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 20, 0, 5, 9, 12, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 6, 0, 7, 0, 7, 13, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 2, 6, 5, 0, 0, 0, 
    
    -- channel=483
    49, 46, 69, 64, 92, 111, 86, 67, 56, 62, 53, 45, 47, 60, 62, 
    47, 49, 73, 57, 115, 132, 132, 120, 79, 82, 97, 108, 112, 118, 112, 
    45, 51, 62, 76, 114, 144, 161, 186, 161, 129, 128, 142, 126, 118, 117, 
    58, 66, 88, 96, 110, 148, 178, 215, 209, 160, 135, 140, 137, 127, 150, 
    116, 130, 133, 79, 116, 155, 168, 175, 218, 206, 190, 176, 183, 206, 216, 
    124, 113, 94, 65, 128, 158, 127, 143, 192, 209, 215, 182, 213, 244, 218, 
    92, 98, 106, 86, 130, 131, 139, 163, 172, 166, 198, 182, 193, 201, 148, 
    100, 124, 132, 137, 140, 158, 181, 197, 168, 138, 169, 177, 168, 154, 164, 
    131, 156, 181, 145, 194, 182, 209, 182, 146, 126, 155, 164, 158, 157, 189, 
    187, 183, 122, 119, 138, 174, 176, 169, 144, 126, 155, 151, 144, 163, 227, 
    137, 128, 22, 102, 104, 126, 137, 152, 165, 146, 159, 159, 166, 222, 228, 
    35, 33, 71, 100, 88, 115, 157, 106, 134, 139, 155, 166, 192, 249, 232, 
    59, 62, 90, 122, 135, 134, 156, 139, 125, 133, 133, 137, 204, 252, 253, 
    102, 125, 134, 147, 174, 203, 167, 173, 157, 132, 115, 117, 178, 250, 256, 
    129, 154, 195, 218, 240, 236, 206, 229, 243, 218, 190, 191, 212, 260, 263, 
    
    -- channel=484
    0, 4, 1, 2, 6, 3, 9, 11, 16, 21, 26, 32, 37, 37, 39, 
    1, 4, 6, 16, 19, 25, 17, 19, 22, 18, 21, 24, 26, 24, 26, 
    6, 6, 26, 25, 29, 35, 36, 37, 23, 7, 6, 10, 17, 17, 24, 
    10, 3, 9, 42, 37, 34, 39, 40, 30, 16, 5, 9, 12, 20, 28, 
    0, 0, 0, 35, 46, 23, 14, 30, 39, 35, 29, 18, 9, 18, 24, 
    0, 0, 0, 35, 23, 13, 12, 23, 29, 38, 40, 24, 18, 13, 18, 
    0, 0, 0, 0, 43, 22, 20, 24, 16, 24, 36, 35, 22, 15, 19, 
    0, 0, 0, 0, 0, 20, 20, 29, 10, 12, 31, 37, 23, 17, 23, 
    0, 0, 0, 0, 0, 0, 0, 22, 10, 7, 22, 33, 27, 32, 37, 
    0, 0, 0, 0, 0, 0, 0, 16, 12, 8, 16, 30, 31, 37, 53, 
    0, 0, 0, 0, 3, 10, 23, 28, 18, 15, 16, 27, 37, 31, 50, 
    0, 0, 0, 0, 23, 40, 20, 22, 27, 20, 15, 15, 39, 34, 37, 
    0, 0, 0, 0, 17, 32, 25, 25, 28, 11, 0, 13, 28, 42, 33, 
    2, 9, 15, 24, 31, 29, 29, 39, 45, 34, 16, 20, 36, 48, 47, 
    24, 32, 41, 51, 48, 34, 38, 46, 53, 51, 47, 44, 48, 58, 55, 
    
    -- channel=485
    16, 8, 7, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    89, 107, 128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    104, 101, 104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    73, 79, 92, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 92, 114, 35, 92, 25, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    152, 201, 235, 211, 88, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    261, 268, 113, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    236, 183, 90, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 49, 35, 18, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=486
    144, 133, 152, 162, 173, 169, 142, 121, 100, 95, 73, 51, 30, 28, 17, 
    139, 128, 145, 120, 157, 173, 163, 130, 96, 97, 85, 81, 81, 93, 93, 
    128, 128, 119, 99, 123, 119, 141, 152, 140, 156, 166, 174, 159, 153, 131, 
    118, 124, 91, 69, 87, 107, 123, 168, 179, 196, 195, 183, 158, 142, 129, 
    180, 225, 230, 72, 87, 158, 177, 157, 172, 169, 186, 184, 191, 194, 187, 
    317, 337, 280, 75, 102, 172, 191, 157, 169, 171, 168, 172, 214, 246, 223, 
    314, 312, 297, 111, 141, 191, 184, 170, 184, 166, 166, 159, 191, 221, 181, 
    284, 307, 320, 281, 158, 137, 186, 191, 208, 183, 158, 143, 164, 156, 152, 
    324, 366, 388, 306, 345, 256, 256, 198, 199, 188, 163, 144, 152, 155, 170, 
    449, 515, 531, 425, 371, 329, 262, 201, 188, 190, 191, 154, 134, 123, 120, 
    573, 554, 321, 304, 232, 236, 178, 190, 203, 196, 197, 155, 132, 157, 129, 
    463, 386, 247, 221, 132, 106, 158, 102, 146, 160, 180, 179, 147, 202, 154, 
    231, 217, 214, 208, 180, 127, 182, 139, 126, 169, 211, 195, 156, 175, 202, 
    175, 187, 201, 187, 168, 173, 134, 161, 135, 159, 203, 163, 164, 164, 184, 
    170, 162, 150, 129, 145, 195, 165, 156, 139, 131, 136, 161, 148, 144, 150, 
    
    -- channel=487
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=488
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 5, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 0, 0, 0, 
    13, 28, 28, 0, 0, 0, 14, 9, 10, 5, 1, 4, 7, 12, 18, 
    20, 13, 0, 0, 0, 1, 0, 0, 8, 8, 11, 0, 7, 21, 18, 
    0, 0, 0, 15, 0, 0, 0, 0, 7, 7, 5, 3, 11, 7, 0, 
    1, 12, 16, 6, 32, 10, 11, 7, 12, 4, 2, 4, 0, 0, 0, 
    17, 27, 46, 57, 36, 39, 10, 17, 3, 0, 4, 3, 0, 0, 0, 
    67, 70, 33, 19, 0, 6, 2, 12, 1, 0, 3, 2, 0, 0, 0, 
    40, 33, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 7, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 8, 18, 
    0, 0, 0, 0, 2, 6, 0, 0, 0, 0, 11, 0, 13, 13, 7, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 5, 8, 
    0, 0, 0, 0, 6, 6, 6, 0, 4, 0, 0, 0, 0, 4, 9, 
    
    -- channel=489
    171, 153, 172, 168, 176, 201, 157, 129, 110, 97, 62, 32, 10, 12, 5, 
    164, 151, 161, 95, 172, 170, 188, 148, 92, 97, 96, 109, 124, 138, 123, 
    139, 139, 94, 96, 107, 126, 133, 157, 194, 230, 218, 211, 174, 148, 102, 
    133, 147, 109, 44, 93, 128, 149, 181, 183, 189, 221, 181, 159, 136, 121, 
    288, 369, 344, 72, 106, 213, 261, 191, 193, 183, 194, 216, 206, 205, 205, 
    413, 411, 323, 70, 148, 225, 213, 195, 210, 193, 192, 190, 218, 248, 221, 
    356, 349, 344, 183, 114, 191, 215, 199, 237, 207, 184, 185, 212, 207, 148, 
    346, 382, 389, 333, 262, 182, 224, 226, 278, 239, 186, 173, 185, 145, 148, 
    416, 481, 559, 443, 489, 355, 309, 232, 246, 236, 214, 183, 182, 164, 105, 
    675, 729, 617, 533, 378, 367, 260, 238, 242, 242, 246, 196, 161, 89, 63, 
    708, 658, 272, 218, 221, 183, 192, 174, 242, 234, 214, 181, 147, 169, 91, 
    440, 305, 281, 260, 124, 97, 203, 107, 123, 181, 240, 223, 133, 176, 145, 
    214, 210, 201, 229, 219, 175, 176, 160, 159, 237, 299, 228, 188, 141, 178, 
    172, 204, 188, 119, 91, 161, 128, 143, 126, 142, 180, 185, 158, 113, 131, 
    136, 79, 75, 77, 98, 168, 153, 101, 87, 93, 89, 102, 91, 84, 89, 
    
    -- channel=490
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=491
    0, 0, 0, 30, 21, 0, 0, 2, 0, 0, 12, 13, 0, 0, 0, 
    0, 0, 5, 26, 0, 54, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    9, 0, 66, 47, 9, 0, 4, 0, 0, 0, 0, 0, 0, 23, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 63, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 2, 
    43, 35, 0, 0, 42, 95, 0, 0, 0, 0, 0, 0, 7, 72, 84, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 122, 
    0, 0, 102, 23, 86, 11, 14, 0, 0, 0, 0, 0, 0, 22, 30, 
    0, 44, 170, 200, 146, 163, 65, 73, 0, 0, 0, 0, 0, 0, 0, 
    364, 326, 57, 0, 0, 12, 0, 0, 34, 0, 0, 0, 0, 33, 0, 
    129, 99, 47, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 26, 19, 
    8, 0, 74, 153, 115, 0, 0, 14, 21, 91, 119, 0, 8, 49, 71, 
    100, 150, 86, 28, 36, 29, 7, 38, 27, 12, 51, 92, 54, 49, 63, 
    
    -- channel=492
    0, 5, 0, 8, 0, 0, 16, 8, 12, 4, 11, 14, 14, 12, 26, 
    0, 5, 0, 19, 0, 0, 0, 6, 23, 12, 26, 30, 34, 37, 44, 
    0, 0, 17, 0, 0, 0, 0, 0, 6, 22, 28, 34, 44, 42, 47, 
    0, 0, 53, 6, 0, 0, 0, 0, 0, 0, 0, 40, 42, 48, 54, 
    10, 13, 55, 66, 0, 0, 0, 16, 0, 0, 0, 4, 46, 76, 77, 
    12, 13, 54, 81, 0, 0, 0, 0, 0, 0, 0, 0, 36, 79, 84, 
    8, 16, 26, 138, 0, 0, 0, 0, 0, 2, 0, 0, 25, 39, 63, 
    5, 17, 31, 49, 116, 14, 22, 0, 0, 0, 0, 0, 0, 22, 57, 
    9, 17, 45, 109, 27, 86, 4, 26, 0, 0, 0, 0, 0, 32, 84, 
    33, 34, 45, 66, 0, 39, 0, 33, 0, 0, 0, 0, 0, 72, 93, 
    29, 46, 142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 61, 113, 
    10, 12, 53, 17, 31, 0, 0, 52, 0, 0, 0, 1, 59, 43, 122, 
    6, 1, 15, 25, 45, 38, 0, 14, 0, 0, 0, 0, 64, 73, 58, 
    15, 19, 27, 50, 54, 44, 39, 11, 3, 0, 0, 0, 27, 86, 66, 
    40, 52, 61, 84, 72, 44, 61, 90, 79, 50, 23, 27, 65, 90, 89, 
    
    -- channel=493
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=494
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 8, 0, 0, 17, 0, 0, 0, 0, 0, 0, 5, 9, 0, 
    0, 0, 0, 11, 0, 2, 7, 6, 24, 14, 0, 0, 0, 0, 0, 
    0, 5, 0, 4, 3, 9, 11, 14, 8, 19, 6, 0, 0, 0, 0, 
    37, 40, 0, 0, 8, 54, 11, 0, 0, 3, 19, 0, 9, 0, 0, 
    24, 6, 0, 0, 1, 75, 0, 0, 6, 0, 0, 23, 23, 0, 0, 
    0, 0, 0, 0, 17, 43, 0, 3, 21, 0, 0, 32, 0, 5, 0, 
    12, 15, 0, 0, 0, 49, 0, 21, 26, 0, 0, 1, 5, 3, 0, 
    29, 44, 13, 0, 0, 0, 9, 0, 23, 0, 0, 0, 24, 0, 0, 
    54, 42, 0, 0, 4, 0, 28, 0, 19, 2, 0, 0, 5, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 39, 0, 24, 20, 12, 0, 0, 34, 0, 
    0, 0, 0, 0, 0, 0, 31, 0, 21, 56, 2, 0, 0, 5, 2, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 28, 12, 0, 0, 0, 14, 
    0, 0, 0, 0, 19, 16, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    
    -- channel=495
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=496
    77, 68, 83, 72, 69, 62, 46, 58, 49, 45, 38, 29, 25, 32, 25, 
    75, 66, 70, 61, 43, 44, 38, 29, 36, 52, 45, 48, 49, 51, 42, 
    67, 67, 35, 46, 26, 16, 12, 20, 48, 69, 65, 60, 53, 48, 35, 
    64, 72, 44, 17, 18, 19, 17, 14, 9, 52, 65, 42, 56, 46, 37, 
    118, 131, 57, 1, 10, 64, 46, 6, 9, 7, 29, 39, 61, 51, 44, 
    140, 137, 77, 7, 34, 74, 37, 21, 26, 8, 0, 31, 56, 57, 45, 
    131, 127, 125, 6, 35, 60, 24, 28, 44, 23, 2, 25, 31, 56, 36, 
    132, 140, 115, 112, 24, 69, 30, 34, 54, 32, 9, 2, 30, 43, 48, 
    148, 179, 193, 99, 124, 45, 86, 16, 52, 44, 23, 3, 33, 26, 3, 
    221, 219, 173, 105, 124, 62, 84, 17, 46, 52, 38, 3, 15, 0, 6, 
    236, 192, 44, 88, 58, 41, 35, 38, 40, 39, 27, 11, 10, 30, 0, 
    135, 131, 93, 67, 7, 18, 62, 0, 40, 48, 53, 28, 0, 45, 1, 
    89, 85, 91, 82, 50, 20, 38, 28, 36, 72, 63, 40, 5, 14, 41, 
    76, 70, 47, 25, 32, 44, 24, 19, 9, 26, 55, 35, 10, 6, 19, 
    32, 20, 19, 5, 23, 38, 19, 4, 0, 3, 10, 9, 0, 0, 0, 
    
    -- channel=497
    93, 89, 89, 84, 115, 153, 120, 105, 96, 94, 86, 82, 85, 90, 99, 
    91, 95, 93, 87, 153, 156, 186, 167, 114, 113, 129, 144, 152, 144, 133, 
    85, 92, 72, 109, 162, 199, 205, 221, 204, 169, 152, 146, 118, 98, 93, 
    100, 107, 130, 130, 191, 213, 230, 237, 209, 163, 163, 139, 117, 116, 135, 
    176, 194, 173, 147, 184, 213, 239, 233, 249, 236, 218, 204, 160, 166, 172, 
    133, 113, 133, 123, 200, 210, 187, 222, 238, 246, 247, 216, 173, 161, 143, 
    84, 88, 124, 152, 116, 146, 206, 228, 226, 224, 240, 226, 179, 129, 93, 
    118, 133, 126, 166, 217, 184, 209, 229, 229, 221, 237, 230, 200, 145, 142, 
    143, 163, 221, 178, 222, 185, 206, 220, 208, 212, 239, 242, 213, 157, 107, 
    215, 178, 82, 151, 127, 178, 164, 223, 217, 213, 233, 241, 204, 141, 134, 
    109, 89, 25, 72, 119, 143, 167, 168, 213, 205, 204, 228, 200, 188, 148, 
    0, 0, 96, 138, 138, 174, 197, 140, 159, 196, 213, 221, 185, 163, 169, 
    60, 68, 85, 121, 166, 172, 153, 184, 198, 212, 209, 200, 216, 162, 172, 
    105, 123, 112, 91, 105, 159, 160, 168, 173, 134, 141, 188, 180, 161, 143, 
    94, 87, 121, 142, 142, 154, 157, 154, 161, 163, 147, 141, 153, 151, 144, 
    
    -- channel=498
    0, 1, 0, 10, 0, 0, 16, 8, 6, 1, 16, 23, 13, 0, 0, 
    0, 1, 0, 20, 0, 0, 8, 5, 20, 0, 0, 0, 0, 0, 0, 
    0, 0, 38, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 15, 32, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 28, 1, 14, 5, 
    0, 0, 7, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 104, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 6, 14, 93, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 52, 
    0, 0, 0, 26, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 8, 0, 0, 0, 0, 0, 0, 69, 
    0, 0, 44, 132, 9, 90, 0, 41, 0, 0, 0, 7, 0, 48, 18, 
    0, 44, 266, 78, 22, 75, 0, 10, 0, 0, 3, 1, 0, 0, 30, 
    148, 148, 75, 29, 60, 0, 0, 36, 0, 0, 0, 0, 27, 0, 47, 
    52, 30, 16, 0, 28, 0, 0, 16, 0, 0, 0, 0, 17, 0, 0, 
    0, 0, 25, 70, 43, 0, 0, 3, 2, 0, 4, 3, 16, 19, 0, 
    41, 63, 35, 22, 0, 0, 7, 36, 18, 2, 0, 17, 41, 7, 14, 
    
    -- channel=499
    110, 112, 109, 104, 155, 179, 146, 126, 118, 126, 125, 124, 126, 122, 122, 
    111, 113, 114, 144, 188, 231, 230, 204, 145, 131, 134, 128, 121, 108, 108, 
    118, 117, 122, 167, 237, 273, 291, 294, 209, 130, 130, 127, 119, 112, 122, 
    126, 120, 117, 182, 275, 282, 290, 297, 283, 220, 185, 166, 120, 117, 133, 
    99, 86, 87, 192, 261, 252, 249, 283, 314, 310, 288, 237, 147, 132, 138, 
    76, 79, 92, 163, 227, 236, 257, 286, 289, 308, 319, 290, 190, 140, 130, 
    83, 84, 89, 110, 175, 232, 268, 289, 264, 269, 306, 304, 226, 151, 126, 
    95, 86, 87, 118, 119, 166, 221, 276, 265, 261, 300, 309, 257, 183, 136, 
    89, 75, 61, 95, 125, 122, 177, 256, 273, 265, 290, 308, 277, 198, 148, 
    26, 12, 31, 95, 158, 153, 195, 264, 277, 267, 279, 307, 282, 193, 147, 
    10, 18, 106, 185, 222, 260, 252, 253, 276, 268, 270, 298, 260, 174, 142, 
    63, 91, 106, 132, 206, 280, 232, 187, 260, 273, 244, 256, 230, 176, 155, 
    115, 112, 115, 119, 139, 172, 212, 221, 247, 256, 221, 253, 233, 182, 168, 
    128, 126, 143, 154, 162, 158, 184, 208, 237, 235, 241, 260, 241, 192, 172, 
    134, 153, 167, 164, 160, 159, 177, 182, 186, 193, 203, 206, 201, 179, 166, 
    
    -- channel=500
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=501
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 8, 0, 15, 
    0, 0, 0, 7, 0, 0, 12, 0, 7, 0, 1, 0, 0, 0, 2, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 37, 
    0, 0, 71, 0, 0, 0, 0, 0, 0, 0, 0, 26, 16, 30, 31, 
    0, 0, 27, 100, 0, 0, 0, 7, 0, 0, 0, 0, 0, 35, 25, 
    0, 0, 143, 83, 0, 0, 0, 10, 0, 0, 0, 0, 0, 31, 44, 
    0, 0, 30, 182, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 0, 64, 152, 0, 1, 0, 0, 2, 3, 0, 0, 0, 31, 
    0, 0, 0, 1, 13, 56, 0, 10, 0, 0, 0, 0, 0, 0, 77, 
    0, 0, 0, 177, 0, 121, 0, 64, 0, 0, 0, 4, 0, 70, 70, 
    0, 11, 256, 31, 0, 40, 0, 7, 0, 0, 0, 10, 0, 38, 71, 
    44, 91, 109, 32, 60, 0, 0, 39, 0, 0, 0, 0, 39, 0, 123, 
    21, 0, 9, 0, 56, 0, 0, 45, 0, 0, 0, 0, 65, 8, 36, 
    0, 0, 0, 52, 54, 28, 3, 0, 0, 0, 0, 0, 18, 58, 5, 
    17, 56, 60, 61, 5, 0, 30, 76, 52, 24, 0, 5, 69, 45, 53, 
    
    -- channel=502
    69, 60, 41, 47, 0, 0, 0, 25, 39, 28, 22, 23, 14, 4, 7, 
    68, 65, 38, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 
    53, 53, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 38, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 84, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    77, 80, 127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 70, 81, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 59, 60, 17, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 58, 107, 44, 45, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    148, 162, 126, 147, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    176, 179, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    125, 82, 72, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 35, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=503
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=504
    0, 4, 0, 0, 6, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 
    0, 1, 0, 14, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 5, 13, 5, 6, 4, 2, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 11, 9, 4, 7, 4, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 31, 13, 0, 1, 20, 2, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 0, 0, 8, 16, 1, 10, 5, 0, 0, 0, 0, 
    0, 0, 0, 35, 3, 5, 8, 4, 0, 13, 1, 9, 8, 0, 0, 
    0, 0, 1, 0, 0, 5, 7, 4, 0, 10, 10, 10, 0, 0, 0, 
    0, 0, 0, 40, 0, 11, 0, 16, 0, 6, 9, 6, 0, 12, 4, 
    0, 0, 10, 0, 0, 0, 0, 16, 0, 6, 6, 11, 10, 11, 0, 
    0, 0, 51, 0, 18, 0, 17, 6, 2, 9, 6, 8, 9, 0, 0, 
    14, 1, 13, 0, 22, 10, 0, 25, 0, 1, 0, 6, 10, 0, 4, 
    4, 2, 0, 0, 0, 19, 0, 0, 3, 2, 0, 12, 11, 0, 0, 
    0, 1, 6, 7, 0, 0, 4, 0, 10, 15, 0, 13, 11, 0, 0, 
    8, 4, 0, 1, 0, 0, 8, 4, 0, 0, 2, 3, 3, 2, 0, 
    
    -- channel=505
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=506
    73, 72, 78, 68, 64, 68, 65, 81, 83, 84, 92, 97, 104, 110, 108, 
    74, 73, 75, 80, 63, 68, 67, 74, 87, 89, 90, 91, 93, 91, 88, 
    76, 78, 70, 93, 71, 75, 70, 69, 89, 73, 68, 66, 71, 72, 77, 
    81, 82, 75, 82, 83, 77, 73, 65, 63, 69, 63, 59, 76, 73, 80, 
    70, 56, 17, 76, 82, 86, 61, 51, 60, 62, 63, 65, 71, 64, 66, 
    32, 22, 14, 67, 85, 74, 46, 54, 64, 58, 60, 71, 65, 57, 56, 
    29, 29, 33, 38, 67, 78, 54, 64, 64, 53, 57, 73, 59, 66, 63, 
    39, 33, 16, 47, 48, 73, 48, 62, 60, 46, 56, 65, 70, 77, 73, 
    33, 27, 8, 0, 15, 12, 50, 44, 60, 49, 54, 59, 75, 67, 70, 
    0, 0, 0, 0, 16, 9, 49, 40, 60, 53, 50, 52, 72, 72, 90, 
    0, 0, 0, 14, 37, 42, 56, 65, 57, 54, 54, 56, 71, 80, 77, 
    0, 3, 28, 51, 48, 79, 84, 65, 73, 70, 60, 52, 65, 80, 65, 
    43, 56, 57, 56, 63, 72, 74, 67, 77, 78, 46, 44, 59, 73, 77, 
    67, 63, 56, 64, 80, 75, 80, 66, 79, 73, 66, 59, 56, 79, 79, 
    66, 75, 82, 83, 91, 77, 67, 76, 85, 85, 86, 78, 78, 85, 86, 
    
    -- channel=507
    94, 79, 109, 103, 100, 99, 74, 59, 38, 26, 3, 0, 0, 0, 0, 
    88, 73, 89, 56, 63, 72, 64, 44, 27, 32, 29, 34, 41, 56, 45, 
    70, 67, 33, 25, 9, 6, 12, 37, 82, 122, 119, 120, 101, 85, 52, 
    60, 74, 34, 0, 0, 0, 17, 48, 64, 101, 124, 100, 101, 76, 60, 
    184, 240, 175, 0, 0, 74, 95, 44, 46, 45, 71, 93, 134, 133, 126, 
    307, 312, 185, 0, 18, 104, 81, 44, 58, 44, 34, 63, 145, 179, 152, 
    279, 274, 251, 63, 45, 89, 59, 54, 88, 62, 31, 53, 105, 144, 94, 
    260, 293, 284, 232, 100, 104, 87, 86, 116, 77, 31, 23, 56, 77, 89, 
    314, 381, 420, 315, 314, 202, 185, 89, 100, 82, 52, 17, 48, 73, 57, 
    519, 570, 506, 347, 287, 207, 179, 89, 88, 92, 84, 24, 26, 20, 31, 
    595, 536, 214, 165, 127, 86, 76, 70, 90, 90, 74, 29, 28, 81, 44, 
    373, 285, 197, 137, 13, 0, 82, 13, 28, 62, 98, 73, 39, 120, 68, 
    161, 149, 153, 158, 104, 53, 74, 40, 31, 103, 133, 90, 63, 85, 112, 
    115, 131, 114, 75, 66, 89, 51, 47, 19, 49, 75, 52, 47, 60, 87, 
    78, 49, 43, 34, 68, 104, 76, 50, 32, 25, 25, 37, 26, 46, 49, 
    
    -- channel=508
    257, 239, 254, 258, 300, 318, 245, 214, 183, 174, 136, 100, 70, 59, 39, 
    251, 235, 247, 194, 301, 332, 337, 260, 168, 167, 142, 137, 140, 150, 141, 
    233, 231, 185, 215, 260, 284, 310, 319, 279, 280, 275, 268, 229, 209, 168, 
    218, 225, 145, 125, 259, 278, 291, 334, 331, 334, 350, 281, 215, 189, 169, 
    310, 385, 382, 159, 248, 367, 392, 338, 357, 349, 368, 349, 272, 239, 234, 
    492, 512, 424, 131, 258, 359, 383, 373, 367, 353, 355, 359, 315, 298, 263, 
    475, 463, 442, 196, 217, 377, 400, 375, 386, 355, 348, 354, 333, 289, 218, 
    448, 465, 480, 418, 266, 225, 333, 374, 440, 403, 355, 339, 336, 239, 196, 
    504, 549, 582, 459, 581, 404, 418, 360, 425, 416, 381, 351, 340, 270, 183, 
    689, 780, 756, 692, 565, 503, 404, 388, 418, 426, 420, 372, 324, 179, 83, 
    831, 796, 430, 436, 431, 410, 372, 348, 420, 416, 392, 353, 279, 219, 95, 
    678, 533, 397, 371, 251, 271, 330, 197, 299, 352, 380, 370, 233, 244, 166, 
    354, 341, 310, 315, 291, 252, 313, 278, 301, 394, 443, 397, 288, 196, 235, 
    264, 287, 298, 239, 185, 223, 202, 261, 258, 307, 386, 367, 295, 177, 186, 
    235, 186, 156, 119, 134, 230, 225, 167, 136, 159, 190, 222, 182, 125, 120, 
    
    -- channel=509
    163, 156, 149, 170, 201, 225, 187, 146, 125, 116, 95, 72, 49, 30, 24, 
    159, 155, 154, 136, 221, 245, 257, 206, 135, 109, 98, 86, 83, 82, 87, 
    151, 150, 145, 132, 215, 233, 259, 262, 200, 175, 181, 181, 159, 149, 130, 
    141, 138, 116, 107, 208, 229, 242, 278, 274, 257, 246, 227, 154, 137, 124, 
    166, 209, 281, 153, 199, 239, 287, 295, 303, 292, 293, 276, 193, 173, 170, 
    297, 327, 343, 144, 185, 232, 313, 311, 296, 302, 309, 286, 238, 220, 206, 
    308, 305, 297, 193, 169, 249, 319, 298, 295, 297, 306, 279, 270, 217, 186, 
    280, 289, 322, 289, 223, 144, 266, 286, 323, 326, 307, 289, 271, 191, 148, 
    306, 324, 357, 336, 383, 315, 283, 302, 320, 330, 314, 306, 267, 221, 170, 
    395, 462, 513, 518, 399, 413, 286, 333, 317, 325, 330, 325, 269, 185, 90, 
    527, 542, 406, 357, 334, 344, 295, 281, 315, 324, 317, 307, 244, 172, 111, 
    487, 402, 300, 268, 230, 227, 230, 186, 232, 272, 285, 301, 228, 176, 163, 
    256, 230, 212, 212, 219, 181, 218, 232, 221, 265, 322, 321, 259, 170, 182, 
    180, 189, 217, 199, 152, 167, 160, 214, 205, 229, 286, 291, 266, 166, 150, 
    179, 159, 138, 117, 104, 165, 182, 160, 132, 141, 152, 187, 172, 124, 118, 
    
    -- channel=510
    36, 30, 28, 46, 29, 26, 26, 12, 6, 0, 0, 0, 0, 0, 0, 
    32, 30, 24, 0, 14, 0, 8, 0, 0, 0, 0, 0, 0, 1, 4, 
    19, 21, 14, 0, 0, 0, 0, 0, 0, 37, 46, 46, 35, 33, 14, 
    9, 14, 24, 0, 0, 0, 0, 0, 0, 1, 33, 42, 30, 27, 10, 
    65, 106, 153, 0, 0, 0, 11, 0, 0, 0, 0, 10, 41, 52, 43, 
    159, 173, 188, 0, 0, 0, 15, 0, 0, 0, 0, 0, 28, 69, 64, 
    153, 154, 157, 92, 0, 0, 16, 0, 0, 2, 0, 0, 14, 38, 43, 
    131, 149, 169, 136, 108, 0, 33, 0, 9, 28, 0, 0, 0, 0, 24, 
    157, 187, 238, 194, 194, 149, 78, 23, 0, 22, 0, 0, 0, 6, 25, 
    282, 328, 329, 302, 151, 181, 54, 38, 0, 14, 14, 0, 0, 0, 0, 
    365, 369, 220, 98, 44, 32, 0, 0, 2, 11, 12, 0, 0, 12, 1, 
    267, 198, 139, 94, 16, 0, 0, 0, 0, 0, 7, 20, 0, 4, 31, 
    89, 75, 71, 71, 65, 15, 0, 1, 0, 0, 50, 30, 18, 0, 19, 
    40, 48, 51, 32, 1, 16, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    33, 8, 0, 0, 0, 11, 12, 2, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=511
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=512
    11, 136, 200, 156, 146, 186, 177, 182, 129, 38, 163, 184, 192, 199, 193, 
    14, 78, 209, 157, 116, 123, 168, 182, 159, 58, 191, 186, 186, 193, 191, 
    17, 35, 204, 148, 145, 64, 102, 151, 139, 129, 174, 195, 183, 187, 183, 
    8, 79, 183, 140, 166, 104, 76, 75, 99, 153, 163, 207, 173, 168, 209, 
    152, 176, 178, 112, 156, 135, 116, 73, 101, 133, 180, 226, 195, 169, 219, 
    186, 186, 188, 135, 158, 132, 100, 80, 95, 119, 157, 241, 210, 181, 212, 
    199, 188, 156, 173, 119, 120, 89, 120, 106, 128, 148, 234, 219, 201, 187, 
    193, 188, 101, 207, 133, 127, 108, 87, 153, 144, 144, 228, 252, 207, 216, 
    173, 173, 133, 163, 151, 138, 101, 75, 160, 128, 150, 108, 199, 196, 252, 
    192, 175, 165, 154, 164, 158, 149, 113, 88, 151, 132, 151, 136, 144, 176, 
    204, 159, 184, 159, 166, 120, 167, 152, 138, 125, 139, 148, 144, 122, 133, 
    205, 167, 195, 164, 154, 139, 164, 153, 141, 103, 158, 139, 151, 124, 113, 
    199, 195, 209, 158, 113, 115, 175, 161, 138, 114, 153, 131, 135, 137, 122, 
    193, 191, 216, 175, 130, 121, 145, 147, 127, 117, 139, 125, 104, 138, 139, 
    186, 191, 193, 180, 146, 138, 127, 141, 101, 126, 127, 129, 111, 130, 137, 
    
    -- channel=513
    42, 8, 108, 98, 89, 91, 90, 76, 82, 72, 33, 86, 104, 94, 103, 
    41, 16, 105, 91, 81, 74, 100, 82, 107, 118, 1, 76, 90, 97, 111, 
    45, 35, 45, 72, 103, 115, 93, 112, 133, 72, 30, 63, 81, 79, 76, 
    0, 0, 0, 85, 103, 117, 69, 77, 75, 54, 93, 58, 98, 100, 65, 
    55, 7, 53, 76, 68, 110, 123, 113, 83, 63, 74, 47, 81, 63, 24, 
    59, 51, 67, 69, 80, 110, 124, 88, 73, 57, 66, 53, 61, 43, 4, 
    45, 52, 97, 94, 71, 74, 112, 82, 90, 64, 61, 51, 60, 57, 5, 
    46, 69, 145, 98, 97, 90, 107, 100, 98, 64, 95, 101, 83, 86, 35, 
    45, 46, 131, 84, 95, 76, 77, 121, 59, 86, 106, 59, 62, 108, 44, 
    37, 29, 91, 94, 77, 118, 121, 87, 60, 86, 113, 101, 66, 90, 68, 
    42, 53, 71, 80, 83, 98, 87, 106, 122, 118, 87, 79, 96, 104, 96, 
    43, 59, 49, 106, 120, 130, 84, 98, 110, 112, 61, 94, 105, 100, 87, 
    40, 40, 30, 95, 144, 124, 119, 109, 123, 104, 79, 91, 111, 103, 86, 
    44, 30, 5, 85, 112, 101, 113, 108, 113, 79, 77, 84, 95, 70, 89, 
    49, 28, 3, 86, 93, 110, 120, 108, 106, 62, 77, 85, 77, 74, 88, 
    
    -- channel=514
    45, 131, 249, 239, 221, 227, 241, 243, 250, 157, 207, 291, 295, 281, 278, 
    48, 87, 211, 242, 273, 225, 230, 261, 262, 183, 284, 291, 290, 287, 287, 
    54, 63, 191, 254, 310, 236, 175, 177, 180, 217, 280, 251, 284, 296, 297, 
    176, 185, 275, 204, 289, 283, 263, 209, 192, 249, 266, 305, 341, 277, 258, 
    227, 273, 245, 183, 275, 281, 262, 196, 193, 231, 259, 315, 308, 215, 210, 
    240, 244, 226, 216, 280, 269, 235, 193, 232, 248, 254, 293, 289, 217, 177, 
    224, 232, 197, 261, 248, 245, 235, 242, 252, 244, 252, 305, 292, 283, 225, 
    203, 230, 244, 316, 272, 267, 241, 253, 233, 224, 231, 185, 274, 267, 243, 
    193, 204, 299, 329, 293, 329, 296, 236, 215, 221, 242, 202, 179, 171, 226, 
    215, 231, 288, 288, 265, 263, 287, 291, 261, 251, 214, 222, 248, 232, 206, 
    237, 211, 268, 297, 294, 247, 255, 277, 260, 225, 197, 248, 259, 218, 202, 
    232, 200, 268, 306, 298, 262, 292, 287, 263, 192, 229, 227, 254, 228, 204, 
    217, 174, 233, 292, 250, 239, 277, 252, 223, 185, 211, 206, 203, 200, 211, 
    204, 154, 186, 282, 266, 323, 250, 215, 188, 163, 199, 198, 176, 200, 222, 
    161, 154, 152, 271, 266, 245, 182, 197, 162, 169, 184, 199, 193, 203, 201, 
    
    -- channel=515
    0, 0, 58, 24, 24, 26, 30, 34, 14, 0, 10, 99, 80, 74, 68, 
    0, 0, 52, 24, 72, 35, 49, 72, 80, 0, 101, 116, 102, 98, 89, 
    0, 0, 23, 41, 135, 35, 0, 27, 10, 0, 127, 119, 125, 126, 115, 
    0, 0, 108, 22, 129, 84, 28, 0, 0, 68, 115, 162, 171, 136, 124, 
    36, 89, 97, 0, 111, 117, 84, 0, 0, 46, 105, 186, 169, 70, 93, 
    90, 94, 92, 21, 109, 104, 53, 0, 33, 57, 96, 184, 169, 81, 55, 
    85, 85, 47, 81, 68, 70, 53, 39, 57, 71, 90, 185, 178, 148, 72, 
    73, 88, 30, 131, 97, 96, 57, 66, 57, 57, 77, 89, 158, 158, 116, 
    58, 57, 85, 127, 122, 142, 104, 38, 42, 22, 74, 0, 64, 62, 121, 
    81, 72, 126, 107, 123, 135, 129, 87, 49, 69, 34, 26, 30, 46, 57, 
    112, 71, 124, 129, 127, 75, 113, 118, 88, 47, 0, 52, 69, 18, 16, 
    111, 62, 134, 152, 142, 72, 116, 106, 95, 0, 41, 41, 75, 30, 0, 
    94, 49, 104, 143, 101, 19, 115, 84, 48, 0, 31, 16, 31, 8, 12, 
    77, 26, 66, 144, 86, 82, 65, 37, 0, 0, 13, 3, 0, 6, 29, 
    32, 21, 26, 141, 106, 81, 0, 5, 0, 0, 0, 6, 0, 10, 12, 
    
    -- channel=516
    9, 40, 118, 112, 120, 120, 128, 126, 118, 97, 69, 143, 141, 147, 142, 
    10, 35, 97, 94, 119, 135, 123, 141, 141, 88, 117, 171, 163, 157, 149, 
    11, 22, 69, 117, 121, 137, 96, 102, 101, 88, 165, 174, 177, 176, 175, 
    90, 51, 152, 146, 113, 132, 124, 100, 81, 104, 156, 170, 186, 193, 177, 
    157, 170, 176, 136, 116, 138, 137, 106, 86, 101, 145, 198, 207, 200, 189, 
    178, 174, 181, 144, 133, 140, 127, 88, 104, 110, 146, 192, 221, 219, 201, 
    192, 174, 157, 133, 138, 119, 127, 97, 126, 126, 142, 194, 218, 216, 209, 
    196, 166, 126, 108, 156, 146, 115, 135, 111, 134, 149, 150, 184, 219, 206, 
    201, 153, 112, 135, 154, 162, 153, 121, 108, 125, 132, 129, 126, 153, 180, 
    202, 176, 158, 157, 163, 160, 147, 138, 154, 124, 124, 105, 114, 130, 140, 
    202, 190, 153, 168, 169, 159, 139, 147, 142, 139, 95, 118, 127, 113, 112, 
    203, 190, 160, 168, 171, 131, 149, 148, 150, 111, 113, 120, 122, 123, 103, 
    202, 191, 171, 168, 157, 79, 134, 143, 128, 107, 109, 110, 110, 98, 109, 
    196, 190, 171, 170, 148, 127, 132, 122, 108, 86, 103, 105, 94, 94, 110, 
    172, 176, 163, 155, 163, 154, 116, 98, 91, 87, 95, 102, 94, 105, 102, 
    
    -- channel=517
    0, 0, 0, 23, 13, 0, 12, 1, 56, 84, 0, 0, 14, 11, 17, 
    0, 0, 0, 0, 33, 36, 0, 0, 28, 124, 0, 29, 35, 24, 26, 
    0, 0, 0, 0, 0, 117, 14, 0, 10, 10, 0, 9, 40, 37, 45, 
    82, 0, 0, 50, 0, 86, 77, 52, 0, 0, 18, 0, 52, 64, 6, 
    77, 0, 28, 96, 0, 30, 65, 85, 0, 0, 0, 0, 54, 96, 0, 
    37, 17, 34, 65, 0, 33, 68, 54, 10, 0, 0, 0, 52, 101, 23, 
    38, 25, 53, 0, 34, 17, 72, 6, 46, 1, 0, 0, 38, 74, 75, 
    50, 15, 92, 0, 64, 33, 59, 35, 0, 12, 21, 0, 0, 56, 32, 
    79, 10, 48, 0, 48, 53, 71, 101, 0, 40, 17, 45, 0, 7, 0, 
    68, 33, 19, 40, 16, 23, 39, 78, 73, 0, 42, 1, 7, 22, 0, 
    43, 67, 0, 40, 39, 81, 0, 21, 66, 51, 6, 0, 9, 43, 11, 
    33, 78, 0, 41, 50, 64, 6, 30, 43, 83, 0, 18, 3, 41, 35, 
    41, 51, 0, 38, 84, 6, 0, 25, 46, 46, 0, 17, 4, 9, 20, 
    47, 47, 0, 21, 91, 30, 30, 17, 31, 17, 0, 9, 31, 0, 5, 
    35, 30, 0, 0, 59, 51, 49, 0, 38, 0, 0, 0, 23, 0, 0, 
    
    -- channel=518
    48, 127, 144, 137, 138, 147, 148, 152, 139, 93, 143, 164, 163, 162, 158, 
    49, 93, 140, 138, 138, 136, 135, 150, 140, 79, 181, 166, 167, 164, 160, 
    50, 65, 149, 150, 149, 107, 111, 116, 108, 124, 173, 158, 162, 168, 169, 
    105, 128, 178, 124, 153, 124, 127, 114, 114, 150, 142, 174, 168, 146, 157, 
    127, 166, 150, 110, 158, 140, 123, 96, 110, 138, 149, 186, 167, 134, 157, 
    146, 152, 141, 124, 151, 134, 115, 103, 122, 139, 149, 182, 169, 140, 148, 
    151, 150, 123, 138, 142, 137, 114, 128, 125, 137, 146, 184, 170, 161, 157, 
    141, 147, 113, 170, 137, 138, 117, 123, 122, 134, 126, 134, 164, 155, 156, 
    132, 144, 143, 175, 144, 160, 145, 109, 144, 122, 127, 120, 147, 117, 161, 
    143, 150, 158, 148, 152, 139, 136, 139, 138, 138, 121, 126, 140, 130, 143, 
    154, 135, 156, 159, 153, 129, 147, 142, 126, 120, 117, 143, 141, 120, 118, 
    154, 126, 166, 155, 148, 126, 154, 148, 134, 102, 141, 129, 135, 121, 115, 
    148, 130, 160, 153, 122, 127, 143, 138, 118, 104, 130, 120, 118, 115, 121, 
    140, 126, 153, 156, 132, 152, 135, 123, 107, 106, 125, 118, 102, 127, 125, 
    125, 126, 138, 153, 140, 131, 104, 115, 95, 112, 117, 117, 113, 123, 122, 
    
    -- channel=519
    0, 0, 0, 9, 0, 0, 0, 0, 17, 74, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 1, 84, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 62, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 39, 0, 21, 31, 21, 0, 0, 0, 0, 0, 17, 0, 
    30, 0, 0, 69, 0, 0, 20, 52, 0, 0, 0, 0, 0, 47, 0, 
    2, 0, 0, 39, 0, 0, 20, 26, 0, 0, 0, 0, 0, 43, 1, 
    3, 0, 34, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 6, 28, 
    19, 0, 57, 0, 22, 0, 14, 10, 0, 3, 0, 0, 0, 4, 0, 
    34, 0, 0, 0, 0, 0, 19, 37, 0, 19, 0, 23, 0, 0, 0, 
    17, 8, 0, 0, 0, 0, 0, 13, 34, 0, 12, 0, 0, 0, 0, 
    0, 33, 0, 0, 0, 32, 0, 0, 15, 24, 0, 0, 0, 17, 3, 
    0, 32, 0, 0, 1, 30, 0, 0, 5, 49, 0, 0, 0, 17, 10, 
    2, 18, 0, 0, 32, 7, 0, 0, 17, 30, 0, 3, 0, 0, 0, 
    12, 19, 0, 0, 30, 7, 0, 0, 18, 11, 0, 0, 16, 0, 0, 
    12, 0, 0, 0, 11, 15, 36, 0, 25, 0, 0, 0, 4, 0, 0, 
    
    -- channel=520
    5, 89, 364, 360, 361, 368, 387, 389, 383, 238, 230, 447, 446, 447, 438, 
    7, 48, 298, 321, 405, 386, 384, 425, 429, 299, 340, 516, 499, 481, 466, 
    11, 23, 229, 338, 427, 413, 275, 299, 315, 312, 456, 507, 532, 539, 535, 
    213, 164, 415, 398, 395, 459, 380, 301, 257, 320, 479, 524, 586, 563, 525, 
    475, 456, 502, 384, 365, 451, 443, 327, 267, 309, 458, 572, 613, 552, 493, 
    510, 492, 509, 413, 419, 442, 398, 291, 319, 333, 432, 566, 639, 592, 506, 
    524, 488, 434, 413, 397, 380, 398, 332, 399, 378, 428, 563, 634, 639, 565, 
    525, 471, 388, 402, 484, 435, 401, 370, 371, 393, 425, 431, 554, 618, 575, 
    528, 420, 423, 433, 504, 520, 466, 400, 322, 364, 412, 328, 334, 436, 503, 
    561, 482, 487, 481, 478, 486, 488, 471, 412, 382, 378, 338, 346, 387, 367, 
    567, 504, 476, 513, 517, 463, 424, 457, 472, 398, 310, 367, 389, 356, 331, 
    556, 516, 472, 533, 524, 440, 458, 462, 455, 351, 330, 366, 391, 371, 316, 
    546, 510, 475, 517, 467, 278, 433, 435, 398, 320, 322, 332, 332, 318, 325, 
    529, 484, 442, 520, 488, 405, 410, 362, 324, 261, 303, 307, 282, 279, 343, 
    457, 458, 399, 479, 497, 453, 347, 303, 268, 240, 282, 305, 290, 301, 311, 
    
    -- channel=521
    133, 49, 0, 0, 0, 0, 0, 0, 0, 6, 57, 0, 0, 0, 0, 
    131, 87, 0, 0, 142, 47, 5, 0, 1, 6, 93, 2, 0, 0, 0, 
    117, 112, 0, 0, 215, 150, 58, 34, 23, 70, 140, 94, 71, 55, 23, 
    37, 82, 78, 12, 201, 186, 108, 65, 78, 134, 160, 155, 171, 149, 117, 
    51, 85, 84, 4, 172, 198, 150, 96, 119, 143, 148, 140, 143, 60, 64, 
    69, 91, 69, 28, 156, 193, 133, 111, 152, 169, 153, 154, 151, 62, 25, 
    38, 45, 0, 39, 119, 175, 157, 161, 174, 184, 171, 146, 153, 130, 66, 
    49, 47, 0, 61, 161, 186, 195, 163, 125, 126, 128, 81, 119, 133, 123, 
    51, 52, 24, 93, 193, 201, 203, 132, 52, 42, 64, 0, 33, 62, 84, 
    79, 90, 120, 118, 164, 204, 223, 177, 66, 60, 13, 0, 0, 8, 10, 
    111, 106, 151, 127, 141, 116, 144, 166, 127, 28, 7, 21, 45, 14, 14, 
    112, 88, 156, 177, 146, 78, 98, 107, 97, 0, 20, 43, 65, 29, 6, 
    96, 53, 119, 187, 103, 2, 67, 51, 34, 3, 23, 34, 48, 24, 13, 
    76, 19, 78, 191, 106, 27, 15, 0, 0, 0, 15, 23, 15, 18, 29, 
    55, 19, 65, 211, 150, 81, 1, 0, 0, 6, 12, 21, 8, 20, 22, 
    
    -- channel=522
    89, 155, 142, 137, 116, 150, 143, 140, 96, 90, 129, 102, 135, 141, 143, 
    92, 135, 145, 139, 46, 85, 112, 108, 97, 73, 113, 84, 106, 121, 129, 
    96, 108, 140, 136, 50, 27, 97, 124, 115, 95, 68, 83, 77, 78, 81, 
    43, 83, 82, 106, 72, 22, 43, 66, 86, 102, 51, 76, 39, 49, 83, 
    67, 88, 70, 90, 81, 45, 46, 64, 84, 92, 65, 74, 50, 66, 112, 
    82, 84, 79, 94, 73, 51, 48, 72, 56, 73, 67, 81, 50, 62, 108, 
    93, 95, 101, 102, 64, 61, 40, 77, 37, 60, 63, 73, 59, 43, 71, 
    91, 103, 89, 106, 48, 50, 42, 55, 76, 84, 70, 132, 97, 60, 81, 
    76, 105, 72, 82, 41, 21, 28, 24, 114, 100, 75, 106, 143, 109, 120, 
    67, 88, 65, 65, 64, 57, 44, 22, 58, 97, 84, 115, 107, 94, 125, 
    71, 74, 70, 55, 60, 49, 79, 69, 48, 81, 113, 99, 90, 92, 108, 
    77, 69, 83, 48, 49, 74, 72, 71, 65, 84, 117, 97, 86, 90, 94, 
    78, 88, 100, 47, 46, 123, 90, 93, 89, 105, 113, 104, 99, 105, 98, 
    82, 100, 125, 51, 41, 89, 84, 111, 111, 119, 110, 107, 100, 117, 100, 
    102, 101, 133, 56, 51, 69, 106, 121, 110, 128, 111, 105, 100, 110, 107, 
    
    -- channel=523
    6, 5, 187, 196, 174, 182, 195, 185, 181, 122, 58, 212, 220, 222, 223, 
    6, 0, 163, 163, 175, 177, 190, 201, 222, 175, 91, 239, 237, 232, 234, 
    11, 9, 96, 149, 187, 216, 155, 169, 196, 131, 182, 231, 242, 237, 239, 
    58, 0, 139, 211, 188, 215, 156, 152, 118, 120, 232, 213, 265, 286, 245, 
    208, 174, 227, 206, 151, 214, 222, 190, 125, 129, 204, 248, 278, 274, 223, 
    237, 224, 251, 188, 190, 220, 219, 139, 136, 127, 191, 243, 290, 274, 224, 
    245, 224, 241, 197, 189, 155, 200, 138, 195, 171, 175, 243, 289, 284, 240, 
    249, 224, 220, 184, 226, 213, 190, 172, 187, 179, 221, 243, 272, 307, 246, 
    256, 192, 200, 196, 224, 224, 198, 211, 145, 179, 206, 163, 171, 244, 227, 
    255, 203, 226, 230, 226, 246, 234, 212, 172, 161, 222, 175, 144, 196, 193, 
    256, 237, 211, 229, 229, 241, 199, 220, 238, 231, 154, 170, 190, 189, 172, 
    253, 252, 203, 248, 260, 232, 209, 219, 231, 201, 143, 188, 194, 187, 165, 
    251, 247, 211, 242, 267, 144, 216, 227, 226, 177, 158, 171, 189, 173, 166, 
    252, 234, 193, 234, 240, 166, 232, 199, 184, 142, 153, 153, 155, 133, 164, 
    229, 216, 176, 220, 235, 232, 206, 174, 165, 104, 146, 152, 143, 144, 167, 
    
    -- channel=524
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=525
    36, 145, 158, 118, 130, 137, 122, 131, 88, 25, 163, 150, 131, 137, 129, 
    37, 102, 183, 134, 153, 133, 172, 174, 157, 56, 190, 184, 162, 155, 148, 
    35, 61, 181, 117, 208, 120, 130, 176, 170, 140, 199, 224, 201, 198, 185, 
    0, 31, 158, 140, 239, 158, 92, 84, 107, 183, 221, 239, 225, 227, 249, 
    140, 174, 197, 106, 199, 204, 168, 111, 131, 175, 227, 258, 243, 193, 234, 
    198, 208, 209, 131, 196, 203, 161, 109, 126, 161, 212, 277, 262, 194, 201, 
    204, 198, 160, 174, 153, 165, 137, 160, 156, 181, 200, 273, 266, 233, 188, 
    203, 206, 94, 209, 177, 195, 164, 144, 198, 174, 201, 276, 310, 259, 251, 
    183, 180, 131, 187, 208, 186, 153, 120, 172, 147, 163, 96, 212, 237, 279, 
    202, 183, 204, 194, 216, 238, 230, 165, 97, 151, 149, 137, 121, 138, 191, 
    229, 187, 227, 196, 201, 164, 214, 212, 184, 146, 143, 142, 157, 130, 134, 
    236, 187, 235, 224, 213, 170, 188, 186, 179, 111, 148, 153, 170, 133, 114, 
    226, 203, 236, 223, 166, 132, 197, 188, 162, 120, 156, 141, 160, 153, 121, 
    216, 191, 224, 236, 160, 123, 165, 155, 131, 118, 136, 128, 108, 139, 139, 
    210, 189, 191, 254, 196, 171, 144, 142, 100, 117, 129, 129, 106, 125, 148, 
    
    -- channel=526
    0, 0, 0, 4, 0, 0, 0, 0, 21, 58, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 26, 0, 23, 24, 13, 0, 0, 0, 0, 0, 17, 0, 
    31, 0, 0, 62, 0, 0, 14, 49, 0, 0, 0, 0, 0, 53, 0, 
    1, 0, 1, 32, 0, 0, 25, 17, 0, 0, 0, 0, 0, 55, 0, 
    3, 0, 21, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 16, 26, 
    18, 0, 56, 0, 9, 0, 4, 0, 0, 0, 0, 0, 0, 9, 0, 
    46, 0, 0, 0, 0, 0, 4, 40, 0, 14, 0, 27, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 14, 24, 0, 8, 0, 0, 0, 0, 
    1, 28, 0, 0, 0, 29, 0, 0, 16, 17, 0, 0, 0, 12, 0, 
    0, 42, 0, 0, 0, 14, 0, 0, 1, 51, 0, 0, 0, 11, 10, 
    4, 24, 0, 0, 34, 0, 0, 0, 16, 25, 0, 0, 0, 0, 0, 
    14, 28, 0, 0, 29, 0, 0, 0, 13, 4, 0, 0, 11, 0, 0, 
    15, 13, 0, 0, 7, 11, 28, 0, 25, 0, 0, 0, 1, 0, 0, 
    
    -- channel=527
    17, 149, 344, 285, 280, 306, 304, 326, 311, 112, 297, 378, 360, 359, 344, 
    19, 78, 322, 287, 365, 276, 326, 368, 342, 181, 412, 425, 396, 384, 367, 
    19, 38, 311, 292, 427, 273, 197, 252, 244, 308, 428, 439, 444, 452, 436, 
    148, 235, 420, 271, 409, 379, 295, 222, 232, 327, 420, 498, 481, 427, 459, 
    384, 415, 416, 246, 382, 387, 346, 215, 247, 298, 421, 532, 507, 392, 420, 
    419, 408, 410, 312, 391, 360, 293, 228, 298, 319, 382, 541, 526, 444, 404, 
    418, 400, 287, 400, 326, 345, 300, 311, 322, 348, 380, 530, 532, 526, 429, 
    399, 386, 251, 443, 377, 364, 337, 279, 360, 310, 341, 342, 518, 487, 493, 
    394, 348, 363, 381, 447, 458, 374, 290, 278, 283, 362, 240, 297, 354, 470, 
    446, 392, 414, 408, 399, 399, 429, 388, 302, 356, 263, 295, 305, 306, 301, 
    468, 376, 445, 425, 443, 334, 389, 388, 377, 269, 272, 318, 330, 266, 259, 
    453, 395, 446, 448, 417, 333, 404, 387, 357, 228, 314, 293, 349, 283, 245, 
    436, 391, 429, 440, 331, 207, 396, 344, 295, 229, 294, 266, 256, 267, 264, 
    411, 365, 397, 463, 370, 340, 304, 285, 237, 196, 267, 252, 209, 256, 300, 
    349, 374, 324, 453, 399, 340, 231, 249, 182, 227, 234, 262, 235, 255, 261, 
    
    -- channel=528
    1, 160, 426, 416, 406, 411, 422, 434, 418, 239, 330, 517, 509, 502, 490, 
    6, 88, 364, 414, 510, 442, 461, 503, 511, 330, 453, 599, 570, 550, 536, 
    11, 39, 295, 417, 592, 493, 348, 383, 394, 401, 551, 608, 632, 633, 618, 
    174, 187, 471, 441, 562, 579, 449, 350, 323, 444, 592, 660, 728, 671, 639, 
    505, 524, 568, 413, 504, 597, 553, 394, 349, 429, 573, 700, 737, 593, 557, 
    579, 572, 574, 464, 543, 577, 499, 369, 402, 448, 549, 699, 748, 620, 519, 
    574, 556, 484, 513, 493, 505, 486, 455, 491, 492, 542, 694, 752, 722, 596, 
    564, 548, 449, 549, 585, 557, 517, 469, 489, 485, 520, 540, 692, 717, 664, 
    550, 486, 528, 569, 638, 652, 587, 476, 414, 447, 491, 367, 427, 518, 606, 
    596, 542, 600, 601, 601, 631, 646, 588, 472, 475, 441, 407, 419, 447, 447, 
    637, 558, 598, 627, 637, 548, 554, 602, 580, 460, 384, 442, 482, 425, 391, 
    628, 556, 593, 675, 652, 557, 572, 581, 558, 397, 405, 447, 491, 441, 369, 
    605, 531, 566, 653, 567, 412, 557, 537, 483, 374, 395, 406, 411, 397, 387, 
    578, 487, 505, 648, 578, 516, 492, 441, 383, 310, 364, 371, 330, 350, 415, 
    497, 463, 437, 620, 609, 536, 405, 370, 303, 290, 336, 365, 338, 358, 382, 
    
    -- channel=529
    0, 0, 225, 245, 225, 230, 250, 248, 260, 168, 77, 275, 289, 290, 287, 
    0, 0, 158, 200, 255, 240, 248, 269, 287, 240, 150, 327, 318, 307, 304, 
    0, 0, 71, 200, 258, 296, 156, 175, 212, 188, 254, 307, 340, 344, 345, 
    130, 39, 223, 277, 227, 314, 254, 194, 145, 156, 306, 314, 382, 383, 327, 
    337, 282, 320, 272, 190, 280, 302, 238, 159, 160, 270, 347, 394, 378, 299, 
    336, 309, 336, 283, 257, 285, 269, 184, 196, 181, 247, 333, 410, 407, 319, 
    340, 307, 289, 271, 235, 209, 271, 198, 264, 225, 245, 329, 406, 427, 364, 
    349, 302, 287, 223, 327, 281, 264, 244, 232, 238, 282, 259, 353, 413, 368, 
    363, 252, 280, 244, 332, 333, 296, 278, 158, 238, 275, 211, 151, 282, 296, 
    377, 309, 311, 311, 287, 309, 322, 307, 265, 236, 251, 215, 210, 252, 207, 
    368, 339, 289, 320, 334, 312, 245, 286, 323, 274, 194, 225, 245, 232, 216, 
    355, 360, 274, 343, 347, 298, 287, 295, 302, 248, 190, 235, 250, 251, 207, 
    352, 344, 285, 330, 323, 140, 271, 281, 271, 220, 191, 212, 211, 202, 207, 
    347, 326, 261, 327, 335, 265, 267, 234, 219, 161, 181, 191, 187, 155, 218, 
    299, 303, 238, 291, 325, 305, 243, 199, 186, 138, 171, 192, 185, 184, 191, 
    
    -- channel=530
    125, 113, 40, 37, 49, 42, 43, 51, 42, 72, 76, 55, 29, 39, 30, 
    123, 118, 54, 33, 59, 67, 52, 59, 47, 48, 107, 57, 39, 33, 26, 
    119, 119, 87, 45, 46, 45, 55, 49, 31, 51, 102, 65, 48, 50, 53, 
    134, 136, 145, 68, 45, 39, 66, 69, 68, 74, 70, 67, 51, 70, 72, 
    96, 117, 94, 64, 66, 41, 43, 52, 67, 68, 79, 80, 62, 92, 108, 
    84, 89, 87, 62, 70, 52, 38, 52, 75, 71, 74, 77, 78, 97, 128, 
    94, 79, 61, 42, 56, 49, 52, 58, 77, 76, 77, 82, 79, 81, 114, 
    100, 69, 6, 43, 62, 59, 50, 61, 59, 85, 71, 81, 61, 75, 92, 
    101, 78, 10, 57, 49, 61, 57, 48, 81, 50, 63, 60, 77, 58, 92, 
    105, 98, 55, 51, 63, 46, 36, 53, 62, 55, 57, 45, 58, 66, 69, 
    95, 91, 64, 55, 58, 57, 60, 42, 42, 59, 51, 61, 49, 45, 62, 
    98, 94, 80, 41, 41, 27, 62, 47, 50, 46, 75, 56, 50, 54, 58, 
    103, 114, 99, 50, 28, 0, 43, 43, 42, 52, 67, 56, 57, 48, 59, 
    102, 119, 113, 61, 45, 31, 56, 42, 47, 63, 71, 60, 62, 68, 60, 
    100, 118, 120, 63, 53, 52, 49, 49, 56, 74, 70, 66, 66, 76, 61, 
    
    -- channel=531
    77, 0, 13, 78, 56, 26, 46, 34, 102, 138, 0, 47, 53, 42, 50, 
    73, 0, 0, 59, 102, 82, 54, 48, 92, 180, 0, 62, 65, 56, 63, 
    74, 37, 0, 44, 86, 188, 87, 48, 95, 59, 24, 44, 76, 68, 72, 
    112, 0, 0, 97, 63, 158, 126, 125, 75, 6, 92, 25, 110, 122, 41, 
    92, 15, 60, 128, 34, 112, 142, 162, 75, 35, 48, 25, 85, 105, 0, 
    64, 49, 68, 86, 68, 117, 154, 116, 92, 49, 53, 9, 73, 92, 10, 
    49, 47, 100, 62, 103, 76, 152, 72, 131, 75, 50, 14, 65, 89, 57, 
    57, 46, 157, 27, 126, 112, 133, 115, 74, 63, 94, 16, 26, 95, 29, 
    86, 36, 117, 65, 107, 120, 132, 181, 13, 84, 92, 80, 0, 62, 0, 
    71, 44, 81, 101, 79, 106, 118, 138, 108, 50, 118, 64, 50, 85, 29, 
    57, 86, 52, 92, 89, 145, 56, 94, 132, 131, 57, 59, 79, 105, 75, 
    48, 97, 23, 107, 124, 130, 71, 95, 112, 137, 20, 83, 79, 99, 95, 
    51, 57, 11, 104, 172, 74, 71, 89, 117, 101, 40, 78, 88, 77, 83, 
    58, 45, 0, 81, 145, 78, 112, 81, 95, 68, 52, 68, 95, 34, 66, 
    49, 33, 0, 63, 111, 115, 109, 73, 108, 23, 60, 64, 79, 53, 67, 
    
    -- channel=532
    32, 168, 0, 0, 0, 0, 0, 0, 0, 0, 89, 0, 0, 0, 0, 
    36, 124, 18, 0, 0, 0, 0, 0, 0, 0, 147, 0, 0, 0, 0, 
    32, 66, 86, 0, 26, 0, 0, 0, 0, 0, 61, 0, 0, 0, 0, 
    0, 70, 106, 0, 52, 0, 0, 0, 0, 87, 0, 18, 0, 0, 0, 
    0, 34, 0, 0, 80, 0, 0, 0, 5, 55, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 0, 5, 48, 13, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 16, 13, 26, 0, 0, 0, 
    0, 0, 0, 48, 0, 0, 0, 0, 0, 1, 0, 17, 0, 0, 0, 
    0, 0, 0, 40, 0, 0, 0, 0, 45, 0, 0, 0, 63, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 13, 13, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    
    -- channel=533
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=534
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 1, 2, 7, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 14, 1, 12, 23, 14, 
    0, 0, 2, 0, 0, 8, 7, 5, 0, 0, 9, 6, 13, 10, 6, 
    6, 5, 10, 0, 1, 12, 7, 0, 0, 0, 8, 9, 15, 8, 4, 
    4, 1, 7, 0, 0, 0, 0, 4, 2, 4, 0, 10, 14, 8, 2, 
    7, 4, 0, 0, 4, 9, 4, 0, 12, 1, 10, 33, 23, 20, 12, 
    7, 0, 0, 0, 6, 1, 0, 2, 0, 0, 2, 0, 1, 17, 15, 
    5, 0, 1, 8, 6, 16, 15, 0, 0, 0, 6, 0, 0, 0, 3, 
    10, 6, 4, 0, 4, 5, 5, 8, 11, 7, 0, 0, 0, 0, 0, 
    11, 10, 1, 10, 11, 13, 0, 2, 6, 0, 0, 0, 1, 0, 0, 
    12, 10, 5, 8, 12, 0, 5, 6, 7, 0, 0, 0, 4, 1, 0, 
    12, 7, 1, 8, 5, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 
    13, 6, 0, 11, 8, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=535
    65, 87, 194, 168, 146, 180, 186, 170, 143, 113, 93, 156, 193, 196, 202, 
    66, 81, 177, 139, 75, 105, 141, 148, 145, 125, 94, 132, 156, 173, 185, 
    71, 76, 127, 137, 65, 81, 97, 126, 136, 95, 84, 103, 113, 116, 124, 
    74, 47, 99, 136, 75, 67, 83, 93, 88, 78, 94, 90, 87, 106, 106, 
    123, 113, 114, 124, 72, 65, 89, 98, 85, 72, 85, 101, 97, 123, 125, 
    124, 112, 126, 127, 87, 74, 90, 76, 74, 64, 79, 95, 97, 129, 136, 
    132, 127, 147, 140, 79, 52, 77, 71, 71, 66, 69, 99, 100, 108, 109, 
    131, 133, 160, 114, 85, 78, 60, 90, 99, 87, 111, 129, 131, 117, 111, 
    131, 112, 118, 91, 76, 62, 54, 78, 97, 121, 128, 142, 116, 137, 130, 
    118, 108, 99, 99, 77, 79, 74, 59, 101, 118, 128, 145, 128, 135, 136, 
    111, 111, 89, 90, 95, 97, 87, 86, 98, 133, 126, 121, 121, 121, 133, 
    111, 121, 87, 83, 100, 113, 107, 103, 111, 127, 126, 120, 120, 127, 124, 
    116, 132, 104, 80, 109, 108, 124, 126, 129, 134, 128, 121, 121, 124, 124, 
    124, 145, 114, 82, 92, 125, 129, 141, 140, 124, 125, 123, 123, 119, 125, 
    128, 145, 114, 79, 88, 115, 141, 146, 139, 129, 123, 126, 121, 126, 124, 
    
    -- channel=536
    12, 0, 161, 188, 189, 175, 191, 183, 177, 169, 50, 197, 209, 214, 214, 
    12, 11, 127, 155, 181, 203, 182, 196, 224, 187, 81, 248, 246, 239, 233, 
    13, 19, 58, 164, 185, 249, 177, 185, 202, 131, 200, 259, 267, 256, 254, 
    98, 0, 124, 230, 173, 226, 176, 164, 127, 124, 244, 224, 276, 308, 263, 
    220, 178, 251, 236, 155, 232, 236, 205, 133, 137, 210, 261, 313, 324, 261, 
    262, 248, 274, 221, 184, 230, 241, 165, 146, 144, 213, 263, 331, 334, 274, 
    280, 252, 271, 204, 227, 196, 227, 132, 202, 178, 203, 258, 326, 320, 293, 
    294, 242, 236, 151, 245, 228, 202, 199, 178, 198, 239, 244, 276, 346, 290, 
    308, 225, 187, 195, 236, 231, 232, 229, 151, 203, 204, 198, 205, 278, 246, 
    298, 235, 233, 241, 257, 274, 244, 225, 216, 174, 223, 171, 154, 201, 218, 
    296, 288, 223, 255, 250, 270, 217, 243, 245, 240, 161, 168, 192, 202, 179, 
    295, 295, 215, 264, 276, 231, 217, 229, 246, 217, 143, 194, 190, 200, 173, 
    296, 290, 228, 267, 293, 166, 220, 237, 238, 191, 159, 181, 194, 173, 174, 
    294, 283, 224, 255, 257, 161, 230, 211, 200, 152, 155, 166, 167, 136, 166, 
    270, 255, 219, 231, 263, 255, 215, 168, 175, 118, 150, 157, 150, 147, 168, 
    
    -- channel=537
    34, 151, 242, 212, 193, 216, 217, 216, 207, 97, 207, 256, 266, 251, 251, 
    37, 90, 219, 219, 223, 172, 211, 218, 214, 135, 253, 226, 237, 246, 255, 
    44, 56, 201, 212, 266, 156, 137, 162, 156, 190, 202, 184, 215, 232, 229, 
    72, 143, 229, 144, 249, 221, 192, 153, 162, 217, 194, 242, 256, 187, 185, 
    160, 197, 165, 111, 229, 219, 206, 141, 164, 194, 203, 226, 210, 106, 125, 
    161, 164, 150, 149, 230, 210, 166, 146, 180, 198, 188, 218, 181, 101, 80, 
    137, 159, 136, 213, 160, 184, 172, 219, 179, 183, 188, 220, 190, 177, 112, 
    114, 173, 200, 299, 202, 190, 192, 187, 195, 168, 161, 162, 202, 163, 148, 
    89, 140, 275, 268, 226, 245, 208, 168, 187, 165, 204, 130, 141, 117, 168, 
    115, 150, 226, 219, 182, 196, 228, 212, 175, 220, 165, 199, 208, 188, 149, 
    141, 114, 206, 216, 221, 157, 204, 213, 207, 166, 170, 212, 216, 174, 174, 
    134, 103, 202, 238, 227, 221, 233, 223, 201, 142, 200, 184, 219, 183, 158, 
    118, 81, 157, 210, 183, 217, 243, 199, 175, 150, 181, 169, 169, 171, 171, 
    110, 60, 114, 207, 202, 286, 198, 175, 154, 132, 169, 161, 142, 172, 192, 
    81, 71, 82, 205, 191, 181, 151, 176, 129, 149, 151, 169, 155, 175, 166, 
    
    -- channel=538
    4, 202, 70, 4, 12, 38, 9, 27, 0, 0, 154, 40, 13, 13, 4, 
    7, 116, 141, 43, 9, 0, 33, 27, 0, 0, 192, 4, 0, 8, 5, 
    6, 45, 207, 42, 75, 0, 11, 67, 7, 21, 86, 30, 0, 6, 0, 
    0, 68, 135, 0, 112, 0, 0, 0, 30, 120, 14, 75, 0, 0, 28, 
    0, 40, 0, 0, 123, 15, 0, 0, 33, 84, 56, 73, 0, 0, 37, 
    0, 6, 0, 0, 68, 6, 0, 0, 18, 61, 48, 98, 0, 0, 0, 
    0, 0, 0, 29, 0, 28, 0, 42, 0, 39, 38, 87, 0, 0, 0, 
    0, 8, 0, 156, 0, 0, 0, 0, 36, 18, 0, 93, 60, 0, 0, 
    0, 19, 0, 85, 0, 0, 0, 0, 95, 0, 8, 0, 134, 3, 88, 
    0, 0, 22, 0, 25, 17, 0, 0, 0, 42, 0, 22, 16, 0, 55, 
    0, 0, 52, 0, 0, 0, 68, 20, 0, 0, 11, 38, 22, 0, 8, 
    0, 0, 85, 5, 0, 0, 32, 2, 0, 0, 71, 7, 31, 0, 0, 
    0, 0, 59, 2, 0, 27, 58, 0, 0, 0, 55, 3, 20, 9, 0, 
    0, 0, 59, 24, 0, 3, 0, 0, 0, 0, 42, 7, 0, 57, 19, 
    0, 0, 33, 61, 0, 0, 0, 18, 0, 40, 20, 17, 0, 33, 25, 
    
    -- channel=539
    0, 93, 381, 357, 322, 365, 379, 371, 365, 178, 227, 415, 443, 437, 435, 
    0, 34, 318, 327, 338, 300, 350, 387, 381, 273, 302, 433, 439, 439, 444, 
    8, 11, 246, 319, 367, 312, 219, 253, 285, 291, 342, 385, 424, 440, 444, 
    142, 131, 328, 322, 352, 376, 311, 249, 221, 272, 376, 419, 468, 425, 405, 
    377, 365, 376, 301, 305, 358, 359, 269, 227, 259, 361, 448, 462, 387, 350, 
    390, 371, 383, 330, 354, 352, 318, 235, 260, 267, 328, 432, 461, 407, 340, 
    386, 372, 335, 373, 301, 284, 303, 295, 314, 299, 317, 435, 461, 467, 385, 
    370, 374, 360, 400, 376, 343, 320, 287, 328, 296, 330, 332, 454, 448, 413, 
    365, 315, 407, 379, 407, 418, 351, 316, 266, 309, 355, 273, 244, 326, 383, 
    394, 354, 400, 399, 354, 366, 398, 376, 315, 332, 322, 323, 317, 331, 293, 
    404, 349, 378, 401, 410, 351, 337, 362, 388, 330, 285, 328, 346, 309, 288, 
    391, 365, 364, 424, 420, 385, 386, 386, 369, 299, 297, 316, 350, 320, 282, 
    379, 351, 356, 399, 369, 271, 382, 367, 338, 279, 288, 289, 284, 291, 287, 
    369, 326, 314, 399, 395, 391, 358, 319, 283, 235, 269, 268, 247, 255, 307, 
    317, 320, 265, 372, 381, 358, 299, 292, 242, 219, 251, 272, 261, 266, 278, 
    
    -- channel=540
    57, 0, 173, 195, 194, 173, 190, 194, 252, 161, 97, 238, 223, 216, 212, 
    54, 0, 121, 170, 288, 224, 217, 238, 248, 251, 149, 296, 268, 246, 238, 
    54, 33, 81, 158, 284, 321, 159, 142, 188, 215, 250, 284, 314, 319, 316, 
    186, 107, 211, 230, 248, 351, 283, 217, 168, 162, 310, 299, 374, 355, 301, 
    321, 262, 296, 254, 202, 300, 309, 252, 179, 177, 276, 320, 370, 336, 241, 
    300, 278, 299, 256, 257, 294, 286, 213, 229, 206, 256, 305, 383, 366, 258, 
    291, 269, 236, 252, 248, 238, 287, 228, 291, 252, 254, 307, 370, 403, 334, 
    292, 258, 256, 219, 323, 295, 297, 243, 251, 223, 268, 190, 316, 365, 331, 
    319, 222, 285, 236, 347, 365, 322, 314, 143, 223, 262, 194, 101, 235, 244, 
    342, 276, 299, 308, 279, 297, 338, 350, 267, 218, 234, 193, 198, 226, 166, 
    335, 302, 288, 315, 324, 310, 241, 278, 329, 245, 186, 210, 232, 222, 188, 
    315, 326, 259, 341, 334, 292, 277, 285, 286, 242, 169, 218, 241, 232, 206, 
    312, 294, 252, 331, 313, 135, 248, 252, 247, 201, 173, 197, 190, 197, 198, 
    304, 270, 212, 327, 342, 248, 244, 203, 189, 154, 167, 179, 179, 147, 205, 
    255, 260, 181, 299, 324, 281, 212, 174, 170, 123, 162, 180, 186, 165, 181, 
    
    -- channel=541
    19, 231, 452, 412, 400, 417, 416, 440, 417, 188, 399, 544, 504, 497, 476, 
    23, 125, 428, 433, 545, 446, 490, 538, 528, 276, 563, 623, 576, 550, 529, 
    27, 59, 393, 434, 666, 467, 347, 404, 399, 428, 637, 653, 661, 667, 643, 
    153, 236, 580, 441, 658, 595, 446, 352, 348, 516, 649, 742, 776, 703, 694, 
    526, 598, 610, 385, 593, 637, 568, 377, 380, 483, 642, 793, 776, 590, 613, 
    614, 617, 609, 453, 619, 617, 498, 361, 443, 499, 602, 799, 797, 624, 558, 
    606, 590, 472, 547, 516, 531, 491, 503, 528, 552, 590, 793, 807, 765, 619, 
    585, 584, 396, 646, 615, 600, 545, 481, 540, 520, 550, 602, 776, 759, 709, 
    560, 517, 539, 629, 685, 710, 609, 470, 460, 440, 528, 337, 481, 540, 687, 
    629, 581, 649, 636, 648, 674, 693, 610, 454, 508, 444, 419, 432, 465, 476, 
    684, 574, 668, 663, 678, 553, 612, 636, 596, 461, 387, 475, 509, 417, 400, 
    675, 573, 679, 721, 685, 561, 617, 613, 573, 362, 449, 465, 528, 438, 365, 
    642, 558, 645, 700, 560, 379, 596, 555, 479, 356, 432, 416, 430, 408, 394, 
    606, 503, 574, 715, 583, 519, 506, 442, 369, 301, 394, 378, 322, 379, 436, 
    517, 493, 485, 704, 631, 544, 388, 381, 283, 304, 353, 382, 339, 382, 403, 
    
    -- channel=542
    6, 0, 0, 36, 0, 0, 5, 0, 112, 207, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 11, 0, 0, 27, 315, 0, 0, 7, 0, 13, 
    0, 0, 0, 0, 0, 248, 10, 0, 42, 0, 0, 0, 0, 0, 0, 
    168, 0, 0, 91, 0, 113, 93, 107, 0, 0, 0, 0, 0, 77, 0, 
    100, 0, 0, 211, 0, 0, 90, 200, 0, 0, 0, 0, 0, 164, 0, 
    0, 0, 16, 76, 0, 0, 141, 67, 0, 0, 0, 0, 0, 157, 0, 
    0, 0, 111, 0, 11, 0, 126, 0, 57, 0, 0, 0, 0, 47, 43, 
    36, 0, 235, 0, 53, 0, 49, 10, 0, 0, 5, 0, 0, 45, 0, 
    136, 0, 49, 0, 0, 0, 32, 226, 0, 23, 10, 81, 0, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 74, 84, 0, 110, 0, 0, 20, 0, 
    0, 72, 0, 0, 0, 147, 0, 0, 95, 135, 0, 0, 0, 78, 0, 
    0, 131, 0, 0, 31, 84, 0, 0, 44, 204, 0, 0, 0, 56, 68, 
    0, 65, 0, 0, 200, 0, 0, 0, 97, 96, 0, 0, 0, 0, 21, 
    26, 68, 0, 0, 150, 0, 61, 19, 73, 18, 0, 0, 69, 0, 0, 
    22, 29, 0, 0, 38, 79, 116, 0, 124, 0, 0, 0, 28, 0, 0, 
    
    -- channel=543
    41, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 41, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 40, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=544
    16, 24, 109, 128, 97, 123, 130, 116, 103, 94, 35, 92, 139, 137, 147, 
    18, 17, 84, 120, 32, 70, 80, 80, 94, 109, 0, 74, 109, 123, 136, 
    25, 17, 41, 111, 27, 58, 77, 83, 101, 61, 2, 44, 59, 61, 73, 
    33, 3, 0, 94, 32, 45, 47, 64, 56, 35, 27, 26, 44, 45, 40, 
    47, 10, 36, 96, 26, 42, 57, 75, 45, 38, 25, 19, 39, 62, 38, 
    49, 44, 46, 80, 33, 43, 69, 69, 25, 25, 24, 16, 25, 40, 35, 
    53, 58, 100, 64, 58, 42, 52, 38, 34, 18, 24, 17, 28, 25, 31, 
    52, 63, 132, 62, 47, 33, 43, 42, 44, 50, 44, 66, 41, 41, 24, 
    46, 57, 96, 72, 33, 18, 32, 58, 65, 84, 56, 86, 73, 74, 30, 
    33, 36, 49, 56, 43, 47, 37, 40, 55, 60, 94, 96, 79, 77, 76, 
    28, 42, 29, 51, 41, 64, 42, 55, 59, 90, 87, 73, 73, 96, 82, 
    30, 42, 21, 44, 58, 88, 50, 65, 66, 106, 60, 79, 64, 84, 87, 
    30, 44, 28, 37, 80, 136, 69, 85, 95, 95, 68, 82, 82, 86, 79, 
    38, 44, 32, 22, 69, 85, 99, 97, 103, 95, 70, 78, 87, 71, 72, 
    51, 36, 44, 13, 46, 71, 103, 97, 102, 68, 78, 73, 80, 67, 79, 
    
    -- channel=545
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=546
    0, 18, 38, 0, 0, 2, 0, 0, 0, 0, 18, 20, 0, 0, 0, 
    0, 0, 74, 0, 7, 0, 5, 9, 1, 0, 54, 1, 0, 0, 0, 
    0, 0, 81, 0, 29, 0, 0, 13, 0, 0, 45, 5, 0, 0, 0, 
    0, 0, 67, 0, 41, 0, 0, 0, 6, 15, 25, 16, 0, 0, 2, 
    0, 17, 6, 0, 40, 0, 0, 0, 7, 4, 22, 34, 0, 0, 4, 
    0, 0, 3, 0, 26, 0, 0, 0, 17, 4, 13, 42, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 4, 13, 0, 40, 0, 0, 0, 
    0, 0, 0, 68, 0, 3, 0, 0, 20, 0, 3, 11, 24, 3, 0, 
    0, 0, 0, 19, 0, 11, 0, 0, 2, 0, 26, 0, 26, 2, 22, 
    0, 0, 6, 1, 1, 1, 0, 0, 0, 11, 0, 6, 0, 8, 11, 
    0, 0, 18, 0, 0, 0, 18, 0, 0, 0, 0, 8, 8, 0, 0, 
    0, 0, 23, 0, 0, 0, 12, 0, 0, 0, 17, 0, 18, 0, 0, 
    0, 0, 9, 2, 0, 0, 30, 0, 0, 0, 17, 0, 3, 0, 0, 
    0, 0, 1, 16, 0, 0, 0, 0, 0, 0, 14, 0, 0, 7, 4, 
    0, 3, 0, 31, 0, 0, 0, 2, 0, 0, 0, 3, 0, 7, 2, 
    
    -- channel=547
    48, 144, 326, 261, 237, 289, 297, 285, 249, 138, 193, 294, 333, 328, 332, 
    51, 89, 309, 229, 168, 174, 221, 244, 233, 152, 232, 243, 277, 298, 310, 
    61, 64, 268, 237, 174, 109, 137, 187, 179, 168, 194, 182, 206, 224, 233, 
    134, 155, 239, 179, 170, 144, 154, 152, 160, 169, 170, 198, 186, 160, 174, 
    191, 194, 188, 146, 180, 142, 153, 119, 142, 140, 176, 209, 185, 158, 179, 
    188, 177, 183, 172, 180, 134, 134, 119, 152, 139, 151, 205, 170, 164, 175, 
    191, 188, 184, 234, 149, 131, 135, 133, 141, 128, 146, 210, 176, 181, 153, 
    172, 189, 220, 279, 153, 131, 120, 138, 167, 139, 152, 166, 198, 174, 159, 
    160, 165, 244, 228, 156, 164, 128, 138, 180, 162, 216, 181, 190, 169, 193, 
    168, 160, 191, 181, 149, 139, 138, 138, 167, 217, 188, 236, 218, 216, 192, 
    165, 137, 173, 181, 181, 143, 171, 154, 166, 189, 189, 220, 209, 187, 197, 
    162, 150, 173, 167, 178, 171, 207, 188, 181, 169, 218, 186, 209, 191, 183, 
    159, 161, 164, 154, 163, 179, 235, 195, 185, 174, 207, 177, 180, 183, 192, 
    158, 163, 155, 161, 167, 239, 211, 202, 191, 163, 200, 182, 170, 193, 206, 
    142, 175, 132, 155, 148, 182, 171, 207, 178, 186, 181, 195, 181, 197, 187, 
    
    -- channel=548
    50, 25, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    51, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    
    -- channel=549
    0, 0, 47, 42, 44, 30, 30, 32, 52, 0, 0, 76, 57, 50, 48, 
    0, 0, 44, 40, 119, 64, 85, 83, 102, 64, 4, 115, 94, 82, 79, 
    0, 0, 0, 12, 160, 134, 47, 68, 94, 60, 90, 134, 143, 138, 125, 
    0, 0, 23, 69, 153, 175, 70, 46, 36, 49, 167, 145, 197, 189, 151, 
    105, 50, 120, 64, 94, 168, 158, 92, 54, 58, 144, 154, 192, 141, 87, 
    122, 112, 133, 68, 121, 161, 143, 65, 73, 64, 117, 167, 198, 142, 69, 
    110, 101, 97, 100, 93, 103, 133, 88, 130, 102, 111, 162, 195, 194, 103, 
    113, 106, 89, 117, 155, 140, 152, 91, 125, 86, 128, 133, 188, 202, 143, 
    115, 71, 126, 103, 179, 170, 135, 144, 40, 66, 120, 4, 47, 142, 121, 
    138, 84, 145, 143, 143, 188, 200, 159, 51, 75, 102, 60, 31, 76, 54, 
    149, 115, 146, 147, 153, 141, 129, 151, 174, 105, 52, 62, 88, 78, 56, 
    141, 132, 122, 189, 185, 147, 122, 133, 139, 82, 32, 80, 108, 77, 50, 
    132, 114, 102, 178, 173, 43, 135, 120, 117, 57, 49, 62, 85, 73, 50, 
    124, 84, 61, 179, 167, 61, 113, 77, 64, 21, 39, 41, 42, 23, 64, 
    98, 78, 30, 175, 159, 132, 83, 55, 36, 0, 31, 45, 31, 28, 56, 
    
    -- channel=550
    0, 141, 404, 356, 344, 375, 378, 377, 329, 166, 261, 432, 444, 439, 435, 
    0, 59, 387, 342, 353, 332, 376, 405, 412, 239, 328, 462, 462, 462, 458, 
    0, 15, 314, 331, 421, 324, 279, 345, 348, 291, 405, 462, 473, 475, 465, 
    72, 93, 337, 344, 425, 391, 281, 251, 249, 326, 445, 477, 514, 488, 479, 
    363, 352, 428, 305, 379, 427, 395, 277, 256, 306, 439, 517, 534, 446, 435, 
    434, 428, 442, 335, 397, 409, 368, 258, 278, 302, 401, 535, 544, 453, 404, 
    443, 425, 402, 403, 362, 355, 345, 302, 349, 335, 386, 531, 549, 520, 422, 
    432, 421, 355, 462, 411, 385, 358, 315, 373, 353, 389, 468, 545, 543, 475, 
    411, 372, 405, 440, 439, 435, 377, 341, 338, 328, 390, 270, 399, 450, 484, 
    444, 382, 443, 432, 445, 470, 451, 394, 304, 361, 371, 348, 314, 361, 380, 
    470, 398, 445, 455, 454, 399, 422, 438, 426, 374, 310, 351, 372, 340, 319, 
    470, 409, 438, 483, 479, 414, 426, 428, 419, 317, 322, 351, 385, 337, 293, 
    452, 418, 422, 467, 428, 336, 451, 423, 390, 296, 329, 319, 347, 327, 306, 
    437, 388, 384, 471, 421, 351, 409, 366, 325, 258, 305, 295, 269, 289, 329, 
    391, 372, 330, 460, 432, 411, 332, 321, 263, 235, 280, 297, 266, 286, 318, 
    
    -- channel=551
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=552
    0, 0, 33, 44, 35, 37, 48, 48, 45, 24, 0, 50, 61, 59, 57, 
    0, 0, 5, 29, 30, 32, 25, 39, 36, 17, 43, 49, 55, 55, 56, 
    0, 0, 0, 43, 26, 21, 0, 0, 0, 11, 40, 25, 41, 51, 55, 
    36, 15, 56, 32, 14, 24, 42, 19, 3, 18, 21, 38, 50, 35, 23, 
    42, 60, 35, 20, 19, 16, 22, 11, 2, 10, 17, 47, 42, 32, 28, 
    34, 32, 27, 33, 31, 20, 10, 3, 19, 19, 18, 32, 41, 39, 29, 
    36, 31, 16, 30, 20, 6, 18, 12, 23, 14, 19, 35, 41, 46, 45, 
    32, 29, 34, 32, 36, 25, 7, 31, 2, 18, 19, 0, 24, 34, 32, 
    31, 17, 36, 51, 29, 45, 38, 13, 11, 23, 22, 28, 0, 0, 17, 
    33, 39, 37, 36, 20, 12, 17, 29, 48, 28, 15, 20, 38, 30, 15, 
    32, 31, 21, 40, 39, 24, 12, 21, 19, 24, 9, 32, 30, 17, 19, 
    30, 25, 27, 34, 35, 18, 39, 33, 27, 12, 27, 21, 23, 27, 17, 
    28, 21, 26, 28, 16, 1, 26, 23, 15, 12, 16, 14, 8, 5, 19, 
    26, 20, 20, 26, 27, 65, 28, 15, 11, 3, 13, 13, 8, 12, 21, 
    10, 17, 16, 14, 25, 28, 9, 12, 6, 10, 9, 15, 15, 21, 10, 
    
    -- channel=553
    0, 106, 440, 399, 378, 407, 423, 436, 418, 185, 290, 508, 509, 504, 488, 
    0, 28, 370, 369, 455, 382, 424, 482, 466, 264, 462, 564, 540, 529, 517, 
    0, 0, 300, 386, 516, 391, 246, 304, 314, 350, 525, 538, 578, 595, 585, 
    175, 190, 509, 390, 482, 489, 401, 293, 265, 380, 523, 608, 649, 583, 564, 
    493, 532, 525, 342, 441, 488, 462, 303, 284, 348, 504, 663, 655, 519, 509, 
    532, 516, 521, 412, 490, 472, 391, 274, 356, 378, 464, 649, 672, 574, 493, 
    531, 500, 398, 491, 407, 395, 396, 375, 422, 417, 455, 646, 674, 671, 554, 
    513, 491, 385, 531, 509, 472, 414, 391, 417, 396, 443, 431, 632, 637, 602, 
    506, 421, 477, 513, 560, 590, 495, 385, 335, 372, 454, 321, 331, 421, 552, 
    558, 500, 539, 531, 502, 509, 539, 499, 421, 438, 365, 370, 389, 409, 378, 
    582, 491, 531, 552, 572, 454, 465, 494, 491, 391, 323, 410, 433, 352, 341, 
    566, 503, 532, 584, 562, 455, 524, 506, 478, 317, 382, 383, 441, 384, 317, 
    545, 485, 513, 558, 456, 272, 500, 456, 397, 306, 357, 340, 334, 328, 337, 
    518, 451, 461, 571, 497, 484, 423, 372, 314, 239, 324, 315, 267, 303, 374, 
    426, 441, 384, 539, 516, 461, 322, 320, 243, 257, 285, 323, 293, 323, 323, 
    
    -- channel=554
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=555
    0, 81, 5, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 65, 105, 41, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 33, 27, 0, 0, 0, 104, 194, 191, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 72, 0, 0, 0, 0, 2, 0, 0, 0, 10, 24, 
    0, 0, 0, 0, 0, 14, 0, 14, 7, 22, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 35, 40, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 21, 0, 1, 0, 0, 0, 0, 36, 15, 49, 313, 109, 33, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 65, 9, 0, 0, 237, 228, 95, 
    0, 0, 0, 0, 30, 119, 26, 0, 0, 0, 64, 12, 0, 0, 122, 
    0, 0, 0, 0, 0, 0, 52, 57, 0, 51, 28, 0, 0, 18, 37, 
    0, 0, 0, 0, 6, 41, 0, 0, 3, 16, 0, 26, 0, 0, 0, 
    0, 0, 7, 0, 54, 149, 43, 66, 82, 43, 29, 38, 115, 70, 0, 
    0, 0, 28, 0, 0, 0, 50, 82, 88, 59, 17, 16, 28, 22, 0, 
    74, 0, 51, 35, 0, 12, 113, 85, 67, 5, 30, 2, 0, 0, 53, 
    
    -- channel=556
    22, 0, 31, 98, 79, 70, 95, 74, 105, 143, 0, 68, 106, 102, 114, 
    22, 0, 0, 67, 47, 85, 44, 45, 76, 157, 0, 68, 93, 96, 105, 
    27, 16, 0, 75, 0, 127, 61, 14, 47, 39, 0, 16, 54, 55, 74, 
    132, 21, 0, 94, 0, 82, 116, 89, 37, 0, 5, 0, 59, 55, 7, 
    76, 22, 33, 125, 0, 36, 75, 107, 27, 9, 0, 0, 41, 84, 0, 
    40, 29, 33, 104, 4, 45, 82, 83, 30, 20, 6, 0, 24, 71, 15, 
    39, 44, 93, 20, 54, 34, 78, 36, 47, 12, 16, 0, 18, 42, 63, 
    47, 45, 166, 0, 70, 41, 53, 81, 0, 48, 38, 0, 0, 27, 15, 
    59, 38, 97, 29, 41, 46, 83, 98, 18, 91, 31, 110, 0, 3, 0, 
    40, 49, 43, 48, 24, 22, 31, 83, 125, 33, 81, 56, 75, 62, 20, 
    21, 62, 0, 56, 43, 91, 0, 40, 70, 87, 59, 49, 54, 88, 61, 
    17, 54, 0, 45, 59, 95, 37, 59, 70, 123, 20, 61, 35, 89, 84, 
    23, 31, 0, 36, 95, 112, 12, 63, 80, 93, 21, 64, 46, 52, 68, 
    34, 35, 0, 6, 100, 118, 73, 67, 80, 76, 31, 60, 80, 31, 48, 
    30, 13, 8, 0, 62, 75, 95, 55, 88, 37, 49, 48, 76, 45, 44, 
    
    -- channel=557
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=558
    0, 181, 49, 0, 0, 10, 0, 9, 0, 0, 147, 28, 0, 0, 0, 
    0, 100, 106, 22, 7, 0, 13, 22, 0, 0, 204, 0, 0, 0, 0, 
    0, 33, 177, 27, 67, 0, 0, 24, 0, 13, 95, 22, 0, 0, 0, 
    0, 97, 152, 0, 99, 0, 0, 0, 12, 111, 13, 79, 0, 0, 27, 
    0, 70, 1, 0, 114, 1, 0, 0, 16, 71, 52, 81, 0, 0, 40, 
    0, 12, 0, 0, 63, 0, 0, 0, 15, 59, 45, 96, 0, 0, 0, 
    0, 0, 0, 24, 0, 14, 0, 34, 0, 36, 39, 93, 5, 0, 0, 
    0, 4, 0, 135, 0, 0, 0, 0, 26, 13, 0, 55, 61, 0, 3, 
    0, 9, 0, 73, 0, 6, 0, 0, 72, 0, 0, 0, 95, 0, 88, 
    0, 0, 15, 0, 16, 0, 0, 0, 0, 31, 0, 1, 17, 0, 38, 
    0, 0, 49, 0, 0, 0, 51, 8, 0, 0, 0, 25, 10, 0, 0, 
    0, 0, 85, 0, 0, 0, 30, 0, 0, 0, 62, 0, 17, 0, 0, 
    0, 0, 64, 0, 0, 0, 35, 0, 0, 0, 39, 0, 0, 0, 0, 
    0, 0, 61, 24, 0, 4, 0, 0, 0, 0, 24, 0, 0, 41, 6, 
    0, 0, 28, 59, 0, 0, 0, 0, 0, 28, 3, 3, 0, 20, 6, 
    
    -- channel=559
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=560
    17, 127, 128, 85, 101, 107, 93, 110, 94, 0, 178, 139, 115, 113, 105, 
    18, 72, 143, 113, 157, 102, 128, 137, 116, 33, 207, 158, 138, 130, 119, 
    15, 33, 176, 104, 203, 84, 83, 112, 96, 141, 178, 182, 170, 175, 162, 
    18, 128, 170, 74, 206, 156, 104, 72, 102, 169, 171, 220, 192, 148, 190, 
    122, 149, 153, 58, 188, 176, 134, 64, 112, 152, 193, 217, 197, 119, 158, 
    146, 154, 143, 101, 168, 156, 113, 98, 125, 155, 172, 233, 201, 129, 126, 
    140, 147, 83, 149, 129, 168, 112, 151, 127, 155, 178, 227, 205, 188, 137, 
    127, 146, 62, 204, 142, 147, 150, 104, 161, 132, 129, 152, 220, 170, 189, 
    109, 135, 150, 167, 189, 186, 150, 103, 138, 104, 132, 60, 140, 138, 199, 
    145, 140, 172, 157, 169, 173, 190, 165, 92, 143, 90, 112, 118, 101, 115, 
    168, 117, 197, 172, 173, 113, 177, 168, 150, 77, 116, 126, 128, 97, 91, 
    165, 118, 198, 189, 162, 129, 163, 155, 134, 69, 128, 111, 141, 97, 86, 
    152, 122, 176, 184, 109, 114, 162, 132, 104, 73, 119, 101, 101, 111, 93, 
    137, 104, 155, 198, 142, 130, 108, 103, 78, 77, 104, 95, 72, 112, 116, 
    118, 114, 115, 208, 158, 121, 73, 91, 49, 92, 92, 100, 86, 95, 105, 
    
    -- channel=561
    67, 66, 193, 167, 145, 180, 192, 194, 207, 107, 133, 203, 215, 216, 213, 
    67, 48, 150, 139, 149, 120, 143, 173, 152, 152, 178, 188, 190, 194, 194, 
    72, 57, 150, 145, 117, 107, 63, 63, 71, 151, 150, 140, 160, 176, 188, 
    210, 215, 224, 128, 88, 143, 168, 129, 113, 102, 129, 161, 154, 130, 145, 
    225, 208, 170, 145, 100, 94, 117, 98, 99, 88, 135, 169, 161, 163, 147, 
    174, 152, 159, 162, 128, 90, 86, 100, 128, 106, 110, 151, 162, 196, 182, 
    173, 160, 117, 168, 102, 95, 103, 117, 122, 113, 115, 156, 162, 199, 198, 
    162, 144, 141, 159, 131, 102, 110, 88, 130, 108, 104, 59, 138, 140, 176, 
    175, 131, 172, 122, 148, 169, 126, 123, 98, 123, 159, 150, 50, 85, 143, 
    194, 168, 137, 145, 98, 68, 107, 151, 156, 153, 112, 152, 166, 151, 92, 
    171, 140, 137, 142, 156, 116, 100, 94, 137, 112, 134, 151, 136, 125, 124, 
    155, 167, 131, 124, 118, 126, 151, 135, 124, 129, 151, 122, 138, 137, 138, 
    160, 168, 142, 116, 94, 55, 132, 117, 112, 122, 129, 118, 87, 116, 136, 
    159, 170, 142, 127, 148, 177, 121, 116, 110, 112, 129, 122, 116, 121, 146, 
    131, 182, 123, 106, 127, 120, 104, 120, 110, 127, 119, 133, 142, 133, 115, 
    
    -- channel=562
    3, 0, 0, 12, 0, 0, 0, 0, 0, 97, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 7, 159, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 110, 38, 0, 54, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 61, 0, 33, 0, 28, 0, 0, 0, 0, 0, 39, 0, 
    10, 0, 0, 124, 0, 0, 38, 109, 0, 0, 0, 0, 0, 93, 0, 
    0, 0, 5, 44, 0, 5, 79, 53, 0, 0, 0, 0, 0, 60, 0, 
    0, 0, 97, 0, 2, 0, 47, 0, 3, 0, 0, 0, 0, 0, 13, 
    27, 0, 112, 0, 17, 0, 30, 0, 0, 0, 9, 1, 0, 27, 0, 
    57, 0, 0, 0, 0, 0, 0, 84, 0, 38, 0, 35, 0, 55, 0, 
    19, 0, 0, 0, 0, 12, 0, 18, 0, 0, 68, 0, 0, 0, 0, 
    0, 42, 0, 0, 0, 77, 0, 0, 44, 69, 3, 0, 0, 50, 4, 
    0, 57, 0, 0, 12, 72, 0, 0, 22, 120, 0, 7, 0, 27, 33, 
    2, 41, 0, 0, 99, 51, 0, 23, 71, 67, 0, 17, 22, 19, 4, 
    24, 41, 0, 0, 61, 0, 39, 30, 60, 46, 0, 0, 46, 0, 0, 
    46, 4, 0, 0, 21, 36, 95, 13, 76, 0, 0, 0, 11, 0, 0, 
    
    -- channel=563
    104, 119, 141, 120, 115, 145, 140, 138, 109, 94, 116, 101, 125, 136, 136, 
    105, 113, 143, 112, 49, 85, 106, 112, 93, 98, 89, 96, 109, 119, 121, 
    106, 104, 143, 108, 29, 41, 87, 108, 109, 102, 69, 99, 85, 86, 92, 
    93, 111, 78, 112, 43, 36, 54, 71, 84, 73, 68, 76, 42, 64, 103, 
    116, 93, 102, 116, 54, 39, 47, 67, 78, 70, 81, 82, 74, 123, 140, 
    113, 106, 113, 116, 56, 40, 57, 79, 59, 58, 70, 93, 88, 131, 164, 
    132, 119, 117, 105, 68, 61, 47, 57, 50, 56, 70, 89, 88, 95, 130, 
    136, 113, 86, 77, 53, 47, 49, 40, 86, 81, 79, 119, 117, 93, 125, 
    135, 118, 62, 51, 53, 28, 26, 46, 97, 102, 85, 118, 126, 138, 139, 
    131, 110, 62, 66, 66, 51, 42, 41, 65, 89, 92, 115, 101, 97, 119, 
    116, 108, 78, 64, 66, 66, 71, 55, 63, 83, 119, 91, 79, 96, 103, 
    118, 123, 80, 44, 49, 67, 70, 66, 67, 106, 107, 91, 80, 92, 105, 
    125, 152, 113, 50, 49, 82, 79, 88, 92, 108, 109, 100, 91, 108, 99, 
    131, 166, 147, 61, 62, 55, 84, 107, 113, 125, 107, 106, 106, 110, 100, 
    148, 167, 152, 62, 64, 77, 108, 114, 116, 127, 113, 107, 110, 102, 106, 
    
    -- channel=564
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=565
    7, 0, 0, 47, 15, 6, 34, 3, 95, 122, 0, 0, 27, 25, 47, 
    0, 0, 0, 3, 0, 1, 0, 0, 16, 252, 0, 0, 23, 21, 39, 
    4, 0, 0, 0, 0, 155, 17, 0, 47, 29, 0, 0, 0, 0, 9, 
    87, 0, 0, 52, 0, 94, 71, 56, 0, 0, 0, 0, 0, 18, 0, 
    78, 0, 0, 163, 0, 0, 56, 134, 0, 0, 0, 0, 0, 108, 0, 
    2, 0, 1, 93, 0, 0, 94, 89, 0, 0, 0, 0, 0, 100, 0, 
    0, 0, 76, 0, 0, 0, 60, 0, 5, 0, 0, 0, 0, 26, 32, 
    18, 0, 184, 0, 17, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 
    74, 0, 68, 0, 11, 0, 11, 134, 0, 67, 0, 87, 0, 19, 0, 
    40, 0, 0, 3, 0, 0, 10, 73, 53, 0, 61, 17, 0, 0, 0, 
    0, 35, 0, 0, 0, 81, 0, 0, 80, 52, 45, 0, 0, 77, 4, 
    0, 76, 0, 0, 4, 96, 0, 0, 24, 171, 0, 8, 0, 53, 72, 
    0, 36, 0, 0, 104, 57, 0, 16, 78, 97, 0, 25, 0, 41, 27, 
    15, 41, 0, 0, 110, 0, 24, 37, 71, 67, 0, 14, 67, 0, 0, 
    31, 20, 0, 0, 36, 37, 102, 23, 97, 0, 0, 0, 51, 0, 0, 
    
    -- channel=566
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 82, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 93, 119, 0, 0, 0, 0, 44, 9, 21, 18, 0, 
    32, 0, 5, 0, 56, 132, 75, 25, 0, 0, 80, 40, 100, 87, 18, 
    41, 16, 26, 0, 25, 91, 87, 51, 17, 1, 42, 42, 73, 29, 0, 
    13, 7, 14, 0, 49, 88, 70, 26, 71, 39, 41, 36, 83, 52, 0, 
    0, 0, 0, 0, 34, 48, 97, 43, 105, 73, 49, 34, 69, 95, 31, 
    0, 0, 0, 0, 94, 94, 105, 72, 28, 6, 43, 0, 10, 69, 34, 
    28, 0, 2, 0, 110, 138, 122, 107, 0, 0, 17, 0, 0, 0, 0, 
    45, 13, 46, 53, 49, 80, 116, 118, 38, 0, 0, 0, 0, 0, 0, 
    46, 45, 45, 54, 67, 65, 20, 49, 75, 0, 0, 0, 0, 0, 0, 
    33, 51, 26, 91, 79, 17, 23, 28, 34, 0, 0, 0, 0, 0, 0, 
    28, 3, 0, 92, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 93, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 87, 76, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=567
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=568
    0, 20, 0, 0, 8, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    0, 32, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 12, 0, 0, 11, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 6, 0, 8, 0, 0, 0, 4, 0, 0, 0, 0, 0, 8, 4, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 2, 0, 0, 0, 7, 4, 
    0, 1, 12, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 13, 
    8, 5, 16, 0, 0, 2, 0, 29, 0, 8, 9, 0, 0, 0, 5, 
    5, 2, 0, 0, 0, 0, 6, 0, 0, 17, 0, 26, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 2, 0, 9, 
    0, 16, 0, 0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 5, 0, 
    4, 0, 0, 0, 0, 19, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    6, 6, 0, 0, 0, 18, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    7, 0, 13, 0, 1, 3, 9, 0, 0, 4, 0, 0, 0, 0, 0, 
    
    -- channel=569
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=570
    121, 123, 28, 27, 16, 26, 16, 23, 25, 27, 96, 5, 0, 0, 0, 
    121, 119, 49, 50, 24, 8, 26, 19, 2, 26, 71, 0, 0, 0, 0, 
    119, 117, 88, 34, 26, 0, 34, 30, 27, 61, 13, 0, 0, 0, 0, 
    55, 113, 37, 4, 40, 0, 19, 33, 53, 57, 0, 10, 0, 0, 0, 
    5, 28, 0, 8, 42, 3, 0, 19, 52, 54, 14, 0, 0, 0, 0, 
    0, 0, 0, 10, 27, 4, 1, 40, 40, 46, 15, 0, 0, 0, 0, 
    0, 0, 0, 22, 10, 22, 0, 54, 14, 34, 15, 0, 0, 0, 0, 
    0, 5, 0, 43, 0, 10, 18, 6, 39, 20, 4, 9, 4, 0, 0, 
    0, 16, 11, 13, 2, 0, 0, 0, 42, 24, 11, 24, 26, 0, 13, 
    0, 6, 0, 0, 0, 0, 2, 5, 0, 24, 6, 32, 38, 13, 20, 
    0, 0, 14, 0, 0, 0, 14, 0, 0, 0, 45, 29, 19, 17, 26, 
    0, 0, 18, 0, 0, 4, 8, 2, 0, 12, 45, 23, 21, 14, 34, 
    0, 0, 19, 0, 0, 36, 6, 1, 2, 25, 41, 31, 22, 38, 31, 
    0, 0, 28, 0, 0, 15, 2, 16, 19, 50, 42, 37, 36, 53, 32, 
    1, 4, 29, 11, 0, 0, 14, 39, 34, 62, 47, 39, 44, 41, 39, 
    
    -- channel=571
    0, 148, 351, 302, 298, 322, 324, 336, 291, 102, 281, 402, 403, 396, 386, 
    0, 46, 314, 309, 351, 301, 336, 375, 366, 157, 395, 446, 433, 425, 414, 
    0, 0, 275, 319, 439, 280, 215, 276, 264, 277, 414, 443, 457, 470, 456, 
    55, 137, 373, 287, 427, 378, 285, 203, 210, 344, 413, 507, 524, 452, 464, 
    331, 381, 400, 234, 391, 416, 363, 212, 226, 311, 419, 535, 528, 383, 408, 
    403, 407, 395, 307, 396, 392, 313, 220, 267, 321, 390, 539, 531, 402, 355, 
    401, 396, 314, 377, 334, 354, 303, 309, 315, 334, 390, 536, 540, 503, 395, 
    381, 395, 291, 448, 394, 374, 333, 311, 337, 332, 350, 391, 524, 498, 470, 
    349, 343, 389, 441, 446, 454, 392, 281, 311, 298, 341, 228, 331, 355, 460, 
    398, 376, 441, 418, 426, 442, 449, 392, 308, 352, 287, 295, 307, 306, 324, 
    441, 362, 441, 450, 452, 349, 405, 426, 388, 295, 268, 325, 346, 281, 265, 
    439, 352, 448, 482, 456, 370, 420, 415, 383, 235, 306, 308, 354, 295, 238, 
    413, 348, 417, 462, 361, 302, 414, 380, 319, 231, 288, 273, 279, 269, 258, 
    386, 312, 366, 466, 385, 389, 340, 305, 249, 194, 255, 250, 202, 253, 292, 
    323, 302, 299, 454, 413, 365, 251, 254, 174, 203, 226, 251, 219, 248, 263, 
    
    -- channel=572
    0, 187, 538, 449, 450, 487, 487, 497, 440, 182, 369, 571, 563, 569, 552, 
    0, 89, 509, 424, 504, 439, 520, 571, 545, 289, 510, 652, 617, 606, 589, 
    0, 26, 424, 416, 591, 444, 337, 435, 445, 414, 605, 674, 679, 682, 662, 
    98, 143, 536, 468, 595, 546, 398, 318, 315, 451, 649, 715, 736, 712, 718, 
    555, 578, 638, 413, 521, 586, 540, 362, 348, 424, 630, 788, 785, 657, 668, 
    651, 635, 662, 481, 564, 568, 487, 327, 395, 432, 579, 806, 826, 712, 643, 
    666, 625, 526, 586, 484, 476, 458, 429, 482, 497, 554, 797, 829, 804, 666, 
    656, 619, 436, 615, 579, 563, 489, 438, 538, 482, 567, 639, 838, 806, 761, 
    643, 539, 515, 562, 650, 640, 529, 443, 427, 452, 545, 380, 499, 631, 745, 
    695, 590, 631, 619, 620, 650, 656, 555, 435, 502, 465, 452, 428, 481, 515, 
    731, 609, 655, 640, 659, 547, 587, 602, 593, 480, 415, 467, 505, 429, 418, 
    722, 637, 650, 687, 669, 545, 604, 588, 573, 395, 449, 466, 528, 450, 381, 
    701, 645, 650, 671, 566, 346, 610, 567, 505, 385, 448, 423, 439, 430, 403, 
    674, 613, 608, 695, 575, 475, 518, 477, 408, 323, 403, 390, 337, 381, 445, 
    597, 600, 516, 684, 620, 558, 429, 414, 321, 326, 365, 397, 349, 383, 417, 
    
    -- channel=573
    0, 18, 336, 337, 320, 344, 357, 351, 328, 202, 146, 375, 400, 405, 404, 
    0, 0, 287, 289, 307, 317, 341, 365, 383, 276, 202, 438, 440, 432, 427, 
    0, 0, 183, 283, 328, 348, 251, 296, 327, 252, 343, 441, 457, 454, 451, 
    99, 23, 267, 364, 319, 369, 270, 239, 204, 226, 409, 418, 475, 496, 460, 
    397, 329, 425, 358, 275, 371, 375, 292, 213, 229, 377, 469, 524, 507, 441, 
    450, 422, 459, 359, 330, 366, 354, 241, 233, 232, 348, 480, 552, 537, 459, 
    471, 429, 419, 367, 332, 301, 336, 244, 315, 292, 334, 467, 549, 550, 479, 
    480, 419, 364, 330, 398, 354, 331, 281, 320, 318, 373, 425, 506, 564, 500, 
    488, 373, 354, 332, 409, 393, 350, 341, 259, 317, 361, 284, 326, 452, 453, 
    500, 398, 403, 405, 407, 432, 411, 365, 310, 314, 353, 308, 272, 338, 341, 
    500, 447, 398, 419, 426, 405, 359, 389, 412, 368, 280, 302, 328, 322, 297, 
    492, 474, 385, 444, 449, 390, 370, 385, 395, 332, 266, 322, 336, 323, 277, 
    488, 478, 404, 435, 435, 247, 383, 392, 378, 300, 281, 296, 309, 294, 284, 
    481, 460, 390, 436, 420, 294, 371, 343, 315, 242, 265, 269, 258, 234, 294, 
    437, 432, 358, 402, 422, 403, 340, 290, 266, 201, 249, 266, 247, 250, 280, 
    
    -- channel=574
    0, 0, 151, 154, 154, 146, 164, 153, 177, 94, 27, 212, 213, 205, 206, 
    0, 0, 101, 123, 196, 173, 168, 188, 216, 162, 76, 253, 246, 234, 230, 
    0, 0, 27, 127, 211, 242, 117, 117, 147, 117, 186, 234, 264, 265, 262, 
    56, 0, 130, 182, 184, 262, 189, 138, 94, 105, 242, 238, 318, 304, 243, 
    220, 171, 231, 186, 146, 242, 247, 174, 101, 110, 210, 263, 322, 277, 192, 
    237, 220, 240, 189, 189, 234, 225, 131, 138, 129, 195, 254, 324, 291, 194, 
    234, 218, 217, 187, 191, 176, 218, 142, 203, 167, 190, 258, 316, 325, 250, 
    236, 212, 229, 169, 254, 221, 212, 189, 171, 170, 208, 181, 257, 322, 257, 
    246, 172, 235, 199, 264, 276, 248, 237, 111, 165, 203, 137, 106, 204, 196, 
    260, 203, 245, 244, 235, 259, 266, 256, 203, 165, 195, 147, 137, 179, 143, 
    264, 237, 222, 262, 262, 254, 197, 234, 263, 211, 122, 156, 183, 173, 141, 
    254, 249, 200, 286, 290, 245, 220, 236, 242, 183, 114, 167, 187, 178, 139, 
    248, 224, 187, 274, 282, 135, 212, 219, 208, 146, 121, 144, 153, 139, 141, 
    240, 200, 145, 262, 277, 199, 209, 170, 150, 92, 112, 123, 119, 91, 146, 
    192, 179, 119, 232, 262, 238, 171, 127, 115, 58, 102, 120, 114, 110, 126, 
    
    -- channel=575
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=576
    159, 162, 142, 116, 132, 122, 143, 159, 181, 181, 178, 186, 148, 179, 153, 
    165, 167, 148, 46, 66, 64, 70, 93, 134, 182, 186, 186, 182, 176, 214, 
    164, 165, 133, 0, 0, 0, 0, 0, 0, 18, 186, 178, 157, 157, 231, 
    163, 153, 124, 0, 49, 59, 0, 0, 0, 0, 48, 194, 156, 142, 162, 
    168, 148, 73, 0, 16, 0, 0, 0, 0, 0, 0, 143, 173, 133, 133, 
    174, 135, 52, 0, 5, 0, 0, 0, 0, 0, 14, 72, 181, 164, 164, 
    139, 92, 83, 0, 0, 0, 0, 0, 0, 0, 1, 67, 136, 166, 177, 
    120, 37, 122, 32, 0, 0, 0, 0, 0, 0, 0, 9, 34, 30, 191, 
    96, 5, 109, 2, 12, 37, 17, 0, 5, 27, 0, 4, 28, 15, 166, 
    100, 0, 87, 0, 16, 0, 3, 51, 14, 20, 9, 16, 41, 0, 127, 
    108, 0, 19, 0, 0, 16, 6, 0, 42, 0, 0, 20, 0, 13, 98, 
    71, 0, 65, 5, 0, 5, 44, 0, 88, 54, 39, 71, 0, 32, 105, 
    44, 0, 8, 23, 0, 0, 4, 7, 19, 136, 74, 0, 0, 21, 84, 
    50, 29, 0, 24, 0, 0, 5, 13, 33, 75, 63, 0, 0, 35, 71, 
    20, 10, 0, 0, 3, 0, 2, 3, 7, 12, 27, 0, 0, 27, 82, 
    
    -- channel=577
    74, 60, 102, 96, 101, 97, 66, 43, 55, 81, 72, 81, 66, 35, 35, 
    100, 96, 124, 140, 153, 160, 153, 170, 172, 111, 70, 87, 94, 69, 43, 
    110, 112, 132, 145, 118, 117, 111, 109, 116, 102, 70, 86, 106, 83, 29, 
    110, 120, 115, 187, 134, 157, 157, 164, 155, 132, 86, 110, 99, 85, 48, 
    113, 126, 150, 195, 139, 144, 186, 159, 159, 146, 152, 96, 94, 96, 52, 
    128, 154, 137, 161, 118, 144, 160, 161, 158, 146, 156, 101, 97, 110, 110, 
    135, 172, 148, 144, 102, 156, 184, 147, 151, 168, 129, 110, 136, 149, 122, 
    171, 159, 116, 156, 159, 124, 121, 148, 145, 131, 138, 138, 121, 134, 118, 
    140, 128, 107, 157, 119, 131, 122, 87, 35, 21, 61, 16, 40, 131, 91, 
    142, 142, 137, 96, 108, 119, 104, 127, 157, 146, 163, 149, 172, 143, 65, 
    143, 150, 85, 103, 83, 87, 69, 108, 97, 110, 111, 79, 111, 118, 52, 
    165, 166, 105, 94, 86, 65, 106, 140, 77, 139, 114, 144, 138, 119, 54, 
    158, 126, 61, 149, 109, 72, 62, 60, 50, 62, 99, 154, 90, 65, 42, 
    148, 172, 152, 151, 117, 99, 47, 52, 69, 100, 147, 195, 81, 58, 66, 
    161, 149, 152, 125, 109, 94, 57, 65, 72, 94, 121, 166, 67, 59, 52, 
    
    -- channel=578
    317, 319, 323, 244, 259, 298, 299, 327, 333, 308, 290, 303, 300, 275, 241, 
    354, 353, 329, 207, 212, 225, 210, 200, 221, 223, 229, 309, 305, 233, 258, 
    354, 354, 322, 221, 268, 315, 314, 304, 276, 235, 249, 332, 294, 205, 207, 
    353, 344, 316, 226, 306, 349, 326, 295, 315, 322, 281, 274, 305, 268, 216, 
    353, 339, 252, 201, 287, 276, 259, 291, 295, 300, 302, 321, 356, 335, 351, 
    343, 316, 296, 221, 197, 256, 256, 238, 232, 255, 240, 263, 337, 355, 356, 
    338, 265, 252, 236, 289, 280, 262, 238, 254, 251, 196, 206, 240, 266, 352, 
    315, 186, 266, 269, 222, 209, 187, 158, 119, 123, 121, 111, 177, 251, 343, 
    331, 212, 276, 115, 221, 220, 259, 253, 296, 320, 308, 287, 333, 287, 335, 
    325, 169, 176, 124, 164, 152, 152, 194, 240, 219, 204, 206, 223, 176, 296, 
    328, 186, 187, 146, 112, 131, 243, 165, 201, 211, 203, 271, 173, 252, 298, 
    327, 133, 157, 248, 134, 94, 100, 66, 159, 195, 244, 225, 109, 131, 245, 
    322, 281, 262, 237, 162, 97, 71, 87, 121, 301, 335, 245, 99, 137, 292, 
    324, 296, 239, 206, 181, 111, 89, 109, 151, 197, 216, 179, 74, 156, 280, 
    299, 290, 253, 161, 160, 122, 117, 129, 142, 168, 198, 169, 99, 146, 308, 
    
    -- channel=579
    163, 168, 170, 73, 94, 101, 114, 154, 192, 173, 161, 169, 132, 131, 81, 
    210, 210, 189, 26, 56, 79, 66, 77, 119, 111, 117, 181, 172, 103, 137, 
    218, 219, 171, 0, 45, 84, 74, 64, 61, 68, 120, 193, 153, 70, 101, 
    216, 212, 154, 3, 130, 148, 115, 107, 107, 108, 122, 167, 139, 102, 69, 
    215, 201, 100, 0, 99, 103, 62, 94, 112, 109, 116, 171, 203, 158, 147, 
    203, 181, 75, 0, 5, 49, 47, 41, 39, 68, 73, 108, 219, 218, 219, 
    177, 96, 67, 0, 43, 57, 43, 7, 38, 54, 0, 50, 130, 153, 220, 
    140, 0, 62, 54, 4, 0, 0, 0, 0, 0, 0, 0, 0, 78, 224, 
    120, 0, 93, 0, 10, 15, 14, 0, 13, 35, 16, 0, 81, 77, 184, 
    132, 0, 4, 0, 0, 0, 0, 23, 46, 53, 34, 33, 70, 0, 135, 
    148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 31, 103, 
    144, 0, 0, 3, 0, 0, 0, 0, 0, 0, 32, 77, 0, 0, 66, 
    129, 2, 21, 42, 0, 0, 0, 0, 0, 114, 113, 22, 0, 0, 94, 
    138, 100, 21, 11, 0, 0, 0, 0, 0, 41, 58, 0, 0, 0, 81, 
    106, 87, 38, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 115, 
    
    -- channel=580
    189, 194, 181, 156, 135, 129, 148, 181, 203, 200, 203, 188, 186, 201, 180, 
    197, 198, 193, 124, 87, 79, 89, 97, 118, 158, 179, 187, 190, 203, 192, 
    196, 196, 175, 114, 21, 53, 49, 59, 51, 80, 143, 181, 192, 178, 181, 
    196, 196, 162, 87, 55, 87, 95, 61, 67, 60, 130, 156, 166, 182, 168, 
    191, 190, 142, 50, 44, 68, 52, 48, 62, 70, 82, 134, 182, 180, 170, 
    162, 180, 117, 56, 14, 29, 40, 33, 33, 48, 57, 91, 160, 196, 196, 
    142, 125, 97, 48, 37, 40, 22, 23, 26, 45, 56, 74, 115, 135, 182, 
    130, 82, 66, 105, 22, 22, 16, 24, 6, 0, 13, 14, 10, 56, 135, 
    130, 82, 95, 36, 26, 53, 48, 39, 64, 75, 83, 73, 82, 75, 108, 
    139, 91, 48, 36, 17, 26, 28, 40, 61, 57, 57, 52, 65, 42, 74, 
    135, 81, 48, 27, 23, 1, 23, 61, 11, 50, 34, 47, 47, 38, 82, 
    119, 79, 14, 51, 40, 25, 26, 2, 37, 52, 63, 93, 40, 25, 45, 
    88, 72, 76, 62, 33, 29, 6, 6, 10, 75, 128, 103, 27, 4, 58, 
    103, 89, 68, 57, 34, 28, 13, 15, 30, 55, 59, 69, 14, 17, 47, 
    80, 76, 73, 38, 31, 22, 23, 22, 23, 28, 38, 24, 25, 15, 55, 
    
    -- channel=581
    63, 51, 68, 85, 37, 34, 39, 29, 24, 53, 52, 36, 85, 39, 71, 
    63, 59, 83, 140, 24, 7, 12, 15, 0, 0, 32, 13, 45, 72, 6, 
    61, 58, 99, 205, 10, 46, 61, 83, 57, 11, 0, 28, 63, 67, 0, 
    61, 70, 76, 217, 0, 37, 112, 61, 67, 59, 25, 0, 65, 84, 20, 
    52, 79, 110, 158, 0, 22, 85, 44, 40, 48, 79, 0, 27, 109, 69, 
    11, 87, 115, 164, 0, 34, 58, 35, 33, 16, 19, 0, 0, 62, 58, 
    12, 96, 36, 114, 40, 39, 70, 49, 19, 35, 45, 0, 0, 0, 24, 
    46, 104, 0, 100, 58, 53, 39, 41, 0, 0, 9, 0, 0, 0, 0, 
    77, 145, 0, 112, 0, 12, 38, 92, 42, 28, 111, 60, 0, 43, 0, 
    86, 174, 0, 83, 0, 35, 0, 0, 47, 11, 42, 24, 17, 75, 0, 
    60, 207, 2, 44, 16, 0, 0, 76, 0, 59, 27, 0, 81, 0, 0, 
    66, 200, 0, 31, 88, 0, 0, 71, 0, 25, 23, 0, 115, 0, 0, 
    51, 170, 26, 31, 83, 51, 0, 0, 0, 0, 69, 140, 59, 0, 0, 
    42, 78, 98, 40, 30, 79, 0, 0, 0, 0, 0, 134, 48, 0, 0, 
    62, 66, 95, 67, 15, 43, 9, 1, 0, 0, 0, 72, 50, 0, 0, 
    
    -- channel=582
    163, 171, 156, 126, 129, 141, 146, 162, 175, 162, 158, 162, 151, 163, 141, 
    171, 172, 152, 90, 98, 100, 104, 102, 110, 129, 144, 167, 160, 139, 161, 
    169, 169, 146, 68, 103, 114, 109, 107, 108, 116, 153, 172, 151, 122, 159, 
    169, 162, 149, 61, 112, 122, 102, 92, 97, 107, 137, 156, 151, 138, 142, 
    168, 156, 113, 52, 106, 102, 77, 91, 96, 104, 101, 163, 176, 158, 174, 
    163, 138, 109, 58, 83, 83, 79, 72, 74, 87, 86, 125, 171, 169, 171, 
    159, 113, 114, 70, 104, 90, 64, 71, 80, 77, 71, 102, 130, 138, 168, 
    132, 81, 128, 93, 74, 68, 67, 47, 38, 42, 40, 44, 80, 113, 172, 
    142, 81, 137, 51, 82, 83, 90, 91, 123, 140, 114, 127, 150, 100, 174, 
    137, 58, 91, 51, 81, 61, 79, 88, 96, 96, 83, 90, 89, 68, 162, 
    142, 54, 90, 61, 58, 66, 103, 64, 98, 82, 79, 118, 72, 88, 158, 
    131, 36, 80, 98, 54, 61, 67, 17, 100, 78, 101, 99, 34, 75, 136, 
    121, 78, 122, 90, 56, 51, 49, 57, 75, 139, 134, 73, 46, 72, 157, 
    125, 107, 78, 75, 71, 42, 59, 66, 78, 117, 99, 49, 39, 89, 139, 
    109, 106, 86, 67, 68, 52, 67, 70, 75, 80, 89, 51, 52, 84, 152, 
    
    -- channel=583
    0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 1, 0, 16, 0, 18, 
    0, 0, 11, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 
    0, 0, 25, 139, 0, 0, 0, 4, 0, 0, 0, 0, 9, 24, 0, 
    0, 0, 16, 146, 0, 0, 41, 0, 0, 0, 0, 0, 0, 30, 0, 
    0, 5, 72, 94, 0, 0, 21, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 21, 57, 106, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 42, 10, 55, 2, 0, 11, 2, 0, 0, 5, 0, 0, 0, 0, 
    1, 81, 0, 57, 12, 0, 0, 17, 0, 0, 6, 0, 0, 0, 0, 
    25, 108, 0, 98, 0, 2, 0, 25, 0, 0, 26, 0, 0, 9, 0, 
    20, 141, 0, 74, 0, 9, 0, 0, 0, 0, 0, 0, 0, 37, 0, 
    0, 153, 0, 18, 15, 0, 0, 59, 0, 22, 0, 0, 68, 0, 0, 
    1, 157, 0, 0, 62, 0, 0, 49, 0, 0, 0, 0, 91, 0, 0, 
    0, 76, 0, 0, 41, 40, 0, 0, 0, 0, 6, 67, 54, 0, 0, 
    0, 11, 42, 0, 1, 50, 0, 0, 0, 0, 0, 56, 45, 0, 0, 
    0, 1, 26, 37, 0, 22, 0, 0, 0, 0, 0, 17, 44, 0, 0, 
    
    -- channel=584
    582, 574, 564, 467, 435, 444, 491, 550, 595, 605, 588, 578, 574, 563, 520, 
    626, 625, 610, 400, 304, 301, 304, 337, 399, 472, 522, 560, 580, 563, 548, 
    623, 622, 583, 345, 194, 265, 265, 274, 248, 279, 433, 577, 564, 496, 490, 
    621, 614, 532, 353, 272, 399, 371, 304, 317, 331, 395, 484, 547, 538, 444, 
    612, 609, 451, 251, 236, 277, 275, 264, 299, 309, 365, 457, 583, 596, 548, 
    546, 576, 413, 237, 119, 196, 212, 191, 191, 219, 261, 328, 524, 624, 623, 
    478, 439, 333, 255, 217, 218, 210, 171, 193, 245, 211, 245, 370, 464, 592, 
    445, 278, 287, 343, 154, 129, 108, 104, 54, 45, 69, 63, 106, 234, 483, 
    466, 295, 295, 168, 160, 228, 241, 230, 262, 295, 333, 274, 288, 302, 406, 
    485, 276, 197, 116, 101, 116, 99, 174, 259, 227, 235, 222, 270, 180, 285, 
    478, 299, 162, 114, 56, 60, 155, 156, 114, 187, 154, 211, 179, 205, 287, 
    441, 235, 129, 219, 126, 38, 61, 66, 117, 229, 263, 295, 133, 102, 191, 
    377, 328, 239, 254, 155, 74, 14, 21, 46, 310, 447, 355, 81, 62, 211, 
    388, 364, 276, 235, 159, 105, 36, 52, 105, 186, 256, 273, 48, 70, 207, 
    344, 328, 299, 168, 134, 103, 75, 78, 86, 113, 154, 186, 68, 67, 231, 
    
    -- channel=585
    228, 218, 230, 172, 203, 224, 241, 260, 259, 237, 208, 217, 203, 174, 164, 
    286, 281, 271, 260, 352, 392, 372, 363, 352, 258, 185, 214, 206, 134, 160, 
    296, 298, 276, 289, 509, 550, 559, 549, 524, 433, 273, 222, 181, 106, 119, 
    294, 292, 282, 363, 553, 525, 564, 658, 635, 616, 414, 246, 196, 136, 96, 
    287, 287, 315, 440, 560, 580, 584, 644, 623, 620, 567, 356, 270, 216, 184, 
    265, 273, 309, 421, 468, 548, 572, 582, 565, 572, 554, 436, 337, 297, 295, 
    231, 206, 208, 336, 509, 575, 596, 532, 554, 540, 406, 375, 335, 318, 308, 
    162, 145, 192, 244, 490, 417, 413, 403, 379, 374, 372, 365, 407, 437, 364, 
    192, 187, 198, 210, 405, 366, 409, 329, 288, 317, 300, 262, 368, 433, 369, 
    237, 218, 214, 220, 339, 329, 340, 394, 384, 422, 415, 401, 411, 364, 392, 
    262, 229, 230, 253, 239, 293, 361, 308, 344, 349, 366, 363, 318, 400, 374, 
    359, 239, 247, 317, 234, 222, 292, 245, 291, 303, 337, 340, 251, 294, 371, 
    430, 345, 306, 348, 290, 202, 188, 206, 235, 352, 342, 309, 221, 255, 402, 
    427, 416, 378, 325, 339, 226, 178, 209, 254, 319, 375, 315, 189, 277, 435, 
    471, 459, 395, 304, 317, 245, 209, 230, 255, 298, 344, 312, 194, 262, 450, 
    
    -- channel=586
    23, 32, 18, 46, 52, 30, 24, 21, 24, 29, 42, 41, 21, 47, 45, 
    9, 10, 4, 29, 27, 22, 36, 36, 43, 56, 67, 46, 43, 56, 78, 
    9, 10, 2, 0, 0, 0, 0, 0, 0, 0, 62, 29, 38, 68, 107, 
    9, 6, 17, 0, 0, 0, 0, 0, 0, 0, 0, 65, 30, 37, 87, 
    15, 3, 24, 0, 0, 0, 0, 0, 0, 0, 0, 10, 23, 0, 21, 
    38, 9, 10, 0, 6, 0, 0, 0, 0, 0, 0, 0, 26, 8, 9, 
    38, 30, 55, 0, 0, 0, 0, 0, 0, 0, 0, 39, 48, 54, 15, 
    47, 66, 77, 23, 0, 0, 0, 2, 34, 32, 27, 48, 40, 11, 23, 
    26, 31, 65, 57, 7, 28, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    14, 24, 66, 59, 40, 23, 40, 58, 0, 12, 0, 8, 7, 8, 53, 
    19, 4, 35, 39, 58, 56, 9, 9, 37, 0, 0, 0, 14, 1, 40, 
    0, 9, 67, 0, 20, 78, 87, 47, 93, 37, 6, 31, 46, 48, 83, 
    0, 0, 12, 0, 8, 45, 77, 73, 70, 37, 0, 0, 48, 63, 52, 
    0, 0, 0, 5, 16, 25, 71, 69, 67, 49, 32, 0, 67, 72, 36, 
    0, 0, 0, 14, 26, 35, 57, 53, 51, 42, 37, 0, 53, 66, 33, 
    
    -- channel=587
    249, 240, 253, 230, 201, 191, 202, 209, 253, 273, 270, 261, 244, 234, 224, 
    278, 276, 291, 239, 177, 170, 168, 203, 230, 238, 252, 247, 272, 273, 235, 
    284, 283, 288, 195, 60, 86, 81, 91, 93, 109, 150, 264, 270, 257, 213, 
    282, 291, 244, 220, 93, 181, 198, 138, 130, 125, 179, 211, 253, 244, 219, 
    281, 290, 261, 147, 106, 129, 141, 121, 137, 132, 168, 177, 255, 268, 191, 
    255, 299, 187, 146, 71, 91, 94, 105, 110, 98, 139, 159, 206, 285, 283, 
    230, 257, 186, 121, 68, 96, 118, 82, 80, 137, 120, 118, 201, 232, 272, 
    253, 193, 108, 212, 81, 72, 47, 65, 76, 69, 58, 79, 87, 102, 195, 
    222, 154, 143, 150, 55, 114, 112, 99, 32, 42, 116, 46, 52, 141, 178, 
    237, 169, 135, 51, 72, 68, 63, 60, 175, 113, 141, 126, 153, 107, 72, 
    229, 171, 78, 62, 32, 35, 31, 92, 49, 92, 68, 57, 100, 69, 87, 
    218, 168, 69, 74, 69, 25, 60, 80, 44, 134, 128, 169, 103, 95, 24, 
    184, 126, 66, 146, 74, 36, 14, 13, 4, 71, 201, 205, 65, 20, 31, 
    170, 195, 145, 149, 82, 66, 10, 11, 38, 123, 129, 187, 30, 14, 49, 
    173, 153, 147, 108, 74, 61, 27, 27, 33, 53, 85, 134, 38, 19, 34, 
    
    -- channel=588
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 5, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=589
    226, 220, 213, 179, 192, 191, 198, 213, 254, 260, 247, 255, 202, 216, 193, 
    258, 258, 240, 159, 203, 222, 230, 262, 289, 301, 256, 257, 254, 227, 249, 
    267, 269, 234, 61, 139, 124, 120, 109, 123, 177, 257, 250, 225, 206, 262, 
    266, 257, 227, 84, 221, 248, 181, 203, 185, 187, 220, 277, 226, 174, 200, 
    270, 249, 205, 116, 196, 211, 183, 193, 209, 215, 199, 256, 265, 197, 153, 
    272, 240, 153, 72, 169, 155, 142, 171, 174, 181, 210, 243, 285, 268, 268, 
    230, 186, 168, 93, 107, 153, 154, 129, 156, 191, 160, 210, 287, 304, 297, 
    195, 121, 179, 110, 139, 99, 85, 96, 135, 132, 108, 156, 194, 194, 311, 
    158, 75, 178, 96, 147, 155, 158, 71, 29, 65, 47, 20, 85, 154, 314, 
    184, 59, 171, 45, 135, 95, 125, 184, 183, 172, 176, 172, 189, 123, 262, 
    204, 47, 86, 68, 58, 104, 97, 53, 160, 79, 97, 116, 67, 130, 226, 
    207, 53, 134, 83, 29, 70, 161, 83, 176, 175, 146, 197, 91, 145, 228, 
    199, 49, 71, 140, 61, 22, 51, 61, 78, 203, 174, 95, 54, 89, 198, 
    192, 186, 121, 129, 109, 39, 38, 57, 97, 202, 202, 104, 36, 100, 206, 
    192, 172, 122, 96, 105, 66, 51, 59, 75, 103, 149, 112, 30, 93, 205, 
    
    -- channel=590
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 22, 
    0, 0, 8, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 
    0, 0, 18, 137, 0, 0, 0, 0, 0, 0, 0, 0, 4, 37, 0, 
    0, 0, 1, 133, 0, 0, 27, 0, 0, 0, 0, 0, 1, 24, 0, 
    0, 2, 47, 84, 0, 0, 6, 0, 0, 0, 0, 0, 0, 24, 0, 
    0, 18, 45, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 69, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 88, 0, 78, 0, 0, 0, 18, 0, 0, 24, 0, 0, 0, 0, 
    14, 122, 0, 63, 0, 3, 0, 0, 0, 0, 0, 0, 0, 24, 0, 
    0, 138, 0, 12, 0, 0, 0, 27, 0, 0, 0, 0, 14, 0, 0, 
    0, 147, 0, 0, 50, 0, 0, 61, 0, 2, 0, 0, 98, 0, 0, 
    0, 86, 0, 0, 39, 23, 0, 0, 0, 0, 0, 77, 36, 0, 0, 
    0, 1, 36, 0, 0, 49, 0, 0, 0, 0, 0, 73, 33, 0, 0, 
    0, 0, 20, 17, 0, 15, 0, 0, 0, 0, 0, 23, 27, 0, 0, 
    
    -- channel=591
    495, 489, 476, 333, 385, 391, 440, 502, 523, 506, 479, 501, 476, 462, 424, 
    529, 530, 486, 217, 252, 277, 245, 263, 348, 417, 438, 499, 489, 425, 500, 
    526, 526, 459, 170, 259, 281, 275, 259, 232, 250, 452, 508, 439, 371, 440, 
    525, 508, 428, 182, 353, 388, 287, 295, 313, 324, 312, 475, 461, 414, 341, 
    523, 498, 290, 155, 294, 255, 244, 263, 288, 296, 337, 443, 523, 490, 484, 
    498, 446, 334, 106, 157, 225, 192, 186, 186, 235, 243, 315, 534, 526, 528, 
    417, 307, 258, 214, 222, 198, 201, 159, 207, 226, 168, 247, 345, 415, 541, 
    356, 128, 331, 241, 154, 132, 118, 84, 54, 62, 58, 64, 163, 242, 536, 
    366, 151, 301, 26, 222, 205, 238, 200, 294, 312, 299, 281, 320, 257, 433, 
    391, 90, 206, 59, 120, 101, 105, 209, 208, 213, 190, 201, 258, 111, 377, 
    402, 123, 143, 105, 36, 101, 220, 56, 211, 153, 168, 286, 79, 267, 309, 
    364, 31, 191, 232, 43, 40, 74, 34, 166, 211, 258, 245, 35, 103, 305, 
    339, 265, 207, 241, 121, 26, 27, 46, 81, 451, 383, 244, 8, 117, 307, 
    353, 294, 207, 206, 151, 48, 50, 75, 136, 194, 261, 164, 18, 133, 294, 
    297, 291, 237, 93, 133, 80, 78, 92, 102, 130, 167, 152, 18, 126, 359, 
    
    -- channel=592
    719, 710, 710, 573, 559, 577, 613, 674, 736, 744, 713, 722, 687, 650, 592, 
    805, 802, 764, 519, 466, 496, 496, 526, 591, 629, 633, 709, 729, 644, 653, 
    815, 814, 752, 444, 407, 485, 496, 483, 453, 457, 597, 731, 692, 567, 578, 
    813, 798, 713, 484, 519, 654, 606, 572, 576, 579, 572, 661, 691, 611, 516, 
    808, 785, 623, 420, 479, 532, 521, 528, 560, 576, 600, 657, 769, 734, 670, 
    759, 745, 586, 376, 323, 435, 437, 427, 426, 461, 499, 557, 746, 816, 816, 
    673, 598, 497, 406, 413, 449, 448, 374, 411, 457, 368, 420, 569, 678, 800, 
    619, 394, 456, 477, 365, 311, 274, 246, 201, 200, 195, 203, 311, 465, 734, 
    618, 384, 443, 265, 333, 384, 416, 359, 359, 409, 426, 343, 433, 494, 656, 
    655, 353, 323, 188, 241, 240, 246, 374, 448, 433, 431, 415, 470, 335, 537, 
    664, 378, 245, 200, 129, 176, 313, 250, 299, 336, 309, 394, 304, 379, 513, 
    653, 310, 252, 333, 172, 101, 186, 143, 247, 370, 409, 448, 227, 224, 428, 
    614, 461, 355, 402, 249, 97, 45, 68, 124, 482, 595, 446, 133, 156, 435, 
    609, 571, 437, 367, 286, 149, 62, 98, 194, 346, 460, 373, 88, 175, 443, 
    572, 543, 455, 278, 246, 174, 123, 140, 170, 232, 319, 305, 104, 165, 469, 
    
    -- channel=593
    372, 359, 366, 309, 291, 284, 321, 361, 381, 391, 383, 368, 380, 354, 343, 
    401, 398, 411, 304, 197, 183, 171, 200, 254, 288, 334, 346, 371, 372, 347, 
    396, 395, 390, 284, 85, 132, 139, 149, 115, 118, 216, 361, 368, 338, 280, 
    394, 399, 334, 304, 143, 258, 267, 183, 192, 199, 214, 272, 351, 369, 278, 
    387, 402, 313, 202, 119, 146, 180, 150, 175, 178, 232, 238, 363, 394, 341, 
    335, 396, 295, 194, 25, 101, 117, 108, 100, 107, 143, 156, 282, 398, 394, 
    283, 297, 204, 189, 132, 122, 151, 99, 119, 170, 137, 126, 197, 276, 372, 
    297, 198, 149, 272, 86, 44, 25, 60, 29, 11, 39, 35, 28, 92, 238, 
    316, 227, 161, 123, 82, 157, 168, 144, 150, 169, 238, 160, 151, 199, 184, 
    322, 228, 109, 94, 31, 62, 15, 71, 158, 102, 126, 108, 158, 103, 79, 
    306, 255, 89, 77, 16, 8, 61, 98, 7, 93, 65, 74, 90, 128, 93, 
    281, 203, 58, 141, 93, 4, 0, 70, 27, 166, 171, 191, 123, 27, 28, 
    229, 249, 124, 168, 111, 49, 1, 0, 0, 169, 320, 302, 59, 14, 42, 
    234, 238, 195, 163, 100, 84, 9, 15, 56, 61, 126, 220, 34, 7, 53, 
    213, 201, 202, 103, 78, 68, 34, 32, 30, 45, 66, 138, 41, 7, 64, 
    
    -- channel=594
    62, 63, 45, 57, 53, 61, 88, 104, 91, 73, 75, 60, 69, 107, 95, 
    44, 46, 44, 32, 24, 13, 14, 14, 20, 60, 73, 54, 53, 88, 91, 
    35, 35, 28, 15, 28, 32, 27, 30, 25, 39, 63, 58, 52, 71, 102, 
    35, 32, 24, 4, 58, 42, 31, 17, 23, 44, 68, 36, 41, 77, 92, 
    32, 33, 18, 0, 41, 25, 0, 26, 28, 24, 23, 55, 44, 37, 57, 
    20, 24, 13, 36, 53, 17, 24, 30, 25, 27, 38, 43, 39, 35, 34, 
    14, 3, 10, 22, 51, 30, 17, 36, 40, 49, 54, 58, 34, 16, 27, 
    7, 11, 20, 30, 19, 27, 41, 54, 67, 61, 66, 74, 38, 7, 29, 
    15, 38, 51, 25, 56, 72, 57, 63, 89, 101, 90, 105, 89, 62, 57, 
    11, 35, 49, 53, 71, 42, 50, 37, 9, 8, 4, 8, 13, 20, 49, 
    11, 29, 77, 61, 83, 78, 61, 75, 42, 45, 42, 42, 61, 44, 71, 
    0, 22, 62, 65, 87, 97, 78, 47, 102, 45, 60, 66, 28, 68, 45, 
    3, 17, 80, 45, 56, 102, 109, 104, 96, 101, 82, 62, 90, 83, 68, 
    18, 12, 27, 50, 60, 80, 112, 108, 96, 64, 6, 21, 82, 91, 55, 
    10, 15, 28, 58, 69, 80, 97, 91, 84, 69, 50, 41, 96, 88, 57, 
    
    -- channel=595
    109, 94, 133, 138, 110, 115, 103, 79, 83, 101, 96, 89, 119, 64, 91, 
    130, 125, 163, 230, 174, 162, 146, 157, 134, 72, 73, 76, 101, 95, 30, 
    134, 133, 181, 301, 179, 214, 215, 235, 220, 145, 5, 100, 125, 108, 0, 
    133, 153, 148, 349, 126, 194, 288, 248, 241, 219, 147, 45, 121, 125, 64, 
    128, 162, 218, 298, 176, 194, 262, 237, 224, 215, 238, 69, 101, 163, 98, 
    106, 187, 198, 315, 147, 211, 238, 227, 223, 196, 194, 114, 48, 135, 133, 
    122, 205, 153, 226, 201, 228, 273, 227, 200, 224, 187, 104, 95, 99, 113, 
    166, 205, 52, 240, 224, 208, 187, 197, 167, 161, 163, 138, 120, 133, 39, 
    171, 216, 74, 229, 130, 148, 177, 208, 121, 104, 207, 133, 112, 188, 39, 
    181, 256, 110, 161, 132, 171, 130, 78, 226, 164, 200, 179, 181, 207, 0, 
    163, 282, 129, 160, 125, 105, 120, 202, 91, 192, 168, 118, 197, 143, 28, 
    199, 291, 89, 160, 187, 92, 74, 186, 16, 155, 161, 141, 208, 133, 0, 
    202, 262, 133, 199, 191, 146, 95, 90, 69, 6, 180, 278, 162, 87, 9, 
    180, 234, 232, 201, 166, 182, 91, 83, 82, 101, 134, 290, 132, 64, 45, 
    221, 213, 237, 198, 151, 152, 109, 110, 109, 121, 128, 226, 140, 77, 23, 
    
    -- channel=596
    0, 0, 0, 0, 0, 0, 0, 22, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 23, 48, 48, 25, 26, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 92, 80, 73, 52, 68, 86, 69, 0, 0, 0, 20, 
    0, 0, 0, 0, 171, 65, 21, 67, 61, 74, 69, 35, 0, 0, 0, 
    0, 0, 0, 0, 136, 105, 16, 89, 86, 87, 20, 93, 1, 0, 0, 
    0, 0, 0, 0, 120, 75, 70, 79, 68, 91, 70, 73, 69, 0, 0, 
    8, 0, 0, 0, 110, 97, 40, 66, 102, 71, 34, 106, 83, 25, 0, 
    0, 0, 43, 0, 49, 20, 58, 40, 56, 51, 50, 75, 109, 103, 103, 
    0, 0, 87, 0, 88, 65, 33, 0, 49, 85, 0, 32, 129, 59, 151, 
    0, 0, 39, 0, 97, 18, 87, 123, 1, 65, 16, 34, 39, 0, 206, 
    0, 0, 42, 0, 42, 71, 84, 14, 93, 12, 35, 72, 0, 64, 181, 
    0, 0, 55, 37, 0, 73, 118, 0, 192, 0, 32, 78, 0, 72, 202, 
    12, 0, 89, 16, 0, 0, 44, 60, 85, 168, 8, 0, 0, 74, 239, 
    43, 0, 0, 0, 30, 0, 43, 67, 91, 129, 46, 0, 0, 131, 196, 
    21, 16, 0, 0, 37, 0, 39, 51, 64, 74, 87, 0, 0, 105, 225, 
    
    -- channel=597
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 22, 9, 14, 23, 0, 0, 0, 
    0, 0, 0, 25, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 19, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 23, 21, 0, 17, 0, 0, 0, 0, 12, 0, 0, 
    0, 8, 0, 0, 17, 31, 34, 30, 18, 0, 0, 0, 15, 18, 0, 
    0, 0, 0, 0, 0, 26, 35, 27, 12, 0, 0, 0, 32, 12, 0, 
    0, 0, 0, 0, 0, 15, 26, 23, 15, 0, 0, 0, 28, 14, 0, 
    
    -- channel=598
    5, 6, 6, 9, 4, 2, 8, 3, 12, 19, 16, 14, 4, 7, 1, 
    16, 15, 16, 18, 21, 21, 21, 33, 38, 40, 15, 10, 17, 20, 10, 
    18, 17, 20, 0, 0, 0, 0, 0, 0, 0, 24, 10, 13, 14, 12, 
    18, 19, 11, 12, 4, 31, 17, 20, 18, 11, 15, 18, 8, 1, 8, 
    18, 16, 28, 11, 14, 17, 21, 19, 19, 19, 18, 18, 18, 7, 0, 
    17, 22, 5, 3, 7, 6, 10, 19, 20, 14, 30, 25, 13, 18, 18, 
    8, 21, 9, 0, 0, 12, 22, 8, 12, 29, 13, 13, 25, 33, 21, 
    19, 9, 0, 10, 9, 0, 0, 4, 18, 14, 6, 22, 10, 12, 24, 
    0, 1, 0, 11, 0, 11, 11, 0, 0, 0, 0, 0, 0, 11, 27, 
    9, 2, 15, 0, 4, 0, 1, 8, 15, 7, 17, 11, 22, 6, 6, 
    8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    15, 15, 3, 0, 0, 0, 8, 8, 0, 16, 6, 16, 10, 8, 0, 
    15, 0, 0, 4, 0, 0, 0, 0, 0, 0, 11, 12, 0, 0, 0, 
    8, 19, 5, 13, 0, 0, 0, 0, 0, 11, 10, 11, 0, 0, 0, 
    15, 11, 3, 7, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 
    
    -- channel=599
    59, 61, 62, 71, 74, 57, 58, 63, 66, 69, 80, 73, 69, 82, 82, 
    46, 46, 58, 48, 17, 1, 0, 14, 38, 64, 85, 77, 78, 101, 101, 
    42, 43, 45, 24, 0, 0, 0, 0, 0, 0, 34, 66, 85, 114, 103, 
    42, 48, 32, 2, 0, 0, 0, 0, 0, 0, 0, 64, 67, 97, 110, 
    46, 48, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 53, 53, 
    55, 62, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 42, 42, 
    56, 63, 56, 4, 0, 0, 0, 0, 0, 0, 0, 0, 22, 39, 49, 
    91, 69, 58, 58, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 5, 
    62, 52, 71, 24, 0, 10, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    51, 48, 55, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 39, 31, 29, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 35, 29, 9, 20, 37, 27, 37, 30, 37, 11, 32, 41, 9, 0, 
    0, 0, 0, 10, 7, 35, 47, 38, 16, 24, 26, 42, 31, 17, 0, 
    0, 0, 0, 13, 1, 30, 44, 37, 37, 5, 0, 24, 42, 16, 0, 
    0, 0, 0, 0, 8, 23, 31, 26, 17, 7, 0, 11, 33, 17, 0, 
    
    -- channel=600
    281, 280, 285, 271, 209, 188, 195, 213, 266, 298, 305, 285, 278, 271, 262, 
    304, 304, 318, 272, 195, 183, 200, 233, 246, 264, 286, 277, 300, 322, 260, 
    316, 315, 311, 261, 67, 101, 100, 120, 125, 164, 182, 273, 310, 303, 251, 
    315, 324, 284, 259, 68, 146, 207, 156, 139, 119, 216, 239, 275, 273, 248, 
    309, 321, 297, 189, 90, 152, 164, 128, 146, 151, 180, 178, 265, 293, 224, 
    273, 324, 211, 182, 71, 102, 122, 114, 121, 125, 149, 174, 230, 316, 314, 
    246, 282, 208, 133, 61, 99, 105, 81, 67, 107, 126, 133, 220, 253, 291, 
    243, 236, 94, 208, 104, 107, 91, 101, 74, 64, 79, 73, 72, 132, 197, 
    227, 175, 131, 183, 51, 94, 79, 75, 33, 32, 87, 43, 54, 127, 150, 
    254, 227, 110, 97, 56, 94, 91, 77, 185, 160, 182, 163, 166, 152, 77, 
    245, 208, 87, 73, 57, 27, 24, 134, 46, 133, 102, 76, 143, 65, 83, 
    234, 236, 38, 74, 90, 44, 78, 94, 28, 117, 110, 163, 143, 99, 37, 
    190, 151, 83, 139, 92, 60, 16, 13, 10, 19, 164, 197, 81, 9, 28, 
    184, 205, 168, 137, 86, 82, 14, 11, 24, 120, 159, 219, 54, 7, 42, 
    187, 168, 168, 123, 79, 66, 36, 35, 41, 61, 91, 123, 58, 17, 35, 
    
    -- channel=601
    220, 216, 233, 160, 209, 239, 233, 244, 231, 209, 188, 215, 200, 171, 137, 
    256, 254, 234, 137, 172, 202, 178, 164, 192, 163, 145, 223, 214, 128, 175, 
    254, 255, 233, 116, 228, 245, 252, 228, 209, 172, 212, 245, 202, 117, 132, 
    254, 244, 225, 149, 294, 307, 233, 233, 251, 269, 185, 226, 219, 185, 134, 
    258, 241, 179, 149, 252, 221, 209, 235, 240, 236, 239, 278, 273, 237, 265, 
    277, 232, 225, 139, 163, 214, 205, 193, 183, 198, 192, 193, 277, 254, 257, 
    274, 204, 204, 188, 253, 233, 231, 201, 238, 229, 152, 178, 198, 229, 263, 
    274, 133, 266, 212, 177, 141, 142, 120, 100, 101, 98, 97, 159, 218, 305, 
    276, 164, 239, 71, 204, 207, 219, 201, 248, 266, 239, 223, 266, 249, 292, 
    252, 99, 173, 91, 146, 117, 119, 205, 170, 179, 157, 162, 205, 121, 276, 
    266, 124, 139, 119, 81, 124, 209, 103, 172, 145, 149, 213, 122, 227, 258, 
    266, 60, 173, 203, 85, 70, 86, 53, 174, 169, 206, 199, 60, 101, 242, 
    266, 215, 210, 194, 127, 63, 60, 74, 102, 310, 266, 177, 61, 129, 266, 
    272, 232, 181, 176, 153, 75, 71, 96, 147, 153, 189, 118, 57, 145, 253, 
    238, 235, 196, 118, 132, 99, 92, 106, 117, 142, 171, 145, 64, 128, 277, 
    
    -- channel=602
    0, 0, 0, 0, 6, 7, 3, 12, 21, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 26, 62, 51, 45, 66, 45, 0, 34, 0, 0, 30, 
    0, 0, 0, 0, 69, 27, 19, 0, 20, 54, 124, 31, 0, 0, 72, 
    0, 0, 0, 0, 151, 50, 0, 13, 4, 23, 22, 102, 0, 0, 0, 
    6, 0, 0, 0, 113, 51, 0, 33, 37, 28, 0, 123, 37, 0, 0, 
    57, 0, 0, 0, 99, 40, 4, 22, 23, 43, 42, 77, 126, 0, 1, 
    52, 0, 2, 0, 34, 26, 0, 3, 47, 26, 0, 94, 119, 79, 32, 
    6, 0, 102, 0, 0, 0, 20, 0, 25, 31, 5, 43, 115, 94, 186, 
    0, 0, 108, 0, 66, 36, 0, 0, 3, 23, 0, 0, 67, 18, 196, 
    0, 0, 87, 0, 82, 0, 65, 115, 0, 58, 10, 34, 56, 0, 228, 
    0, 0, 13, 0, 0, 63, 61, 0, 116, 0, 10, 71, 0, 42, 169, 
    0, 0, 95, 0, 0, 29, 101, 0, 182, 0, 21, 64, 0, 77, 213, 
    16, 0, 28, 11, 0, 0, 12, 30, 57, 192, 0, 0, 0, 62, 218, 
    33, 0, 0, 0, 1, 0, 9, 32, 62, 137, 71, 0, 0, 107, 183, 
    3, 0, 0, 0, 12, 0, 4, 18, 34, 50, 75, 0, 0, 85, 212, 
    
    -- channel=603
    431, 423, 427, 336, 352, 365, 390, 422, 445, 446, 425, 435, 425, 394, 367, 
    471, 469, 454, 279, 225, 224, 208, 233, 296, 345, 371, 423, 437, 390, 407, 
    466, 465, 442, 234, 149, 186, 186, 177, 147, 146, 321, 446, 417, 350, 343, 
    465, 457, 395, 256, 226, 343, 269, 201, 226, 237, 242, 370, 425, 401, 321, 
    464, 455, 317, 180, 186, 172, 196, 179, 202, 210, 253, 347, 461, 459, 428, 
    439, 438, 340, 153, 77, 142, 131, 124, 122, 137, 167, 220, 395, 467, 467, 
    393, 350, 277, 216, 172, 157, 164, 121, 150, 196, 150, 172, 269, 356, 463, 
    402, 217, 287, 299, 117, 80, 49, 51, 35, 32, 28, 41, 90, 162, 387, 
    399, 243, 268, 119, 142, 191, 225, 202, 221, 250, 290, 223, 236, 239, 335, 
    398, 180, 187, 82, 79, 76, 50, 129, 200, 141, 150, 145, 202, 111, 226, 
    390, 224, 124, 96, 28, 54, 144, 74, 112, 114, 99, 171, 88, 183, 222, 
    352, 140, 139, 187, 77, 15, 23, 52, 92, 212, 226, 219, 98, 65, 156, 
    303, 263, 176, 210, 116, 33, 9, 16, 33, 296, 378, 286, 44, 64, 175, 
    302, 286, 205, 194, 123, 69, 24, 39, 97, 133, 187, 191, 26, 65, 173, 
    260, 247, 220, 113, 101, 75, 53, 58, 64, 88, 123, 156, 35, 62, 191, 
    
    -- channel=604
    385, 368, 380, 311, 304, 322, 357, 378, 386, 392, 368, 367, 396, 339, 346, 
    419, 416, 419, 326, 263, 261, 232, 253, 285, 304, 318, 342, 364, 344, 317, 
    413, 411, 418, 346, 258, 311, 322, 333, 287, 239, 257, 371, 354, 312, 242, 
    412, 414, 366, 391, 266, 389, 394, 357, 368, 370, 316, 278, 372, 356, 253, 
    404, 418, 338, 322, 272, 280, 333, 325, 333, 333, 387, 308, 388, 434, 371, 
    349, 404, 354, 314, 162, 266, 276, 263, 260, 258, 270, 266, 320, 416, 413, 
    304, 323, 235, 290, 283, 279, 326, 262, 265, 308, 248, 201, 241, 298, 400, 
    305, 219, 198, 309, 229, 209, 165, 171, 127, 127, 131, 114, 142, 206, 304, 
    341, 278, 189, 185, 202, 222, 289, 303, 269, 281, 373, 285, 257, 293, 264, 
    363, 266, 166, 163, 127, 174, 118, 141, 278, 204, 236, 219, 249, 214, 167, 
    345, 323, 166, 168, 99, 110, 205, 179, 141, 205, 192, 218, 176, 244, 183, 
    354, 269, 145, 248, 187, 70, 48, 165, 62, 247, 268, 222, 204, 113, 111, 
    338, 390, 215, 263, 227, 128, 76, 78, 79, 242, 389, 379, 136, 113, 140, 
    326, 342, 300, 254, 203, 182, 87, 93, 126, 140, 214, 316, 113, 89, 168, 
    331, 328, 319, 204, 176, 165, 120, 122, 122, 138, 156, 251, 123, 98, 177, 
    
    -- channel=605
    771, 764, 754, 573, 608, 638, 693, 766, 830, 808, 765, 786, 722, 708, 629, 
    868, 865, 811, 493, 519, 557, 537, 575, 664, 696, 688, 780, 782, 662, 730, 
    874, 874, 789, 375, 489, 557, 554, 528, 504, 503, 694, 809, 722, 571, 655, 
    871, 850, 740, 443, 657, 767, 659, 646, 653, 665, 627, 747, 726, 633, 552, 
    867, 832, 627, 396, 598, 594, 566, 609, 639, 650, 659, 765, 850, 764, 710, 
    824, 780, 588, 350, 402, 495, 483, 486, 482, 524, 568, 622, 848, 875, 876, 
    724, 590, 505, 395, 490, 517, 502, 423, 488, 541, 404, 495, 657, 750, 879, 
    644, 334, 514, 485, 402, 318, 293, 257, 235, 233, 213, 247, 385, 517, 865, 
    631, 337, 515, 217, 403, 444, 481, 387, 412, 484, 474, 398, 531, 552, 795, 
    672, 270, 389, 144, 310, 248, 282, 430, 484, 467, 450, 446, 527, 321, 658, 
    699, 301, 275, 209, 133, 225, 380, 232, 378, 338, 330, 457, 285, 441, 615, 
    691, 204, 325, 384, 149, 124, 235, 112, 351, 413, 476, 517, 163, 283, 523, 
    664, 428, 404, 459, 239, 88, 68, 102, 164, 646, 680, 460, 115, 207, 565, 
    668, 612, 434, 415, 319, 128, 86, 135, 253, 443, 507, 352, 64, 251, 559, 
    621, 585, 475, 283, 283, 177, 147, 172, 208, 277, 375, 319, 88, 231, 605, 
    
    -- channel=606
    0, 0, 21, 101, 0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 37, 
    0, 0, 74, 273, 18, 0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 
    0, 0, 108, 455, 0, 0, 0, 33, 0, 0, 0, 0, 42, 108, 0, 
    0, 20, 16, 506, 0, 0, 137, 0, 0, 0, 0, 0, 20, 105, 0, 
    0, 49, 169, 323, 0, 0, 86, 0, 0, 0, 41, 0, 0, 118, 0, 
    0, 116, 130, 365, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 186, 24, 180, 0, 0, 86, 18, 0, 1, 32, 0, 0, 0, 0, 
    54, 243, 0, 228, 42, 63, 0, 69, 5, 0, 19, 0, 0, 0, 0, 
    78, 273, 0, 295, 0, 0, 0, 127, 0, 0, 154, 0, 0, 0, 0, 
    96, 392, 0, 147, 0, 59, 0, 0, 100, 0, 42, 0, 0, 124, 0, 
    12, 459, 0, 86, 17, 0, 0, 159, 0, 76, 2, 0, 118, 0, 0, 
    35, 499, 0, 0, 203, 0, 0, 217, 0, 22, 0, 0, 270, 0, 0, 
    0, 293, 0, 65, 159, 127, 0, 0, 0, 0, 31, 360, 146, 0, 0, 
    0, 98, 170, 105, 23, 207, 0, 0, 0, 0, 0, 397, 107, 0, 0, 
    25, 28, 160, 139, 10, 94, 0, 0, 0, 0, 0, 203, 111, 0, 0, 
    
    -- channel=607
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 3, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 30, 25, 11, 0, 0, 0, 2, 2, 0, 
    0, 0, 0, 0, 0, 0, 24, 18, 3, 0, 0, 0, 7, 3, 0, 
    0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 8, 3, 0, 
    
    -- channel=608
    14, 14, 24, 54, 31, 25, 0, 0, 0, 10, 20, 22, 18, 7, 19, 
    14, 12, 26, 66, 14, 1, 21, 29, 15, 5, 30, 18, 30, 37, 15, 
    18, 18, 35, 67, 0, 0, 0, 0, 0, 0, 0, 18, 44, 51, 21, 
    19, 21, 39, 61, 0, 0, 0, 0, 0, 0, 0, 16, 40, 38, 43, 
    21, 26, 50, 39, 0, 0, 0, 0, 0, 0, 0, 0, 8, 28, 19, 
    34, 41, 43, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 18, 
    52, 84, 77, 44, 0, 0, 0, 0, 0, 0, 0, 0, 7, 28, 11, 
    77, 113, 43, 52, 0, 2, 2, 3, 10, 11, 9, 6, 0, 0, 0, 
    66, 77, 25, 116, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    53, 79, 32, 47, 4, 15, 8, 0, 25, 11, 19, 15, 1, 38, 0, 
    47, 78, 20, 23, 24, 11, 0, 19, 1, 19, 2, 0, 43, 0, 0, 
    28, 83, 13, 0, 24, 12, 19, 46, 0, 24, 0, 1, 64, 22, 0, 
    11, 8, 0, 6, 11, 20, 14, 10, 10, 0, 0, 9, 37, 4, 0, 
    0, 20, 17, 11, 3, 23, 11, 4, 0, 7, 20, 37, 34, 0, 0, 
    1, 0, 4, 35, 3, 16, 10, 6, 6, 7, 9, 28, 29, 0, 0, 
    
    -- channel=609
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=610
    0, 0, 2, 0, 2, 1, 8, 18, 23, 1, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 13, 21, 0, 0, 24, 17, 0, 18, 2, 0, 10, 
    0, 0, 0, 0, 20, 10, 0, 0, 1, 9, 35, 20, 0, 0, 14, 
    0, 2, 0, 0, 55, 14, 0, 0, 0, 0, 5, 37, 0, 0, 0, 
    0, 0, 0, 0, 51, 0, 0, 2, 3, 0, 5, 35, 15, 0, 0, 
    13, 0, 0, 0, 12, 3, 0, 0, 0, 3, 0, 2, 39, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 4, 18, 0, 20, 38, 5, 18, 
    10, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 72, 
    0, 0, 48, 0, 18, 0, 0, 0, 6, 0, 3, 5, 22, 0, 45, 
    0, 0, 43, 0, 22, 0, 5, 0, 0, 0, 0, 0, 27, 0, 32, 
    0, 0, 4, 0, 0, 0, 6, 0, 26, 0, 0, 24, 0, 17, 4, 
    0, 0, 29, 11, 0, 0, 9, 0, 37, 0, 17, 31, 0, 29, 3, 
    0, 0, 1, 34, 0, 0, 0, 1, 0, 84, 9, 0, 0, 4, 34, 
    5, 0, 0, 26, 0, 0, 0, 0, 13, 47, 1, 0, 0, 20, 20, 
    0, 0, 0, 0, 2, 0, 0, 1, 1, 6, 12, 0, 0, 19, 41, 
    
    -- channel=611
    144, 141, 151, 107, 136, 144, 135, 149, 145, 139, 137, 149, 139, 154, 121, 
    134, 135, 136, 12, 28, 21, 5, 12, 53, 89, 119, 164, 150, 137, 168, 
    126, 128, 110, 0, 0, 0, 0, 0, 0, 0, 117, 167, 154, 135, 159, 
    127, 125, 94, 0, 28, 10, 0, 0, 0, 0, 1, 152, 147, 170, 138, 
    133, 128, 17, 0, 0, 0, 0, 0, 0, 0, 0, 106, 146, 143, 179, 
    152, 123, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 140, 126, 130, 
    159, 102, 102, 31, 0, 0, 0, 0, 0, 0, 0, 12, 63, 80, 137, 
    172, 60, 159, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 146, 
    160, 49, 164, 0, 27, 35, 10, 15, 115, 99, 83, 106, 97, 19, 92, 
    129, 3, 104, 0, 13, 0, 0, 12, 0, 0, 0, 0, 21, 0, 66, 
    128, 6, 76, 29, 10, 13, 30, 0, 33, 5, 9, 56, 0, 50, 40, 
    73, 0, 75, 78, 5, 17, 8, 0, 69, 37, 56, 69, 0, 22, 38, 
    35, 31, 61, 66, 5, 24, 33, 32, 32, 158, 92, 62, 0, 37, 50, 
    51, 25, 6, 52, 14, 11, 46, 48, 51, 42, 23, 27, 8, 48, 21, 
    0, 0, 17, 0, 19, 17, 39, 41, 33, 31, 26, 32, 11, 44, 55, 
    
    -- channel=612
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 12, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 28, 14, 17, 20, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 35, 42, 33, 21, 0, 0, 0, 26, 14, 0, 
    0, 0, 0, 0, 0, 19, 38, 33, 17, 0, 0, 0, 35, 13, 0, 
    0, 0, 0, 0, 0, 13, 24, 19, 11, 0, 0, 0, 30, 9, 0, 
    
    -- channel=613
    198, 176, 208, 150, 157, 162, 168, 166, 197, 218, 193, 205, 186, 144, 136, 
    248, 244, 257, 177, 186, 201, 186, 223, 245, 211, 174, 196, 210, 167, 149, 
    257, 257, 260, 146, 158, 181, 174, 172, 171, 150, 154, 211, 198, 148, 113, 
    255, 259, 218, 224, 205, 274, 252, 267, 253, 244, 180, 197, 205, 162, 91, 
    253, 263, 215, 210, 203, 210, 254, 243, 251, 239, 265, 201, 226, 224, 143, 
    236, 267, 183, 165, 123, 182, 193, 198, 197, 191, 219, 180, 221, 258, 256, 
    199, 214, 143, 149, 132, 192, 232, 166, 180, 226, 143, 132, 203, 242, 266, 
    196, 112, 104, 152, 158, 109, 90, 99, 88, 81, 76, 81, 112, 151, 243, 
    180, 100, 92, 103, 115, 129, 151, 109, 40, 48, 109, 31, 67, 170, 197, 
    208, 100, 111, 10, 74, 74, 59, 103, 191, 156, 181, 162, 201, 125, 111, 
    213, 131, 40, 43, 0, 31, 62, 50, 82, 90, 90, 91, 76, 121, 93, 
    238, 114, 70, 89, 22, 0, 33, 69, 28, 142, 138, 159, 70, 81, 53, 
    233, 159, 46, 166, 73, 0, 0, 0, 0, 118, 190, 189, 9, 5, 55, 
    215, 236, 167, 156, 95, 32, 0, 0, 9, 104, 170, 204, 0, 0, 91, 
    231, 211, 186, 99, 75, 37, 0, 0, 9, 46, 93, 159, 0, 0, 88, 
    
    -- channel=614
    486, 474, 485, 396, 383, 391, 398, 422, 493, 516, 496, 510, 454, 453, 396, 
    542, 541, 531, 317, 314, 324, 333, 386, 438, 469, 462, 513, 521, 470, 470, 
    554, 556, 514, 220, 197, 226, 202, 194, 214, 268, 422, 519, 499, 424, 455, 
    553, 545, 476, 258, 289, 373, 298, 279, 273, 274, 335, 500, 488, 433, 378, 
    554, 540, 395, 210, 259, 269, 266, 253, 284, 281, 313, 443, 521, 487, 425, 
    541, 524, 334, 162, 179, 199, 202, 199, 208, 231, 280, 335, 520, 555, 556, 
    488, 434, 356, 211, 146, 208, 190, 154, 180, 231, 188, 259, 427, 496, 559, 
    455, 281, 324, 288, 168, 142, 130, 118, 106, 99, 98, 116, 183, 270, 535, 
    417, 206, 324, 188, 171, 216, 202, 149, 143, 166, 176, 131, 202, 255, 458, 
    441, 181, 263, 52, 146, 113, 138, 211, 285, 266, 268, 259, 304, 183, 334, 
    452, 185, 152, 91, 49, 89, 129, 104, 189, 171, 159, 210, 159, 185, 297, 
    421, 152, 170, 170, 53, 33, 137, 69, 170, 230, 236, 306, 90, 180, 236, 
    371, 193, 163, 261, 97, 23, 5, 18, 52, 290, 337, 249, 46, 68, 229, 
    364, 354, 231, 237, 145, 52, 10, 32, 84, 263, 308, 253, 11, 84, 235, 
    334, 299, 254, 158, 130, 75, 43, 57, 78, 125, 194, 200, 20, 79, 250, 
    
    -- channel=615
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 22, 18, 35, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=616
    42, 44, 38, 22, 21, 33, 39, 60, 53, 36, 38, 32, 43, 43, 34, 
    41, 42, 37, 9, 0, 0, 0, 0, 0, 0, 14, 31, 30, 24, 30, 
    36, 36, 25, 16, 0, 0, 0, 0, 0, 0, 0, 39, 35, 18, 11, 
    35, 33, 21, 0, 0, 9, 14, 0, 0, 0, 7, 0, 27, 43, 27, 
    34, 33, 6, 0, 0, 0, 0, 0, 0, 0, 0, 9, 41, 41, 63, 
    23, 25, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 36, 36, 
    24, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    21, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 14, 17, 0, 0, 0, 0, 0, 40, 54, 45, 44, 42, 8, 1, 
    26, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 23, 0, 0, 0, 0, 0, 0, 21, 48, 19, 0, 0, 1, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=617
    632, 628, 615, 452, 483, 502, 558, 647, 680, 652, 623, 629, 610, 594, 527, 
    690, 690, 653, 343, 315, 327, 300, 322, 422, 497, 531, 624, 626, 551, 600, 
    683, 683, 611, 285, 244, 314, 312, 301, 256, 271, 498, 644, 588, 477, 512, 
    681, 667, 555, 290, 388, 490, 404, 338, 366, 381, 401, 550, 585, 556, 444, 
    677, 657, 423, 202, 314, 298, 285, 298, 336, 347, 401, 536, 674, 639, 625, 
    627, 608, 445, 175, 121, 226, 215, 197, 188, 238, 260, 344, 620, 684, 685, 
    543, 424, 337, 253, 273, 247, 234, 180, 237, 283, 204, 272, 404, 502, 681, 
    497, 208, 364, 377, 148, 101, 73, 63, 11, 4, 22, 28, 119, 256, 603, 
    516, 250, 376, 49, 205, 256, 290, 235, 342, 388, 396, 335, 391, 343, 503, 
    527, 182, 215, 62, 95, 84, 71, 200, 256, 220, 205, 203, 287, 121, 379, 
    529, 215, 161, 94, 7, 44, 206, 91, 143, 154, 142, 262, 92, 275, 350, 
    488, 104, 152, 268, 61, 1, 25, 0, 153, 248, 304, 322, 51, 65, 269, 
    422, 341, 272, 284, 124, 9, 0, 0, 27, 480, 532, 363, 1, 67, 315, 
    448, 384, 265, 244, 154, 40, 1, 34, 126, 197, 265, 216, 0, 97, 293, 
    372, 355, 300, 110, 122, 60, 47, 61, 73, 111, 164, 152, 1, 80, 356, 
    
    -- channel=618
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=619
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 130, 201, 223, 282, 362, 332, 203, 70, 0, 1, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 38, 0, 1, 49, 76, 
    0, 0, 9, 25, 0, 0, 0, 51, 0, 0, 0, 126, 0, 0, 22, 
    0, 0, 182, 124, 44, 125, 132, 55, 61, 55, 0, 0, 0, 0, 0, 
    65, 58, 0, 0, 175, 49, 51, 135, 150, 103, 189, 125, 20, 0, 0, 
    60, 148, 150, 0, 0, 37, 51, 25, 32, 87, 87, 154, 281, 267, 18, 
    88, 208, 26, 0, 121, 28, 48, 113, 256, 231, 184, 288, 259, 163, 86, 
    0, 0, 29, 277, 3, 63, 0, 0, 0, 0, 0, 0, 0, 0, 117, 
    0, 41, 192, 0, 153, 82, 169, 193, 166, 197, 228, 204, 199, 152, 83, 
    6, 0, 0, 0, 50, 88, 0, 11, 100, 0, 3, 0, 72, 0, 26, 
    49, 111, 90, 0, 0, 73, 317, 171, 174, 111, 0, 163, 149, 248, 104, 
    43, 0, 0, 28, 0, 0, 27, 24, 8, 0, 0, 0, 54, 0, 0, 
    0, 67, 0, 61, 24, 0, 0, 0, 0, 233, 223, 88, 24, 14, 28, 
    64, 6, 0, 84, 45, 0, 0, 0, 0, 45, 137, 87, 0, 9, 0, 
    
    -- channel=620
    41, 39, 49, 89, 35, 37, 26, 15, 5, 22, 33, 18, 63, 25, 55, 
    36, 34, 53, 140, 1, 0, 5, 0, 0, 0, 9, 0, 26, 48, 0, 
    34, 32, 67, 201, 0, 19, 39, 56, 31, 0, 0, 14, 55, 56, 0, 
    35, 39, 68, 175, 0, 3, 83, 4, 15, 22, 20, 0, 52, 74, 42, 
    30, 48, 99, 120, 0, 9, 32, 1, 1, 13, 26, 0, 11, 79, 75, 
    4, 59, 117, 153, 0, 8, 31, 8, 6, 0, 0, 0, 0, 37, 33, 
    32, 96, 68, 114, 42, 26, 35, 36, 6, 0, 41, 0, 0, 0, 0, 
    72, 146, 0, 102, 40, 55, 38, 40, 6, 6, 20, 0, 0, 0, 0, 
    105, 178, 0, 129, 0, 27, 44, 97, 62, 63, 101, 75, 22, 50, 0, 
    87, 198, 0, 122, 0, 42, 0, 0, 38, 3, 24, 10, 0, 82, 0, 
    62, 208, 42, 58, 48, 0, 12, 100, 0, 68, 31, 0, 103, 5, 0, 
    56, 205, 0, 42, 112, 19, 0, 72, 0, 29, 18, 0, 141, 0, 0, 
    40, 156, 57, 10, 86, 75, 21, 12, 10, 0, 60, 105, 94, 2, 0, 
    31, 57, 92, 16, 35, 92, 29, 17, 1, 0, 0, 87, 79, 0, 0, 
    41, 46, 72, 71, 20, 57, 38, 26, 20, 11, 0, 47, 88, 0, 0, 
    
    -- channel=621
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=622
    0, 5, 0, 0, 0, 11, 23, 49, 47, 0, 0, 11, 0, 9, 0, 
    0, 2, 0, 0, 0, 14, 2, 0, 15, 23, 0, 35, 0, 0, 42, 
    0, 0, 0, 0, 53, 22, 9, 0, 0, 28, 105, 33, 0, 0, 69, 
    0, 0, 0, 0, 135, 42, 0, 0, 0, 19, 18, 80, 0, 0, 0, 
    5, 0, 0, 0, 87, 29, 0, 11, 15, 15, 0, 103, 42, 0, 3, 
    42, 0, 0, 0, 63, 14, 0, 0, 0, 22, 13, 59, 113, 0, 0, 
    31, 0, 0, 0, 29, 4, 0, 0, 26, 6, 0, 63, 73, 40, 32, 
    0, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 9, 77, 58, 158, 
    0, 0, 91, 0, 57, 17, 1, 0, 34, 59, 0, 16, 92, 6, 178, 
    0, 0, 41, 0, 56, 0, 26, 78, 0, 9, 0, 0, 5, 0, 215, 
    0, 0, 1, 0, 0, 36, 61, 0, 93, 0, 0, 67, 0, 40, 165, 
    0, 0, 61, 4, 0, 8, 58, 0, 150, 0, 13, 32, 0, 30, 199, 
    0, 0, 28, 0, 0, 0, 0, 14, 44, 204, 0, 0, 0, 47, 213, 
    12, 0, 0, 0, 0, 0, 0, 23, 52, 98, 25, 0, 0, 90, 173, 
    0, 0, 0, 0, 0, 0, 0, 6, 18, 27, 43, 0, 0, 69, 209, 
    
    -- channel=623
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=624
    205, 198, 194, 127, 165, 179, 187, 201, 212, 208, 186, 212, 184, 174, 156, 
    227, 228, 196, 75, 137, 168, 160, 164, 190, 203, 183, 215, 202, 148, 199, 
    231, 232, 194, 34, 196, 190, 189, 170, 168, 173, 238, 220, 168, 124, 187, 
    231, 214, 198, 55, 240, 239, 156, 209, 210, 225, 178, 235, 200, 142, 122, 
    233, 210, 121, 94, 207, 191, 172, 200, 208, 209, 207, 251, 235, 195, 198, 
    236, 180, 147, 54, 158, 176, 155, 157, 160, 182, 181, 211, 278, 231, 233, 
    202, 131, 129, 118, 149, 159, 155, 138, 164, 157, 117, 164, 206, 229, 253, 
    149, 52, 197, 67, 132, 124, 120, 84, 78, 90, 74, 80, 156, 184, 304, 
    156, 53, 153, 30, 164, 128, 151, 122, 143, 161, 118, 126, 165, 150, 281, 
    170, 10, 125, 31, 107, 81, 102, 168, 136, 158, 140, 148, 159, 97, 273, 
    188, 26, 85, 63, 41, 102, 156, 28, 178, 100, 124, 186, 67, 167, 224, 
    186, 0, 134, 125, 20, 37, 89, 42, 135, 127, 141, 130, 26, 95, 245, 
    200, 119, 107, 128, 72, 14, 31, 48, 84, 251, 164, 69, 16, 99, 224, 
    197, 167, 115, 108, 103, 27, 38, 59, 86, 143, 180, 67, 22, 104, 226, 
    184, 178, 129, 71, 93, 58, 53, 65, 78, 100, 128, 99, 17, 98, 254, 
    
    -- channel=625
    149, 144, 131, 92, 117, 129, 169, 194, 155, 139, 131, 134, 173, 165, 169, 
    121, 123, 110, 15, 0, 0, 0, 0, 0, 44, 106, 119, 122, 138, 166, 
    101, 99, 95, 33, 0, 0, 3, 1, 0, 0, 84, 136, 109, 120, 121, 
    102, 95, 70, 10, 0, 29, 0, 0, 0, 0, 0, 68, 132, 169, 115, 
    100, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 123, 164, 202, 
    81, 75, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 102, 102, 
    59, 34, 18, 59, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 
    78, 0, 91, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 
    111, 72, 62, 0, 14, 24, 47, 102, 190, 181, 204, 204, 125, 27, 19, 
    94, 17, 19, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    74, 64, 44, 37, 4, 9, 67, 0, 0, 0, 0, 57, 0, 56, 7, 
    18, 0, 52, 89, 48, 8, 0, 0, 0, 27, 59, 0, 0, 0, 0, 
    3, 125, 70, 25, 50, 50, 44, 39, 32, 164, 142, 102, 14, 46, 9, 
    15, 0, 11, 26, 15, 49, 69, 61, 58, 0, 0, 0, 39, 30, 0, 
    0, 0, 17, 0, 12, 43, 58, 51, 32, 6, 0, 20, 43, 33, 22, 
    
    -- channel=626
    0, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 22, 203, 33, 0, 35, 68, 18, 0, 9, 0, 0, 55, 0, 
    0, 0, 62, 241, 0, 0, 0, 0, 0, 0, 0, 0, 23, 74, 0, 
    0, 5, 38, 276, 0, 0, 78, 11, 0, 0, 0, 0, 10, 20, 2, 
    0, 19, 155, 212, 0, 0, 85, 0, 0, 0, 4, 0, 0, 16, 0, 
    0, 66, 83, 201, 0, 0, 27, 33, 42, 0, 29, 0, 0, 0, 0, 
    0, 143, 66, 111, 0, 0, 45, 21, 0, 3, 48, 0, 0, 0, 0, 
    39, 212, 0, 90, 65, 61, 35, 68, 78, 72, 61, 50, 0, 0, 0, 
    19, 168, 0, 275, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 
    44, 247, 0, 111, 0, 52, 4, 0, 79, 13, 79, 45, 13, 133, 0, 
    10, 265, 0, 42, 39, 0, 0, 97, 0, 56, 7, 0, 132, 0, 0, 
    24, 318, 0, 0, 101, 0, 0, 168, 0, 40, 0, 0, 217, 23, 0, 
    13, 81, 0, 1, 71, 59, 4, 0, 0, 0, 0, 108, 117, 0, 0, 
    0, 66, 91, 36, 16, 103, 0, 0, 0, 0, 2, 184, 85, 0, 0, 
    33, 19, 60, 111, 11, 55, 0, 0, 0, 0, 0, 107, 74, 0, 0, 
    
    -- channel=627
    39, 42, 24, 55, 48, 31, 36, 33, 33, 48, 60, 55, 55, 79, 91, 
    9, 12, 12, 12, 0, 0, 0, 3, 12, 71, 91, 51, 52, 100, 103, 
    5, 6, 4, 0, 0, 0, 0, 0, 0, 0, 64, 31, 48, 105, 134, 
    6, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 56, 49, 69, 99, 
    9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 31, 
    16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 5, 
    5, 14, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 14, 
    7, 40, 45, 0, 0, 0, 0, 0, 0, 2, 4, 14, 0, 0, 0, 
    0, 21, 21, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 41, 49, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 27, 28, 44, 32, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 14, 44, 0, 27, 58, 46, 61, 34, 27, 0, 0, 48, 23, 11, 
    0, 0, 0, 0, 9, 53, 77, 68, 58, 7, 0, 0, 46, 46, 0, 
    0, 0, 0, 0, 0, 42, 76, 63, 37, 4, 0, 0, 71, 36, 0, 
    0, 0, 0, 3, 11, 38, 56, 46, 34, 14, 0, 0, 57, 40, 0, 
    
    -- channel=628
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=629
    0, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 36, 
    0, 0, 9, 178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 
    0, 0, 60, 292, 0, 0, 0, 0, 0, 0, 0, 0, 1, 74, 0, 
    0, 0, 33, 307, 0, 0, 33, 0, 0, 0, 0, 0, 40, 42, 0, 
    0, 6, 88, 244, 0, 0, 60, 0, 0, 0, 5, 0, 0, 80, 0, 
    0, 40, 143, 200, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 131, 35, 185, 0, 0, 33, 0, 0, 0, 13, 0, 0, 0, 0, 
    23, 196, 0, 78, 41, 65, 1, 27, 1, 15, 4, 0, 0, 0, 0, 
    48, 223, 0, 242, 0, 0, 11, 106, 0, 0, 62, 0, 0, 0, 0, 
    71, 269, 0, 160, 0, 48, 0, 0, 40, 0, 27, 0, 0, 117, 0, 
    11, 347, 0, 68, 15, 0, 0, 48, 0, 41, 6, 0, 71, 0, 0, 
    8, 354, 0, 0, 125, 0, 0, 214, 0, 49, 0, 0, 269, 0, 0, 
    0, 238, 0, 0, 131, 69, 0, 0, 0, 0, 0, 150, 106, 0, 0, 
    0, 45, 113, 12, 11, 147, 0, 0, 0, 0, 0, 207, 118, 0, 0, 
    3, 15, 75, 86, 0, 78, 0, 0, 0, 0, 0, 130, 87, 0, 0, 
    
    -- channel=630
    146, 129, 152, 88, 107, 132, 154, 173, 161, 144, 115, 114, 144, 92, 96, 
    183, 178, 191, 168, 199, 215, 172, 169, 172, 108, 72, 104, 106, 68, 52, 
    181, 181, 189, 235, 305, 361, 369, 382, 337, 242, 95, 127, 103, 49, 0, 
    179, 189, 156, 301, 305, 336, 391, 424, 421, 404, 257, 82, 115, 104, 10, 
    169, 192, 186, 300, 331, 329, 370, 402, 387, 375, 392, 184, 160, 179, 131, 
    124, 185, 196, 305, 207, 321, 352, 340, 325, 322, 301, 208, 150, 181, 180, 
    99, 114, 70, 208, 331, 351, 401, 330, 336, 351, 235, 166, 133, 125, 179, 
    78, 44, 37, 184, 270, 225, 202, 211, 155, 148, 165, 137, 153, 204, 159, 
    129, 123, 62, 76, 206, 185, 247, 238, 210, 212, 283, 211, 226, 263, 136, 
    155, 148, 73, 102, 134, 171, 129, 135, 230, 201, 219, 202, 227, 186, 106, 
    153, 187, 109, 130, 83, 97, 191, 173, 117, 184, 188, 185, 141, 234, 113, 
    228, 173, 84, 210, 145, 58, 47, 118, 50, 160, 206, 171, 129, 99, 66, 
    259, 304, 180, 223, 188, 101, 53, 60, 55, 174, 259, 289, 94, 87, 130, 
    259, 267, 250, 208, 186, 140, 55, 68, 99, 107, 160, 255, 69, 84, 159, 
    291, 293, 279, 164, 161, 126, 86, 98, 102, 123, 140, 202, 81, 85, 177, 
    
    -- channel=631
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=632
    0, 3, 0, 15, 0, 0, 0, 0, 1, 0, 5, 0, 0, 4, 3, 
    0, 0, 0, 31, 0, 0, 15, 3, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 33, 0, 0, 0, 0, 0, 11, 0, 0, 5, 10, 0, 
    0, 0, 5, 0, 0, 0, 8, 0, 0, 0, 37, 0, 0, 0, 19, 
    0, 0, 21, 1, 0, 16, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 9, 16, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 19, 11, 0, 0, 0, 
    0, 27, 0, 0, 0, 0, 0, 4, 0, 0, 4, 3, 0, 6, 0, 
    0, 29, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 46, 0, 36, 0, 4, 2, 10, 0, 0, 0, 0, 0, 18, 0, 
    0, 24, 1, 0, 13, 0, 0, 31, 0, 0, 0, 0, 9, 0, 18, 
    0, 51, 0, 0, 22, 14, 8, 0, 0, 0, 0, 0, 49, 0, 13, 
    0, 1, 11, 0, 3, 11, 0, 0, 0, 0, 0, 0, 23, 0, 2, 
    0, 0, 7, 0, 0, 9, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    
    -- channel=633
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=634
    0, 0, 0, 0, 16, 18, 20, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 38, 31, 19, 12, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 88, 58, 61, 52, 52, 36, 33, 0, 0, 0, 10, 
    0, 0, 0, 0, 71, 39, 19, 43, 43, 51, 5, 6, 0, 0, 8, 
    0, 0, 0, 33, 74, 45, 44, 54, 43, 47, 29, 18, 0, 0, 0, 
    0, 0, 15, 23, 95, 73, 50, 66, 66, 59, 50, 45, 0, 0, 0, 
    0, 0, 17, 57, 81, 61, 66, 75, 80, 62, 61, 60, 21, 5, 0, 
    0, 10, 67, 10, 72, 68, 67, 60, 91, 104, 79, 95, 110, 59, 19, 
    0, 27, 46, 45, 89, 65, 83, 80, 75, 78, 57, 74, 68, 40, 50, 
    0, 4, 69, 76, 102, 78, 84, 81, 43, 45, 39, 50, 38, 53, 83, 
    0, 14, 69, 87, 90, 116, 107, 39, 111, 47, 66, 78, 39, 82, 78, 
    0, 3, 109, 70, 69, 103, 92, 90, 103, 74, 64, 28, 67, 80, 112, 
    23, 31, 58, 46, 72, 84, 118, 120, 120, 94, 27, 7, 82, 124, 107, 
    15, 15, 30, 48, 77, 76, 116, 115, 109, 76, 51, 4, 98, 121, 105, 
    26, 33, 26, 59, 82, 88, 104, 103, 101, 90, 76, 58, 91, 117, 103, 
    
    -- channel=635
    503, 500, 495, 363, 380, 401, 418, 475, 525, 518, 495, 515, 465, 453, 390, 
    569, 569, 525, 266, 276, 306, 307, 326, 392, 428, 434, 520, 514, 422, 475, 
    577, 578, 501, 186, 241, 287, 284, 261, 251, 279, 438, 531, 479, 360, 426, 
    576, 554, 488, 199, 361, 426, 335, 325, 333, 348, 361, 493, 482, 407, 343, 
    575, 542, 362, 176, 298, 316, 278, 298, 330, 342, 349, 484, 556, 494, 483, 
    556, 498, 359, 134, 174, 234, 225, 215, 214, 262, 283, 363, 569, 578, 580, 
    494, 372, 322, 207, 226, 245, 214, 176, 222, 240, 176, 260, 398, 478, 582, 
    422, 200, 348, 252, 172, 134, 118, 80, 49, 48, 52, 64, 175, 296, 570, 
    425, 178, 330, 75, 202, 219, 235, 165, 224, 273, 221, 198, 300, 292, 505, 
    438, 123, 196, 33, 110, 84, 109, 239, 248, 257, 233, 233, 275, 147, 427, 
    459, 128, 130, 57, 6, 62, 179, 68, 189, 158, 154, 254, 118, 233, 379, 
    431, 60, 137, 194, 7, 0, 85, 0, 174, 204, 239, 280, 35, 98, 338, 
    397, 227, 204, 226, 74, 0, 0, 0, 37, 381, 377, 205, 0, 58, 335, 
    404, 345, 224, 183, 128, 0, 0, 6, 82, 222, 295, 150, 0, 89, 324, 
    350, 324, 243, 99, 101, 28, 12, 29, 56, 110, 182, 123, 0, 71, 370, 
    
    -- channel=636
    724, 717, 700, 543, 563, 557, 614, 692, 775, 780, 751, 760, 695, 696, 629, 
    795, 796, 759, 418, 424, 440, 428, 496, 612, 708, 699, 756, 761, 705, 742, 
    801, 801, 718, 271, 245, 279, 265, 253, 244, 340, 647, 754, 706, 631, 695, 
    798, 784, 655, 297, 411, 532, 403, 377, 377, 376, 487, 719, 696, 632, 567, 
    798, 769, 521, 239, 348, 353, 336, 325, 377, 387, 444, 630, 778, 711, 628, 
    757, 728, 472, 156, 183, 245, 223, 239, 246, 292, 350, 470, 754, 802, 801, 
    640, 534, 422, 249, 207, 241, 246, 176, 236, 323, 255, 363, 575, 684, 826, 
    582, 286, 429, 374, 180, 122, 77, 93, 92, 83, 80, 131, 222, 334, 761, 
    540, 246, 434, 127, 235, 278, 302, 191, 221, 269, 291, 212, 295, 336, 637, 
    588, 193, 321, 65, 145, 123, 133, 270, 344, 300, 306, 297, 380, 181, 474, 
    599, 209, 172, 106, 22, 82, 179, 81, 221, 159, 164, 270, 95, 279, 402, 
    552, 142, 214, 233, 42, 32, 139, 67, 219, 331, 332, 401, 115, 167, 346, 
    476, 278, 210, 325, 124, 1, 0, 13, 45, 496, 522, 360, 20, 85, 331, 
    481, 440, 288, 291, 179, 50, 4, 37, 136, 310, 381, 287, 0, 108, 329, 
    421, 390, 315, 144, 158, 81, 48, 64, 85, 137, 221, 211, 0, 99, 372, 
    
    -- channel=637
    462, 452, 457, 398, 353, 326, 355, 384, 451, 497, 493, 482, 459, 449, 426, 
    499, 498, 507, 358, 258, 244, 251, 312, 371, 425, 466, 463, 493, 504, 468, 
    506, 505, 489, 278, 61, 91, 85, 98, 103, 166, 333, 467, 483, 463, 435, 
    504, 509, 431, 307, 104, 230, 225, 159, 151, 146, 252, 414, 454, 446, 381, 
    498, 506, 397, 201, 101, 145, 176, 117, 153, 157, 221, 307, 453, 479, 387, 
    452, 499, 307, 153, 34, 77, 86, 84, 92, 104, 168, 223, 399, 507, 505, 
    385, 403, 287, 166, 46, 73, 90, 44, 57, 126, 117, 157, 312, 407, 483, 
    382, 275, 201, 273, 70, 37, 19, 42, 26, 12, 30, 41, 56, 140, 363, 
    363, 220, 204, 186, 51, 129, 112, 86, 60, 68, 140, 70, 81, 158, 266, 
    390, 236, 173, 66, 40, 61, 45, 92, 201, 162, 188, 170, 215, 126, 138, 
    380, 244, 79, 57, 2, 1, 16, 78, 43, 102, 70, 81, 107, 85, 121, 
    336, 220, 80, 91, 50, 0, 47, 75, 39, 171, 160, 221, 117, 84, 62, 
    262, 184, 82, 178, 77, 16, 0, 0, 0, 136, 279, 265, 36, 0, 42, 
    253, 266, 186, 175, 80, 52, 0, 0, 22, 133, 205, 251, 13, 0, 55, 
    231, 207, 195, 110, 68, 47, 7, 6, 13, 39, 84, 149, 10, 0, 56, 
    
    -- channel=638
    307, 297, 316, 251, 220, 229, 244, 263, 299, 318, 304, 299, 303, 265, 246, 
    352, 349, 357, 244, 175, 174, 167, 197, 226, 237, 250, 289, 309, 285, 244, 
    357, 355, 353, 239, 112, 174, 173, 182, 163, 150, 184, 308, 312, 249, 188, 
    356, 359, 309, 277, 143, 258, 262, 219, 225, 216, 225, 238, 299, 284, 191, 
    348, 360, 279, 200, 142, 177, 208, 192, 208, 205, 248, 234, 313, 345, 282, 
    303, 355, 253, 194, 54, 135, 160, 140, 141, 147, 171, 179, 269, 358, 356, 
    274, 286, 197, 159, 125, 155, 174, 121, 122, 167, 121, 107, 192, 253, 334, 
    277, 174, 125, 220, 115, 97, 68, 73, 25, 13, 30, 14, 32, 131, 250, 
    278, 178, 132, 109, 76, 111, 134, 136, 108, 116, 185, 112, 125, 183, 194, 
    298, 182, 87, 39, 22, 57, 30, 61, 178, 136, 159, 137, 171, 119, 96, 
    286, 208, 60, 40, 0, 0, 55, 92, 32, 115, 87, 104, 107, 102, 105, 
    283, 181, 26, 107, 54, 0, 0, 30, 0, 118, 140, 156, 79, 34, 23, 
    249, 225, 106, 157, 83, 1, 0, 0, 0, 99, 250, 243, 17, 0, 42, 
    242, 252, 189, 146, 77, 43, 0, 0, 0, 69, 142, 217, 0, 0, 61, 
    232, 217, 205, 98, 55, 30, 0, 0, 0, 29, 69, 130, 0, 0, 63, 
    
    -- channel=639
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
