library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    24, 47, 31, 33, 25, 40, 36, 44, 27, 0, 8, 25, 40, 42, 39, 
    28, 59, 29, 33, 25, 27, 19, 16, 19, 15, 0, 8, 11, 16, 27, 
    0, 0, 33, 43, 20, 34, 52, 44, 9, 0, 7, 18, 3, 0, 32, 
    48, 0, 27, 29, 18, 15, 12, 0, 0, 0, 50, 14, 48, 16, 0, 
    32, 0, 18, 0, 0, 0, 55, 42, 29, 0, 27, 28, 14, 33, 0, 
    0, 0, 50, 15, 47, 48, 65, 43, 52, 0, 5, 53, 0, 18, 21, 
    11, 2, 25, 92, 0, 0, 0, 25, 56, 0, 47, 37, 8, 4, 15, 
    0, 50, 0, 32, 0, 0, 25, 20, 59, 0, 38, 55, 0, 4, 61, 
    0, 0, 21, 0, 0, 40, 66, 15, 0, 25, 17, 66, 25, 39, 2, 
    12, 0, 59, 0, 12, 0, 6, 25, 0, 3, 35, 30, 0, 0, 16, 
    0, 0, 64, 0, 2, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 43, 8, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 
    30, 19, 0, 0, 1, 183, 14, 10, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 34, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 135, 167, 21, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 11, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 95, 90, 0, 72, 3, 2, 0, 35, 14, 
    0, 0, 0, 0, 0, 153, 0, 0, 0, 36, 62, 109, 58, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 63, 71, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    134, 0, 0, 0, 191, 117, 99, 80, 0, 0, 0, 0, 0, 0, 0, 
    0, 116, 0, 46, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 89, 95, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 89, 
    0, 0, 13, 110, 26, 33, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    46, 32, 54, 35, 37, 39, 40, 45, 37, 13, 17, 40, 36, 23, 19, 
    40, 36, 58, 28, 66, 0, 0, 0, 1, 21, 0, 0, 13, 37, 12, 
    0, 99, 43, 34, 59, 11, 0, 0, 33, 61, 0, 0, 0, 33, 27, 
    0, 98, 4, 54, 0, 72, 0, 0, 0, 151, 0, 0, 0, 0, 111, 
    0, 0, 0, 240, 0, 30, 0, 0, 0, 232, 0, 0, 0, 0, 81, 
    0, 0, 0, 112, 68, 84, 0, 0, 0, 302, 0, 0, 8, 0, 0, 
    43, 0, 6, 0, 91, 99, 0, 0, 0, 189, 0, 0, 0, 2, 0, 
    17, 0, 0, 0, 128, 67, 0, 0, 0, 135, 0, 0, 40, 0, 18, 
    0, 0, 0, 0, 7, 56, 0, 0, 44, 0, 0, 0, 47, 30, 31, 
    0, 0, 0, 61, 0, 106, 109, 0, 0, 3, 0, 0, 26, 45, 4, 
    0, 0, 0, 251, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 42, 0, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 63, 216, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 250, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    
    -- channel=3
    1, 0, 0, 0, 3, 0, 0, 4, 7, 0, 0, 0, 0, 0, 1, 
    6, 0, 0, 0, 0, 0, 5, 0, 0, 55, 28, 83, 86, 0, 0, 
    0, 0, 3, 5, 5, 80, 53, 167, 37, 0, 0, 0, 0, 44, 0, 
    15, 82, 12, 8, 3, 62, 0, 0, 0, 0, 0, 0, 8, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 35, 0, 0, 0, 42, 
    0, 0, 0, 1, 75, 0, 0, 12, 0, 0, 0, 8, 0, 0, 0, 
    21, 0, 57, 0, 11, 0, 0, 0, 0, 0, 7, 35, 50, 2, 0, 
    0, 6, 25, 16, 0, 0, 0, 0, 0, 0, 0, 74, 0, 0, 8, 
    0, 0, 0, 0, 0, 99, 113, 29, 0, 130, 59, 3, 49, 21, 0, 
    0, 0, 0, 85, 0, 0, 52, 0, 23, 0, 0, 10, 0, 0, 0, 
    9, 5, 31, 18, 0, 0, 0, 0, 0, 29, 52, 0, 0, 50, 51, 
    30, 0, 0, 0, 0, 156, 177, 170, 54, 0, 0, 0, 7, 9, 0, 
    0, 46, 23, 0, 98, 0, 0, 0, 6, 0, 0, 0, 0, 0, 1, 
    0, 0, 11, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 16, 156, 30, 7, 0, 0, 0, 2, 0, 18, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 51, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 6, 160, 0, 0, 0, 0, 0, 0, 
    74, 0, 0, 0, 0, 120, 9, 10, 0, 0, 12, 0, 80, 0, 0, 
    128, 0, 0, 0, 0, 0, 0, 20, 2, 0, 25, 38, 13, 0, 0, 
    79, 0, 29, 0, 0, 21, 50, 0, 42, 0, 0, 52, 0, 25, 0, 
    67, 0, 0, 25, 0, 0, 0, 10, 44, 0, 98, 61, 0, 15, 0, 
    0, 75, 0, 57, 0, 0, 94, 0, 104, 0, 82, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 189, 46, 0, 0, 11, 13, 0, 18, 0, 
    0, 0, 35, 0, 0, 86, 0, 0, 0, 100, 0, 129, 0, 0, 0, 
    0, 0, 68, 0, 41, 0, 0, 0, 0, 69, 189, 20, 0, 0, 21, 
    0, 0, 112, 0, 0, 0, 14, 136, 139, 56, 0, 0, 0, 0, 15, 
    53, 0, 1, 0, 376, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 89, 156, 0, 18, 0, 0, 0, 0, 0, 25, 18, 0, 
    15, 0, 0, 199, 15, 0, 0, 0, 0, 0, 3, 2, 0, 0, 152, 
    42, 0, 0, 85, 43, 0, 26, 0, 0, 0, 9, 0, 0, 10, 82, 
    
    -- channel=5
    66, 86, 79, 88, 88, 69, 84, 92, 95, 71, 62, 55, 73, 81, 90, 
    87, 80, 69, 94, 60, 151, 100, 104, 64, 30, 69, 50, 20, 35, 87, 
    126, 0, 86, 97, 72, 0, 141, 23, 0, 0, 29, 28, 83, 0, 49, 
    181, 0, 75, 71, 150, 5, 78, 39, 40, 0, 133, 0, 77, 69, 0, 
    102, 0, 112, 0, 105, 10, 95, 107, 71, 0, 22, 100, 30, 99, 0, 
    0, 12, 140, 67, 0, 0, 165, 50, 166, 0, 106, 101, 0, 46, 61, 
    0, 121, 22, 184, 0, 0, 31, 100, 114, 0, 109, 86, 1, 0, 59, 
    23, 64, 0, 110, 0, 0, 131, 16, 83, 0, 99, 88, 0, 0, 50, 
    59, 0, 161, 0, 73, 0, 39, 77, 0, 67, 0, 103, 0, 3, 48, 
    26, 0, 196, 0, 36, 0, 0, 82, 3, 26, 101, 0, 0, 13, 79, 
    0, 0, 152, 0, 248, 16, 0, 9, 110, 67, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 133, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 62, 109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 184, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 61, 51, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 95, 0, 0, 0, 0, 52, 0, 
    16, 168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 76, 
    0, 0, 0, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 90, 84, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 74, 0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 128, 43, 22, 7, 0, 0, 0, 8, 8, 0, 
    0, 0, 0, 34, 0, 38, 0, 0, 40, 0, 0, 41, 0, 0, 0, 
    0, 0, 0, 0, 27, 16, 0, 0, 0, 161, 85, 38, 48, 0, 0, 
    14, 0, 0, 0, 0, 0, 107, 181, 139, 0, 0, 0, 0, 23, 19, 
    133, 135, 67, 0, 0, 30, 0, 0, 3, 3, 1, 0, 0, 0, 0, 
    0, 53, 101, 0, 51, 0, 0, 0, 0, 0, 0, 0, 4, 26, 0, 
    0, 0, 114, 79, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 21, 0, 11, 72, 23, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 20, 36, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 22, 0, 30, 0, 26, 15, 0, 
    60, 18, 0, 0, 0, 0, 13, 23, 35, 0, 5, 19, 16, 39, 0, 
    24, 44, 0, 0, 0, 0, 47, 0, 77, 0, 25, 14, 0, 25, 20, 
    7, 122, 0, 0, 0, 0, 13, 13, 46, 0, 38, 35, 17, 16, 6, 
    34, 88, 0, 0, 0, 0, 21, 0, 0, 0, 32, 37, 0, 0, 0, 
    84, 68, 83, 13, 0, 0, 0, 39, 0, 0, 0, 6, 0, 0, 0, 
    56, 56, 121, 41, 16, 0, 0, 73, 1, 0, 19, 4, 0, 0, 0, 
    68, 36, 103, 0, 166, 64, 49, 61, 75, 65, 86, 115, 121, 80, 80, 
    106, 67, 32, 38, 141, 129, 132, 127, 155, 152, 177, 186, 204, 204, 204, 
    249, 105, 0, 120, 126, 174, 175, 168, 175, 186, 205, 211, 207, 202, 225, 
    260, 219, 34, 191, 150, 172, 191, 174, 176, 194, 218, 219, 231, 242, 252, 
    258, 241, 205, 145, 166, 166, 166, 171, 182, 210, 214, 200, 205, 275, 259, 
    
    -- channel=8
    213, 227, 225, 226, 225, 213, 235, 253, 225, 169, 136, 149, 174, 199, 196, 
    221, 242, 238, 234, 223, 232, 192, 181, 129, 61, 39, 48, 76, 132, 180, 
    132, 144, 234, 242, 243, 214, 111, 51, 23, 59, 28, 16, 44, 47, 150, 
    47, 102, 206, 230, 193, 110, 90, 28, 28, 42, 58, 47, 18, 25, 104, 
    0, 93, 167, 127, 110, 103, 64, 34, 34, 37, 55, 39, 34, 24, 58, 
    0, 43, 147, 212, 81, 53, 93, 47, 50, 61, 44, 4, 22, 15, 22, 
    0, 76, 72, 183, 142, 84, 61, 45, 25, 85, 15, 16, 27, 21, 40, 
    0, 14, 8, 89, 107, 66, 34, 42, 29, 130, 50, 21, 13, 52, 104, 
    0, 0, 0, 34, 63, 51, 45, 55, 18, 131, 38, 14, 37, 104, 185, 
    22, 13, 0, 32, 0, 27, 27, 61, 33, 20, 13, 0, 37, 163, 162, 
    5, 11, 0, 18, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    102, 118, 103, 99, 100, 97, 115, 143, 126, 112, 104, 101, 77, 78, 91, 
    98, 117, 116, 110, 102, 0, 34, 117, 147, 0, 0, 0, 20, 80, 71, 
    111, 154, 112, 121, 128, 194, 52, 12, 0, 0, 0, 0, 0, 0, 59, 
    0, 0, 75, 119, 75, 4, 0, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 109, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 74, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 62, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    35, 36, 25, 36, 35, 28, 33, 36, 37, 44, 24, 17, 18, 26, 42, 
    38, 38, 28, 40, 30, 80, 2, 29, 21, 28, 40, 28, 19, 39, 46, 
    47, 38, 39, 40, 45, 96, 15, 17, 2, 44, 20, 0, 40, 22, 56, 
    73, 46, 53, 35, 43, 6, 66, 0, 29, 13, 10, 15, 25, 28, 45, 
    0, 86, 0, 0, 53, 0, 0, 0, 41, 0, 24, 0, 38, 42, 0, 
    0, 52, 0, 0, 73, 0, 40, 7, 75, 13, 0, 0, 31, 17, 0, 
    0, 109, 0, 66, 78, 0, 68, 0, 54, 68, 0, 3, 17, 37, 17, 
    0, 43, 0, 75, 13, 64, 0, 4, 27, 56, 9, 21, 17, 26, 0, 
    0, 1, 0, 52, 0, 0, 24, 72, 7, 51, 83, 0, 21, 47, 41, 
    0, 0, 18, 25, 9, 0, 0, 99, 0, 3, 10, 19, 49, 52, 25, 
    102, 0, 23, 0, 0, 0, 0, 0, 0, 0, 34, 23, 11, 61, 52, 
    67, 0, 0, 64, 46, 0, 29, 22, 26, 35, 43, 35, 39, 35, 29, 
    39, 26, 0, 104, 0, 18, 25, 26, 37, 40, 40, 35, 33, 20, 24, 
    37, 31, 0, 139, 12, 20, 26, 29, 20, 23, 32, 49, 33, 40, 61, 
    24, 35, 25, 115, 47, 44, 35, 16, 24, 34, 38, 24, 29, 59, 40, 
    
    -- channel=11
    78, 89, 79, 82, 77, 84, 90, 86, 75, 78, 69, 65, 61, 63, 51, 
    73, 86, 83, 89, 75, 130, 89, 96, 60, 29, 41, 42, 46, 55, 61, 
    99, 60, 87, 84, 86, 145, 62, 13, 0, 63, 84, 33, 41, 24, 63, 
    57, 41, 93, 84, 98, 33, 90, 25, 29, 70, 87, 59, 19, 3, 37, 
    51, 140, 89, 33, 172, 98, 113, 45, 36, 0, 98, 51, 33, 8, 4, 
    64, 169, 96, 85, 187, 100, 147, 59, 46, 70, 138, 38, 41, 18, 0, 
    35, 202, 83, 76, 109, 116, 198, 85, 65, 126, 108, 44, 26, 39, 42, 
    95, 144, 46, 84, 47, 203, 123, 96, 49, 122, 102, 53, 33, 75, 30, 
    141, 168, 75, 103, 71, 70, 66, 78, 42, 87, 105, 23, 9, 40, 80, 
    160, 159, 112, 83, 106, 18, 35, 135, 72, 77, 26, 0, 32, 93, 82, 
    179, 155, 115, 111, 150, 94, 148, 161, 72, 0, 0, 0, 30, 62, 48, 
    132, 137, 100, 251, 251, 45, 51, 40, 21, 10, 22, 21, 26, 37, 29, 
    32, 96, 78, 302, 38, 21, 24, 16, 9, 8, 12, 30, 48, 30, 33, 
    23, 25, 101, 221, 22, 23, 20, 20, 13, 21, 27, 38, 17, 38, 87, 
    33, 22, 42, 72, 13, 21, 27, 15, 24, 33, 30, 7, 27, 81, 16, 
    
    -- channel=12
    0, 7, 8, 3, 0, 16, 0, 0, 11, 0, 0, 0, 0, 0, 1, 
    10, 26, 11, 0, 8, 172, 0, 33, 0, 30, 32, 14, 0, 0, 12, 
    21, 0, 11, 0, 14, 0, 0, 0, 31, 90, 0, 0, 0, 0, 30, 
    0, 163, 0, 20, 53, 0, 66, 0, 0, 18, 0, 0, 0, 0, 30, 
    0, 142, 0, 4, 133, 0, 0, 0, 0, 53, 0, 0, 22, 0, 17, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 300, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 60, 105, 0, 0, 0, 204, 0, 0, 0, 37, 0, 
    0, 0, 0, 0, 17, 131, 0, 0, 0, 112, 0, 0, 6, 0, 0, 
    0, 0, 0, 41, 13, 0, 0, 62, 0, 0, 39, 0, 0, 8, 63, 
    0, 0, 0, 32, 0, 0, 0, 44, 0, 0, 0, 0, 74, 85, 0, 
    71, 0, 0, 235, 0, 61, 97, 0, 0, 0, 46, 95, 37, 0, 0, 
    0, 0, 0, 186, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 28, 0, 
    0, 84, 0, 0, 0, 197, 0, 0, 0, 47, 0, 0, 0, 19, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 0, 0, 0, 0, 146, 
    0, 15, 0, 59, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 
    0, 45, 0, 0, 346, 0, 0, 0, 0, 146, 0, 0, 54, 0, 0, 
    0, 0, 4, 0, 215, 0, 89, 0, 0, 190, 0, 0, 0, 4, 0, 
    0, 25, 0, 0, 62, 212, 0, 7, 0, 135, 0, 0, 54, 7, 0, 
    0, 14, 0, 97, 0, 95, 17, 0, 45, 0, 182, 0, 29, 67, 0, 
    0, 0, 0, 77, 0, 0, 0, 0, 0, 42, 0, 34, 68, 2, 0, 
    180, 0, 0, 133, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    256, 58, 0, 81, 0, 0, 60, 61, 7, 0, 0, 0, 0, 0, 0, 
    0, 139, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 130, 67, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 256, 0, 50, 48, 0, 0, 0, 0, 0, 11, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    144, 139, 147, 151, 146, 131, 156, 171, 155, 116, 90, 102, 113, 121, 127, 
    154, 153, 154, 152, 158, 102, 118, 110, 57, 42, 0, 0, 32, 110, 125, 
    55, 124, 161, 160, 159, 77, 57, 21, 34, 0, 0, 0, 0, 38, 98, 
    0, 50, 145, 159, 102, 90, 20, 0, 0, 22, 0, 0, 0, 0, 70, 
    0, 0, 105, 159, 23, 0, 0, 0, 0, 34, 0, 0, 0, 0, 5, 
    0, 0, 110, 47, 6, 18, 0, 0, 0, 44, 0, 0, 0, 0, 0, 
    0, 0, 94, 98, 0, 37, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 55, 54, 17, 0, 0, 20, 0, 0, 0, 0, 0, 71, 
    0, 0, 0, 0, 17, 0, 18, 0, 32, 0, 47, 0, 0, 55, 94, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 26, 0, 0, 2, 75, 106, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 9, 0, 0, 0, 45, 11, 14, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 8, 0, 11, 0, 0, 0, 3, 46, 43, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 5, 3, 18, 19, 6, 24, 0, 32, 0, 0, 0, 
    80, 82, 101, 91, 77, 63, 59, 46, 47, 61, 45, 38, 33, 17, 0, 
    47, 0, 48, 49, 54, 49, 53, 54, 65, 69, 65, 22, 9, 41, 0, 
    42, 24, 93, 91, 58, 47, 28, 281, 247, 199, 144, 136, 36, 0, 0, 
    58, 43, 47, 57, 46, 43, 101, 398, 310, 174, 47, 0, 0, 0, 0, 
    54, 26, 18, 28, 37, 29, 19, 134, 55, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 76, 12, 46, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    266, 209, 0, 0, 0, 0, 0, 0, 0, 0, 76, 174, 212, 83, 0, 
    0, 0, 0, 70, 51, 212, 224, 174, 77, 0, 0, 0, 0, 0, 0, 
    287, 270, 98, 0, 0, 0, 0, 0, 0, 14, 118, 186, 136, 186, 116, 
    5, 0, 61, 79, 0, 0, 0, 15, 152, 62, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 45, 0, 0, 0, 0, 43, 119, 187, 109, 
    140, 211, 214, 191, 163, 104, 59, 24, 38, 3, 79, 40, 0, 0, 1, 
    213, 188, 239, 299, 340, 346, 306, 260, 215, 186, 123, 67, 0, 0, 0, 
    17, 18, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 12, 12, 0, 
    0, 59, 113, 57, 6, 6, 213, 142, 105, 144, 228, 120, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 59, 96, 139, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 59, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 34, 0, 0, 0, 
    0, 70, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 131, 0, 
    0, 0, 0, 0, 0, 0, 49, 49, 65, 0, 0, 0, 0, 72, 0, 
    0, 105, 10, 45, 0, 0, 0, 14, 70, 0, 0, 0, 15, 0, 97, 
    163, 0, 0, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    369, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 34, 0, 26, 54, 83, 39, 34, 0, 0, 0, 4, 21, 0, 27, 
    0, 121, 0, 0, 0, 55, 74, 0, 0, 0, 0, 0, 20, 15, 44, 
    0, 43, 24, 0, 0, 8, 324, 94, 109, 80, 65, 58, 26, 30, 43, 
    0, 0, 9, 0, 0, 1, 192, 115, 102, 76, 39, 31, 0, 37, 34, 
    0, 0, 0, 0, 0, 0, 50, 23, 38, 71, 4, 0, 10, 23, 25, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 15, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 18, 13, 0, 4, 50, 63, 0, 0, 0, 
    232, 182, 16, 0, 0, 1, 0, 0, 0, 0, 0, 0, 64, 58, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 33, 0, 0, 0, 0, 
    118, 165, 66, 0, 0, 155, 244, 340, 105, 0, 0, 0, 0, 0, 5, 
    17, 0, 104, 119, 99, 0, 0, 0, 120, 236, 262, 204, 158, 82, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 
    0, 0, 36, 55, 82, 99, 113, 141, 91, 59, 54, 51, 0, 0, 0, 
    200, 199, 182, 143, 106, 72, 32, 7, 4, 29, 35, 36, 83, 27, 0, 
    0, 0, 0, 0, 0, 0, 18, 153, 180, 147, 91, 0, 0, 10, 11, 
    0, 11, 67, 32, 0, 0, 24, 0, 0, 0, 0, 146, 59, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 142, 63, 0, 0, 0, 0, 
    12, 0, 4, 9, 13, 18, 38, 146, 59, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 54, 16, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 119, 124, 78, 0, 0, 
    0, 0, 24, 43, 0, 258, 178, 136, 54, 0, 0, 0, 0, 0, 0, 
    88, 36, 0, 0, 68, 28, 0, 0, 0, 27, 133, 165, 101, 178, 0, 
    0, 0, 0, 0, 0, 0, 0, 148, 53, 0, 0, 0, 0, 0, 0, 
    0, 61, 0, 0, 22, 55, 25, 65, 11, 147, 65, 169, 159, 130, 0, 
    210, 119, 95, 66, 37, 0, 19, 0, 0, 0, 39, 1, 0, 0, 0, 
    48, 0, 45, 73, 100, 114, 120, 128, 107, 99, 48, 2, 0, 0, 0, 
    49, 0, 28, 53, 40, 0, 0, 0, 0, 0, 0, 0, 80, 0, 0, 
    67, 8, 24, 43, 10, 11, 0, 1, 43, 116, 187, 0, 0, 0, 0, 
    117, 10, 12, 16, 9, 9, 0, 0, 169, 0, 0, 0, 0, 0, 0, 
    92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 55, 0, 36, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 2, 0, 76, 0, 0, 
    0, 0, 0, 0, 60, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 53, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 0, 71, 76, 28, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 
    89, 0, 0, 38, 30, 15, 0, 27, 31, 43, 16, 0, 0, 0, 0, 
    208, 22, 9, 25, 21, 18, 0, 49, 64, 12, 0, 0, 0, 0, 0, 
    148, 50, 32, 28, 26, 20, 0, 0, 2, 0, 1, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 29, 72, 66, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 62, 26, 0, 0, 0, 0, 0, 0, 0, 82, 87, 69, 128, 0, 
    0, 0, 0, 31, 30, 239, 328, 296, 201, 0, 0, 0, 0, 0, 0, 
    92, 114, 92, 46, 0, 0, 0, 0, 0, 24, 150, 193, 247, 137, 137, 
    122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 3, 15, 46, 32, 78, 201, 108, 196, 206, 189, 216, 110, 14, 
    148, 175, 115, 113, 65, 36, 0, 0, 0, 0, 0, 5, 0, 34, 0, 
    0, 0, 0, 32, 90, 141, 168, 194, 143, 106, 77, 27, 0, 0, 0, 
    45, 95, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 
    0, 0, 17, 14, 0, 0, 107, 163, 109, 114, 107, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 33, 71, 126, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    57, 56, 56, 56, 55, 56, 55, 55, 51, 61, 63, 55, 56, 56, 56, 
    56, 56, 56, 57, 56, 57, 55, 56, 62, 98, 56, 51, 56, 57, 57, 
    51, 52, 55, 57, 55, 62, 53, 83, 72, 98, 47, 40, 55, 55, 57, 
    73, 71, 58, 53, 55, 92, 39, 88, 100, 127, 123, 68, 70, 65, 61, 
    69, 28, 56, 44, 54, 75, 55, 65, 75, 95, 96, 82, 61, 7, 67, 
    106, 104, 83, 24, 56, 24, 24, 26, 34, 113, 114, 110, 142, 73, 65, 
    79, 29, 46, 53, 136, 125, 104, 101, 60, 69, 55, 45, 33, 62, 24, 
    18, 132, 52, 21, 74, 112, 100, 108, 71, 88, 107, 102, 92, 102, 87, 
    0, 101, 88, 67, 76, 89, 81, 92, 98, 94, 109, 111, 90, 84, 90, 
    85, 98, 116, 120, 126, 131, 160, 143, 137, 138, 136, 130, 118, 95, 81, 
    49, 70, 81, 67, 52, 55, 103, 99, 116, 114, 109, 105, 105, 93, 53, 
    23, 0, 51, 50, 25, 9, 109, 166, 146, 132, 106, 85, 44, 34, 24, 
    27, 2, 0, 0, 5, 7, 0, 0, 0, 0, 0, 0, 0, 16, 35, 
    67, 4, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 13, 17, 40, 
    31, 5, 9, 10, 6, 10, 0, 0, 0, 0, 0, 9, 13, 28, 47, 
    
    -- channel=24
    18, 20, 20, 20, 20, 20, 20, 24, 25, 17, 13, 18, 21, 20, 21, 
    18, 20, 20, 21, 20, 20, 20, 22, 17, 9, 0, 11, 21, 20, 21, 
    18, 20, 22, 22, 22, 20, 11, 11, 0, 0, 0, 2, 19, 21, 20, 
    0, 0, 13, 23, 24, 34, 12, 1, 0, 0, 0, 3, 0, 6, 14, 
    0, 0, 0, 24, 19, 8, 31, 6, 11, 0, 0, 0, 0, 0, 6, 
    0, 7, 45, 3, 4, 0, 0, 0, 0, 0, 0, 0, 7, 24, 1, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 4, 39, 0, 0, 18, 32, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 9, 17, 7, 0, 15, 0, 0, 0, 0, 9, 41, 23, 19, 
    20, 24, 27, 13, 6, 17, 87, 153, 181, 161, 122, 61, 27, 34, 16, 
    7, 17, 21, 13, 14, 14, 111, 276, 223, 106, 60, 69, 35, 15, 9, 
    0, 35, 25, 19, 24, 18, 56, 95, 60, 99, 70, 21, 18, 14, 9, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 70, 71, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 57, 18, 0, 0, 84, 48, 11, 43, 98, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 53, 308, 339, 113, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    21, 0, 36, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 21, 5, 0, 0, 3, 0, 
    0, 0, 5, 0, 68, 0, 30, 24, 1, 0, 0, 0, 0, 0, 0, 
    0, 63, 0, 17, 16, 0, 0, 3, 0, 0, 5, 17, 11, 19, 0, 
    0, 42, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 6, 0, 3, 0, 0, 0, 0, 
    15, 24, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 19, 6, 5, 14, 0, 35, 4, 14, 0, 0, 0, 0, 0, 2, 
    30, 28, 17, 5, 22, 30, 0, 0, 0, 0, 0, 0, 0, 14, 25, 
    56, 36, 29, 24, 32, 34, 0, 0, 0, 0, 0, 19, 26, 24, 37, 
    49, 56, 61, 57, 47, 47, 9, 0, 0, 11, 24, 38, 38, 28, 33, 
    
    -- channel=27
    235, 236, 236, 236, 236, 237, 236, 238, 234, 237, 236, 236, 236, 236, 237, 
    236, 237, 237, 237, 236, 237, 236, 236, 239, 244, 208, 229, 236, 236, 238, 
    235, 236, 237, 237, 237, 242, 231, 246, 204, 172, 187, 212, 239, 238, 239, 
    229, 234, 241, 239, 241, 256, 215, 210, 163, 158, 146, 209, 240, 239, 241, 
    152, 153, 227, 234, 238, 227, 230, 228, 225, 233, 230, 201, 189, 169, 241, 
    137, 159, 242, 212, 231, 217, 205, 210, 201, 213, 163, 153, 145, 188, 236, 
    131, 120, 176, 150, 225, 35, 29, 62, 172, 244, 229, 205, 192, 202, 177, 
    0, 120, 90, 158, 167, 128, 161, 218, 170, 131, 98, 84, 92, 117, 163, 
    3, 204, 150, 198, 226, 237, 239, 176, 153, 165, 166, 172, 156, 146, 126, 
    157, 136, 144, 144, 142, 138, 134, 104, 121, 78, 93, 61, 57, 69, 86, 
    0, 0, 7, 5, 17, 24, 47, 48, 52, 32, 19, 17, 20, 61, 85, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 88, 65, 87, 
    0, 0, 0, 0, 0, 0, 42, 102, 90, 91, 77, 34, 47, 83, 127, 
    0, 0, 0, 0, 0, 0, 0, 92, 40, 0, 11, 71, 81, 97, 145, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 83, 75, 91, 111, 152, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 144, 0, 
    0, 0, 0, 0, 0, 0, 0, 48, 145, 0, 0, 0, 0, 0, 0, 
    0, 231, 0, 0, 0, 13, 132, 0, 0, 0, 0, 0, 0, 35, 49, 
    375, 0, 44, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 48, 6, 5, 9, 38, 175, 90, 66, 80, 104, 143, 0, 0, 18, 
    0, 39, 0, 0, 8, 39, 98, 0, 0, 0, 0, 0, 37, 18, 39, 
    0, 37, 41, 21, 36, 38, 84, 56, 0, 0, 105, 106, 0, 4, 0, 
    0, 44, 57, 45, 53, 55, 84, 36, 121, 135, 22, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 60, 55, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 
    133, 189, 126, 0, 0, 0, 0, 0, 0, 0, 0, 20, 76, 176, 0, 
    0, 0, 0, 0, 22, 65, 133, 114, 82, 0, 0, 0, 0, 0, 0, 
    123, 208, 172, 0, 0, 0, 0, 0, 16, 3, 14, 28, 117, 43, 124, 
    173, 0, 0, 140, 69, 0, 0, 0, 24, 16, 0, 0, 0, 0, 0, 
    33, 50, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 30, 52, 60, 
    109, 104, 119, 114, 87, 87, 40, 2, 58, 0, 49, 27, 11, 6, 15, 
    63, 125, 104, 156, 194, 213, 193, 164, 122, 88, 81, 52, 39, 0, 8, 
    0, 125, 0, 0, 0, 12, 43, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 103, 31, 0, 0, 345, 99, 16, 1, 12, 77, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 14, 61, 13, 24, 0, 0, 0, 0, 28, 
    0, 0, 0, 0, 0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 8, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 21, 0, 0, 0, 0, 
    1, 2, 0, 0, 0, 0, 0, 0, 31, 16, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 
    4, 0, 0, 9, 3, 0, 0, 0, 0, 82, 0, 16, 0, 0, 0, 
    31, 2, 26, 0, 24, 5, 0, 6, 0, 0, 0, 0, 0, 42, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 3, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 64, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 15, 
    0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 16, 0, 1, 7, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 17, 7, 40, 
    0, 0, 0, 0, 0, 20, 18, 0, 0, 2, 6, 0, 27, 17, 14, 
    33, 34, 12, 0, 0, 0, 0, 7, 0, 0, 19, 16, 19, 10, 16, 
    21, 8, 0, 0, 0, 0, 0, 13, 0, 34, 21, 29, 9, 9, 44, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 82, 34, 71, 30, 48, 3, 8, 0, 
    32, 3, 58, 42, 35, 6, 1, 0, 171, 122, 115, 273, 157, 89, 116, 
    169, 137, 148, 179, 174, 173, 118, 83, 0, 0, 0, 0, 0, 41, 116, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 94, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 85, 94, 2, 0, 0, 0, 
    7, 97, 28, 0, 8, 53, 49, 0, 0, 0, 0, 0, 0, 0, 76, 
    0, 0, 0, 29, 0, 0, 0, 43, 58, 0, 0, 8, 102, 125, 93, 
    0, 0, 0, 34, 112, 45, 33, 63, 1, 64, 127, 105, 49, 27, 53, 
    21, 8, 21, 10, 0, 0, 67, 4, 25, 34, 50, 50, 5, 26, 10, 
    55, 111, 119, 78, 122, 118, 14, 0, 67, 64, 0, 24, 28, 0, 0, 
    120, 102, 53, 27, 31, 49, 46, 26, 0, 0, 17, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 29, 29, 8, 4, 0, 0, 0, 46, 
    
    -- channel=34
    0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 68, 2, 0, 0, 0, 0, 0, 0, 0, 119, 5, 0, 0, 24, 
    0, 92, 30, 0, 0, 0, 0, 1, 57, 0, 170, 65, 0, 0, 26, 
    0, 115, 21, 44, 0, 9, 0, 0, 0, 0, 0, 48, 123, 0, 99, 
    0, 39, 0, 36, 12, 34, 27, 0, 0, 0, 0, 34, 80, 0, 40, 
    0, 29, 0, 31, 0, 0, 0, 0, 0, 0, 97, 0, 0, 0, 0, 
    0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 53, 6, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 23, 0, 0, 0, 
    0, 0, 52, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 7, 
    4, 0, 0, 0, 0, 21, 0, 0, 95, 0, 0, 0, 0, 0, 0, 
    40, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 99, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 101, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 7, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 68, 266, 239, 325, 57, 0, 0, 
    69, 54, 147, 97, 89, 57, 69, 26, 0, 0, 0, 0, 0, 90, 118, 
    38, 0, 0, 57, 19, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 59, 35, 101, 44, 63, 44, 40, 22, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 36, 4, 61, 110, 
    0, 0, 101, 0, 0, 0, 49, 86, 20, 0, 0, 0, 13, 0, 0, 
    126, 0, 0, 10, 76, 0, 0, 0, 0, 0, 0, 0, 0, 30, 70, 
    0, 0, 0, 0, 0, 0, 23, 162, 121, 0, 0, 68, 0, 3, 0, 
    9, 16, 37, 132, 92, 0, 0, 0, 0, 57, 0, 33, 37, 0, 26, 
    0, 0, 0, 0, 15, 119, 50, 0, 0, 39, 12, 0, 0, 5, 0, 
    75, 80, 33, 0, 0, 0, 42, 49, 0, 0, 7, 0, 2, 0, 0, 
    0, 3, 19, 26, 5, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 0, 176, 0, 0, 0, 0, 0, 
    58, 0, 1, 0, 17, 0, 23, 13, 163, 0, 0, 0, 0, 47, 26, 
    51, 40, 13, 33, 35, 60, 22, 101, 0, 38, 16, 0, 23, 0, 0, 
    0, 0, 44, 0, 0, 0, 0, 27, 0, 0, 0, 0, 1, 0, 144, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 124, 109, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 107, 0, 0, 0, 0, 0, 
    5, 99, 0, 0, 19, 48, 0, 0, 0, 0, 0, 0, 0, 0, 94, 
    0, 0, 18, 21, 0, 0, 0, 85, 53, 0, 0, 25, 124, 93, 3, 
    0, 0, 0, 69, 84, 0, 50, 5, 0, 38, 111, 55, 46, 35, 88, 
    0, 0, 38, 0, 0, 0, 131, 70, 7, 0, 71, 48, 0, 30, 10, 
    16, 107, 126, 86, 65, 0, 0, 9, 86, 27, 0, 14, 65, 0, 2, 
    24, 0, 0, 0, 36, 52, 9, 0, 0, 82, 11, 17, 1, 0, 0, 
    7, 0, 0, 0, 0, 0, 21, 41, 0, 61, 16, 0, 1, 0, 108, 
    
    -- channel=37
    6, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 28, 0, 0, 179, 0, 0, 7, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 61, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 104, 0, 
    0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 0, 136, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 0, 143, 68, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 25, 0, 
    0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 8, 14, 0, 17, 
    0, 0, 39, 0, 0, 0, 6, 9, 0, 0, 0, 0, 11, 7, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 28, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 4, 0, 12, 
    10, 0, 0, 0, 0, 0, 0, 15, 0, 62, 0, 3, 0, 0, 51, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 17, 41, 0, 60, 111, 0, 0, 0, 
    34, 32, 56, 74, 16, 0, 0, 0, 0, 0, 0, 0, 195, 103, 112, 
    90, 50, 2, 52, 80, 94, 82, 55, 42, 8, 23, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 7, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 16, 0, 0, 0, 0, 
    28, 66, 0, 0, 12, 40, 0, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 7, 0, 0, 0, 0, 63, 126, 0, 0, 6, 71, 39, 13, 
    33, 0, 0, 69, 94, 62, 0, 0, 0, 57, 71, 19, 36, 32, 21, 
    0, 0, 0, 0, 0, 0, 134, 93, 0, 0, 40, 0, 0, 0, 0, 
    77, 122, 149, 104, 17, 0, 0, 14, 49, 1, 0, 6, 10, 0, 0, 
    0, 0, 0, 14, 40, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 23, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    180, 102, 142, 123, 121, 87, 83, 98, 72, 76, 51, 61, 66, 85, 50, 
    149, 69, 92, 86, 87, 64, 73, 77, 58, 119, 0, 45, 55, 70, 40, 
    114, 28, 48, 52, 55, 49, 79, 28, 16, 145, 1, 18, 52, 42, 30, 
    68, 0, 16, 0, 5, 13, 31, 79, 86, 85, 86, 14, 0, 12, 0, 
    37, 25, 32, 2, 0, 0, 18, 82, 96, 115, 95, 42, 4, 76, 0, 
    95, 52, 110, 59, 113, 90, 129, 129, 102, 110, 45, 68, 101, 20, 39, 
    117, 93, 95, 98, 111, 148, 161, 156, 156, 135, 58, 24, 44, 0, 38, 
    137, 134, 135, 151, 151, 153, 155, 148, 117, 116, 22, 7, 28, 83, 81, 
    143, 120, 109, 146, 155, 146, 141, 125, 85, 109, 57, 52, 57, 48, 9, 
    160, 139, 151, 147, 143, 138, 123, 101, 55, 86, 75, 76, 57, 51, 27, 
    153, 162, 152, 132, 106, 106, 157, 97, 43, 75, 72, 73, 66, 53, 58, 
    120, 139, 181, 121, 124, 96, 100, 88, 79, 78, 73, 78, 75, 66, 48, 
    88, 102, 102, 96, 90, 79, 77, 79, 73, 76, 70, 55, 68, 56, 56, 
    70, 61, 67, 61, 64, 62, 70, 73, 51, 91, 60, 58, 57, 57, 57, 
    46, 45, 57, 59, 63, 66, 69, 58, 24, 80, 56, 52, 55, 52, 50, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 6, 9, 6, 6, 17, 2, 18, 6, 
    0, 0, 0, 0, 11, 8, 18, 15, 11, 20, 0, 20, 11, 27, 17, 
    0, 0, 10, 16, 43, 20, 36, 15, 0, 5, 0, 2, 19, 42, 31, 
    2, 0, 42, 44, 62, 50, 31, 29, 0, 0, 0, 0, 0, 38, 44, 
    0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 39, 72, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 68, 57, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 42, 13, 28, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 22, 15, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 12, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 
    0, 0, 0, 3, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    18, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 5, 0, 0, 9, 0, 35, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 26, 0, 35, 0, 0, 46, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 2, 21, 2, 25, 24, 0, 28, 7, 0, 
    0, 0, 15, 7, 0, 0, 0, 41, 0, 22, 7, 0, 0, 55, 0, 
    34, 0, 34, 0, 49, 7, 20, 6, 11, 36, 0, 15, 11, 121, 0, 
    31, 0, 4, 0, 14, 3, 21, 0, 29, 41, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 20, 0, 0, 0, 0, 60, 
    0, 0, 0, 0, 0, 0, 20, 32, 4, 16, 0, 0, 0, 0, 10, 
    0, 10, 4, 0, 1, 18, 13, 5, 0, 18, 0, 3, 4, 8, 0, 
    7, 6, 6, 1, 5, 6, 59, 1, 0, 48, 13, 22, 35, 26, 52, 
    50, 7, 55, 8, 28, 38, 12, 0, 14, 40, 45, 47, 47, 36, 31, 
    19, 4, 17, 1, 27, 38, 26, 35, 34, 42, 42, 24, 32, 30, 33, 
    32, 28, 44, 37, 40, 43, 44, 54, 24, 45, 33, 28, 31, 37, 39, 
    38, 38, 50, 48, 50, 46, 51, 46, 19, 23, 37, 21, 34, 34, 53, 
    
    -- channel=43
    175, 122, 199, 206, 225, 214, 236, 243, 233, 252, 231, 241, 230, 253, 228, 
    185, 129, 205, 209, 234, 215, 240, 242, 229, 260, 161, 242, 235, 259, 229, 
    188, 119, 199, 205, 239, 208, 239, 207, 202, 205, 149, 220, 233, 243, 229, 
    180, 111, 207, 197, 220, 201, 203, 196, 148, 77, 74, 96, 161, 222, 189, 
    98, 77, 108, 130, 140, 144, 129, 140, 62, 68, 47, 32, 93, 162, 107, 
    27, 31, 74, 21, 80, 71, 95, 79, 62, 57, 32, 133, 143, 153, 52, 
    64, 42, 37, 47, 93, 85, 93, 66, 76, 93, 127, 177, 149, 131, 16, 
    61, 65, 75, 108, 133, 143, 148, 149, 145, 149, 109, 141, 141, 49, 48, 
    101, 89, 88, 136, 155, 144, 131, 115, 118, 110, 116, 138, 134, 124, 138, 
    40, 76, 119, 126, 98, 120, 140, 146, 101, 138, 141, 152, 123, 85, 46, 
    81, 104, 117, 109, 117, 106, 136, 42, 37, 136, 115, 80, 49, 12, 30, 
    81, 91, 103, 30, 35, 109, 104, 47, 47, 57, 47, 15, 9, 0, 0, 
    63, 82, 67, 41, 42, 36, 23, 32, 31, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 2, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    32, 2, 0, 0, 46, 2, 4, 0, 0, 0, 21, 87, 0, 17, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 29, 20, 63, 0, 0, 0, 0, 
    0, 15, 70, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 142, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 0, 0, 
    0, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 10, 22, 
    0, 13, 8, 11, 14, 16, 0, 0, 20, 0, 3, 0, 6, 7, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 0, 0, 0, 20, 0, 0, 44, 0, 0, 0, 0, 
    0, 0, 12, 0, 9, 0, 0, 63, 27, 0, 125, 53, 0, 24, 0, 
    0, 0, 12, 15, 21, 0, 20, 0, 0, 99, 5, 95, 342, 71, 49, 
    109, 9, 91, 123, 105, 105, 66, 76, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 255, 0, 
    8, 0, 2, 0, 41, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 76, 50, 0, 0, 0, 
    0, 23, 45, 30, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 72, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 11, 0, 0, 0, 6, 12, 
    23, 0, 0, 0, 64, 67, 0, 0, 4, 87, 19, 29, 5, 3, 10, 
    117, 3, 0, 0, 0, 74, 45, 0, 0, 28, 15, 2, 9, 0, 1, 
    84, 36, 84, 3, 22, 67, 39, 0, 4, 22, 8, 0, 0, 2, 0, 
    40, 69, 40, 36, 17, 17, 16, 20, 25, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 60, 0, 8, 0, 0, 4, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 19, 0, 1, 7, 2, 1, 5, 3, 1, 0, 0, 0, 
    0, 0, 0, 189, 165, 157, 155, 154, 158, 132, 130, 103, 0, 0, 0, 
    0, 0, 11, 139, 99, 63, 118, 80, 50, 52, 36, 24, 0, 0, 0, 
    0, 0, 78, 179, 127, 120, 106, 140, 139, 184, 156, 127, 57, 0, 0, 
    0, 0, 0, 2, 0, 0, 1, 10, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 27, 46, 25, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 78, 24, 10, 17, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 132, 36, 35, 37, 20, 60, 34, 10, 0, 0, 0, 
    0, 0, 0, 56, 61, 39, 54, 0, 0, 30, 4, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 11, 0, 0, 0, 0, 25, 9, 
    1, 33, 17, 4, 0, 3, 3, 4, 34, 29, 33, 35, 39, 55, 52, 
    50, 70, 68, 48, 41, 47, 44, 37, 27, 22, 19, 16, 17, 2, 0, 
    31, 25, 24, 14, 21, 30, 25, 13, 20, 18, 8, 3, 0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 88, 181, 176, 148, 161, 153, 146, 99, 0, 0, 0, 
    0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 251, 183, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 35, 221, 113, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 198, 301, 223, 98, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 77, 63, 12, 0, 67, 241, 350, 329, 204, 56, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    201, 222, 247, 263, 281, 178, 103, 136, 163, 49, 87, 15, 79, 113, 93, 
    0, 0, 0, 0, 0, 0, 0, 72, 116, 144, 163, 187, 204, 216, 225, 
    114, 128, 114, 84, 69, 62, 51, 48, 24, 16, 7, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 
    
    -- channel=50
    25, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 48, 86, 49, 91, 60, 60, 65, 120, 9, 0, 0, 
    20, 0, 0, 57, 0, 13, 5, 62, 1, 0, 2, 52, 58, 0, 0, 
    0, 0, 0, 18, 7, 11, 0, 16, 17, 0, 2, 0, 106, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 132, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 150, 117, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 88, 111, 109, 38, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 29, 16, 11, 0, 137, 102, 111, 50, 0, 
    2, 0, 0, 0, 0, 0, 0, 74, 0, 0, 0, 0, 60, 0, 0, 
    63, 24, 25, 31, 50, 0, 34, 81, 0, 0, 8, 0, 0, 0, 7, 
    6, 0, 0, 0, 0, 0, 10, 38, 0, 23, 19, 37, 38, 15, 50, 
    5, 4, 0, 8, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 
    
    -- channel=51
    0, 0, 36, 35, 37, 57, 72, 77, 74, 91, 72, 76, 51, 0, 0, 
    0, 0, 0, 52, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 88, 75, 88, 43, 84, 121, 132, 129, 94, 119, 6, 4, 
    0, 0, 0, 0, 19, 24, 52, 33, 0, 30, 39, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 8, 
    0, 100, 181, 169, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 24, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 124, 81, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 45, 3, 0, 76, 237, 200, 0, 0, 0, 0, 
    1, 0, 0, 62, 51, 5, 231, 126, 0, 106, 8, 182, 68, 33, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    115, 123, 110, 96, 83, 86, 64, 54, 35, 27, 26, 4, 13, 38, 56, 
    11, 16, 18, 11, 17, 41, 21, 25, 38, 33, 0, 0, 28, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 16, 31, 0, 16, 18, 22, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 152, 0, 11, 31, 79, 48, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 241, 31, 0, 0, 11, 44, 15, 96, 90, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    154, 177, 191, 186, 192, 178, 172, 124, 104, 52, 92, 51, 96, 37, 31, 
    10, 0, 0, 30, 31, 34, 52, 66, 89, 86, 104, 91, 97, 119, 100, 
    32, 0, 0, 0, 2, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 194, 
    
    -- channel=53
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 0, 16, 0, 0, 14, 2, 0, 0, 0, 0, 
    0, 0, 36, 44, 0, 0, 17, 0, 0, 30, 0, 9, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 46, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 219, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 280, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 65, 82, 219, 12, 0, 88, 57, 62, 45, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 9, 16, 1, 9, 7, 0, 0, 
    31, 10, 11, 6, 15, 7, 21, 3, 23, 21, 17, 22, 0, 0, 11, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 52, 26, 32, 44, 49, 54, 57, 0, 0, 0, 
    0, 0, 0, 84, 18, 5, 21, 23, 31, 11, 14, 13, 41, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 90, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 249, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 124, 209, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 132, 285, 159, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 19, 0, 0, 0, 64, 276, 305, 145, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    228, 259, 270, 275, 282, 329, 303, 200, 148, 195, 149, 182, 80, 69, 110, 
    0, 10, 25, 62, 68, 84, 92, 80, 97, 117, 117, 118, 132, 124, 103, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    
    -- channel=55
    87, 117, 123, 77, 76, 90, 91, 74, 84, 82, 86, 81, 68, 77, 75, 
    103, 128, 123, 11, 0, 0, 0, 0, 0, 0, 0, 0, 82, 79, 78, 
    101, 133, 117, 0, 5, 0, 0, 0, 0, 7, 0, 0, 45, 90, 85, 
    112, 131, 116, 0, 0, 3, 2, 0, 2, 8, 0, 29, 0, 92, 94, 
    129, 131, 119, 120, 89, 85, 87, 84, 87, 85, 74, 64, 92, 105, 103, 
    114, 119, 84, 116, 121, 114, 108, 109, 111, 111, 103, 105, 106, 101, 102, 
    99, 151, 130, 7, 15, 92, 104, 108, 104, 106, 97, 102, 101, 99, 95, 
    95, 117, 99, 142, 40, 0, 28, 89, 97, 94, 92, 99, 105, 106, 108, 
    89, 91, 88, 82, 123, 15, 0, 0, 0, 56, 78, 104, 103, 101, 105, 
    81, 76, 84, 99, 98, 0, 0, 2, 15, 24, 0, 0, 5, 57, 95, 
    78, 82, 83, 122, 84, 150, 81, 13, 105, 66, 100, 83, 42, 77, 76, 
    23, 35, 30, 26, 20, 35, 38, 49, 71, 79, 77, 83, 99, 96, 84, 
    44, 60, 63, 51, 44, 45, 45, 44, 54, 43, 46, 40, 40, 47, 36, 
    5, 10, 17, 4, 3, 8, 8, 3, 7, 5, 1, 6, 7, 9, 24, 
    0, 9, 13, 6, 3, 14, 18, 4, 15, 14, 7, 0, 6, 54, 56, 
    
    -- channel=56
    0, 0, 0, 4, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 
    0, 0, 0, 82, 115, 103, 101, 102, 102, 97, 86, 57, 12, 0, 0, 
    0, 0, 0, 41, 86, 86, 98, 90, 66, 76, 66, 56, 35, 0, 0, 
    0, 0, 12, 81, 73, 59, 60, 87, 75, 87, 96, 93, 37, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 25, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 38, 50, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 2, 0, 2, 0, 9, 18, 37, 51, 26, 0, 0, 0, 0, 0, 
    20, 0, 0, 8, 0, 59, 41, 9, 47, 2, 44, 35, 24, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 19, 16, 17, 23, 19, 17, 23, 19, 22, 20, 21, 21, 12, 0, 
    26, 21, 19, 23, 22, 30, 31, 33, 34, 28, 26, 25, 8, 0, 12, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 77, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 108, 106, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 9, 7, 0, 9, 26, 0, 0, 0, 0, 0, 
    11, 0, 0, 3, 0, 0, 29, 0, 14, 0, 28, 6, 26, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 17, 13, 32, 24, 23, 26, 41, 37, 39, 40, 32, 40, 76, 
    0, 23, 28, 31, 33, 27, 27, 31, 37, 36, 36, 43, 48, 114, 107, 
    
    -- channel=59
    150, 178, 156, 151, 150, 169, 168, 156, 159, 161, 170, 163, 163, 196, 195, 
    153, 180, 187, 156, 167, 156, 157, 156, 168, 169, 164, 142, 192, 199, 198, 
    150, 173, 201, 117, 157, 146, 141, 136, 153, 174, 163, 165, 185, 205, 200, 
    152, 168, 193, 132, 137, 142, 140, 154, 148, 161, 152, 168, 146, 195, 193, 
    167, 171, 168, 180, 150, 148, 140, 155, 161, 151, 154, 161, 189, 193, 190, 
    184, 192, 160, 159, 168, 162, 170, 177, 171, 169, 171, 184, 191, 190, 190, 
    191, 152, 129, 135, 141, 172, 190, 198, 195, 194, 190, 193, 193, 197, 194, 
    201, 202, 176, 124, 80, 124, 166, 195, 202, 193, 190, 189, 190, 188, 186, 
    211, 212, 210, 196, 95, 42, 78, 136, 159, 175, 171, 192, 193, 190, 186, 
    214, 212, 211, 236, 75, 6, 18, 27, 46, 70, 89, 150, 157, 170, 184, 
    203, 206, 208, 182, 73, 49, 13, 38, 102, 21, 43, 28, 95, 153, 181, 
    178, 186, 180, 175, 170, 143, 127, 148, 159, 136, 148, 139, 154, 154, 156, 
    66, 68, 67, 60, 59, 51, 50, 67, 75, 68, 68, 70, 74, 78, 62, 
    21, 32, 28, 17, 18, 9, 9, 9, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 2, 0, 2, 0, 0, 0, 0, 43, 68, 
    
    -- channel=60
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 46, 0, 24, 0, 22, 23, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 62, 102, 197, 111, 0, 152, 63, 212, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 
    0, 0, 0, 8, 0, 28, 20, 24, 7, 23, 11, 5, 7, 156, 0, 
    
    -- channel=61
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 95, 87, 50, 69, 57, 68, 65, 59, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 
    17, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 153, 243, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 234, 168, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 12, 56, 262, 211, 56, 9, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 66, 46, 0, 0, 68, 246, 279, 184, 48, 0, 
    58, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 25, 0, 0, 
    172, 101, 110, 124, 132, 140, 54, 38, 91, 28, 45, 31, 0, 57, 71, 
    0, 0, 0, 0, 0, 0, 0, 13, 33, 65, 61, 85, 94, 84, 89, 
    0, 56, 58, 38, 24, 23, 25, 23, 20, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 20, 0, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 45, 
    0, 0, 0, 0, 0, 14, 32, 10, 33, 16, 16, 0, 0, 0, 8, 
    0, 0, 0, 0, 17, 8, 19, 22, 28, 32, 23, 0, 12, 0, 13, 
    0, 0, 0, 0, 0, 45, 3, 32, 19, 42, 31, 0, 46, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 11, 28, 24, 25, 25, 53, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 26, 46, 41, 51, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 39, 26, 45, 35, 35, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 10, 46, 24, 63, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 24, 39, 46, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 
    
    -- channel=65
    0, 0, 0, 0, 1, 0, 0, 0, 18, 22, 0, 0, 0, 26, 0, 
    0, 0, 0, 0, 0, 27, 23, 0, 0, 0, 0, 0, 0, 0, 0, 
    81, 32, 0, 16, 0, 0, 0, 0, 7, 67, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 76, 0, 0, 0, 0, 0, 0, 50, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 46, 
    19, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 69, 
    0, 0, 48, 23, 72, 0, 0, 0, 0, 0, 0, 0, 74, 74, 0, 
    0, 65, 17, 4, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    160, 118, 0, 0, 0, 0, 26, 147, 99, 0, 0, 0, 0, 34, 4, 
    0, 224, 130, 0, 0, 0, 0, 0, 0, 16, 0, 25, 98, 0, 0, 
    2, 0, 126, 99, 0, 0, 0, 0, 57, 70, 133, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 0, 0, 113, 0, 63, 0, 26, 0, 190, 0, 58, 0, 
    0, 0, 0, 0, 0, 56, 0, 83, 0, 6, 0, 211, 0, 38, 0, 
    0, 19, 0, 0, 0, 66, 0, 0, 36, 0, 0, 205, 0, 0, 0, 
    0, 33, 0, 0, 65, 0, 0, 0, 80, 0, 0, 99, 0, 0, 0, 
    0, 89, 0, 0, 131, 0, 0, 103, 0, 0, 0, 115, 0, 0, 0, 
    0, 109, 0, 0, 0, 0, 0, 25, 0, 0, 0, 148, 0, 0, 0, 
    0, 38, 68, 0, 0, 26, 7, 0, 0, 31, 40, 36, 0, 0, 0, 
    0, 31, 22, 0, 0, 12, 41, 4, 0, 0, 4, 64, 0, 0, 0, 
    0, 0, 0, 0, 64, 0, 54, 10, 0, 0, 0, 45, 0, 11, 0, 
    0, 0, 0, 3, 0, 73, 39, 1, 7, 0, 15, 0, 0, 0, 57, 
    0, 37, 0, 0, 5, 0, 95, 0, 0, 0, 10, 0, 0, 25, 0, 
    7, 0, 0, 17, 0, 29, 28, 0, 3, 0, 0, 0, 0, 74, 0, 
    25, 122, 0, 0, 0, 22, 0, 0, 143, 0, 0, 0, 0, 143, 0, 
    0, 119, 142, 0, 0, 0, 0, 0, 71, 8, 6, 0, 0, 74, 18, 
    0, 0, 165, 141, 0, 0, 0, 0, 0, 21, 21, 0, 0, 0, 85, 
    
    -- channel=67
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 48, 37, 
    15, 0, 0, 0, 0, 0, 25, 34, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 12, 0, 0, 38, 0, 0, 0, 22, 18, 5, 0, 0, 0, 
    31, 31, 2, 0, 59, 0, 0, 81, 66, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 58, 24, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 14, 29, 0, 0, 0, 0, 32, 0, 0, 0, 0, 
    0, 3, 16, 0, 0, 0, 0, 60, 59, 0, 0, 27, 0, 0, 0, 
    18, 16, 16, 0, 0, 95, 35, 0, 0, 44, 78, 0, 0, 0, 58, 
    0, 0, 0, 10, 24, 0, 0, 0, 22, 89, 18, 0, 18, 0, 0, 
    0, 9, 6, 0, 0, 49, 0, 0, 16, 0, 28, 0, 0, 51, 75, 
    8, 0, 0, 0, 45, 0, 43, 0, 0, 35, 4, 30, 5, 21, 0, 
    56, 0, 0, 32, 0, 68, 0, 0, 15, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 4, 0, 0, 0, 6, 0, 0, 33, 0, 70, 0, 
    0, 77, 27, 0, 0, 0, 34, 31, 40, 0, 0, 0, 0, 0, 87, 
    0, 0, 68, 0, 0, 0, 0, 62, 1, 0, 0, 40, 75, 128, 0, 
    
    -- channel=68
    0, 0, 0, 0, 117, 0, 15, 0, 36, 0, 40, 0, 168, 0, 0, 
    0, 0, 52, 0, 102, 5, 21, 0, 10, 0, 64, 0, 55, 0, 35, 
    46, 0, 0, 43, 64, 0, 0, 58, 0, 120, 0, 0, 22, 0, 0, 
    59, 0, 8, 0, 0, 0, 51, 112, 0, 0, 0, 0, 34, 0, 177, 
    37, 0, 19, 57, 0, 0, 116, 0, 31, 0, 0, 0, 8, 0, 222, 
    111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 51, 0, 188, 
    0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 40, 0, 112, 
    0, 0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 194, 
    0, 0, 63, 16, 0, 0, 0, 0, 0, 0, 0, 0, 31, 139, 0, 
    0, 70, 11, 0, 35, 48, 0, 0, 0, 0, 0, 0, 70, 0, 0, 
    141, 0, 8, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 
    56, 0, 0, 0, 0, 0, 22, 179, 0, 0, 33, 0, 54, 2, 0, 
    55, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 217, 0, 0, 
    118, 0, 0, 0, 0, 0, 0, 0, 15, 6, 140, 3, 0, 0, 0, 
    
    -- channel=69
    49, 31, 11, 1, 122, 0, 50, 0, 9, 0, 111, 0, 268, 0, 17, 
    0, 16, 24, 3, 112, 0, 0, 0, 47, 0, 106, 0, 241, 0, 70, 
    47, 27, 20, 0, 91, 0, 0, 38, 0, 60, 12, 0, 156, 12, 73, 
    73, 0, 43, 91, 0, 0, 93, 55, 0, 89, 0, 0, 73, 13, 188, 
    63, 0, 172, 16, 0, 9, 162, 0, 8, 0, 58, 0, 37, 14, 252, 
    84, 0, 0, 173, 0, 0, 34, 0, 51, 15, 35, 0, 84, 0, 278, 
    94, 0, 0, 46, 46, 24, 48, 14, 20, 5, 14, 13, 22, 0, 201, 
    63, 0, 0, 16, 82, 0, 0, 16, 49, 38, 23, 0, 151, 0, 142, 
    0, 0, 0, 0, 0, 201, 0, 3, 41, 14, 10, 8, 36, 8, 172, 
    6, 1, 55, 0, 25, 0, 64, 23, 0, 69, 16, 50, 130, 47, 0, 
    110, 0, 82, 0, 0, 104, 0, 28, 53, 18, 34, 38, 68, 0, 2, 
    0, 44, 145, 0, 38, 0, 0, 11, 0, 62, 44, 40, 75, 0, 0, 
    0, 0, 100, 96, 89, 0, 0, 58, 0, 37, 0, 78, 112, 0, 26, 
    126, 0, 0, 29, 123, 54, 12, 88, 0, 0, 29, 64, 137, 0, 0, 
    133, 129, 0, 0, 25, 109, 89, 42, 11, 0, 0, 44, 103, 0, 0, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 34, 0, 39, 0, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 75, 0, 0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 78, 0, 0, 0, 
    0, 25, 11, 0, 0, 0, 38, 29, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 17, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 0, 0, 
    0, 0, 15, 20, 9, 0, 0, 6, 0, 0, 0, 0, 39, 96, 0, 
    0, 23, 0, 0, 15, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    34, 200, 0, 0, 0, 65, 32, 62, 147, 0, 0, 0, 0, 36, 0, 
    0, 23, 165, 18, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 
    0, 0, 10, 140, 63, 0, 0, 0, 0, 80, 154, 43, 0, 0, 0, 
    
    -- channel=71
    37, 0, 29, 40, 67, 0, 25, 0, 1, 0, 48, 0, 84, 0, 4, 
    17, 0, 31, 45, 39, 0, 8, 0, 21, 0, 43, 0, 75, 0, 51, 
    19, 0, 30, 22, 19, 0, 11, 27, 2, 29, 10, 0, 67, 29, 51, 
    45, 14, 32, 39, 0, 0, 27, 0, 0, 22, 5, 0, 47, 29, 111, 
    35, 6, 99, 0, 0, 3, 51, 0, 9, 0, 9, 0, 17, 44, 119, 
    16, 0, 37, 72, 10, 0, 0, 0, 3, 0, 0, 0, 17, 36, 109, 
    27, 11, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 69, 
    23, 7, 18, 26, 2, 0, 0, 0, 0, 0, 0, 0, 19, 17, 46, 
    7, 19, 0, 3, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 57, 
    29, 2, 24, 16, 23, 0, 0, 0, 0, 0, 0, 0, 17, 30, 0, 
    56, 0, 26, 12, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 50, 
    0, 30, 24, 5, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 
    58, 0, 0, 0, 2, 0, 0, 16, 0, 0, 0, 0, 0, 0, 11, 
    44, 26, 0, 0, 0, 10, 10, 6, 0, 0, 0, 0, 13, 28, 0, 
    
    -- channel=72
    23, 0, 24, 0, 0, 6, 15, 0, 25, 0, 6, 2, 50, 25, 0, 
    6, 0, 0, 0, 0, 26, 0, 0, 4, 8, 11, 27, 32, 27, 26, 
    1, 0, 0, 0, 0, 16, 22, 9, 0, 0, 8, 29, 37, 8, 2, 
    0, 30, 14, 17, 0, 45, 15, 0, 26, 0, 69, 42, 21, 9, 33, 
    0, 24, 5, 0, 18, 27, 25, 0, 37, 32, 38, 0, 36, 0, 3, 
    0, 23, 0, 0, 59, 61, 26, 69, 38, 52, 40, 34, 27, 0, 8, 
    0, 33, 0, 3, 63, 108, 98, 121, 76, 82, 77, 98, 23, 3, 0, 
    0, 9, 0, 8, 92, 63, 101, 88, 113, 123, 108, 72, 85, 20, 0, 
    0, 16, 0, 0, 34, 70, 98, 90, 124, 107, 75, 109, 41, 22, 0, 
    0, 0, 0, 5, 32, 24, 82, 102, 80, 112, 77, 92, 79, 19, 0, 
    9, 16, 3, 7, 0, 36, 68, 101, 93, 76, 101, 98, 75, 4, 18, 
    0, 103, 53, 25, 0, 11, 101, 107, 81, 66, 119, 102, 83, 34, 0, 
    23, 13, 42, 45, 38, 11, 61, 87, 52, 85, 103, 96, 90, 0, 0, 
    29, 22, 23, 33, 49, 46, 45, 25, 57, 104, 91, 83, 52, 0, 0, 
    7, 38, 33, 42, 31, 45, 33, 57, 46, 66, 74, 38, 14, 45, 71, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 37, 32, 0, 0, 0, 0, 0, 0, 
    0, 77, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 30, 6, 0, 0, 0, 0, 0, 4, 49, 0, 0, 0, 0, 
    
    -- channel=74
    134, 55, 154, 138, 138, 90, 136, 69, 160, 116, 164, 47, 206, 112, 83, 
    88, 49, 147, 136, 79, 109, 122, 71, 158, 115, 175, 57, 195, 111, 152, 
    109, 88, 112, 81, 44, 106, 162, 157, 112, 109, 190, 52, 187, 133, 170, 
    153, 175, 118, 78, 8, 220, 236, 86, 133, 62, 202, 143, 194, 121, 204, 
    94, 176, 165, 82, 60, 155, 147, 77, 205, 159, 195, 102, 170, 121, 181, 
    37, 162, 145, 83, 209, 76, 0, 94, 114, 118, 123, 72, 160, 143, 169, 
    62, 145, 100, 126, 28, 5, 0, 39, 17, 0, 0, 0, 108, 139, 120, 
    81, 137, 88, 133, 59, 0, 20, 1, 0, 0, 0, 0, 18, 120, 82, 
    85, 114, 78, 111, 32, 0, 0, 0, 0, 1, 0, 0, 0, 23, 100, 
    101, 70, 104, 138, 135, 45, 0, 0, 0, 0, 0, 14, 49, 94, 89, 
    117, 134, 112, 149, 88, 75, 59, 0, 0, 0, 0, 12, 34, 38, 183, 
    56, 156, 179, 145, 158, 82, 46, 11, 0, 0, 8, 0, 34, 68, 171, 
    104, 113, 157, 187, 169, 138, 49, 10, 0, 0, 4, 0, 50, 11, 212, 
    168, 86, 175, 174, 195, 204, 193, 128, 32, 10, 0, 0, 31, 125, 143, 
    172, 153, 116, 180, 161, 174, 231, 225, 98, 29, 9, 8, 68, 166, 216, 
    
    -- channel=75
    29, 0, 11, 0, 0, 0, 15, 0, 58, 26, 47, 0, 96, 0, 0, 
    25, 0, 23, 16, 0, 0, 0, 0, 36, 27, 42, 18, 81, 17, 58, 
    63, 11, 10, 12, 0, 0, 7, 48, 2, 29, 23, 29, 142, 60, 92, 
    2, 16, 53, 1, 0, 56, 80, 0, 17, 0, 65, 75, 151, 88, 130, 
    7, 75, 81, 25, 0, 69, 27, 0, 58, 57, 111, 40, 123, 103, 83, 
    0, 78, 93, 14, 77, 73, 30, 81, 82, 78, 64, 52, 122, 94, 65, 
    1, 58, 75, 116, 89, 76, 60, 92, 81, 84, 72, 93, 86, 93, 43, 
    22, 48, 74, 120, 110, 49, 94, 112, 91, 88, 99, 113, 126, 91, 23, 
    29, 72, 68, 74, 121, 94, 103, 109, 130, 130, 111, 118, 126, 64, 4, 
    91, 54, 42, 72, 71, 115, 98, 137, 133, 152, 105, 123, 86, 37, 11, 
    70, 44, 31, 42, 59, 54, 127, 160, 153, 142, 111, 112, 84, 23, 110, 
    27, 136, 81, 57, 79, 69, 141, 163, 135, 118, 133, 128, 94, 60, 72, 
    124, 134, 143, 108, 72, 95, 135, 145, 86, 118, 150, 105, 102, 0, 90, 
    68, 41, 111, 139, 121, 84, 97, 50, 72, 144, 126, 120, 49, 33, 3, 
    61, 0, 39, 126, 153, 126, 112, 107, 92, 113, 126, 48, 10, 20, 126, 
    
    -- channel=76
    36, 0, 117, 6, 0, 114, 29, 0, 5, 0, 0, 42, 0, 16, 28, 
    0, 0, 0, 14, 0, 63, 0, 62, 0, 28, 0, 101, 0, 146, 4, 
    0, 0, 0, 0, 0, 102, 101, 22, 0, 0, 58, 57, 0, 0, 35, 
    0, 160, 1, 0, 0, 143, 0, 0, 172, 0, 123, 87, 0, 0, 0, 
    0, 137, 0, 0, 96, 0, 0, 153, 6, 82, 17, 0, 0, 0, 0, 
    0, 113, 0, 0, 142, 0, 0, 74, 0, 0, 0, 99, 0, 0, 0, 
    0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 3, 0, 
    0, 30, 22, 0, 20, 0, 17, 16, 0, 19, 16, 0, 0, 0, 0, 
    0, 28, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 50, 0, 0, 0, 24, 0, 0, 0, 0, 0, 21, 17, 
    0, 75, 0, 0, 20, 0, 75, 0, 0, 0, 0, 0, 0, 0, 65, 
    0, 154, 0, 37, 0, 0, 27, 0, 0, 0, 30, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 0, 0, 0, 159, 0, 
    0, 39, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 207, 
    
    -- channel=77
    0, 0, 0, 0, 0, 49, 0, 0, 9, 25, 0, 29, 0, 88, 0, 
    0, 0, 0, 0, 0, 70, 60, 0, 0, 0, 0, 37, 0, 0, 0, 
    0, 3, 0, 0, 0, 1, 0, 0, 53, 0, 134, 13, 0, 0, 0, 
    0, 58, 0, 0, 0, 24, 0, 0, 37, 0, 97, 0, 69, 0, 0, 
    0, 155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 3, 0, 0, 
    0, 198, 31, 0, 24, 0, 0, 0, 0, 0, 44, 0, 0, 43, 0, 
    0, 71, 81, 0, 0, 0, 0, 0, 11, 0, 0, 0, 39, 0, 0, 
    0, 56, 0, 11, 0, 0, 13, 3, 0, 0, 0, 82, 0, 27, 0, 
    0, 0, 0, 36, 43, 0, 5, 0, 0, 0, 19, 0, 55, 0, 0, 
    0, 0, 0, 36, 2, 263, 0, 0, 0, 0, 0, 0, 0, 0, 44, 
    0, 70, 0, 86, 0, 0, 181, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 18, 0, 36, 0, 0, 0, 0, 0, 0, 0, 
    23, 240, 0, 0, 0, 100, 0, 0, 121, 0, 49, 0, 0, 6, 0, 
    0, 80, 270, 25, 0, 0, 0, 0, 0, 20, 0, 0, 0, 1, 0, 
    0, 0, 159, 186, 33, 0, 0, 0, 0, 61, 63, 0, 0, 0, 98, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    9, 26, 19, 21, 0, 51, 24, 44, 41, 57, 25, 76, 0, 29, 47, 
    14, 46, 21, 16, 6, 19, 16, 56, 36, 39, 24, 65, 22, 38, 0, 
    10, 51, 31, 3, 17, 46, 55, 27, 36, 0, 65, 62, 13, 31, 46, 
    14, 46, 14, 2, 54, 64, 73, 34, 54, 38, 25, 90, 29, 32, 0, 
    22, 35, 0, 18, 68, 63, 6, 92, 43, 73, 66, 112, 40, 11, 0, 
    5, 31, 38, 11, 52, 64, 59, 22, 55, 68, 59, 102, 43, 18, 0, 
    28, 13, 43, 45, 49, 27, 54, 10, 45, 28, 27, 26, 56, 40, 16, 
    28, 32, 29, 35, 17, 8, 30, 57, 20, 22, 15, 24, 0, 31, 0, 
    44, 29, 22, 32, 21, 17, 8, 15, 0, 17, 50, 2, 15, 4, 25, 
    17, 10, 28, 42, 7, 40, 5, 0, 23, 0, 24, 12, 0, 12, 71, 
    0, 69, 36, 23, 38, 10, 46, 0, 0, 2, 2, 23, 16, 33, 5, 
    84, 29, 63, 52, 28, 38, 7, 19, 0, 7, 0, 15, 49, 36, 61, 
    11, 94, 100, 98, 57, 62, 7, 0, 37, 11, 0, 1, 12, 55, 66, 
    3, 42, 114, 125, 94, 82, 79, 52, 30, 0, 19, 9, 0, 81, 67, 
    22, 37, 65, 115, 112, 91, 96, 74, 75, 13, 0, 20, 46, 20, 95, 
    
    -- channel=80
    128, 39, 122, 116, 136, 132, 148, 114, 119, 84, 113, 113, 121, 93, 121, 
    61, 86, 117, 121, 127, 132, 145, 152, 159, 86, 103, 121, 124, 127, 122, 
    69, 79, 96, 111, 107, 129, 148, 123, 137, 130, 102, 129, 135, 134, 118, 
    88, 61, 102, 95, 109, 140, 152, 122, 116, 154, 131, 134, 141, 127, 128, 
    65, 82, 93, 98, 116, 94, 111, 106, 117, 133, 101, 107, 98, 107, 123, 
    60, 107, 90, 83, 83, 23, 32, 40, 105, 87, 106, 130, 76, 103, 117, 
    0, 66, 66, 80, 55, 16, 106, 108, 42, 37, 108, 108, 69, 100, 112, 
    135, 34, 85, 60, 15, 73, 78, 56, 42, 59, 97, 80, 59, 83, 97, 
    172, 44, 76, 47, 35, 88, 112, 92, 95, 76, 147, 115, 40, 57, 119, 
    190, 49, 46, 120, 21, 25, 177, 107, 137, 110, 112, 99, 56, 25, 122, 
    170, 81, 66, 197, 52, 82, 154, 134, 163, 81, 74, 114, 73, 14, 123, 
    186, 129, 82, 128, 133, 139, 117, 123, 83, 66, 54, 33, 92, 57, 117, 
    159, 176, 102, 74, 69, 122, 175, 161, 117, 85, 83, 67, 40, 109, 66, 
    155, 144, 159, 100, 140, 150, 146, 195, 144, 131, 139, 110, 117, 94, 126, 
    199, 143, 190, 147, 141, 167, 150, 167, 156, 179, 153, 150, 152, 150, 121, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 5, 0, 0, 96, 14, 0, 1, 35, 5, 0, 1, 
    4, 0, 0, 0, 0, 8, 33, 0, 0, 0, 0, 0, 0, 0, 14, 
    6, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 24, 53, 38, 25, 164, 131, 203, 199, 45, 0, 0, 0, 
    0, 0, 0, 41, 137, 34, 33, 0, 13, 42, 0, 0, 0, 0, 0, 
    0, 28, 66, 26, 28, 207, 115, 172, 95, 31, 77, 0, 0, 42, 0, 
    15, 0, 2, 0, 0, 0, 0, 28, 13, 7, 2, 55, 12, 109, 14, 
    0, 0, 15, 40, 0, 1, 0, 0, 0, 0, 0, 0, 6, 0, 72, 
    10, 17, 12, 30, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 18, 11, 14, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 42, 36, 45, 18, 35, 29, 81, 0, 50, 33, 8, 33, 67, 0, 
    43, 0, 70, 30, 31, 34, 30, 54, 0, 18, 61, 53, 56, 7, 46, 
    0, 13, 51, 52, 44, 35, 3, 86, 47, 0, 48, 27, 46, 54, 44, 
    25, 22, 36, 69, 39, 67, 33, 56, 76, 47, 55, 0, 19, 63, 47, 
    59, 39, 35, 58, 37, 44, 10, 1, 0, 98, 86, 0, 64, 44, 40, 
    285, 2, 20, 28, 32, 104, 0, 2, 0, 69, 0, 0, 49, 44, 56, 
    179, 157, 0, 0, 90, 11, 8, 0, 0, 2, 0, 0, 40, 33, 31, 
    0, 207, 0, 58, 83, 0, 38, 41, 0, 0, 0, 0, 100, 28, 0, 
    17, 180, 0, 19, 0, 124, 0, 57, 48, 31, 0, 0, 152, 106, 0, 
    0, 193, 0, 0, 174, 104, 0, 40, 0, 17, 2, 0, 136, 175, 0, 
    0, 176, 0, 0, 60, 55, 33, 102, 0, 27, 21, 31, 89, 237, 0, 
    53, 63, 42, 0, 0, 41, 52, 0, 0, 1, 0, 43, 117, 151, 4, 
    85, 51, 52, 86, 0, 10, 56, 0, 0, 0, 0, 5, 52, 71, 59, 
    0, 146, 0, 115, 0, 29, 78, 0, 35, 6, 21, 32, 8, 53, 0, 
    37, 58, 28, 71, 42, 10, 49, 44, 41, 56, 63, 63, 33, 0, 88, 
    
    -- channel=83
    30, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 26, 68, 0, 0, 
    0, 0, 3, 8, 0, 0, 0, 0, 20, 38, 13, 0, 0, 0, 13, 
    0, 13, 0, 0, 0, 3, 3, 17, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 16, 20, 40, 7, 
    0, 0, 0, 29, 4, 0, 14, 18, 23, 0, 0, 0, 0, 0, 0, 
    96, 82, 77, 0, 23, 2, 0, 0, 0, 0, 9, 73, 0, 0, 0, 
    0, 0, 0, 0, 46, 0, 12, 0, 19, 9, 2, 21, 23, 10, 0, 
    13, 1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 133, 0, 0, 0, 0, 13, 58, 34, 3, 0, 
    41, 48, 0, 0, 0, 0, 0, 0, 0, 59, 35, 0, 0, 0, 0, 
    0, 4, 0, 43, 123, 190, 76, 113, 3, 0, 11, 0, 0, 0, 0, 
    1, 0, 15, 0, 0, 0, 0, 0, 106, 53, 0, 45, 55, 2, 0, 
    0, 26, 43, 0, 0, 0, 29, 0, 0, 0, 36, 30, 0, 81, 109, 
    0, 26, 0, 3, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 0, 22, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 2, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    49, 0, 0, 0, 0, 1, 0, 0, 7, 0, 0, 117, 0, 17, 0, 
    0, 0, 0, 0, 15, 0, 58, 99, 52, 0, 26, 81, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 67, 34, 0, 0, 0, 
    11, 0, 0, 1, 0, 0, 0, 0, 0, 0, 29, 73, 0, 0, 65, 
    0, 0, 0, 58, 0, 0, 45, 62, 35, 160, 237, 10, 0, 0, 76, 
    6, 0, 0, 188, 21, 18, 91, 0, 120, 43, 0, 6, 0, 0, 117, 
    7, 0, 30, 191, 0, 11, 0, 0, 130, 58, 36, 0, 0, 0, 110, 
    21, 0, 0, 0, 83, 0, 0, 123, 0, 0, 34, 0, 0, 7, 0, 
    0, 0, 0, 13, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 43, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 
    0, 0, 0, 0, 0, 0, 0, 17, 7, 0, 0, 0, 0, 2, 0, 
    
    -- channel=85
    110, 47, 55, 68, 89, 68, 81, 31, 108, 18, 31, 63, 26, 0, 81, 
    68, 105, 52, 61, 64, 79, 99, 75, 136, 45, 0, 7, 29, 70, 23, 
    100, 51, 61, 51, 61, 68, 114, 31, 80, 157, 19, 68, 33, 27, 45, 
    73, 19, 57, 40, 65, 75, 76, 84, 30, 62, 58, 118, 46, 16, 28, 
    0, 38, 65, 55, 62, 72, 71, 85, 87, 8, 46, 182, 20, 25, 32, 
    0, 55, 36, 58, 54, 0, 106, 0, 124, 5, 69, 105, 0, 34, 16, 
    0, 0, 59, 92, 6, 20, 54, 148, 21, 37, 119, 83, 0, 33, 27, 
    79, 0, 76, 0, 0, 58, 65, 11, 20, 51, 190, 98, 0, 18, 79, 
    77, 0, 50, 65, 57, 0, 130, 20, 32, 16, 114, 67, 0, 0, 232, 
    97, 0, 39, 304, 0, 0, 131, 25, 144, 43, 47, 80, 0, 0, 306, 
    99, 0, 46, 216, 16, 0, 18, 0, 90, 62, 12, 4, 0, 0, 229, 
    33, 44, 0, 148, 63, 57, 41, 108, 60, 16, 34, 0, 0, 0, 21, 
    43, 24, 46, 0, 129, 95, 36, 108, 101, 65, 61, 22, 0, 15, 0, 
    81, 0, 83, 28, 79, 49, 0, 120, 49, 70, 67, 47, 79, 38, 40, 
    33, 38, 69, 30, 68, 51, 51, 40, 56, 45, 40, 27, 61, 90, 16, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 
    55, 0, 0, 0, 0, 0, 0, 0, 0, 22, 12, 0, 18, 19, 0, 
    91, 0, 0, 0, 0, 0, 0, 105, 101, 0, 0, 0, 24, 0, 0, 
    0, 88, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 16, 0, 0, 0, 0, 0, 0, 0, 9, 41, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 68, 97, 127, 137, 0, 0, 0, 0, 
    0, 0, 0, 0, 283, 75, 58, 37, 0, 0, 0, 0, 27, 0, 0, 
    0, 7, 0, 0, 0, 0, 74, 0, 157, 14, 31, 77, 0, 64, 0, 
    34, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 16, 85, 
    0, 0, 0, 129, 28, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 14, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    137, 204, 195, 203, 209, 217, 197, 183, 132, 103, 115, 123, 110, 129, 98, 
    163, 184, 190, 215, 223, 219, 227, 234, 191, 103, 111, 118, 146, 147, 116, 
    162, 170, 200, 210, 215, 227, 230, 216, 206, 172, 171, 156, 156, 137, 142, 
    105, 179, 196, 207, 218, 231, 222, 209, 199, 209, 196, 158, 144, 143, 142, 
    131, 168, 198, 212, 214, 210, 165, 174, 177, 192, 171, 131, 121, 135, 141, 
    84, 188, 186, 194, 185, 136, 131, 100, 118, 155, 147, 72, 102, 124, 137, 
    155, 133, 165, 168, 136, 171, 121, 136, 130, 133, 106, 67, 84, 121, 131, 
    159, 153, 155, 132, 151, 144, 181, 158, 120, 127, 105, 62, 71, 135, 109, 
    167, 176, 140, 117, 168, 122, 152, 155, 136, 112, 64, 51, 80, 135, 86, 
    187, 158, 117, 113, 64, 142, 118, 187, 177, 71, 57, 104, 104, 135, 93, 
    187, 156, 131, 71, 124, 59, 90, 166, 69, 71, 57, 74, 121, 131, 91, 
    163, 187, 127, 122, 161, 142, 164, 141, 45, 25, 26, 45, 77, 124, 111, 
    191, 187, 164, 119, 116, 174, 163, 147, 109, 83, 65, 65, 98, 86, 123, 
    178, 153, 161, 160, 124, 159, 191, 179, 142, 141, 139, 162, 146, 155, 136, 
    174, 209, 174, 179, 169, 204, 193, 167, 183, 160, 184, 186, 176, 170, 146, 
    
    -- channel=89
    0, 0, 59, 58, 59, 75, 82, 46, 16, 28, 16, 0, 0, 4, 0, 
    6, 30, 41, 39, 65, 52, 71, 80, 45, 8, 37, 46, 25, 14, 11, 
    0, 23, 31, 66, 54, 70, 68, 99, 64, 0, 0, 0, 54, 59, 9, 
    0, 12, 49, 59, 58, 100, 101, 93, 103, 69, 26, 24, 51, 32, 32, 
    31, 8, 26, 45, 57, 84, 19, 0, 17, 125, 67, 30, 46, 52, 36, 
    70, 0, 0, 28, 70, 0, 0, 71, 43, 27, 37, 33, 42, 42, 41, 
    0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 43, 
    0, 43, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 30, 8, 17, 137, 118, 153, 144, 37, 0, 0, 0, 
    36, 27, 0, 0, 187, 23, 31, 0, 0, 42, 0, 0, 19, 0, 0, 
    29, 58, 0, 0, 0, 145, 137, 188, 161, 41, 58, 47, 0, 69, 0, 
    67, 19, 4, 0, 0, 0, 0, 28, 4, 6, 0, 28, 52, 90, 45, 
    47, 45, 0, 78, 0, 39, 17, 0, 0, 0, 0, 0, 0, 8, 51, 
    62, 82, 44, 33, 50, 0, 42, 32, 0, 0, 0, 0, 0, 0, 26, 
    29, 0, 26, 6, 0, 9, 77, 89, 58, 47, 40, 35, 13, 18, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 25, 20, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 26, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    33, 75, 74, 86, 78, 75, 54, 38, 34, 0, 13, 9, 0, 32, 11, 
    108, 111, 64, 91, 95, 85, 73, 68, 36, 0, 12, 24, 39, 41, 12, 
    120, 107, 93, 99, 104, 100, 91, 73, 65, 19, 37, 25, 45, 32, 34, 
    59, 113, 102, 105, 118, 102, 105, 76, 89, 83, 52, 47, 24, 27, 41, 
    71, 104, 109, 101, 116, 108, 93, 94, 85, 88, 77, 70, 24, 37, 42, 
    0, 94, 124, 121, 104, 87, 138, 135, 68, 71, 87, 8, 20, 20, 37, 
    72, 88, 146, 127, 74, 166, 96, 65, 88, 98, 65, 0, 0, 17, 34, 
    43, 89, 139, 102, 133, 148, 118, 143, 142, 133, 101, 6, 0, 42, 29, 
    64, 88, 138, 94, 182, 93, 161, 126, 124, 120, 49, 0, 0, 73, 49, 
    68, 93, 151, 114, 83, 126, 90, 101, 84, 0, 0, 0, 0, 77, 100, 
    98, 84, 146, 34, 0, 30, 31, 95, 29, 0, 0, 0, 0, 82, 121, 
    64, 98, 85, 59, 20, 0, 21, 26, 0, 0, 0, 0, 0, 48, 81, 
    78, 84, 88, 95, 74, 68, 50, 30, 0, 0, 0, 0, 0, 0, 72, 
    97, 70, 95, 53, 71, 52, 87, 69, 28, 27, 0, 22, 8, 28, 38, 
    60, 99, 73, 71, 56, 99, 85, 73, 64, 41, 59, 70, 65, 58, 28, 
    
    -- channel=92
    0, 133, 0, 44, 1, 16, 0, 14, 0, 0, 14, 22, 30, 65, 0, 
    7, 0, 0, 1, 18, 23, 6, 30, 0, 0, 34, 4, 33, 6, 0, 
    0, 27, 7, 0, 8, 0, 5, 7, 4, 19, 109, 9, 24, 0, 25, 
    0, 0, 0, 11, 0, 0, 0, 0, 6, 0, 0, 0, 0, 52, 16, 
    0, 33, 0, 0, 0, 1, 0, 62, 0, 25, 0, 0, 37, 0, 8, 
    41, 0, 66, 0, 0, 62, 0, 0, 0, 43, 0, 0, 38, 9, 27, 
    224, 0, 0, 0, 0, 34, 0, 4, 144, 67, 0, 0, 32, 46, 20, 
    0, 114, 0, 0, 42, 0, 0, 16, 0, 0, 0, 0, 0, 95, 0, 
    20, 91, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 84, 93, 0, 
    0, 108, 0, 0, 0, 0, 0, 131, 0, 0, 16, 74, 64, 127, 0, 
    0, 24, 0, 0, 116, 0, 0, 19, 0, 0, 0, 0, 78, 81, 0, 
    0, 65, 0, 29, 0, 88, 98, 0, 0, 14, 13, 38, 30, 18, 0, 
    33, 0, 13, 0, 0, 0, 42, 7, 23, 42, 51, 79, 102, 0, 92, 
    18, 0, 0, 0, 0, 51, 51, 0, 26, 35, 33, 110, 52, 99, 0, 
    0, 100, 0, 39, 1, 30, 9, 0, 0, 0, 39, 25, 2, 0, 53, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 28, 0, 0, 0, 
    0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 2, 1, 0, 
    121, 0, 5, 0, 0, 10, 0, 79, 0, 0, 0, 0, 59, 0, 5, 
    36, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 128, 0, 5, 0, 0, 0, 12, 0, 0, 0, 0, 8, 15, 0, 
    0, 19, 0, 0, 75, 8, 0, 63, 71, 59, 63, 0, 23, 63, 0, 
    0, 99, 0, 0, 441, 0, 0, 93, 0, 0, 0, 0, 39, 130, 0, 
    0, 35, 13, 0, 0, 146, 86, 125, 49, 0, 32, 91, 0, 176, 0, 
    0, 0, 69, 0, 0, 0, 0, 0, 0, 24, 7, 14, 77, 8, 178, 
    0, 16, 0, 158, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 56, 
    0, 37, 0, 0, 48, 0, 33, 0, 0, 0, 0, 0, 0, 0, 65, 
    38, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    79, 62, 55, 56, 63, 62, 71, 53, 29, 16, 10, 6, 25, 12, 11, 
    70, 68, 79, 62, 69, 81, 70, 64, 48, 19, 16, 24, 13, 1, 27, 
    27, 77, 70, 79, 72, 83, 72, 85, 87, 45, 37, 13, 0, 24, 15, 
    63, 47, 72, 79, 78, 83, 71, 69, 66, 71, 47, 35, 11, 22, 16, 
    39, 66, 69, 70, 93, 54, 39, 38, 26, 58, 61, 17, 30, 13, 12, 
    109, 22, 76, 68, 65, 100, 0, 12, 25, 22, 4, 14, 14, 21, 17, 
    12, 76, 33, 33, 79, 24, 60, 6, 18, 5, 0, 0, 9, 25, 4, 
    0, 48, 30, 46, 47, 56, 50, 25, 16, 9, 0, 0, 20, 26, 0, 
    30, 15, 31, 23, 5, 59, 18, 24, 27, 3, 0, 5, 32, 24, 0, 
    0, 44, 8, 0, 56, 8, 31, 42, 0, 2, 15, 0, 15, 42, 0, 
    4, 27, 0, 0, 0, 1, 12, 0, 28, 0, 0, 18, 7, 35, 0, 
    24, 0, 27, 60, 16, 36, 9, 0, 0, 8, 0, 0, 31, 9, 39, 
    30, 14, 10, 56, 57, 0, 22, 20, 5, 0, 0, 9, 0, 10, 0, 
    0, 30, 16, 11, 29, 23, 13, 10, 32, 14, 31, 25, 26, 22, 0, 
    34, 2, 25, 25, 23, 7, 17, 23, 14, 25, 27, 30, 24, 15, 41, 
    
    -- channel=96
    350, 341, 344, 342, 346, 329, 314, 311, 287, 266, 263, 221, 75, 132, 230, 
    342, 326, 341, 353, 339, 316, 306, 291, 280, 265, 224, 142, 133, 151, 259, 
    265, 318, 325, 320, 303, 303, 301, 282, 272, 265, 56, 77, 130, 182, 240, 
    297, 304, 301, 299, 304, 312, 306, 276, 252, 193, 88, 98, 238, 252, 272, 
    300, 316, 316, 311, 307, 250, 201, 239, 215, 160, 70, 41, 192, 248, 249, 
    318, 317, 309, 302, 271, 171, 0, 0, 0, 0, 0, 57, 38, 186, 239, 
    314, 321, 307, 274, 112, 48, 88, 117, 120, 0, 0, 137, 12, 72, 169, 
    316, 313, 208, 110, 79, 46, 50, 62, 0, 0, 0, 59, 121, 40, 50, 
    319, 251, 62, 41, 34, 3, 0, 0, 0, 0, 33, 251, 157, 0, 0, 
    284, 26, 47, 18, 75, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    143, 0, 86, 32, 69, 1, 0, 0, 1, 141, 3, 0, 0, 3, 119, 
    173, 34, 17, 62, 18, 0, 0, 0, 118, 39, 55, 0, 11, 85, 95, 
    147, 27, 0, 54, 0, 0, 0, 0, 110, 1, 53, 7, 0, 116, 66, 
    155, 46, 0, 10, 0, 7, 4, 26, 132, 0, 85, 65, 35, 84, 41, 
    136, 74, 43, 19, 5, 10, 24, 44, 49, 2, 37, 73, 39, 32, 19, 
    
    -- channel=97
    8, 35, 40, 48, 43, 39, 35, 25, 46, 136, 45, 0, 22, 19, 2, 
    0, 0, 30, 32, 24, 19, 20, 12, 12, 1, 0, 0, 6, 0, 0, 
    62, 81, 30, 20, 16, 3, 6, 0, 0, 0, 0, 0, 0, 0, 4, 
    18, 6, 6, 0, 0, 0, 0, 0, 0, 0, 82, 59, 41, 57, 15, 
    5, 8, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    11, 1, 5, 7, 0, 0, 0, 0, 74, 103, 0, 0, 31, 0, 0, 
    0, 6, 11, 0, 0, 153, 216, 252, 150, 0, 0, 0, 0, 66, 0, 
    8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 119, 0, 0, 0, 
    14, 0, 0, 11, 76, 63, 0, 0, 0, 0, 38, 33, 0, 0, 0, 
    0, 0, 0, 4, 43, 25, 0, 0, 0, 203, 137, 0, 0, 0, 75, 
    0, 286, 0, 18, 3, 0, 0, 0, 163, 217, 252, 194, 63, 128, 262, 
    41, 0, 0, 0, 0, 0, 0, 0, 60, 0, 0, 147, 5, 110, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 158, 95, 25, 
    0, 36, 171, 155, 311, 436, 453, 465, 232, 42, 52, 15, 172, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 72, 15, 0, 0, 0, 
    
    -- channel=98
    174, 157, 155, 164, 133, 135, 138, 107, 140, 64, 81, 91, 0, 52, 57, 
    157, 119, 114, 133, 123, 113, 114, 99, 101, 90, 107, 1, 0, 86, 62, 
    112, 100, 110, 106, 113, 103, 103, 95, 98, 121, 52, 0, 6, 61, 44, 
    95, 113, 110, 104, 115, 114, 104, 84, 86, 110, 0, 92, 74, 80, 69, 
    103, 118, 118, 111, 131, 107, 79, 94, 73, 0, 0, 25, 7, 58, 78, 
    118, 116, 106, 103, 147, 122, 23, 19, 58, 8, 0, 0, 106, 0, 62, 
    119, 113, 89, 129, 103, 77, 0, 0, 0, 331, 1, 0, 0, 0, 26, 
    122, 110, 143, 37, 0, 66, 0, 0, 0, 62, 0, 0, 0, 84, 0, 
    114, 157, 11, 31, 0, 54, 270, 53, 0, 0, 0, 0, 35, 91, 0, 
    203, 133, 0, 40, 0, 116, 372, 0, 0, 0, 96, 0, 0, 0, 0, 
    343, 66, 0, 0, 0, 88, 290, 0, 0, 0, 81, 249, 0, 0, 0, 
    169, 71, 0, 0, 46, 61, 238, 0, 0, 0, 0, 286, 0, 0, 13, 
    131, 38, 0, 0, 83, 0, 51, 0, 0, 68, 0, 48, 61, 0, 37, 
    78, 63, 0, 26, 107, 73, 71, 57, 0, 89, 0, 0, 15, 0, 22, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 1, 26, 
    
    -- channel=99
    0, 0, 0, 2, 7, 15, 16, 10, 13, 111, 34, 0, 0, 35, 0, 
    48, 12, 8, 21, 21, 16, 15, 13, 9, 0, 43, 13, 17, 0, 0, 
    0, 46, 33, 20, 21, 12, 14, 9, 0, 0, 0, 0, 6, 0, 0, 
    33, 10, 0, 2, 0, 0, 12, 18, 1, 0, 33, 74, 0, 5, 13, 
    0, 0, 0, 0, 0, 0, 0, 51, 189, 185, 63, 0, 4, 9, 0, 
    0, 0, 0, 1, 21, 114, 0, 0, 0, 0, 0, 18, 29, 0, 5, 
    0, 0, 0, 14, 0, 0, 162, 243, 160, 219, 15, 0, 35, 4, 3, 
    0, 0, 10, 0, 86, 0, 7, 207, 197, 0, 0, 0, 0, 30, 28, 
    0, 42, 96, 68, 0, 76, 118, 0, 0, 5, 26, 254, 149, 0, 0, 
    42, 0, 0, 24, 10, 0, 0, 13, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 66, 61, 0, 0, 208, 188, 47, 0, 0, 52, 
    6, 48, 0, 10, 14, 0, 5, 0, 0, 16, 37, 42, 2, 6, 18, 
    25, 0, 1, 75, 71, 62, 47, 75, 0, 0, 10, 0, 0, 11, 1, 
    1, 0, 0, 0, 0, 20, 18, 37, 0, 0, 81, 25, 86, 40, 0, 
    0, 44, 150, 22, 1, 13, 21, 29, 34, 37, 0, 3, 0, 0, 0, 
    
    -- channel=100
    0, 0, 0, 1, 19, 11, 0, 19, 8, 57, 0, 0, 153, 0, 0, 
    0, 0, 33, 10, 9, 9, 0, 1, 0, 0, 0, 60, 12, 0, 0, 
    65, 43, 0, 11, 0, 0, 0, 0, 0, 0, 16, 83, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 214, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 135, 269, 289, 0, 165, 0, 0, 0, 
    0, 0, 0, 0, 0, 175, 86, 65, 0, 0, 0, 39, 64, 51, 0, 
    0, 0, 0, 0, 11, 0, 65, 0, 0, 0, 0, 388, 10, 0, 0, 
    0, 0, 44, 0, 199, 0, 0, 0, 66, 0, 71, 32, 0, 0, 0, 
    0, 0, 220, 0, 101, 0, 0, 0, 0, 257, 115, 0, 0, 0, 74, 
    0, 370, 47, 50, 0, 0, 0, 0, 197, 93, 0, 0, 105, 88, 315, 
    22, 0, 0, 129, 0, 0, 0, 0, 344, 0, 0, 0, 0, 277, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 187, 0, 0, 0, 9, 176, 0, 
    0, 29, 157, 119, 167, 206, 217, 223, 207, 0, 66, 64, 91, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 3, 114, 36, 0, 0, 0, 
    
    -- channel=101
    128, 144, 135, 142, 155, 136, 116, 139, 86, 66, 94, 60, 86, 0, 80, 
    122, 141, 132, 125, 113, 106, 96, 107, 89, 97, 55, 87, 77, 0, 87, 
    93, 98, 93, 96, 80, 87, 86, 89, 86, 59, 46, 67, 43, 34, 103, 
    73, 70, 75, 84, 76, 81, 88, 99, 82, 64, 100, 0, 60, 77, 87, 
    66, 73, 74, 84, 62, 78, 65, 56, 52, 160, 116, 0, 85, 83, 72, 
    72, 77, 84, 83, 34, 0, 0, 8, 0, 0, 108, 245, 0, 139, 67, 
    72, 77, 100, 44, 17, 0, 26, 13, 17, 0, 0, 452, 14, 0, 48, 
    69, 85, 7, 59, 70, 0, 36, 46, 0, 0, 0, 186, 222, 0, 27, 
    79, 23, 27, 0, 60, 0, 0, 0, 0, 0, 115, 212, 0, 0, 0, 
    0, 0, 246, 0, 79, 0, 0, 0, 0, 0, 0, 181, 0, 0, 59, 
    0, 0, 231, 60, 49, 0, 0, 0, 161, 85, 0, 0, 28, 53, 110, 
    0, 0, 30, 99, 0, 0, 0, 0, 309, 16, 37, 0, 0, 172, 37, 
    0, 0, 0, 86, 0, 0, 0, 0, 320, 0, 118, 0, 0, 161, 0, 
    13, 0, 0, 1, 0, 0, 0, 0, 106, 0, 25, 66, 0, 47, 0, 
    21, 38, 3, 73, 4, 15, 18, 25, 29, 0, 48, 81, 17, 14, 0, 
    
    -- channel=102
    0, 0, 18, 27, 27, 22, 29, 17, 0, 5, 0, 3, 11, 82, 0, 
    14, 0, 20, 26, 34, 27, 20, 9, 0, 0, 0, 0, 0, 0, 0, 
    80, 49, 38, 20, 3, 0, 0, 0, 0, 0, 7, 111, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 28, 260, 356, 429, 0, 0, 139, 0, 0, 
    0, 0, 0, 1, 8, 73, 0, 0, 0, 0, 0, 0, 0, 93, 54, 
    0, 0, 13, 0, 0, 26, 0, 0, 0, 0, 0, 102, 31, 0, 0, 
    0, 0, 0, 65, 34, 0, 41, 4, 41, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 52, 101, 0, 0, 155, 426, 4, 0, 0, 0, 
    53, 259, 42, 0, 8, 0, 0, 0, 0, 37, 0, 264, 55, 38, 103, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 36, 0, 18, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 69, 9, 
    0, 41, 109, 178, 161, 235, 270, 266, 258, 0, 0, 0, 0, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 115, 31, 0, 0, 0, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 138, 77, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 43, 17, 14, 0, 85, 218, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 33, 83, 61, 92, 113, 132, 70, 0, 31, 
    0, 0, 0, 0, 57, 1, 0, 80, 78, 84, 161, 48, 0, 17, 50, 
    0, 0, 116, 30, 32, 0, 0, 107, 102, 75, 0, 120, 90, 95, 80, 
    0, 0, 157, 72, 11, 34, 4, 113, 182, 48, 23, 0, 121, 99, 43, 
    0, 29, 132, 66, 19, 61, 34, 109, 186, 49, 40, 0, 97, 122, 0, 
    0, 33, 109, 76, 58, 129, 96, 111, 181, 24, 94, 14, 43, 63, 0, 
    0, 0, 56, 32, 22, 19, 18, 20, 60, 43, 62, 37, 13, 12, 0, 
    0, 13, 57, 86, 51, 58, 50, 44, 27, 0, 45, 16, 9, 6, 0, 
    
    -- channel=104
    489, 470, 472, 462, 437, 403, 390, 362, 332, 277, 266, 201, 105, 81, 204, 
    424, 393, 393, 379, 351, 324, 322, 302, 285, 273, 233, 152, 56, 149, 235, 
    308, 297, 296, 302, 293, 288, 292, 288, 280, 267, 150, 18, 109, 213, 243, 
    260, 276, 283, 281, 291, 299, 299, 297, 279, 234, 77, 48, 210, 253, 243, 
    270, 288, 289, 287, 287, 269, 250, 246, 227, 167, 16, 69, 184, 228, 233, 
    288, 287, 286, 282, 262, 180, 87, 47, 36, 0, 16, 30, 8, 154, 210, 
    290, 288, 280, 246, 164, 93, 25, 0, 20, 0, 26, 0, 16, 34, 118, 
    284, 281, 195, 139, 50, 36, 31, 26, 37, 67, 0, 0, 10, 24, 65, 
    282, 230, 97, 0, 2, 0, 0, 46, 2, 0, 39, 0, 74, 24, 50, 
    246, 134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 7, 
    165, 22, 0, 2, 0, 0, 0, 0, 6, 0, 12, 0, 0, 0, 0, 
    174, 0, 0, 0, 0, 6, 0, 0, 0, 7, 0, 6, 0, 0, 0, 
    113, 3, 0, 0, 0, 0, 18, 0, 0, 0, 1, 5, 11, 0, 42, 
    123, 39, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 24, 0, 22, 
    105, 44, 0, 0, 0, 0, 0, 1, 5, 8, 0, 0, 12, 12, 11, 
    
    -- channel=105
    340, 406, 456, 480, 469, 431, 415, 380, 350, 295, 251, 204, 103, 71, 142, 
    441, 379, 397, 417, 389, 342, 329, 305, 270, 236, 177, 102, 0, 4, 163, 
    353, 353, 331, 312, 285, 250, 251, 233, 223, 206, 109, 0, 0, 66, 170, 
    240, 238, 232, 229, 232, 236, 205, 184, 174, 169, 49, 0, 101, 201, 216, 
    208, 238, 241, 241, 240, 218, 169, 145, 0, 0, 0, 0, 104, 190, 195, 
    232, 236, 234, 238, 216, 21, 0, 0, 13, 5, 0, 0, 62, 25, 165, 
    238, 234, 244, 213, 109, 81, 37, 39, 55, 0, 0, 0, 0, 66, 91, 
    237, 238, 144, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    240, 179, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    211, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    196, 100, 0, 0, 0, 0, 0, 0, 0, 0, 19, 60, 0, 0, 11, 
    196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 9, 
    52, 0, 0, 0, 67, 148, 166, 166, 53, 0, 0, 0, 39, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 32, 0, 40, 0, 101, 24, 0, 43, 0, 
    0, 0, 0, 0, 0, 0, 13, 26, 43, 37, 0, 61, 0, 0, 41, 
    0, 0, 0, 0, 51, 21, 0, 82, 0, 0, 48, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 48, 39, 0, 25, 0, 28, 106, 0, 19, 38, 0, 21, 0, 
    0, 0, 148, 9, 14, 74, 0, 0, 90, 29, 31, 0, 30, 50, 0, 
    0, 0, 119, 0, 35, 49, 46, 0, 45, 15, 22, 0, 107, 0, 4, 
    0, 0, 63, 0, 25, 18, 10, 0, 22, 32, 35, 22, 71, 12, 19, 
    0, 0, 34, 64, 37, 46, 45, 36, 39, 28, 21, 0, 40, 36, 35, 
    
    -- channel=107
    90, 91, 111, 99, 90, 73, 75, 54, 46, 48, 24, 0, 6, 0, 0, 
    85, 82, 77, 61, 53, 40, 44, 30, 23, 15, 3, 6, 0, 0, 2, 
    67, 49, 35, 28, 21, 20, 22, 20, 18, 8, 54, 0, 0, 23, 19, 
    10, 9, 13, 12, 16, 23, 29, 33, 34, 27, 16, 0, 12, 15, 7, 
    11, 12, 15, 17, 21, 43, 60, 47, 31, 73, 0, 0, 32, 13, 3, 
    12, 14, 18, 19, 11, 20, 112, 146, 176, 123, 119, 25, 0, 38, 0, 
    15, 20, 23, 3, 54, 69, 81, 5, 0, 0, 226, 104, 0, 13, 0, 
    19, 18, 0, 43, 32, 5, 1, 0, 6, 166, 212, 206, 0, 0, 17, 
    20, 0, 27, 12, 32, 0, 0, 221, 240, 219, 250, 11, 0, 5, 129, 
    0, 97, 52, 0, 0, 0, 0, 210, 184, 236, 148, 99, 131, 145, 159, 
    0, 146, 63, 6, 0, 0, 23, 180, 248, 0, 32, 107, 164, 148, 29, 
    0, 0, 85, 0, 0, 36, 70, 185, 138, 0, 0, 0, 98, 76, 0, 
    0, 0, 76, 0, 0, 57, 153, 167, 99, 0, 5, 0, 86, 0, 0, 
    0, 0, 61, 0, 46, 86, 98, 99, 17, 7, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    
    -- channel=108
    99, 42, 52, 25, 16, 23, 36, 15, 45, 0, 8, 37, 15, 0, 38, 
    31, 52, 12, 31, 32, 28, 44, 33, 42, 41, 59, 51, 0, 92, 51, 
    11, 0, 19, 27, 41, 50, 51, 56, 60, 50, 168, 0, 15, 115, 45, 
    42, 53, 50, 48, 62, 58, 75, 83, 80, 85, 0, 0, 41, 18, 25, 
    60, 54, 48, 48, 58, 100, 53, 23, 78, 171, 24, 45, 48, 41, 47, 
    58, 53, 51, 48, 56, 117, 233, 83, 0, 0, 105, 0, 0, 37, 38, 
    55, 48, 52, 42, 188, 0, 0, 0, 0, 47, 122, 0, 3, 0, 0, 
    44, 43, 70, 118, 0, 38, 0, 110, 306, 390, 0, 0, 0, 0, 222, 
    48, 49, 38, 0, 0, 0, 0, 253, 0, 0, 0, 0, 76, 252, 55, 
    24, 409, 0, 17, 0, 58, 105, 0, 0, 0, 0, 0, 124, 0, 0, 
    174, 0, 0, 0, 0, 125, 211, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 1, 52, 0, 68, 161, 115, 0, 0, 46, 0, 43, 0, 0, 0, 
    62, 23, 34, 0, 181, 125, 142, 0, 0, 53, 15, 33, 51, 0, 33, 
    70, 46, 0, 0, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 44, 
    52, 0, 5, 104, 47, 60, 48, 32, 25, 50, 0, 0, 42, 43, 56, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 3, 0, 0, 94, 2, 9, 0, 52, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 4, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 159, 0, 0, 138, 0, 0, 
    0, 0, 0, 0, 0, 10, 94, 48, 116, 78, 224, 0, 0, 173, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 115, 9, 48, 81, 91, 0, 2, 0, 0, 53, 0, 15, 
    0, 0, 0, 18, 0, 52, 16, 98, 0, 20, 255, 0, 0, 0, 0, 
    0, 279, 0, 0, 0, 0, 0, 26, 0, 0, 37, 506, 0, 0, 0, 
    46, 0, 152, 0, 0, 73, 54, 0, 0, 0, 0, 83, 102, 0, 0, 
    25, 33, 158, 0, 0, 0, 0, 0, 0, 62, 0, 0, 287, 0, 26, 
    0, 86, 138, 4, 149, 258, 255, 240, 156, 52, 61, 0, 134, 13, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 132, 12, 0, 0, 0, 2, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    155, 154, 165, 172, 154, 132, 127, 116, 87, 58, 77, 49, 0, 38, 34, 
    137, 132, 102, 91, 79, 69, 67, 69, 62, 61, 39, 4, 7, 19, 30, 
    61, 50, 62, 45, 55, 49, 44, 62, 56, 60, 0, 0, 21, 34, 29, 
    45, 45, 42, 43, 51, 44, 44, 51, 64, 37, 0, 36, 50, 36, 45, 
    31, 37, 39, 38, 42, 42, 35, 23, 26, 0, 0, 0, 1, 40, 40, 
    36, 33, 36, 37, 21, 22, 14, 0, 0, 0, 0, 0, 30, 0, 29, 
    37, 34, 23, 27, 5, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 
    37, 25, 26, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    24, 7, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 18, 24, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 18, 12, 15, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 27, 45, 
    0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 38, 46, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 61, 48, 
    0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 54, 
    0, 0, 5, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 44, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 117, 
    0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 95, 
    0, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 96, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 67, 
    9, 0, 0, 45, 78, 52, 0, 0, 0, 0, 0, 0, 0, 74, 61, 
    20, 65, 89, 88, 74, 46, 27, 82, 71, 44, 3, 17, 61, 91, 99, 
    
    -- channel=113
    0, 0, 0, 10, 16, 0, 1, 1, 0, 0, 5, 5, 0, 0, 0, 
    0, 0, 0, 13, 0, 48, 3, 8, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 42, 20, 15, 0, 27, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 56, 7, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 35, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 
    10, 3, 0, 0, 9, 44, 0, 0, 0, 0, 0, 0, 6, 20, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 87, 
    0, 0, 51, 0, 72, 0, 17, 0, 0, 0, 0, 0, 0, 23, 0, 
    0, 8, 158, 155, 108, 136, 52, 15, 0, 0, 3, 0, 0, 0, 0, 
    263, 236, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 3, 0, 
    72, 72, 30, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 58, 120, 81, 0, 0, 6, 14, 77, 84, 0, 9, 12, 34, 
    72, 111, 54, 3, 0, 2, 0, 17, 5, 0, 40, 65, 35, 15, 16, 
    
    -- channel=114
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 34, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 0, 0, 0, 7, 43, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 3, 24, 30, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 0, 0, 0, 6, 25, 0, 8, 0, 1, 
    0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 17, 40, 14, 0, 
    0, 0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 48, 0, 17, 0, 
    0, 0, 0, 0, 0, 40, 0, 14, 0, 0, 0, 0, 0, 8, 0, 
    1, 11, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 2, 0, 
    0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 2, 6, 0, 0, 0, 67, 0, 
    0, 0, 0, 0, 0, 0, 30, 0, 7, 55, 0, 0, 0, 39, 18, 
    0, 2, 0, 0, 41, 0, 22, 0, 21, 48, 2, 0, 0, 26, 65, 
    0, 7, 16, 13, 83, 30, 0, 4, 32, 14, 45, 22, 0, 42, 36, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 21, 
    0, 0, 0, 44, 0, 0, 0, 0, 4, 15, 35, 17, 0, 0, 0, 
    0, 0, 0, 0, 24, 0, 14, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 75, 51, 22, 50, 37, 0, 7, 1, 0, 2, 5, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 29, 27, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 8, 10, 15, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 10, 0, 0, 0, 94, 4, 0, 0, 0, 0, 0, 0, 40, 19, 
    0, 59, 76, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 22, 0, 0, 0, 0, 0, 0, 22, 14, 
    0, 0, 123, 206, 0, 33, 0, 0, 0, 0, 0, 27, 0, 0, 0, 
    0, 128, 0, 0, 65, 43, 0, 34, 100, 52, 0, 0, 0, 0, 0, 
    28, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    39, 0, 0, 0, 55, 1, 19, 0, 0, 0, 5, 2, 0, 0, 0, 
    0, 8, 48, 10, 0, 0, 0, 0, 4, 3, 9, 0, 3, 0, 0, 
    
    -- channel=116
    0, 0, 0, 25, 0, 0, 2, 0, 1, 4, 12, 20, 6, 0, 0, 
    0, 0, 0, 0, 16, 16, 18, 9, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 58, 1, 0, 0, 8, 0, 0, 0, 0, 0, 0, 28, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 34, 38, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 93, 16, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 30, 39, 0, 0, 0, 8, 0, 0, 7, 57, 
    0, 0, 0, 6, 37, 0, 0, 0, 0, 7, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 6, 0, 13, 96, 
    0, 0, 126, 124, 61, 128, 0, 9, 0, 0, 0, 20, 3, 13, 0, 
    0, 28, 185, 2, 26, 90, 7, 24, 0, 4, 25, 0, 0, 0, 18, 
    246, 106, 0, 75, 23, 0, 0, 25, 0, 0, 0, 0, 14, 0, 0, 
    0, 40, 0, 0, 18, 8, 52, 0, 0, 0, 0, 13, 4, 0, 0, 
    0, 0, 50, 84, 0, 0, 0, 3, 5, 14, 34, 0, 27, 4, 0, 
    73, 65, 0, 0, 0, 0, 0, 2, 0, 0, 0, 14, 7, 0, 6, 
    
    -- channel=117
    5, 13, 0, 0, 11, 32, 30, 18, 27, 24, 21, 26, 25, 12, 31, 
    6, 27, 2, 0, 44, 0, 62, 43, 17, 21, 27, 32, 25, 26, 38, 
    3, 12, 28, 12, 42, 45, 36, 42, 9, 36, 29, 38, 23, 31, 38, 
    7, 8, 103, 0, 38, 59, 52, 37, 44, 0, 19, 49, 28, 36, 40, 
    0, 0, 163, 86, 29, 6, 66, 87, 68, 56, 21, 47, 20, 46, 47, 
    0, 0, 154, 47, 69, 0, 40, 97, 70, 71, 85, 14, 0, 43, 50, 
    0, 0, 22, 229, 0, 0, 90, 55, 40, 82, 87, 9, 55, 14, 47, 
    0, 0, 29, 0, 201, 0, 92, 29, 30, 93, 87, 66, 49, 5, 36, 
    0, 0, 24, 71, 116, 182, 59, 70, 18, 70, 86, 88, 12, 29, 67, 
    0, 0, 0, 213, 0, 150, 0, 114, 29, 43, 70, 99, 37, 90, 54, 
    0, 32, 138, 14, 16, 38, 46, 17, 41, 42, 67, 94, 51, 72, 58, 
    0, 0, 76, 61, 121, 19, 8, 104, 0, 7, 43, 92, 62, 0, 134, 
    1, 0, 0, 10, 71, 87, 0, 89, 14, 0, 68, 59, 121, 32, 29, 
    3, 8, 26, 37, 14, 45, 30, 39, 42, 0, 0, 68, 74, 51, 12, 
    31, 33, 39, 52, 0, 22, 69, 68, 52, 52, 13, 29, 76, 41, 49, 
    
    -- channel=118
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 21, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 120, 32, 0, 0, 0, 0, 0, 0, 11, 10, 
    0, 0, 0, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 86, 91, 30, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 35, 64, 0, 80, 0, 0, 0, 0, 0, 0, 0, 
    173, 64, 65, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    25, 16, 0, 0, 49, 0, 20, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 17, 32, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 
    35, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    
    -- channel=119
    26, 24, 11, 12, 0, 0, 0, 11, 19, 13, 12, 14, 12, 7, 13, 
    26, 31, 16, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 3, 4, 
    20, 23, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 19, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 27, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 20, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 18, 27, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 14, 21, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 15, 47, 6, 23, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 45, 8, 74, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 69, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 27, 20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    3, 5, 15, 15, 35, 50, 42, 24, 13, 18, 16, 11, 15, 21, 20, 
    3, 8, 25, 4, 56, 65, 69, 78, 40, 30, 42, 43, 45, 51, 48, 
    5, 9, 16, 30, 54, 81, 99, 102, 81, 62, 53, 64, 49, 47, 49, 
    12, 21, 35, 45, 59, 82, 91, 114, 132, 85, 70, 76, 58, 53, 70, 
    31, 37, 67, 26, 55, 66, 83, 96, 118, 126, 114, 96, 99, 99, 105, 
    42, 31, 27, 7, 60, 83, 65, 71, 98, 107, 123, 104, 112, 116, 98, 
    19, 20, 18, 48, 42, 50, 69, 90, 92, 83, 104, 101, 106, 92, 59, 
    30, 37, 49, 16, 90, 66, 88, 95, 86, 72, 89, 104, 93, 83, 70, 
    44, 53, 48, 45, 81, 103, 82, 94, 75, 61, 79, 91, 85, 82, 108, 
    46, 58, 29, 32, 55, 79, 83, 83, 77, 63, 77, 83, 86, 92, 104, 
    27, 28, 7, 24, 45, 58, 75, 50, 81, 77, 87, 83, 90, 112, 118, 
    2, 0, 0, 31, 40, 47, 63, 74, 57, 62, 66, 89, 106, 123, 120, 
    0, 21, 25, 41, 36, 62, 85, 60, 64, 58, 66, 66, 116, 139, 115, 
    31, 50, 68, 82, 84, 90, 86, 86, 80, 73, 46, 54, 93, 126, 131, 
    66, 82, 95, 107, 117, 117, 104, 117, 128, 113, 105, 101, 110, 134, 133, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 22, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 20, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 5, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 
    0, 0, 0, 0, 2, 41, 12, 24, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 38, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 41, 30, 
    0, 0, 0, 31, 38, 0, 0, 0, 2, 23, 20, 0, 0, 60, 68, 
    0, 45, 42, 30, 44, 21, 0, 32, 48, 27, 33, 54, 49, 74, 81, 
    
    -- channel=122
    55, 50, 39, 38, 68, 105, 79, 56, 51, 62, 49, 46, 47, 36, 35, 
    56, 62, 66, 4, 120, 132, 140, 122, 56, 54, 49, 43, 36, 23, 19, 
    59, 66, 56, 52, 144, 172, 188, 177, 97, 55, 47, 43, 13, 13, 13, 
    63, 65, 55, 66, 182, 196, 181, 178, 150, 129, 95, 68, 17, 16, 15, 
    44, 43, 117, 12, 163, 178, 176, 162, 193, 185, 174, 145, 39, 0, 0, 
    22, 24, 116, 0, 146, 174, 173, 189, 194, 180, 199, 190, 64, 0, 0, 
    23, 17, 40, 3, 89, 115, 178, 192, 192, 170, 201, 175, 116, 32, 5, 
    39, 23, 41, 2, 50, 51, 127, 155, 193, 189, 195, 202, 191, 78, 19, 
    29, 10, 30, 0, 107, 77, 104, 115, 195, 200, 201, 223, 194, 85, 0, 
    0, 0, 0, 82, 93, 163, 83, 124, 205, 199, 198, 216, 188, 66, 0, 
    0, 10, 0, 144, 144, 161, 149, 108, 182, 182, 168, 202, 153, 54, 0, 
    9, 17, 4, 76, 105, 178, 168, 67, 178, 184, 164, 179, 90, 18, 0, 
    40, 41, 32, 30, 46, 53, 107, 130, 155, 163, 186, 173, 113, 13, 19, 
    39, 36, 45, 21, 0, 40, 34, 109, 93, 118, 161, 168, 148, 4, 0, 
    23, 5, 5, 0, 0, 17, 28, 0, 0, 39, 50, 60, 39, 0, 0, 
    
    -- channel=123
    35, 30, 32, 44, 44, 37, 34, 19, 12, 9, 0, 0, 0, 0, 0, 
    32, 30, 38, 0, 46, 40, 34, 19, 2, 0, 0, 0, 0, 0, 0, 
    26, 26, 32, 0, 14, 11, 21, 17, 4, 38, 39, 45, 34, 33, 18, 
    17, 18, 0, 0, 0, 5, 8, 29, 33, 43, 51, 47, 26, 21, 9, 
    35, 67, 128, 0, 0, 24, 46, 34, 34, 30, 40, 42, 41, 36, 35, 
    123, 136, 127, 0, 0, 36, 55, 38, 37, 31, 34, 29, 51, 61, 57, 
    123, 118, 103, 28, 35, 41, 51, 32, 45, 41, 35, 20, 52, 59, 45, 
    100, 109, 138, 73, 41, 9, 50, 37, 60, 57, 32, 25, 38, 21, 19, 
    117, 124, 139, 125, 148, 124, 81, 47, 53, 56, 39, 29, 24, 36, 35, 
    188, 237, 252, 214, 144, 150, 76, 51, 49, 54, 53, 36, 21, 11, 0, 
    261, 276, 128, 118, 88, 71, 58, 33, 53, 56, 53, 29, 15, 17, 4, 
    225, 156, 87, 75, 30, 1, 19, 14, 22, 25, 47, 49, 17, 30, 18, 
    79, 69, 56, 61, 44, 21, 39, 21, 15, 26, 79, 60, 33, 26, 30, 
    36, 50, 64, 45, 10, 27, 2, 36, 9, 32, 52, 37, 43, 11, 22, 
    46, 24, 4, 0, 0, 34, 31, 8, 0, 1, 5, 19, 5, 0, 5, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 13, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 14, 44, 58, 63, 39, 
    0, 0, 0, 0, 0, 0, 0, 4, 35, 51, 15, 19, 0, 0, 0, 
    0, 0, 0, 9, 0, 27, 37, 23, 2, 0, 0, 0, 0, 0, 0, 
    77, 96, 58, 0, 26, 52, 41, 0, 12, 2, 0, 0, 5, 8, 27, 
    0, 0, 0, 0, 23, 87, 0, 0, 25, 0, 17, 0, 12, 0, 0, 
    0, 0, 0, 0, 51, 0, 0, 0, 27, 0, 0, 19, 8, 0, 0, 
    0, 0, 0, 0, 0, 98, 12, 20, 25, 0, 0, 18, 11, 0, 5, 
    0, 0, 23, 19, 14, 38, 25, 0, 0, 0, 0, 0, 15, 4, 0, 
    95, 42, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 1, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 33, 9, 
    0, 0, 0, 0, 0, 0, 59, 0, 0, 0, 27, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 13, 30, 21, 0, 0, 30, 6, 
    0, 3, 0, 0, 0, 15, 0, 1, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 28, 25, 10, 0, 0, 21, 4, 0, 0, 18, 16, 
    
    -- channel=125
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 2, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 12, 0, 14, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 5, 0, 75, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 20, 6, 0, 0, 
    0, 0, 7, 0, 67, 70, 0, 0, 1, 0, 0, 0, 0, 25, 0, 
    0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 
    0, 0, 0, 0, 0, 0, 35, 0, 5, 0, 0, 0, 21, 0, 0, 
    0, 0, 0, 0, 72, 40, 38, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 150, 36, 84, 0, 35, 3, 0, 0, 0, 0, 0, 0, 
    34, 79, 0, 0, 0, 23, 42, 0, 76, 24, 0, 0, 0, 47, 0, 
    43, 11, 13, 0, 0, 0, 33, 0, 0, 1, 0, 0, 0, 0, 55, 
    4, 0, 0, 13, 28, 33, 0, 37, 0, 12, 117, 0, 0, 0, 13, 
    0, 23, 31, 0, 0, 37, 0, 0, 0, 3, 22, 47, 5, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 0, 24, 52, 19, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 54, 94, 91, 66, 19, 4, 12, 17, 15, 0, 0, 
    0, 0, 0, 30, 90, 125, 136, 160, 100, 14, 15, 12, 5, 0, 0, 
    3, 0, 0, 46, 126, 132, 150, 158, 126, 96, 60, 33, 3, 1, 16, 
    14, 8, 0, 52, 123, 120, 112, 134, 166, 158, 149, 111, 33, 30, 31, 
    0, 0, 0, 44, 87, 106, 108, 142, 145, 162, 161, 149, 84, 29, 15, 
    0, 0, 0, 0, 58, 94, 124, 147, 121, 126, 150, 166, 88, 25, 0, 
    0, 0, 0, 45, 0, 67, 86, 140, 127, 119, 149, 154, 114, 51, 33, 
    0, 0, 2, 14, 26, 0, 68, 109, 128, 124, 144, 154, 137, 84, 8, 
    0, 0, 0, 0, 36, 19, 65, 122, 134, 131, 139, 154, 139, 61, 26, 
    0, 0, 0, 50, 97, 99, 116, 125, 133, 133, 118, 153, 136, 55, 19, 
    0, 0, 32, 6, 40, 140, 115, 16, 109, 140, 113, 114, 105, 60, 26, 
    12, 0, 0, 18, 40, 41, 57, 90, 105, 134, 81, 115, 101, 55, 55, 
    17, 19, 20, 20, 38, 45, 51, 85, 104, 90, 97, 122, 109, 67, 45, 
    7, 16, 45, 43, 43, 34, 54, 59, 56, 63, 75, 79, 73, 52, 33, 
    
    -- channel=128
    48, 0, 36, 36, 10, 19, 25, 2, 49, 47, 0, 11, 38, 23, 41, 
    47, 0, 28, 41, 1, 0, 0, 0, 27, 110, 0, 0, 8, 19, 34, 
    51, 20, 0, 26, 0, 47, 37, 16, 46, 28, 0, 0, 0, 0, 0, 
    53, 12, 0, 0, 0, 45, 26, 43, 39, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 0, 10, 28, 54, 26, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 51, 60, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 18, 17, 24, 35, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 108, 0, 0, 0, 34, 5, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 88, 0, 0, 0, 0, 72, 0, 25, 20, 36, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 18, 11, 8, 37, 50, 18, 10, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 30, 26, 43, 4, 12, 49, 18, 
    0, 0, 0, 0, 0, 44, 0, 4, 13, 72, 0, 17, 19, 29, 48, 
    0, 0, 0, 0, 63, 101, 8, 15, 44, 47, 6, 27, 24, 45, 35, 
    0, 0, 0, 0, 39, 26, 18, 39, 51, 44, 15, 31, 52, 16, 24, 
    0, 0, 0, 0, 0, 10, 40, 41, 62, 18, 26, 28, 43, 6, 25, 
    
    -- channel=129
    0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 64, 104, 97, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 197, 42, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 173, 141, 32, 
    0, 0, 0, 0, 18, 66, 0, 0, 0, 0, 48, 0, 0, 0, 91, 
    0, 0, 0, 0, 0, 0, 24, 15, 0, 43, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 72, 0, 28, 44, 1, 0, 0, 69, 17, 0, 
    0, 0, 4, 0, 0, 0, 35, 39, 39, 17, 0, 0, 2, 0, 0, 
    39, 0, 25, 0, 0, 0, 54, 31, 29, 0, 1, 0, 0, 0, 20, 
    
    -- channel=130
    0, 315, 33, 0, 0, 30, 0, 19, 0, 0, 238, 0, 0, 6, 0, 
    0, 199, 63, 101, 0, 0, 24, 27, 0, 0, 230, 0, 0, 0, 0, 
    1, 64, 154, 84, 42, 0, 0, 43, 0, 50, 21, 6, 0, 0, 0, 
    0, 111, 49, 0, 99, 0, 0, 0, 0, 173, 0, 81, 0, 0, 37, 
    0, 55, 0, 0, 102, 0, 0, 0, 9, 126, 31, 43, 0, 0, 51, 
    0, 8, 0, 0, 42, 0, 0, 0, 0, 82, 40, 61, 0, 0, 0, 
    0, 1, 0, 0, 0, 20, 0, 81, 0, 14, 46, 61, 0, 0, 0, 
    0, 18, 0, 109, 0, 0, 0, 0, 21, 57, 0, 128, 89, 0, 16, 
    0, 19, 0, 87, 0, 0, 0, 0, 137, 21, 0, 0, 139, 0, 128, 
    0, 5, 0, 0, 3, 0, 0, 0, 0, 19, 0, 0, 49, 0, 70, 
    0, 0, 28, 0, 0, 0, 41, 27, 0, 0, 39, 13, 0, 0, 0, 
    0, 0, 80, 0, 0, 0, 9, 0, 0, 0, 74, 0, 0, 0, 0, 
    0, 0, 81, 0, 0, 140, 1, 0, 0, 0, 42, 8, 0, 12, 0, 
    0, 0, 101, 0, 0, 39, 0, 0, 0, 30, 14, 7, 0, 70, 0, 
    0, 0, 90, 24, 0, 0, 0, 10, 0, 71, 20, 0, 0, 20, 18, 
    
    -- channel=131
    0, 19, 0, 0, 14, 0, 0, 0, 0, 34, 46, 0, 0, 0, 0, 
    0, 5, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 16, 6, 0, 
    0, 0, 61, 31, 0, 0, 64, 45, 4, 7, 0, 40, 0, 0, 0, 
    90, 126, 0, 0, 0, 0, 0, 9, 42, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 38, 15, 0, 0, 1, 6, 0, 0, 0, 18, 13, 
    0, 0, 0, 0, 0, 0, 16, 62, 0, 6, 13, 7, 0, 0, 7, 
    0, 5, 8, 0, 104, 136, 12, 0, 0, 0, 38, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 49, 0, 3, 0, 0, 5, 21, 35, 0, 0, 28, 153, 54, 0, 
    0, 0, 0, 0, 47, 10, 0, 0, 7, 0, 0, 3, 0, 0, 41, 
    0, 0, 4, 15, 0, 3, 39, 6, 0, 0, 27, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 7, 
    0, 0, 0, 3, 19, 137, 0, 0, 0, 0, 0, 0, 0, 5, 3, 
    0, 0, 3, 0, 0, 0, 0, 11, 12, 28, 3, 9, 10, 16, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 4, 5, 6, 0, 4, 0, 3, 
    
    -- channel=132
    7, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 46, 29, 0, 51, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 59, 0, 0, 0, 10, 0, 0, 0, 0, 0, 58, 0, 
    0, 0, 0, 71, 0, 0, 0, 92, 0, 0, 0, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 2, 33, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 77, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 3, 103, 0, 16, 0, 
    8, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 43, 0, 0, 0, 103, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 38, 0, 0, 0, 50, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 66, 0, 0, 0, 41, 18, 0, 0, 37, 0, 0, 
    0, 4, 0, 0, 0, 0, 72, 0, 12, 1, 0, 0, 3, 0, 0, 
    21, 0, 0, 0, 0, 0, 83, 12, 51, 0, 0, 0, 0, 0, 0, 
    
    -- channel=133
    18, 0, 18, 39, 45, 4, 46, 17, 106, 142, 0, 7, 42, 38, 51, 
    12, 0, 0, 0, 22, 18, 0, 3, 34, 173, 0, 25, 36, 34, 44, 
    12, 0, 0, 0, 0, 156, 0, 0, 23, 0, 0, 0, 12, 12, 29, 
    172, 0, 0, 56, 0, 67, 102, 70, 0, 0, 8, 0, 0, 50, 0, 
    90, 0, 21, 105, 0, 0, 53, 104, 0, 0, 0, 0, 10, 98, 0, 
    26, 0, 34, 76, 0, 0, 80, 24, 23, 0, 0, 0, 10, 135, 11, 
    25, 0, 45, 45, 15, 0, 74, 0, 36, 0, 0, 0, 0, 63, 47, 
    43, 0, 172, 0, 28, 19, 0, 62, 0, 0, 40, 0, 0, 38, 0, 
    118, 0, 41, 0, 8, 17, 29, 121, 0, 37, 43, 120, 0, 0, 0, 
    68, 0, 0, 14, 0, 0, 0, 39, 126, 0, 43, 16, 7, 34, 0, 
    16, 66, 0, 0, 1, 80, 0, 0, 51, 76, 0, 0, 10, 40, 16, 
    0, 105, 0, 0, 29, 12, 0, 0, 41, 104, 0, 1, 2, 56, 58, 
    22, 53, 0, 0, 115, 0, 0, 0, 47, 64, 0, 4, 0, 3, 35, 
    36, 75, 0, 0, 73, 38, 20, 25, 48, 1, 0, 15, 47, 0, 8, 
    19, 68, 0, 0, 28, 60, 54, 15, 79, 0, 0, 14, 39, 0, 0, 
    
    -- channel=134
    0, 59, 9, 0, 0, 12, 0, 0, 0, 0, 33, 0, 0, 0, 0, 
    0, 15, 41, 3, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 26, 66, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 60, 0, 0, 200, 116, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 78, 
    0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    13, 0, 0, 1, 0, 0, 49, 29, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    18, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 32, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 25, 73, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    66, 0, 0, 0, 3, 52, 38, 24, 0, 0, 27, 0, 13, 26, 0, 
    0, 0, 0, 0, 0, 23, 32, 30, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 18, 39, 1, 39, 0, 0, 0, 11, 19, 0, 
    0, 0, 0, 0, 25, 6, 53, 0, 43, 21, 0, 0, 0, 25, 0, 
    0, 0, 0, 0, 23, 38, 27, 39, 0, 0, 14, 0, 0, 16, 0, 
    13, 0, 0, 0, 28, 55, 52, 67, 0, 0, 7, 0, 0, 0, 0, 
    2, 0, 3, 8, 3, 15, 29, 39, 35, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 6, 7, 34, 0, 0, 17, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 17, 22, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 31, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    13, 56, 144, 116, 92, 114, 132, 115, 99, 69, 50, 139, 152, 154, 157, 
    13, 37, 141, 84, 49, 58, 73, 100, 106, 50, 101, 101, 118, 128, 136, 
    18, 31, 113, 106, 49, 37, 58, 66, 60, 28, 95, 56, 65, 68, 81, 
    97, 45, 128, 74, 60, 21, 54, 72, 55, 53, 64, 56, 55, 69, 54, 
    51, 96, 78, 59, 74, 34, 43, 46, 44, 42, 47, 91, 60, 61, 78, 
    71, 68, 76, 51, 71, 37, 49, 19, 55, 41, 51, 67, 51, 56, 76, 
    78, 72, 85, 93, 72, 22, 39, 17, 51, 50, 35, 83, 56, 48, 48, 
    64, 72, 96, 104, 38, 54, 6, 63, 51, 43, 68, 49, 64, 69, 38, 
    69, 66, 76, 97, 28, 56, 39, 47, 66, 58, 89, 105, 87, 48, 61, 
    52, 54, 73, 67, 56, 37, 22, 28, 81, 72, 90, 92, 85, 96, 101, 
    52, 52, 53, 60, 53, 64, 65, 46, 39, 99, 59, 89, 91, 70, 77, 
    55, 57, 64, 43, 62, 45, 87, 68, 73, 59, 93, 75, 82, 72, 76, 
    57, 58, 67, 52, 83, 49, 93, 78, 75, 65, 89, 67, 77, 64, 85, 
    58, 64, 59, 46, 45, 91, 104, 88, 74, 59, 89, 73, 68, 81, 76, 
    47, 69, 48, 46, 42, 69, 64, 88, 78, 69, 76, 78, 70, 87, 80, 
    
    -- channel=137
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 16, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    20, 0, 21, 0, 0, 0, 0, 0, 10, 0, 0, 6, 0, 0, 0, 
    14, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    10, 0, 72, 0, 0, 0, 0, 0, 0, 0, 56, 20, 5, 4, 0, 
    33, 0, 88, 0, 0, 0, 0, 2, 4, 0, 41, 0, 0, 20, 10, 
    41, 10, 46, 0, 3, 0, 0, 0, 0, 0, 15, 46, 17, 44, 48, 
    40, 15, 58, 0, 3, 0, 0, 0, 20, 0, 0, 63, 39, 79, 91, 
    52, 12, 0, 32, 2, 0, 9, 0, 12, 6, 0, 48, 32, 54, 32, 
    53, 2, 0, 22, 0, 0, 0, 0, 8, 0, 2, 0, 15, 64, 22, 
    89, 16, 0, 0, 0, 5, 0, 25, 0, 0, 58, 0, 19, 45, 28, 
    84, 7, 0, 0, 2, 0, 0, 0, 0, 2, 1, 0, 0, 13, 0, 
    60, 35, 19, 0, 0, 0, 10, 0, 0, 12, 0, 0, 0, 0, 0, 
    51, 81, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    60, 89, 30, 0, 33, 0, 18, 0, 0, 0, 7, 0, 0, 0, 0, 
    54, 89, 38, 28, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    42, 108, 23, 28, 0, 7, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    
    -- channel=139
    0, 0, 145, 119, 127, 124, 131, 123, 110, 59, 29, 169, 161, 159, 158, 
    0, 0, 142, 85, 133, 130, 137, 148, 166, 67, 98, 187, 184, 178, 173, 
    0, 0, 80, 100, 165, 146, 97, 132, 128, 61, 182, 185, 196, 196, 188, 
    0, 0, 152, 139, 161, 154, 100, 92, 74, 97, 194, 181, 220, 232, 186, 
    136, 138, 181, 105, 143, 173, 170, 108, 83, 90, 169, 220, 236, 195, 175, 
    178, 171, 192, 111, 159, 172, 153, 67, 107, 97, 158, 223, 242, 205, 166, 
    183, 165, 165, 151, 141, 118, 155, 85, 144, 129, 144, 222, 239, 228, 166, 
    185, 165, 141, 164, 177, 163, 131, 146, 126, 124, 169, 188, 211, 258, 186, 
    186, 135, 147, 170, 173, 184, 157, 149, 103, 102, 168, 88, 147, 180, 181, 
    188, 146, 187, 179, 185, 209, 182, 144, 130, 135, 150, 115, 91, 145, 144, 
    198, 176, 172, 186, 186, 174, 168, 175, 174, 171, 79, 126, 146, 118, 120, 
    200, 181, 173, 207, 216, 151, 169, 168, 180, 106, 107, 128, 151, 126, 90, 
    194, 176, 160, 202, 211, 70, 187, 167, 154, 100, 114, 107, 137, 100, 107, 
    186, 163, 133, 203, 172, 128, 167, 135, 117, 57, 105, 95, 86, 82, 115, 
    153, 152, 110, 192, 179, 183, 125, 107, 89, 56, 83, 100, 73, 101, 104, 
    
    -- channel=140
    18, 95, 49, 0, 0, 0, 0, 0, 0, 0, 59, 17, 0, 0, 0, 
    23, 74, 84, 0, 0, 0, 0, 0, 0, 0, 220, 0, 0, 0, 0, 
    23, 44, 113, 27, 19, 0, 0, 0, 0, 0, 107, 0, 0, 0, 0, 
    76, 148, 258, 0, 0, 0, 0, 0, 1, 51, 0, 7, 0, 0, 0, 
    0, 92, 0, 0, 73, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 24, 0, 0, 0, 51, 28, 0, 5, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 82, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 48, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 25, 0, 
    
    -- channel=141
    0, 78, 62, 0, 0, 0, 0, 0, 0, 0, 95, 0, 0, 0, 0, 
    0, 0, 220, 2, 0, 0, 17, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 259, 0, 63, 0, 0, 100, 47, 6, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 118, 0, 0, 0, 18, 25, 25, 17, 0, 0, 16, 
    0, 0, 0, 0, 79, 0, 0, 0, 11, 0, 84, 0, 0, 0, 0, 
    0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 97, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 
    0, 0, 0, 210, 0, 0, 18, 0, 91, 0, 0, 194, 69, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 50, 0, 177, 122, 104, 
    0, 0, 0, 0, 0, 30, 4, 0, 0, 5, 0, 24, 0, 0, 0, 
    0, 0, 46, 0, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 2, 0, 24, 0, 0, 
    0, 0, 6, 0, 0, 0, 83, 0, 0, 0, 27, 0, 30, 20, 0, 
    0, 0, 1, 14, 0, 0, 0, 0, 0, 0, 24, 0, 0, 6, 0, 
    0, 0, 0, 70, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=143
    0, 30, 45, 15, 7, 50, 38, 42, 6, 0, 53, 15, 39, 48, 47, 
    0, 0, 32, 28, 0, 0, 21, 20, 0, 0, 20, 9, 21, 36, 35, 
    0, 0, 35, 21, 0, 0, 0, 2, 0, 25, 0, 22, 9, 10, 9, 
    0, 52, 0, 3, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 23, 
    47, 8, 11, 8, 0, 0, 0, 0, 0, 0, 2, 1, 0, 20, 45, 
    26, 14, 18, 34, 0, 0, 0, 0, 0, 0, 0, 21, 7, 34, 62, 
    37, 37, 18, 10, 0, 0, 0, 0, 0, 0, 0, 8, 19, 22, 38, 
    40, 30, 0, 0, 0, 0, 0, 0, 1, 7, 0, 36, 27, 0, 56, 
    24, 27, 0, 0, 0, 0, 0, 0, 18, 7, 0, 0, 19, 36, 65, 
    43, 30, 0, 0, 0, 0, 0, 0, 0, 21, 0, 22, 20, 0, 0, 
    31, 7, 4, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 6, 
    27, 20, 4, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    29, 49, 27, 0, 0, 7, 0, 0, 0, 5, 7, 4, 0, 8, 0, 
    33, 53, 58, 0, 0, 0, 0, 3, 7, 18, 2, 4, 0, 8, 12, 
    39, 53, 62, 0, 0, 0, 4, 4, 0, 30, 4, 6, 6, 3, 0, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 18, 18, 8, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 118, 84, 76, 63, 66, 69, 6, 0, 0, 0, 0, 0, 
    0, 0, 7, 132, 3, 9, 41, 60, 63, 30, 0, 0, 0, 0, 0, 
    0, 0, 5, 145, 34, 23, 96, 60, 45, 33, 45, 0, 0, 1, 0, 
    0, 5, 75, 117, 72, 97, 89, 78, 89, 73, 53, 2, 0, 0, 0, 
    15, 81, 77, 140, 15, 59, 94, 79, 45, 24, 40, 0, 0, 0, 0, 
    61, 100, 57, 62, 117, 155, 142, 120, 103, 115, 98, 64, 65, 44, 0, 
    38, 77, 6, 134, 68, 20, 46, 87, 36, 0, 34, 19, 0, 20, 0, 
    50, 94, 55, 87, 54, 95, 70, 28, 83, 74, 89, 86, 67, 112, 0, 
    34, 125, 53, 91, 76, 79, 64, 69, 105, 120, 120, 100, 100, 72, 0, 
    41, 130, 70, 60, 73, 41, 37, 144, 0, 52, 36, 0, 114, 73, 0, 
    66, 129, 0, 80, 99, 68, 56, 55, 49, 0, 0, 68, 73, 60, 0, 
    36, 76, 97, 81, 71, 96, 52, 40, 11, 4, 70, 142, 90, 24, 0, 
    65, 64, 88, 88, 71, 82, 52, 56, 57, 65, 63, 138, 68, 42, 0, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 87, 84, 135, 199, 167, 93, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 17, 
    0, 0, 101, 21, 0, 62, 31, 4, 6, 0, 0, 0, 0, 0, 0, 
    3, 18, 0, 10, 123, 0, 3, 75, 93, 59, 121, 90, 0, 0, 0, 
    19, 90, 88, 0, 0, 0, 0, 0, 0, 8, 27, 63, 163, 116, 0, 
    46, 142, 0, 0, 72, 41, 39, 85, 201, 181, 131, 216, 173, 68, 0, 
    0, 0, 7, 185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 
    0, 18, 100, 0, 104, 25, 115, 56, 116, 100, 132, 112, 83, 89, 0, 
    0, 0, 0, 0, 30, 38, 0, 33, 63, 15, 5, 0, 70, 0, 0, 
    0, 68, 0, 0, 0, 48, 236, 82, 87, 22, 0, 96, 69, 199, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 
    0, 22, 0, 16, 0, 0, 0, 0, 0, 185, 101, 48, 0, 0, 0, 
    10, 0, 0, 46, 11, 0, 0, 0, 0, 15, 88, 33, 0, 0, 0, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 49, 22, 14, 38, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 113, 0, 0, 0, 90, 
    0, 0, 0, 0, 108, 44, 0, 0, 0, 0, 0, 66, 0, 0, 10, 
    0, 0, 0, 0, 23, 44, 0, 0, 0, 35, 0, 81, 16, 0, 0, 
    45, 0, 0, 0, 98, 0, 0, 0, 0, 11, 15, 90, 89, 0, 0, 
    28, 0, 8, 0, 10, 0, 0, 0, 23, 0, 0, 96, 87, 100, 5, 
    0, 0, 141, 0, 0, 0, 0, 0, 25, 44, 0, 59, 143, 91, 124, 
    0, 0, 65, 0, 51, 50, 37, 0, 0, 36, 0, 0, 26, 0, 245, 
    0, 0, 3, 0, 56, 0, 44, 179, 0, 17, 0, 0, 0, 0, 329, 
    0, 0, 0, 0, 1, 80, 62, 0, 123, 0, 0, 16, 0, 8, 293, 
    0, 0, 60, 0, 0, 37, 131, 0, 218, 21, 0, 0, 0, 4, 386, 
    0, 0, 0, 0, 0, 0, 2, 25, 101, 154, 0, 0, 0, 80, 309, 
    0, 0, 0, 0, 0, 0, 0, 30, 67, 92, 59, 0, 0, 122, 275, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 31, 60, 0, 0, 83, 273, 
    
    -- channel=147
    0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 25, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 12, 84, 67, 29, 53, 129, 161, 9, 0, 0, 2, 26, 
    0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 9, 44, 22, 0, 0, 
    0, 0, 0, 15, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 89, 45, 32, 0, 29, 60, 11, 73, 63, 0, 0, 
    36, 35, 51, 22, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 
    0, 74, 8, 0, 47, 197, 218, 57, 0, 38, 25, 0, 54, 99, 50, 
    0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 55, 121, 0, 54, 158, 128, 147, 25, 112, 62, 
    2, 0, 22, 0, 37, 34, 3, 16, 157, 167, 163, 164, 144, 0, 0, 
    0, 20, 0, 0, 0, 0, 57, 23, 0, 0, 0, 0, 0, 104, 76, 
    14, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 126, 41, 8, 0, 10, 
    9, 6, 2, 27, 0, 0, 0, 1, 14, 28, 30, 25, 0, 11, 32, 
    
    -- channel=148
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 199, 89, 32, 54, 120, 79, 19, 0, 0, 0, 11, 0, 
    0, 0, 22, 97, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 
    0, 0, 0, 213, 0, 24, 111, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 188, 92, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 42, 0, 154, 0, 0, 0, 23, 23, 0, 21, 0, 0, 0, 0, 
    0, 103, 10, 0, 0, 13, 46, 7, 0, 109, 63, 0, 25, 2, 0, 
    61, 153, 0, 146, 27, 0, 0, 3, 99, 69, 14, 96, 0, 0, 0, 
    0, 95, 0, 232, 0, 34, 2, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 153, 54, 0, 65, 0, 0, 0, 101, 0, 26, 0, 20, 38, 0, 
    0, 152, 0, 0, 8, 0, 0, 88, 0, 0, 0, 0, 67, 0, 0, 
    0, 221, 0, 0, 73, 15, 28, 64, 0, 44, 0, 71, 102, 99, 0, 
    0, 0, 0, 24, 0, 36, 13, 0, 0, 0, 46, 149, 110, 0, 0, 
    0, 55, 0, 81, 0, 47, 0, 0, 0, 73, 0, 126, 7, 0, 0, 
    3, 0, 0, 113, 0, 18, 0, 0, 0, 0, 0, 70, 41, 0, 0, 
    
    -- channel=149
    0, 0, 28, 30, 0, 0, 0, 0, 0, 0, 3, 0, 55, 0, 48, 
    0, 0, 34, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 
    0, 0, 16, 239, 0, 0, 0, 0, 0, 0, 0, 0, 28, 82, 0, 
    0, 4, 0, 185, 0, 0, 14, 0, 0, 0, 0, 0, 5, 81, 0, 
    0, 16, 2, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 20, 
    0, 41, 64, 136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 32, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 58, 0, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 109, 0, 1, 0, 0, 0, 25, 29, 0, 126, 52, 0, 0, 0, 
    37, 175, 0, 96, 0, 19, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 190, 17, 47, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 
    0, 218, 0, 45, 99, 0, 0, 86, 0, 0, 0, 0, 139, 0, 0, 
    0, 201, 0, 21, 88, 67, 0, 0, 0, 0, 23, 220, 40, 0, 0, 
    0, 0, 74, 19, 0, 113, 1, 0, 0, 0, 0, 197, 51, 0, 0, 
    0, 0, 63, 0, 0, 34, 3, 0, 0, 0, 0, 51, 48, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 13, 7, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 58, 81, 106, 116, 167, 200, 167, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 0, 0, 0, 12, 
    0, 0, 0, 0, 68, 165, 0, 9, 0, 21, 0, 38, 0, 0, 0, 
    0, 0, 33, 43, 4, 0, 64, 10, 22, 25, 0, 45, 0, 0, 0, 
    8, 0, 0, 0, 4, 0, 0, 27, 14, 0, 57, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 79, 21, 94, 165, 75, 76, 94, 182, 7, 
    8, 0, 74, 0, 0, 0, 0, 0, 77, 63, 7, 125, 89, 0, 56, 
    0, 12, 0, 61, 12, 119, 117, 0, 0, 0, 0, 0, 0, 11, 125, 
    0, 0, 95, 0, 28, 0, 0, 127, 0, 0, 0, 0, 50, 0, 51, 
    0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 116, 0, 0, 0, 47, 117, 111, 178, 15, 50, 98, 0, 82, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 89, 18, 0, 0, 17, 0, 
    0, 0, 0, 3, 1, 0, 0, 0, 51, 0, 44, 0, 6, 0, 22, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 37, 0, 0, 0, 
    
    -- channel=151
    47, 43, 66, 21, 29, 26, 33, 49, 48, 34, 29, 22, 49, 13, 27, 
    57, 55, 73, 63, 88, 91, 48, 45, 46, 4, 0, 28, 24, 9, 0, 
    58, 58, 69, 152, 151, 185, 177, 200, 177, 118, 0, 40, 34, 15, 0, 
    57, 77, 47, 171, 112, 105, 191, 193, 191, 161, 121, 0, 28, 35, 0, 
    51, 76, 73, 153, 152, 146, 166, 180, 168, 158, 190, 27, 40, 78, 42, 
    23, 77, 80, 184, 81, 158, 169, 160, 155, 158, 122, 78, 32, 59, 58, 
    29, 46, 20, 98, 154, 151, 197, 149, 136, 149, 98, 51, 28, 0, 56, 
    30, 16, 0, 113, 144, 140, 117, 118, 73, 71, 83, 58, 61, 85, 25, 
    44, 45, 29, 7, 102, 46, 90, 110, 105, 74, 150, 112, 108, 103, 0, 
    65, 88, 24, 53, 60, 96, 69, 16, 128, 94, 108, 102, 107, 86, 0, 
    55, 91, 66, 80, 44, 28, 85, 108, 53, 116, 119, 111, 58, 120, 0, 
    95, 105, 15, 118, 80, 35, 10, 62, 0, 49, 96, 69, 61, 55, 0, 
    110, 171, 85, 129, 104, 61, 31, 32, 10, 38, 102, 176, 43, 31, 14, 
    109, 120, 134, 111, 90, 82, 32, 30, 34, 46, 57, 172, 34, 27, 27, 
    128, 134, 148, 68, 83, 64, 46, 54, 51, 60, 62, 110, 42, 39, 48, 
    
    -- channel=152
    27, 41, 41, 18, 22, 16, 18, 35, 51, 31, 42, 32, 22, 50, 27, 
    20, 22, 24, 0, 0, 0, 0, 0, 0, 0, 22, 46, 42, 43, 52, 
    19, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 56, 49, 41, 44, 
    19, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 23, 45, 66, 
    22, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 26, 34, 
    26, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 21, 
    47, 19, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    74, 6, 5, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 79, 0, 0, 0, 0, 0, 4, 0, 17, 18, 27, 0, 2, 
    23, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 10, 0, 10, 0, 
    0, 0, 10, 11, 0, 0, 0, 0, 0, 10, 21, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    
    -- channel=153
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=154
    0, 0, 10, 0, 0, 0, 0, 0, 10, 12, 9, 3, 0, 29, 8, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 24, 13, 1, 35, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 0, 27, 47, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 23, 0, 41, 0, 0, 0, 
    0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    211, 205, 224, 165, 155, 148, 154, 182, 224, 228, 224, 215, 188, 197, 153, 
    242, 241, 255, 138, 144, 149, 136, 166, 203, 197, 188, 226, 227, 210, 192, 
    249, 251, 232, 103, 49, 86, 68, 77, 86, 116, 149, 231, 234, 185, 172, 
    248, 258, 193, 127, 123, 149, 146, 120, 115, 103, 168, 205, 192, 200, 154, 
    244, 253, 189, 75, 111, 119, 103, 106, 125, 111, 144, 183, 223, 210, 166, 
    224, 256, 114, 83, 36, 65, 84, 78, 76, 91, 112, 119, 219, 248, 250, 
    208, 185, 131, 38, 53, 82, 82, 49, 64, 111, 67, 100, 186, 196, 241, 
    206, 95, 79, 155, 50, 28, 29, 44, 22, 0, 23, 29, 31, 94, 218, 
    176, 60, 138, 24, 50, 74, 46, 16, 25, 24, 62, 24, 69, 116, 161, 
    185, 78, 98, 0, 33, 20, 32, 51, 114, 102, 105, 95, 143, 40, 87, 
    190, 57, 44, 7, 0, 0, 0, 57, 12, 56, 42, 48, 44, 54, 73, 
    187, 63, 22, 54, 0, 0, 33, 0, 48, 57, 89, 165, 0, 60, 16, 
    148, 59, 63, 122, 10, 0, 0, 0, 0, 100, 152, 151, 0, 0, 46, 
    164, 152, 95, 111, 39, 0, 0, 0, 2, 99, 101, 138, 0, 0, 40, 
    137, 121, 116, 37, 33, 0, 0, 0, 0, 22, 60, 69, 0, 0, 55, 
    
    -- channel=156
    0, 0, 0, 0, 0, 0, 0, 64, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 24, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 130, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 11, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 72, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 106, 0, 41, 0, 0, 0, 205, 182, 64, 170, 234, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 
    0, 0, 34, 0, 0, 0, 44, 0, 0, 0, 0, 43, 0, 85, 0, 
    0, 0, 0, 94, 0, 21, 0, 0, 131, 0, 0, 34, 0, 0, 41, 
    0, 0, 123, 0, 0, 0, 12, 17, 7, 284, 8, 0, 0, 14, 147, 
    0, 0, 0, 0, 0, 0, 34, 57, 82, 0, 0, 0, 0, 98, 52, 
    0, 0, 0, 0, 0, 0, 17, 33, 20, 9, 0, 0, 0, 65, 171, 
    
    -- channel=157
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 44, 100, 54, 128, 178, 104, 13, 0, 0, 0, 11, 
    0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 160, 0, 0, 0, 76, 
    0, 0, 0, 0, 147, 32, 0, 7, 0, 0, 0, 174, 0, 0, 0, 
    0, 0, 0, 0, 131, 0, 11, 17, 15, 0, 0, 94, 0, 0, 0, 
    53, 0, 0, 0, 131, 26, 0, 24, 38, 26, 118, 19, 134, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 44, 0, 52, 156, 162, 1, 
    3, 0, 109, 0, 0, 0, 31, 4, 97, 98, 46, 93, 143, 44, 269, 
    0, 0, 2, 0, 45, 32, 0, 0, 0, 0, 0, 0, 0, 0, 152, 
    0, 0, 208, 0, 123, 0, 38, 117, 0, 72, 45, 70, 171, 0, 130, 
    0, 0, 0, 0, 0, 104, 0, 0, 164, 0, 0, 22, 0, 0, 0, 
    0, 0, 230, 0, 0, 0, 121, 16, 154, 0, 3, 67, 0, 176, 87, 
    1, 0, 0, 66, 0, 0, 0, 8, 0, 191, 0, 0, 0, 39, 20, 
    0, 0, 0, 92, 0, 0, 0, 0, 0, 135, 140, 0, 0, 44, 48, 
    0, 0, 0, 0, 14, 0, 0, 0, 0, 14, 60, 120, 0, 40, 52, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 6, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 3, 46, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
