library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    517, 513, 519, 522, 520, 524, 525, 532, 531, 513, 504, 510, 529, 552, 559, 562, 548, 524, 502, 487, 478, 476, 480, 489, 494, 512, 529, 546, 553, 550, 
    537, 530, 535, 530, 523, 523, 526, 532, 523, 479, 469, 496, 522, 541, 540, 529, 521, 489, 453, 428, 425, 434, 446, 461, 468, 485, 510, 534, 545, 545, 
    534, 530, 540, 537, 528, 525, 530, 532, 513, 404, 393, 448, 489, 499, 500, 500, 485, 430, 377, 340, 336, 352, 389, 411, 432, 455, 478, 502, 525, 537, 
    504, 493, 510, 528, 531, 532, 539, 540, 521, 394, 373, 413, 462, 482, 475, 470, 449, 362, 294, 248, 248, 279, 316, 350, 397, 430, 446, 460, 494, 521, 
    483, 470, 473, 504, 530, 541, 544, 548, 536, 434, 423, 417, 435, 456, 445, 443, 398, 298, 226, 206, 225, 251, 274, 304, 364, 411, 430, 430, 467, 505, 
    453, 444, 438, 473, 524, 546, 543, 540, 535, 500, 461, 403, 395, 414, 386, 374, 350, 270, 196, 198, 248, 278, 278, 307, 362, 405, 422, 417, 445, 488, 
    412, 374, 367, 429, 506, 536, 522, 493, 496, 473, 403, 328, 319, 348, 336, 330, 330, 290, 219, 210, 265, 305, 315, 332, 359, 397, 432, 428, 430, 468, 
    305, 257, 266, 369, 479, 515, 442, 344, 334, 346, 293, 245, 258, 309, 322, 328, 346, 334, 253, 226, 253, 296, 334, 343, 355, 373, 425, 449, 435, 446, 
    195, 123, 171, 318, 448, 502, 351, 170, 140, 190, 181, 190, 231, 285, 325, 336, 372, 366, 249, 206, 210, 273, 324, 324, 333, 350, 401, 448, 442, 441, 
    124, 54, 98, 279, 423, 505, 351, 116, 28, 107, 130, 155, 213, 271, 313, 333, 399, 343, 184, 158, 164, 251, 310, 310, 306, 321, 363, 420, 430, 441, 
    97, 32, 69, 251, 401, 508, 428, 202, 96, 145, 144, 120, 181, 244, 297, 299, 391, 287, 118, 114, 146, 255, 307, 307, 301, 310, 329, 369, 392, 438, 
    95, 22, 86, 246, 379, 486, 520, 312, 209, 190, 161, 81, 127, 205, 258, 270, 358, 225, 83, 102, 165, 271, 313, 323, 311, 304, 297, 325, 349, 429, 
    83, 14, 108, 251, 358, 449, 536, 387, 289, 197, 137, 65, 100, 157, 204, 246, 333, 189, 83, 107, 175, 255, 302, 316, 310, 290, 269, 295, 337, 418, 
    54, 10, 111, 241, 311, 385, 491, 404, 314, 137, 47, 46, 105, 154, 199, 249, 318, 206, 116, 126, 188, 260, 307, 310, 295, 265, 257, 305, 361, 426, 
    26, 0, 66, 211, 244, 294, 390, 402, 310, 126, 42, 85, 159, 206, 233, 274, 325, 243, 194, 184, 200, 252, 314, 313, 286, 266, 282, 349, 404, 452, 
    0, 0, 5, 166, 201, 212, 269, 351, 306, 187, 120, 180, 236, 266, 286, 284, 296, 288, 317, 260, 235, 284, 345, 349, 321, 297, 321, 382, 422, 463, 
    0, 0, 0, 111, 176, 166, 179, 283, 285, 296, 247, 258, 293, 272, 294, 281, 258, 281, 351, 316, 297, 328, 381, 385, 371, 351, 378, 414, 449, 481, 
    0, 0, 0, 66, 175, 151, 152, 193, 227, 331, 299, 297, 277, 209, 245, 269, 232, 270, 319, 315, 345, 388, 415, 381, 375, 362, 402, 433, 467, 493, 
    0, 0, 0, 43, 162, 141, 105, 141, 210, 319, 290, 283, 198, 120, 165, 233, 250, 289, 307, 336, 379, 408, 408, 344, 340, 334, 392, 438, 461, 473, 
    3, 0, 0, 50, 168, 128, 26, 26, 121, 237, 211, 183, 83, 18, 61, 163, 221, 300, 342, 362, 360, 351, 326, 271, 251, 246, 286, 325, 340, 345, 
    0, 0, 0, 55, 160, 77, 0, 0, 0, 99, 125, 75, 7, 0, 18, 109, 184, 263, 314, 312, 280, 256, 213, 188, 165, 149, 156, 186, 193, 197, 
    0, 0, 0, 29, 111, 0, 0, 0, 0, 36, 73, 65, 47, 48, 62, 106, 141, 199, 217, 200, 169, 147, 123, 104, 86, 73, 66, 84, 89, 89, 
    0, 0, 0, 10, 43, 0, 0, 0, 0, 71, 106, 118, 121, 124, 128, 140, 141, 151, 143, 123, 107, 98, 82, 63, 51, 42, 40, 50, 50, 47, 
    0, 0, 0, 4, 0, 0, 0, 0, 66, 116, 127, 132, 135, 144, 143, 141, 138, 134, 120, 99, 85, 74, 56, 34, 30, 31, 32, 30, 15, 0, 
    24, 19, 3, 25, 0, 0, 0, 46, 112, 117, 103, 108, 115, 123, 129, 134, 131, 123, 107, 85, 62, 41, 28, 19, 21, 27, 12, 0, 0, 0, 
    15, 38, 42, 37, 0, 0, 0, 93, 122, 115, 91, 100, 115, 122, 124, 124, 116, 103, 84, 66, 44, 18, 6, 14, 27, 21, 0, 0, 0, 0, 
    5, 29, 48, 38, 0, 0, 0, 96, 118, 104, 81, 90, 101, 114, 120, 117, 101, 84, 67, 54, 36, 20, 19, 27, 28, 0, 0, 0, 0, 0, 
    4, 17, 32, 44, 0, 0, 49, 107, 131, 114, 84, 79, 81, 96, 104, 101, 87, 73, 59, 54, 50, 46, 43, 30, 5, 0, 0, 0, 36, 53, 
    7, 20, 28, 43, 51, 34, 110, 135, 151, 134, 112, 100, 90, 96, 96, 91, 72, 51, 43, 52, 61, 69, 57, 18, 0, 0, 0, 0, 61, 78, 
    17, 35, 45, 46, 74, 94, 126, 154, 165, 152, 143, 131, 128, 134, 123, 103, 73, 40, 31, 50, 69, 86, 60, 3, 0, 0, 0, 12, 59, 92, 
    
    
    others => 0);
end gold_package;
