library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    174, 174, 112, 165, 0, 32, 0, 109, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 78, 0, 0, 6, 89, 5, 88, 50, 50, 0, 161, 63, 68, 812, 370, 192, 154, 921, 191, 41, 0, 1072, 0, 0, 0, 1094, 0, 0, 0, 316, 124, 26, 21, 265, 117, 47, 99, 166, 31, 40, 97, 0, 23, 0, 158, 27, 35, 3, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 277, 252, 344, 4, 462, 292, 386, 57, 866, 784, 959, 1204, 443, 558, 1184, 1304, 0, 0, 0, 19, 0, 92, 95, 0, 0, 76, 12, 1, 612, 445, 463, 482, 349, 369, 248, 370, 67, 126, 101, 281, 0, 0, 0, 106, 0, 0, 0, 0, 770, 711, 625, 346, 570, 516, 433, 136, 564, 388, 675, 859, 0, 0, 406, 349, 912, 812, 445, 374, 779, 667, 341, 285, 506, 336, 152, 198, 93, 0, 0, 0, 225, 347, 259, 540, 287, 247, 217, 599, 121, 319, 145, 600, 0, 134, 0, 738, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 90, 206, 59, 535, 564, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 465, 359, 361, 391, 804, 742, 997, 1147, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 0, 0, 10, 133, 196, 23, 0, 57, 153, 101, 0, 0, 0, 179, 128, 91, 208, 0, 0, 0, 126, 157, 199, 78, 529, 370, 360, 178, 953, 856, 683, 807, 828, 719, 1036, 1228, 503, 0, 0, 0, 756, 0, 0, 0, 1078, 0, 0, 0, 1340, 0, 19, 4, 522, 381, 224, 279, 323, 195, 68, 93, 0, 0, 0, 0, 147, 0, 0, 0, 241, 160, 115, 0, 616, 80, 27, 0, 898, 0, 157, 278, 790, 302, 535, 574, 0, 0, 0, 0, 722, 166, 145, 0, 1188, 474, 652, 713, 1334, 655, 1163, 1215, 267, 169, 336, 166, 628, 297, 375, 155, 618, 463, 413, 663, 605, 654, 424, 774, 34, 118, 62, 136, 0, 22, 12, 86, 0, 104, 180, 84, 23, 0, 0, 0, 140, 151, 131, 128, 74, 62, 80, 45, 0, 111, 7, 88, 0, 0, 0, 0, 273, 330, 267, 238, 160, 150, 88, 109, 4, 159, 47, 275, 0, 0, 0, 11, 350, 327, 187, 343, 31, 74, 61, 269, 0, 0, 0, 155, 0, 0, 0, 0, 351, 245, 149, 122, 189, 59, 8, 82, 40, 0, 0, 36, 0, 0, 0, 0, 304, 106, 41, 0, 598, 154, 0, 0, 882, 53, 42, 197, 958, 0, 129, 156, 0, 0, 0, 0, 125, 0, 0, 0, 581, 289, 229, 334, 829, 710, 1194, 1327, 87, 51, 62, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 904, 878, 598, 564, 483, 512, 269, 386, 0, 0, 0, 101, 0, 0, 0, 0, 0, 0, 0, 100, 0, 16, 0, 66, 0, 22, 149, 112, 315, 350, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 607, 460, 381, 388, 430, 384, 255, 298, 35, 92, 58, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 239, 81, 74, 0, 611, 530, 618, 573, 750, 845, 1018, 1057, 166, 92, 124, 11, 139, 85, 84, 1, 129, 50, 137, 139, 203, 106, 71, 0, 0, 0, 0, 0, 0, 0, 10, 26, 6, 0, 0, 0, 1257, 1314, 1106, 1189, 107, 0, 105, 0, 934, 211, 150, 0, 1217, 559, 870, 904, 1403, 903, 1146, 1220, 628, 538, 378, 203, 430, 343, 198, 132, 275, 198, 230, 395, 0, 0, 0, 0, 0, 287, 296, 781, 312, 339, 615, 999, 228, 723, 334, 1632, 83, 941, 0, 2184, 525, 597, 393, 461, 294, 417, 411, 429, 0, 263, 244, 124, 0, 0, 0, 0, 144, 9, 14, 54, 90, 47, 59, 92, 84, 62, 0, 37, 98, 59, 0, 340, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1473, 1368, 1304, 1434, 43, 0, 0, 0, 80, 80, 32, 0, 118, 129, 134, 63, 232, 245, 98, 66, 38, 0, 0, 0, 346, 0, 0, 0, 788, 0, 0, 0, 994, 0, 204, 226, 761, 726, 500, 551, 387, 449, 235, 326, 0, 12, 0, 61, 0, 0, 0, 0, 278, 280, 164, 143, 0, 40, 0, 66, 0, 0, 0, 16, 0, 0, 0, 0, 570, 470, 403, 280, 614, 412, 365, 82, 374, 482, 349, 687, 0, 0, 242, 350, 272, 191, 230, 0, 421, 236, 176, 77, 660, 563, 760, 807, 389, 591, 785, 713, 74, 119, 51, 353, 0, 62, 64, 196, 0, 0, 0, 27, 26, 0, 0, 0, 93, 0, 36, 0, 93, 0, 0, 0, 143, 0, 4, 52, 0, 11, 16, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 706, 688, 418, 349, 424, 425, 136, 306, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 116, 0, 0, 0, 0, 1452, 1332, 1077, 1205, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 141, 111, 160, 131, 189, 131, 174, 201, 53, 221, 514, 416, 427, 517, 0, 161, 120, 438, 205, 205, 309, 497, 110, 409, 278, 829, 52, 506, 0, 1064, 0, 0, 0, 0, 130, 0, 0, 0, 453, 40, 126, 167, 741, 615, 941, 1077, 444, 222, 316, 27, 474, 267, 326, 0, 632, 70, 96, 217, 660, 45, 179, 125, 418, 141, 276, 26, 374, 165, 316, 113, 458, 0, 272, 239, 285, 189, 348, 129, 0, 0, 18, 0, 80, 0, 0, 0, 99, 0, 61, 178, 84, 0, 119, 105, 
    
    
    others => 0);
end ifmap_package;
