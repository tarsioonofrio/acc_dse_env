library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -14779, -6268, 2153, -18975, -719, 17228, 6543, 28779, 15072, 26517, 18611, 2851, -3368, -35807, -8963, 11843, 

    -- weights
    -- filter=0 channel=0
    53, 59, 5, 34, 27, 18, 50, 3, 63,
    -- filter=0 channel=1
    74, 50, 0, 19, 78, 31, 51, 33, 49,
    -- filter=0 channel=2
    -60, -16, -28, -16, -70, -82, 14, -15, -73,
    -- filter=1 channel=0
    -45, -15, -18, 41, 6, -5, 19, 47, -46,
    -- filter=1 channel=1
    -16, 0, 24, -21, -27, -35, 26, -38, -49,
    -- filter=1 channel=2
    -14, -6, 23, 19, -10, 14, -6, -13, 40,
    -- filter=2 channel=0
    -15, 15, -26, 41, 34, -9, 30, 54, 61,
    -- filter=2 channel=1
    -53, 28, 11, -39, -24, -36, -24, -19, 15,
    -- filter=2 channel=2
    -32, -49, 49, -51, -56, 52, 45, -34, -28,
    -- filter=3 channel=0
    -14, 22, -39, -45, 1, 18, 0, -2, 45,
    -- filter=3 channel=1
    19, 29, -32, 43, 44, 38, 30, 33, 25,
    -- filter=3 channel=2
    75, 9, 45, 8, 62, 53, 9, 83, -9,
    -- filter=4 channel=0
    99, 93, -1, 39, 28, -10, -69, -81, -19,
    -- filter=4 channel=1
    79, 84, 39, 7, -11, -24, -59, -102, -85,
    -- filter=4 channel=2
    91, 1, -5, -12, 24, 0, 6, -59, -40,
    -- filter=5 channel=0
    26, 35, 67, -27, 42, 7, -33, 10, -13,
    -- filter=5 channel=1
    32, 1, -6, 29, -14, 30, -47, -2, -8,
    -- filter=5 channel=2
    -15, 11, 14, -29, -49, 13, -6, -59, -79,
    -- filter=6 channel=0
    36, 110, 38, 59, 56, 48, -23, -52, -45,
    -- filter=6 channel=1
    30, 28, 58, -26, -14, -44, -81, -48, -68,
    -- filter=6 channel=2
    10, -8, 71, -5, -9, -16, -52, -28, -45,
    -- filter=7 channel=0
    -33, -60, -8, -41, -19, -43, -77, -1, 25,
    -- filter=7 channel=1
    100, 69, 15, 52, 93, 91, 75, 91, 39,
    -- filter=7 channel=2
    -25, -49, -65, -70, -67, -22, -4, -68, -74,
    -- filter=8 channel=0
    -16, -84, -44, 31, -98, -132, 17, -27, -97,
    -- filter=8 channel=1
    47, -67, -72, 20, 2, -83, 16, -22, -9,
    -- filter=8 channel=2
    57, 65, 64, 76, 75, 44, 87, 63, 24,
    -- filter=9 channel=0
    1, 33, -10, -37, -51, -47, 1, 24, -21,
    -- filter=9 channel=1
    61, 78, 39, -18, 54, 76, 18, 16, 30,
    -- filter=9 channel=2
    8, -34, 14, 1, -75, -57, -73, -65, -52,
    -- filter=10 channel=0
    3, -17, -7, -4, 0, -49, -41, -36, -65,
    -- filter=10 channel=1
    37, 15, 29, 0, -25, 7, -48, -35, -15,
    -- filter=10 channel=2
    41, 46, 4, -31, 51, 42, -36, -37, 44,
    -- filter=11 channel=0
    -7, 31, -36, -32, -31, -43, -48, -5, 21,
    -- filter=11 channel=1
    38, 30, -31, 15, 15, -18, 1, -18, 29,
    -- filter=11 channel=2
    -45, 22, -44, -40, 22, 35, 4, -20, -24,
    -- filter=12 channel=0
    -41, -7, 33, -47, 8, 18, -71, 3, -52,
    -- filter=12 channel=1
    64, 48, 43, 43, 39, 75, -15, -2, 66,
    -- filter=12 channel=2
    21, 21, 55, -31, 28, 28, 41, 0, -45,
    -- filter=13 channel=0
    36, 15, 40, -31, 41, 49, 32, -29, -5,
    -- filter=13 channel=1
    -68, -4, -75, 33, -2, -31, -40, 10, -79,
    -- filter=13 channel=2
    54, 20, 53, 113, 84, 87, 74, 55, 27,
    -- filter=14 channel=0
    39, -9, 25, -31, -21, 14, -26, 47, -19,
    -- filter=14 channel=1
    -28, 8, 40, 7, -37, -11, -10, 38, 1,
    -- filter=14 channel=2
    -17, -48, 24, -11, -22, -45, 41, 42, -30,
    -- filter=15 channel=0
    57, 83, 39, 27, 102, 115, 79, 107, 108,
    -- filter=15 channel=1
    -44, -51, -42, 25, -59, -61, 44, 16, 21,
    -- filter=15 channel=2
    -87, -84, -103, -26, -59, -14, -49, -42, -62,

    others => 0);
end iwght_package;
