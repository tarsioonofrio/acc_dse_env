library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 126, 276, 171, 3, 65, 0, 0, 0, 177, 193, 129, 0, 186, 0, 27, 60, 81, 0, 0, 38, 0, 0, 0, 136, 81, 129, 0, 265, 152, 203, 31, 81, 0, 0, 33, 65, 294, 124, 124, 181, 0, 0, 36, 72, 174, 0, 0, 142, 328, 0, 90, 0, 0, 78, 0, 368, 0, 0, 0, 0, 0, 213, 0, 0, 38, 101, 105, 0, 188, 0, 77, 0, 31, 41, 0, 77, 57, 0, 75, 0, 69, 0, 102, 0, 100, 0, 0, 0, 204, 73, 65, 48, 190, 208, 0, 156, 225, 0, 0, 0, 0, 0, 0, 0, 0, 15, 76, 0, 234, 0, 0, 0, 0, 0, 237, 0, 181, 37, 239, 199, 120, 0, 0, 153, 37, 41, 0, 11, 0, 196, 21, 56, 0, 196, 111, 28, 0, 60, 193, 0, 117, 0, 114, 484, 137, 136, 2, 0, 150, 211, 0, 76, 83, 0, 0, 0, 0, 0, 158, 171, 0, 0, 185, 182, 0, 0, 231, 0, 0, 419, 0, 0, 0, 0, 0, 97, 0, 0, 4, 0, 0, 38, 48, 0, 422, 3, 0, 407, 80, 0, 38, 17, 149, 121, 0, 0, 125, 163, 319, 161, 0, 24, 58, 0, 41, 71, 80, 0, 146, 0, 129, 0, 111, 43, 0, 32, 0, 44, 0, 0, 0, 0, 17, 70, 95, 0, 265, 155, 0, 0, 0, 69, 276, 64, 379, 279, 0, 0, 0, 0, 20, 29, 158, 328, 0, 0, 171, 0, 419, 0, 175, 0, 0, 100, 0, 0, 2, 79, 0, 0, 0, 0, 0, 51, 0, 0, 0, 123, 19, 0, 15, 85, 97, 0, 0, 80, 158, 300, 0, 146, 0, 18, 397, 0, 0, 245, 0, 445, 0, 41, 0, 0, 177, 0, 187, 9, 0, 0, 0, 0, 0, 276, 0, 137, 84, 234, 19, 2, 98, 121, 188, 147, 139, 159, 212, 0, 326, 0, 219, 17, 0, 0, 104, 51, 0, 0, 322, 0, 20, 0, 346, 243, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 66, 0, 23, 0, 94, 0, 131, 0, 0, 33, 267, 58, 137, 0, 26, 0, 92, 0, 0, 0, 0, 462, 38, 201, 0, 0, 256, 0, 0, 135, 312, 0, 0, 0, 0, 0, 238, 271, 0, 0, 141, 0, 102, 0, 50, 37, 184, 171, 15, 0, 0, 0, 10, 164, 0, 207, 85, 0, 41, 75, 56, 0, 0, 0, 0, 0, 68, 44, 26, 92, 22, 36, 297, 0, 88, 38, 0, 0, 40, 177, 59, 75, 0, 35, 341, 0, 79, 48, 142, 179, 157, 112, 0, 151, 274, 0, 106, 64, 17, 0, 146, 1, 0, 2, 22, 0, 124, 0, 41, 0, 0, 0, 214, 61, 129, 4, 83, 0, 0, 428, 0, 0, 0, 227, 0, 0, 0, 0, 0, 0, 60, 237, 318, 43, 120, 0, 141, 194, 129, 200, 28, 126, 0, 107, 16, 0, 0, 0, 0, 18, 0, 0, 372, 211, 71, 128, 0, 0, 0, 64, 32, 0, 0, 0, 67, 0, 0, 0, 0, 155, 169, 224, 0, 128, 0, 0, 108, 0, 239, 107, 0, 0, 0, 91, 93, 75, 0, 3, 43, 29, 20, 425, 0, 9, 0, 5, 0, 0, 113, 45, 0, 228, 0, 13, 39, 0, 0, 25, 0, 54, 79, 169, 95, 0, 36, 1, 81, 0, 34, 92, 97, 0, 171, 0, 297, 321, 90, 10, 0, 48, 0, 0, 34, 201, 253, 0, 406, 0, 253, 110, 0, 0, 280, 230, 0, 0, 0, 14, 23, 0, 0, 0, 0, 0, 227, 63, 321, 35, 0, 0, 0, 0, 0, 30, 66, 18, 0, 0, 87, 168, 103, 0, 0, 0, 46, 0, 0, 0, 49, 0, 15, 0, 269, 179, 132, 96, 83, 27, 0, 119, 39, 288, 285, 355, 0, 0, 0, 0, 0, 71, 0, 64, 0, 0, 58, 73, 36, 28, 0, 23, 26, 0, 65, 306, 0, 82, 45, 64, 106, 154, 69, 0, 0, 103, 0, 91, 134, 228, 0, 287, 0, 0, 11, 146, 31, 130, 0, 285, 0, 102, 141, 70, 0, 0, 230, 109, 0, 0, 27, 0, 0, 0, 80, 29, 0, 0, 124, 0, 0, 202, 84, 0, 23, 0, 0, 176, 61, 78, 0, 221, 0, 143, 367, 157, 0, 0, 14, 248, 0, 0, 94, 0, 0, 122, 208, 0, 314, 370, 5, 323, 115, 17, 115, 116, 176, 0, 0, 43, 0, 73, 0, 43, 0, 181, 0, 105, 280, 326, 50, 0, 257, 163, 83, 0, 36, 203, 177, 45, 0, 124, 152, 0, 0, 74, 77, 125, 0, 0, 55, 97, 0, 148, 39, 21, 4, 0, 32, 16, 21, 0, 57, 176, 0, 139, 3, 0, 284, 0, 0, 55, 301, 0, 0, 0, 94, 161, 0, 0, 63, 0, 58, 0, 0, 0, 0, 0, 0, 0, 100, 168, 0, 49, 0, 286, 0, 39, 96, 0, 0, 0, 178, 287, 0, 64, 84, 95, 0, 0, 0, 125, 134, 132, 0, 0, 0, 145, 0, 57, 118, 62, 0, 0, 0, 41, 0, 343, 0, 0, 0, 103, 0, 0, 0, 0, 273, 0, 141, 0, 0, 213, 0, 106, 43, 62, 180, 101, 0, 0, 11, 63, 98, 0, 0, 91, 210, 332, 0, 153, 25, 45, 215, 0, 0, 225, 20, 195, 106, 244, 9, 269, 75, 128, 17, 100, 162, 171, 0, 0, 50, 39, 0, 0, 17, 0, 23, 214, 0, 31, 218, 10, 0, 288, 0, 45, 60, 43, 82, 2, 43, 0, 0, 98, 364, 0, 0, 0, 0, 0, 12, 0, 0, 188, 0, 23, 10, 0, 0, 0, 0, 217, 0, 54, 9, 49, 40, 0, 36, 0, 296, 0, 0, 0, 112, 132, 0, 32, 0, 204, 206, 0, 0, 58, 222, 0, 13, 175, 30, 150, 332, 0, 180, 221, 0, 0, 0, 0, 0, 52, 207, 2, 0, 0, 47, 128, 0, 0, 0, 7, 0, 24, 0, 0, 0, 146, 0, 19, 190, 104, 252, 230, 76, 54, 0, 21, 25, 0, 0, 0, 321, 77, 241, 0, 250, 115, 0, 21, 212, 0, 17, 0, 283, 0, 114, 0, 0, 70, 343, 282, 162, 130, 0, 0, 89, 213, 94, 13, 91, 0, 123, 47, 455, 248, 112, 82, 0, 0, 55, 0, 83, 161, 0, 68, 0, 0, 57, 0, 5, 91, 75, 0, 108, 0, 0, 152, 0, 0, 0, 0, 132, 0, 35, 0, 265, 0, 0, 48, 394, 0, 0, 0, 176, 0, 71, 42, 0, 55, 0, 67, 77, 222, 44, 119, 39, 122, 0, 3, 0, 128, 18, 0, 0, 0, 94, 62, 214, 29, 0, 0, 176, 4, 0, 0, 35, 99, 119, 0, 11, 0, 80, 2, 146, 174, 0, 246, 6, 26, 118, 190, 0, 0, 64, 0, 0, 0, 342, 0, 61, 68, 0, 66, 0, 0, 141, 0, 0, 0, 221, 0, 40, 0, 142, 108, 85, 0, 339, 0, 157, 66, 122, 114, 115, 47, 89, 107, 0, 0, 243, 201, 0, 321, 5, 90, 34, 89, 104, 194, 0, 0, 19, 124, 22, 0, 0, 121, 68, 0, 0, 0, 5, 618, 127, 0, 0, 177, 56, 417, 0, 26, 0, 0, 184, 26, 230, 32, 4, 119, 0, 41, 0, 0, 0, 198, 305, 0, 56, 220, 22, 0, 113, 46, 0, 15, 0, 30, 49, 30, 262, 7, 0, 0, 186, 115, 0, 0, 0, 0, 0, 0, 76, 0, 0, 47, 38, 344, 0, 0, 23, 0, 130, 135, 0, 0, 0, 0, 22, 0, 64, 59, 0, 169, 397, 0, 0, 0, 32, 0, 62, 0, 95, 86, 0, 0, 0, 0, 117, 128, 97, 109, 91, 196, 60, 579, 0, 0, 0, 0, 176, 208, 65, 167, 0, 304, 273, 313, 0, 0, 0, 230, 118, 0, 0, 0, 0, 122, 0, 0, 0, 85, 0, 84, 82, 0, 0, 0, 0, 71, 0, 365, 10, 33, 108, 117, 0, 159, 8, 259, 45, 0, 0, 0, 22, 239, 78, 173, 234, 186, 0, 0, 0, 0, 181, 255, 0, 0, 10, 0, 0, 56, 0, 191, 0, 0, 182, 0, 14, 47, 85, 65, 95, 0, 147, 187, 0, 0, 0, 0, 86, 6, 0, 46, 0, 0, 0, 0, 0, 0, 186, 0, 0, 0, 410, 0, 110, 0, 26, 0, 0, 30, 0, 0, 0, 0, 79, 0, 0, 0, 0, 45, 0, 0, 85, 472, 0, 141, 0, 200, 0, 123, 30, 0, 0, 83, 30, 38, 111, 0, 0, 0, 73, 0, 9, 0, 62, 63, 0, 180, 80, 89, 232, 0, 0, 221, 43, 6, 0, 87, 121, 0, 98, 232, 79, 197, 80, 0, 35, 17, 160, 0, 165, 0, 95, 0, 81, 0, 0, 0, 0, 2, 0, 0, 0, 0, 121, 47, 0, 308, 146, 0, 0, 0, 130, 89, 0, 0, 92, 330, 95, 43, 149, 0, 0, 0, 0, 16, 0, 0, 0, 0, 65, 0, 397, 109, 0, 62, 0, 223, 148, 117, 0, 332, 89, 0, 131, 92, 0, 382, 96, 0, 0, 19, 82, 200, 141, 0, 0, 0, 121, 0, 228, 255, 21, 0, 52, 0, 167, 346, 143, 56, 0, 53, 0, 0, 0, 53, 0, 242, 115, 107, 288, 0, 41, 0, 107, 72, 30, 0, 0, 0, 162, 115, 53, 0, 0, 0, 190, 0, 382, 0, 235, 0, 0, 0, 161, 141, 284, 0, 136, 0, 52, 21, 33, 112, 0, 0, 52, 0, 88, 0, 0, 232, 100, 85, 0, 0, 26, 0, 4, 0, 0, 0, 75, 0, 10, 0, 424, 102, 0, 286, 0, 0, 0, 0, 316, 53, 81, 218, 150, 0, 235, 254, 0, 0, 187, 9, 26, 164, 19, 0, 0, 108, 0, 0, 0, 21, 229, 0, 0, 161, 0, 268, 91, 0, 160, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 169, 0, 0, 326, 0, 0, 0, 0, 0, 67, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167, 0, 0, 0, 0, 0, 0, 184, 33, 75, 201, 0, 201, 0, 0, 113, 0, 0, 26, 218, 273, 340, 416, 715, 65, 96, 0, 0, 0, 0, 146, 77, 0, 0, 185, 155, 103, 0, 0, 84, 13, 0, 6, 122, 68, 28, 0, 0, 0, 0, 0, 117, 0, 293, 0, 0, 50, 0, 0, 16, 0, 0, 0, 67, 321, 0, 298, 0, 115, 94, 0, 288, 119, 132, 0, 0, 57, 0, 0, 118, 0, 0, 0, 22, 269, 62, 276, 24, 0, 0, 0, 0, 61, 99, 0, 150, 112, 116, 174, 15, 0, 102, 200, 153, 274, 0, 49, 0, 114, 25, 0, 0, 0, 120, 0, 25, 100, 0, 162, 35, 84, 99, 122, 126, 70, 204, 257, 0, 187, 0, 256, 0, 0, 230, 0, 144, 159, 87, 28, 14, 253, 0, 38, 0, 0, 115, 28, 23, 57, 38, 39, 108, 19, 0, 132, 0, 75, 153, 0, 0, 92, 0, 0, 0, 441, 243, 71, 0, 379, 0, 0, 0, 0, 0, 0, 84, 0, 82, 0, 65, 0, 0, 199, 244, 0, 0, 77, 0, 142, 188, 91, 0, 9, 225, 0, 0, 0, 0, 325, 46, 83, 0, 0, 0, 168, 0, 0, 0, 63, 0, 0, 56, 0, 98, 38, 0, 0, 0, 0, 202, 0, 121, 467, 69, 93, 345, 56, 193, 138, 311, 0, 206, 92, 139, 87, 113, 0, 0, 464, 139, 0, 9, 476, 61, 0, 0, 0, 89, 0, 78, 75, 37, 0, 0, 0, 22, 84, 134, 0, 105, 0, 189, 159, 0, 0, 0, 150, 0, 95, 70, 136, 64, 235, 65, 87, 0, 63, 0, 261, 0, 187, 184, 0, 0, 0, 0, 239, 225, 0, 60, 0, 0, 39, 0, 0, 98, 385, 73, 0, 0, 31, 311, 0, 162, 0, 59, 105, 51, 0, 0, 108, 57, 0, 84, 0, 0, 22, 351, 0, 32, 108, 0, 121, 16, 0, 371, 0, 43, 0, 28, 0, 0, 250, 83, 279, 0, 0, 69, 38, 0, 208, 62, 0, 104, 248, 238, 0, 25, 89, 0, 0, 0, 0, 0, 175, 20, 0, 0, 274, 89, 7, 0, 0, 0, 294, 19, 69, 76, 0, 0, 124, 0, 0, 0, 88, 0, 0, 380, 14, 19, 153, 0, 0, 0, 0, 0, 24, 72, 137, 0, 111, 173, 0, 295, 319, 0, 0, 44, 406, 190, 0, 187, 0, 0, 0, 86, 0, 90, 63, 38, 62, 0, 51, 0, 0, 0, 139, 131, 0, 26, 0, 60, 98, 0, 0, 139, 0, 0, 0, 151, 119, 0, 0, 121, 130, 0, 19, 119, 0, 235, 0, 0, 154, 94, 100, 28, 0, 11, 0, 57, 218, 19, 313, 52, 0, 146, 33, 68, 0, 0, 0, 250, 0, 0, 0, 0, 63, 152, 89, 119, 0, 9, 0, 57, 18, 152, 149, 0, 124, 27, 81, 0, 0, 127, 0, 101, 397, 0, 8, 0, 0, 131, 0, 48, 0, 90, 0, 77, 5, 10, 0, 2, 0, 0, 0, 39, 0, 67, 0, 322, 248, 267, 100, 0, 0, 0, 0, 84, 159, 9, 0, 0, 0, 0, 0, 178, 0, 0, 0, 0, 0, 0, 0, 385, 93, 329, 111, 17, 205, 0, 0, 0, 70, 74, 0, 308, 86, 0, 0, 27, 0, 2, 0, 0, 0, 28, 243, 0, 25, 0, 41, 132, 0, 47, 121, 69, 0, 0, 0, 47, 136, 0, 293, 0, 0, 267, 0, 0, 30, 322, 0, 237, 141, 0, 0, 119, 0, 0, 320, 202, 0, 0, 40, 138, 0, 310, 0, 9, 91, 32, 0, 0, 0, 0, 116, 0, 0, 0, 63, 0, 205, 114, 191, 0, 148, 337, 103, 48, 0, 151, 0, 26, 0, 0, 77, 0, 0, 132, 0, 109, 0, 161, 0, 0, 0, 3, 0, 235, 
    
    
    others => 0);
end ifmap_package;
