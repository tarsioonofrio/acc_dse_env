library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 59, 29, 46, 38, 35, 35, 32, 31, 26, 24, 25, 23, 29, 44, 41, 35, 31, 30, 40, 48, 51, 58, 66, 65, 57, 46, 33, 25, 11, 3, 0, 0, 14, 0, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 13, 14, 11, 0, 0, 0, 0, 19, 36, 35, 24, 8, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 31, 33, 24, 10, 0, 0, 0, 0, 0, 0, 0, 22, 18, 0, 0, 0, 2, 20, 4, 24, 13, 0, 0, 0, 0, 0, 20, 43, 24, 0, 0, 7, 24, 14, 5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 25, 8, 0, 0, 0, 19, 2, 38, 40, 4, 0, 0, 0, 0, 0, 34, 47, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 9, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 13, 22, 0, 0, 0, 9, 0, 0, 0, 0, 12, 27, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 59, 9, 0, 0, 0, 4, 0, 0, 0, 0, 34, 23, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 1, 0, 0, 0, 0, 0, 0, 0, 0, 25, 55, 3, 11, 0, 0, 0, 0, 0, 11, 46, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 15, 32, 0, 0, 0, 0, 0, 0, 64, 130, 81, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 18, 0, 0, 0, 0, 0, 0, 0, 102, 101, 30, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 4, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 18, 0, 0, 32, 56, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 18, 0, 0, 1, 27, 0, 0, 0, 12, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 12, 0, 0, 24, 40, 25, 0, 0, 0, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 73, 59, 42, 32, 35, 30, 0, 0, 0, 33, 47, 10, 0, 0, 9, 21, 20, 14, 0, 0, 0, 15, 6, 0, 0, 0, 0, 0, 2, 0, 0, 0, 71, 105, 70, 22, 4, 0, 0, 0, 0, 25, 71, 50, 26, 5, 10, 17, 21, 5, 0, 0, 0, 14, 27, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 45, 27, 0, 0, 0, 0, 0, 0, 0, 4, 43, 36, 2, 0, 0, 0, 0, 0, 0, 0, 10, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 20, 0, 0, 0, 0, 3, 12, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 7, 78, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 53, 29, 4, 0, 0, 0, 0, 0, 0, 0, 0, 18, 2, 84, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 8, 79, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 48, 58, 77, 52, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 75, 80, 32, 0, 0, 0, 0, 0, 0, 21, 20, 36, 66, 84, 96, 103, 83, 44, 28, 16, 13, 16, 23, 23, 20, 21, 23, 28, 15, 0, 0, 0, 49, 75, 91, 57, 6, 0, 0, 0, 1, 56, 35, 4, 1, 8, 25, 37, 37, 27, 26, 29, 29, 23, 21, 21, 19, 17, 19, 24, 15, 0, 0, 0, 13, 6, 58, 94, 35, 15, 0, 0, 16, 60, 43, 15, 7, 8, 12, 19, 24, 24, 24, 23, 22, 19, 15, 13, 13, 15, 19, 21, 9, 0, 0, 17, 19, 0, 12, 47, 38, 42, 0, 0, 20, 45, 33, 22, 17, 19, 22, 22, 21, 19, 19, 18, 17, 16, 14, 14, 18, 26, 30, 26, 6, 0, 0, 20, 46, 0, 0, 0, 17, 67, 29, 12, 26, 26, 23, 18, 14, 14, 18, 20, 21, 20, 19, 19, 19, 22, 25, 26, 29, 30, 29, 22, 7, 0, 5, 19, 49, 13, 0, 0, 0, 38, 102, 73, 42, 24, 24, 20, 13, 8, 10, 17, 22, 23, 22, 22, 22, 25, 31, 36, 34, 27, 19, 14, 8, 0, 21, 19, 48, 14, 13, 0, 0, 1, 99, 98, 55, 34, 34, 33, 26, 17, 12, 12, 14, 15, 15, 15, 17, 22, 28, 32, 28, 17, 3, 0, 0, 0, 6, 14, 48, 8, 13, 0, 0, 0, 32, 58, 32, 22, 27, 33, 35, 31, 25, 22, 17, 11, 5, 0, 1, 8, 11, 9, 10, 0, 0, 0, 1, 0, 0, 9, 68, 47, 42, 41, 40, 31, 34, 49, 36, 33, 36, 38, 42, 44, 43, 47, 49, 49, 47, 42, 39, 38, 35, 33, 41, 48, 47, 47, 43, 30, 25, 0, 41, 55, 43, 43, 43, 40, 33, 33, 24, 19, 20, 22, 23, 22, 22, 26, 36, 50, 62, 62, 54, 44, 40, 47, 65, 90, 93, 79, 52, 35, 37, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 49, 64, 43, 43, 38, 38, 42, 43, 41, 35, 41, 43, 34, 31, 34, 32, 29, 28, 31, 34, 34, 32, 35, 38, 41, 42, 41, 35, 0, 0, 0, 46, 57, 78, 54, 55, 47, 49, 55, 58, 53, 37, 48, 63, 41, 29, 36, 40, 41, 34, 38, 44, 43, 37, 36, 42, 48, 53, 53, 51, 4, 0, 0, 48, 59, 79, 54, 62, 55, 53, 58, 64, 53, 33, 51, 76, 42, 18, 30, 38, 38, 34, 36, 46, 40, 29, 29, 32, 44, 49, 55, 58, 18, 0, 0, 38, 55, 75, 49, 66, 67, 58, 58, 66, 55, 30, 48, 85, 52, 9, 11, 27, 34, 15, 11, 40, 34, 14, 8, 25, 40, 41, 44, 49, 25, 5, 0, 27, 43, 65, 41, 72, 79, 63, 56, 64, 59, 37, 52, 74, 51, 5, 2, 8, 13, 0, 0, 23, 26, 3, 2, 21, 32, 31, 39, 31, 15, 14, 0, 10, 29, 48, 15, 63, 86, 68, 53, 58, 66, 43, 27, 32, 38, 0, 0, 0, 14, 0, 0, 14, 52, 16, 5, 11, 31, 12, 24, 21, 0, 8, 9, 0, 29, 6, 10, 68, 89, 75, 49, 38, 66, 34, 6, 1, 29, 5, 0, 0, 31, 22, 0, 14, 77, 45, 9, 2, 18, 2, 0, 20, 0, 0, 18, 0, 32, 0, 27, 91, 95, 72, 37, 11, 76, 59, 0, 0, 31, 13, 0, 1, 30, 36, 0, 8, 69, 51, 6, 0, 0, 0, 0, 4, 0, 0, 13, 0, 15, 1, 48, 109, 104, 67, 28, 0, 50, 86, 7, 2, 45, 21, 0, 0, 8, 32, 0, 0, 53, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 59, 125, 107, 67, 20, 0, 20, 127, 61, 20, 61, 21, 0, 0, 0, 10, 0, 0, 36, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 70, 129, 107, 72, 37, 0, 18, 129, 97, 21, 66, 34, 0, 0, 0, 0, 0, 0, 41, 27, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 71, 113, 93, 73, 60, 0, 5, 111, 105, 40, 58, 46, 0, 0, 0, 0, 0, 0, 54, 32, 11, 7, 15, 8, 4, 2, 0, 0, 0, 0, 0, 0, 60, 99, 57, 58, 78, 26, 15, 86, 94, 70, 58, 60, 0, 15, 0, 0, 0, 0, 57, 29, 1, 0, 20, 19, 11, 21, 0, 0, 0, 0, 0, 0, 44, 82, 18, 23, 88, 61, 27, 46, 65, 86, 83, 73, 40, 54, 47, 0, 0, 5, 58, 30, 0, 0, 15, 26, 33, 60, 18, 8, 0, 0, 0, 0, 20, 72, 0, 4, 90, 87, 28, 8, 26, 86, 115, 87, 67, 85, 74, 33, 0, 22, 43, 39, 1, 1, 15, 38, 69, 96, 50, 18, 0, 0, 0, 0, 0, 63, 0, 0, 70, 110, 50, 2, 15, 82, 118, 88, 79, 81, 71, 67, 51, 41, 40, 49, 23, 11, 23, 47, 86, 111, 51, 9, 0, 0, 0, 0, 0, 49, 3, 0, 38, 112, 73, 25, 23, 79, 100, 67, 81, 58, 48, 65, 89, 60, 36, 44, 39, 14, 28, 51, 83, 105, 42, 1, 0, 0, 0, 0, 0, 30, 14, 0, 0, 89, 81, 36, 30, 47, 63, 23, 57, 33, 13, 39, 89, 57, 32, 36, 21, 4, 22, 52, 81, 103, 45, 7, 0, 0, 0, 36, 0, 20, 24, 0, 0, 50, 52, 0, 2, 16, 38, 1, 33, 30, 0, 16, 59, 55, 31, 12, 0, 0, 17, 50, 78, 103, 47, 11, 0, 0, 0, 68, 0, 26, 36, 0, 0, 0, 33, 0, 0, 5, 12, 0, 0, 20, 0, 0, 21, 15, 0, 0, 0, 0, 5, 39, 70, 87, 37, 6, 0, 0, 0, 58, 14, 46, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 37, 0, 0, 0, 0, 0, 8, 10, 63, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 35, 26, 26, 24, 22, 21, 20, 23, 23, 20, 20, 26, 28, 27, 23, 21, 20, 16, 13, 14, 18, 21, 22, 20, 17, 13, 9, 0, 0, 17, 27, 77, 81, 68, 69, 69, 63, 59, 58, 65, 63, 46, 51, 69, 69, 63, 58, 58, 54, 42, 30, 30, 40, 49, 55, 56, 52, 45, 34, 21, 0, 14, 21, 64, 76, 68, 72, 73, 66, 61, 61, 72, 66, 28, 33, 63, 69, 68, 66, 58, 40, 7, 0, 0, 0, 15, 31, 40, 48, 50, 37, 23, 0, 12, 34, 84, 104, 99, 98, 97, 90, 87, 92, 114, 116, 65, 54, 80, 89, 86, 75, 65, 46, 0, 0, 0, 0, 0, 3, 28, 53, 66, 60, 42, 0, 16, 34, 80, 108, 105, 97, 93, 89, 87, 95, 126, 133, 83, 41, 47, 47, 46, 35, 41, 45, 2, 0, 0, 0, 0, 0, 0, 24, 62, 67, 50, 0, 15, 17, 48, 92, 97, 84, 85, 88, 86, 82, 105, 110, 68, 5, 0, 0, 0, 1, 22, 45, 19, 0, 0, 0, 0, 0, 0, 0, 37, 73, 66, 0, 17, 0, 0, 51, 69, 59, 76, 89, 90, 61, 54, 65, 44, 0, 0, 0, 0, 0, 10, 55, 44, 0, 0, 0, 0, 0, 0, 0, 9, 69, 84, 0, 22, 0, 0, 20, 9, 21, 63, 89, 91, 38, 0, 29, 32, 0, 0, 0, 0, 0, 0, 53, 67, 0, 0, 0, 0, 0, 0, 0, 0, 44, 92, 1, 23, 0, 0, 0, 0, 0, 54, 89, 112, 61, 0, 17, 39, 0, 0, 0, 0, 0, 0, 42, 72, 0, 0, 0, 0, 0, 0, 0, 0, 12, 83, 18, 17, 0, 0, 8, 0, 0, 41, 92, 158, 147, 54, 50, 56, 0, 0, 0, 0, 0, 0, 33, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 11, 7, 0, 0, 15, 0, 0, 22, 84, 169, 193, 89, 45, 45, 0, 0, 0, 0, 0, 0, 34, 77, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 14, 0, 0, 15, 56, 134, 165, 88, 21, 46, 0, 0, 0, 0, 0, 0, 55, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 29, 28, 103, 142, 95, 49, 47, 7, 0, 0, 0, 0, 8, 72, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 15, 59, 108, 91, 64, 37, 11, 0, 0, 0, 0, 15, 76, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 35, 1, 10, 67, 89, 88, 52, 13, 0, 0, 0, 0, 7, 69, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 7, 0, 0, 27, 0, 0, 39, 93, 118, 75, 9, 0, 0, 0, 0, 4, 52, 60, 13, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 7, 11, 2, 19, 0, 0, 17, 7, 0, 1, 66, 89, 57, 0, 0, 0, 0, 0, 1, 24, 32, 14, 0, 0, 0, 0, 7, 10, 0, 0, 8, 0, 13, 27, 8, 22, 0, 0, 2, 12, 0, 0, 3, 35, 38, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 11, 18, 9, 17, 35, 0, 14, 47, 8, 9, 0, 0, 0, 12, 0, 0, 0, 0, 15, 7, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 8, 23, 28, 37, 43, 0, 9, 64, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 29, 27, 24, 25, 0, 0, 72, 8, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 17, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 32, 0, 0, 0, 0, 22, 13, 0, 0, 35, 50, 37, 54, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 69, 15, 0, 0, 0, 37, 42, 13, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 58, 30, 18, 0, 31, 35, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 29, 25, 25, 9, 47, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 7, 17, 13, 36, 82, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 12, 53, 114, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 103, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 57, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 56, 89, 101, 89, 62, 24, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 28, 49, 45, 31, 27, 61, 96, 121, 121, 96, 61, 18, 0, 0, 0, 3, 0, 4, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 60, 107, 129, 114, 51, 0, 0, 0, 0, 1, 50, 91, 82, 52, 6, 0, 0, 0, 36, 92, 89, 38, 0, 0, 0, 0, 27, 34, 0, 0, 0, 62, 119, 142, 141, 97, 10, 0, 0, 0, 0, 0, 0, 45, 92, 80, 39, 0, 0, 0, 68, 175, 179, 106, 34, 2, 0, 0, 32, 76, 82, 57, 13, 16, 55, 58, 53, 32, 0, 0, 0, 0, 0, 0, 0, 24, 100, 100, 73, 0, 0, 0, 12, 111, 148, 60, 23, 5, 0, 0, 0, 65, 109, 53, 0, 0, 0, 0, 0, 25, 1, 0, 0, 0, 0, 0, 0, 29, 96, 121, 91, 16, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 66, 75, 11, 0, 0, 3, 10, 2, 9, 55, 124, 114, 44, 25, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 92, 98, 28, 0, 0, 0, 0, 0, 0, 0, 87, 131, 72, 78, 51, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 90, 63, 0, 0, 0, 0, 0, 0, 0, 0, 27, 110, 88, 88, 64, 0, 0, 0, 0, 0, 0, 44, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 61, 62, 50, 0, 0, 0, 0, 0, 0, 6, 88, 49, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 13, 8, 0, 0, 0, 0, 0, 16, 23, 0, 0, 0, 0, 2, 0, 0, 68, 57, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 34, 8, 0, 32, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 33, 0, 0, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 0, 14, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 53, 26, 0, 0, 0, 11, 32, 0, 0, 0, 0, 0, 0, 50, 67, 65, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 84, 58, 24, 0, 0, 0, 33, 0, 0, 0, 0, 1, 58, 93, 95, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 107, 91, 42, 0, 0, 0, 0, 0, 0, 0, 24, 80, 119, 122, 113, 69, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 80, 94, 111, 106, 98, 83, 62, 44, 25, 37, 13, 15, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 53, 41, 32, 27, 22, 23, 21, 31, 49, 22, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 16, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 81, 111, 107, 76, 48, 22, 12, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 126, 107, 34, 0, 0, 0, 0, 0, 0, 0, 0, 28, 35, 28, 22, 13, 7, 8, 9, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 78, 60, 34, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 27, 61, 65, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 28, 73, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 40, 108, 46, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 0, 0, 39, 44, 0, 0, 1, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 3, 21, 18, 19, 18, 20, 20, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 21, 26, 35, 32, 34, 38, 33, 28, 36, 46, 46, 48, 50, 53, 57, 54, 45, 31, 17, 10, 14, 24, 35, 40, 21, 0, 0, 0, 14, 27, 35, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 18, 5, 0, 0, 34, 0, 0, 0, 0, 0, 95, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 21, 24, 0, 0, 21, 29, 0, 0, 0, 0, 96, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 81, 7, 0, 0, 0, 0, 0, 16, 63, 0, 0, 0, 22, 0, 0, 0, 0, 86, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 20, 89, 19, 0, 9, 0, 0, 0, 0, 89, 18, 0, 0, 0, 28, 0, 0, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 25, 92, 12, 16, 22, 0, 0, 0, 13, 104, 46, 0, 0, 0, 26, 3, 0, 0, 44, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 11, 0, 0, 15, 95, 0, 18, 39, 0, 0, 0, 61, 125, 59, 0, 0, 0, 0, 12, 0, 0, 22, 0, 0, 0, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 10, 98, 0, 11, 52, 0, 0, 0, 99, 119, 43, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 7, 115, 0, 0, 0, 0, 0, 0, 0, 0, 10, 86, 0, 12, 49, 0, 0, 0, 106, 102, 37, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 47, 156, 0, 0, 0, 0, 0, 0, 0, 0, 22, 35, 0, 14, 23, 0, 0, 0, 65, 75, 32, 0, 0, 0, 0, 0, 0, 0, 63, 0, 0, 0, 38, 201, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 9, 0, 0, 0, 0, 4, 61, 48, 0, 0, 0, 0, 0, 0, 0, 82, 0, 0, 0, 4, 218, 19, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 61, 53, 0, 0, 0, 0, 0, 0, 0, 98, 0, 0, 0, 0, 191, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 48, 0, 0, 0, 0, 0, 0, 0, 111, 0, 0, 0, 0, 144, 155, 0, 0, 1, 54, 0, 0, 0, 0, 0, 25, 55, 0, 0, 0, 0, 0, 35, 28, 0, 0, 0, 0, 0, 0, 0, 115, 0, 0, 0, 0, 105, 186, 0, 0, 0, 107, 56, 0, 0, 0, 0, 21, 106, 0, 0, 0, 6, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 122, 0, 0, 0, 0, 85, 190, 0, 0, 0, 97, 87, 0, 0, 0, 0, 18, 141, 26, 0, 0, 19, 26, 0, 0, 0, 0, 0, 0, 0, 0, 30, 120, 0, 0, 0, 0, 68, 154, 0, 0, 0, 128, 131, 1, 0, 0, 0, 16, 124, 84, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 110, 0, 0, 0, 0, 52, 85, 0, 0, 0, 188, 203, 53, 0, 0, 0, 41, 103, 86, 32, 3, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 50, 91, 0, 0, 0, 0, 23, 0, 0, 0, 38, 249, 222, 74, 0, 0, 0, 20, 47, 42, 19, 3, 0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 45, 89, 0, 0, 0, 0, 0, 0, 0, 0, 165, 243, 139, 44, 0, 2, 4, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 34, 99, 0, 2, 0, 0, 0, 0, 0, 10, 242, 177, 51, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 46, 122, 0, 0, 39, 6, 0, 0, 0, 93, 259, 123, 2, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 0, 0, 60, 131, 0, 0, 44, 38, 0, 0, 0, 116, 239, 83, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 9, 14, 58, 114, 0, 0, 31, 34, 23, 0, 0, 105, 194, 58, 0, 0, 0, 9, 12, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 27, 27, 55, 85, 0, 0, 34, 23, 38, 0, 0, 55, 118, 38, 0, 0, 0, 9, 16, 9, 0, 0, 0, 4, 20, 23, 16, 0, 0, 0, 0, 38, 67, 50, 57, 70, 0, 0, 34, 12, 27, 28, 4, 17, 46, 22, 1, 0, 0, 4, 9, 0, 0, 0, 0, 0, 21, 29, 20, 0, 0, 0, 0, 41, 69, 40, 43, 51, 0, 0, 21, 0, 0, 6, 0, 2, 14, 6, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 14, 15, 6, 0, 0, 0, 0, 38, 43, 13, 9, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 43, 0, 9, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 3, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 46, 0, 26, 15, 0, 0, 0, 0, 0, 12, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 76, 32, 0, 25, 20, 0, 0, 0, 0, 4, 27, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 0, 0, 0, 56, 0, 0, 18, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 16, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 37, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 32, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 0, 0, 26, 0, 0, 0, 17, 55, 22, 0, 0, 4, 0, 0, 0, 0, 0, 0, 29, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 32, 0, 67, 0, 0, 4, 52, 117, 122, 5, 0, 30, 0, 0, 0, 0, 0, 0, 36, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 63, 50, 91, 0, 0, 27, 61, 140, 171, 62, 18, 54, 0, 0, 0, 0, 0, 0, 70, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 117, 71, 69, 81, 0, 0, 27, 19, 77, 143, 70, 35, 46, 0, 0, 0, 0, 0, 6, 113, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 117, 66, 68, 70, 0, 0, 14, 0, 3, 80, 64, 57, 51, 0, 0, 0, 0, 0, 30, 130, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 123, 75, 56, 58, 0, 0, 2, 0, 0, 31, 75, 96, 69, 0, 0, 0, 0, 0, 37, 117, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 140, 96, 46, 54, 0, 0, 0, 0, 0, 8, 94, 124, 83, 3, 0, 0, 0, 0, 31, 62, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 162, 121, 41, 70, 0, 0, 0, 0, 0, 0, 91, 110, 67, 0, 0, 0, 0, 0, 20, 20, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 180, 147, 48, 84, 0, 0, 0, 23, 0, 0, 43, 70, 39, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 190, 173, 57, 81, 7, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 183, 188, 56, 67, 25, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 195, 56, 52, 18, 0, 0, 70, 30, 0, 0, 0, 0, 43, 53, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 159, 208, 83, 58, 15, 0, 0, 116, 100, 0, 0, 0, 49, 105, 115, 79, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 13, 0, 0, 0, 0, 162, 202, 133, 97, 35, 0, 44, 168, 144, 16, 0, 9, 101, 141, 136, 101, 41, 0, 0, 0, 0, 0, 0, 0, 7, 14, 10, 0, 0, 0, 0, 0, 162, 201, 159, 147, 77, 33, 109, 204, 123, 22, 0, 30, 82, 107, 97, 66, 27, 0, 0, 0, 0, 8, 18, 30, 39, 38, 32, 28, 22, 11, 21, 0, 125, 184, 155, 162, 130, 111, 182, 187, 47, 0, 0, 0, 2, 14, 14, 11, 7, 4, 6, 13, 24, 33, 37, 43, 49, 54, 55, 56, 56, 47, 55, 0, 79, 128, 115, 142, 156, 165, 232, 143, 0, 0, 0, 0, 10, 15, 16, 19, 20, 19, 20, 25, 34, 43, 49, 55, 61, 66, 70, 75, 79, 74, 79, 0, 77, 97, 72, 112, 158, 196, 259, 128, 0, 0, 0, 27, 37, 29, 24, 26, 28, 30, 33, 39, 46, 56, 67, 75, 74, 70, 70, 77, 87, 94, 97, 0, 84, 99, 46, 87, 149, 204, 253, 130, 0, 0, 14, 49, 51, 37, 25, 24, 30, 37, 43, 50, 57, 65, 72, 77, 74, 66, 63, 73, 90, 92, 85, 0, 87, 105, 49, 68, 132, 173, 197, 113, 0, 0, 27, 55, 63, 55, 44, 39, 41, 45, 49, 54, 55, 57, 62, 68, 72, 73, 76, 82, 81, 59, 40, 0, 99, 126, 72, 78, 100, 119, 114, 78, 21, 8, 35, 58, 70, 72, 66, 60, 66, 75, 80, 77, 68, 63, 66, 71, 90, 116, 124, 107, 78, 49, 33, 0, 95, 132, 96, 96, 93, 80, 68, 52, 29, 25, 43, 59, 68, 71, 72, 75, 87, 98, 108, 109, 94, 82, 77, 85, 116, 162, 170, 139, 98, 66, 48, 0, 86, 128, 109, 107, 104, 91, 77, 67, 59, 55, 61, 68, 72, 74, 77, 81, 88, 99, 108, 112, 102, 94, 96, 108, 132, 151, 153, 129, 99, 77, 63, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 40, 30, 29, 24, 19, 18, 19, 23, 31, 36, 34, 26, 24, 27, 23, 17, 12, 13, 21, 30, 31, 31, 29, 27, 24, 21, 21, 25, 37, 53, 6, 0, 72, 66, 68, 58, 53, 55, 55, 58, 60, 50, 40, 33, 36, 48, 49, 47, 52, 57, 65, 65, 63, 63, 70, 75, 71, 66, 61, 58, 72, 86, 23, 0, 60, 53, 59, 54, 52, 57, 59, 59, 54, 28, 9, 0, 8, 38, 59, 69, 78, 77, 57, 27, 11, 5, 17, 35, 51, 63, 72, 69, 79, 94, 28, 0, 58, 54, 62, 59, 57, 60, 63, 58, 56, 40, 37, 37, 41, 64, 87, 96, 88, 68, 34, 0, 0, 0, 0, 0, 8, 38, 66, 78, 84, 96, 28, 0, 80, 73, 90, 83, 68, 64, 64, 59, 56, 64, 85, 84, 69, 59, 51, 49, 47, 31, 0, 0, 0, 0, 0, 0, 0, 15, 41, 70, 90, 99, 30, 0, 76, 50, 67, 81, 73, 74, 74, 77, 76, 79, 89, 74, 50, 20, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 10, 29, 52, 87, 103, 34, 0, 13, 0, 0, 34, 56, 75, 79, 81, 80, 66, 46, 34, 20, 0, 0, 0, 0, 14, 17, 4, 0, 4, 0, 7, 14, 7, 12, 35, 74, 106, 36, 0, 0, 0, 0, 0, 28, 63, 62, 38, 0, 0, 0, 0, 0, 0, 0, 0, 14, 38, 47, 35, 6, 4, 0, 0, 9, 0, 0, 19, 53, 104, 45, 0, 0, 0, 0, 0, 10, 54, 55, 15, 0, 0, 0, 0, 0, 0, 0, 0, 20, 28, 29, 2, 0, 0, 0, 0, 0, 0, 0, 2, 26, 89, 60, 0, 0, 0, 0, 0, 0, 45, 62, 35, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 60, 49, 0, 0, 0, 0, 0, 0, 36, 66, 56, 47, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 16, 0, 0, 0, 0, 0, 3, 42, 52, 37, 63, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 22, 4, 0, 0, 0, 0, 0, 0, 49, 61, 41, 50, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 12, 0, 0, 0, 0, 0, 0, 30, 50, 34, 33, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 46, 21, 0, 0, 0, 0, 0, 0, 0, 26, 25, 21, 2, 0, 0, 0, 0, 1, 11, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 37, 69, 26, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 27, 27, 11, 21, 22, 32, 23, 3, 0, 15, 26, 11, 2, 0, 10, 24, 31, 27, 28, 45, 76, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 52, 50, 34, 18, 17, 0, 0, 0, 2, 23, 33, 38, 36, 34, 33, 33, 30, 27, 42, 77, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 15, 51, 37, 0, 0, 0, 0, 0, 0, 0, 24, 47, 48, 22, 14, 11, 10, 18, 42, 78, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 10, 8, 0, 0, 0, 0, 0, 0, 28, 47, 51, 35, 20, 7, 0, 0, 1, 19, 50, 80, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 33, 13, 0, 0, 0, 0, 0, 0, 13, 37, 57, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 88, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 115, 56, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 154, 98, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 185, 143, 79, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 190, 168, 104, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 169, 173, 116, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 131, 155, 111, 57, 0, 0, 0, 0, 0, 0, 0, 0, 24, 36, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 137, 99, 46, 0, 49, 104, 66, 0, 0, 4, 50, 106, 115, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 138, 100, 44, 13, 148, 254, 242, 162, 92, 81, 72, 70, 66, 46, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 114, 139, 128, 65, 59, 193, 268, 236, 134, 54, 14, 0, 0, 5, 11, 1, 0, 0, 0, 3, 21, 35, 46, 55, 61, 60, 48, 46, 10, 29, 0, 20, 105, 115, 101, 49, 94, 197, 209, 136, 37, 0, 0, 0, 2, 9, 13, 12, 10, 14, 25, 36, 46, 59, 77, 92, 96, 89, 79, 90, 53, 58, 0, 15, 90, 83, 54, 5, 97, 181, 169, 66, 2, 0, 21, 35, 34, 33, 32, 29, 27, 32, 43, 55, 69, 88, 107, 113, 104, 95, 101, 140, 104, 85, 0, 19, 73, 64, 36, 20, 125, 163, 123, 32, 0, 33, 59, 57, 49, 43, 40, 39, 42, 51, 65, 82, 99, 113, 118, 105, 90, 98, 135, 186, 144, 101, 0, 39, 73, 51, 46, 62, 144, 158, 105, 27, 21, 61, 74, 66, 57, 50, 47, 49, 56, 68, 82, 96, 110, 114, 100, 78, 78, 114, 158, 183, 127, 80, 8, 60, 94, 56, 55, 75, 123, 123, 83, 31, 34, 70, 83, 82, 73, 65, 62, 64, 72, 81, 90, 96, 100, 95, 83, 82, 108, 145, 158, 141, 75, 45, 34, 98, 137, 98, 80, 94, 120, 104, 70, 39, 52, 82, 101, 105, 97, 88, 90, 99, 112, 121, 123, 116, 108, 104, 113, 148, 188, 197, 165, 120, 57, 35, 61, 122, 161, 141, 119, 110, 116, 98, 70, 51, 65, 87, 105, 115, 115, 113, 114, 123, 143, 154, 149, 136, 124, 126, 153, 203, 245, 230, 183, 129, 65, 28, 91, 131, 153, 147, 138, 122, 111, 96, 78, 65, 69, 77, 82, 84, 84, 87, 99, 119, 142, 155, 151, 137, 127, 136, 168, 211, 228, 208, 168, 124, 67, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 4, 6, 0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 18, 56, 18, 0, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 22, 0, 0, 0, 0, 0, 0, 4, 0, 13, 61, 65, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 43, 14, 0, 0, 0, 0, 0, 17, 3, 0, 43, 77, 39, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 46, 39, 9, 0, 0, 0, 0, 26, 27, 0, 12, 63, 80, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 44, 58, 30, 0, 0, 0, 0, 44, 44, 0, 0, 47, 89, 62, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 41, 58, 44, 0, 0, 0, 0, 64, 49, 0, 0, 16, 68, 80, 13, 8, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 41, 38, 0, 0, 0, 0, 72, 51, 0, 0, 0, 29, 57, 36, 56, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 18, 0, 0, 0, 6, 71, 55, 3, 0, 0, 0, 11, 12, 63, 84, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 54, 13, 0, 0, 0, 0, 0, 35, 81, 0, 0, 0, 0, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 54, 4, 0, 0, 0, 0, 0, 0, 70, 0, 0, 0, 0, 102, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 41, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 111, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 38, 0, 0, 0, 0, 0, 0, 0, 67, 0, 0, 0, 0, 102, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 10, 29, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 76, 105, 0, 0, 0, 15, 13, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 6, 19, 8, 0, 0, 0, 0, 0, 0, 0, 78, 0, 0, 0, 0, 43, 91, 0, 0, 0, 42, 47, 0, 0, 0, 0, 0, 76, 41, 0, 0, 9, 44, 38, 15, 0, 0, 0, 0, 0, 0, 10, 87, 0, 0, 0, 0, 5, 45, 0, 0, 0, 58, 93, 27, 0, 0, 0, 0, 91, 90, 57, 32, 31, 47, 56, 57, 49, 23, 0, 0, 0, 0, 65, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 175, 110, 23, 0, 0, 31, 107, 126, 115, 95, 93, 103, 121, 132, 129, 113, 87, 70, 71, 86, 162, 151, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 222, 158, 85, 63, 51, 70, 116, 145, 152, 158, 163, 173, 181, 185, 183, 178, 173, 172, 173, 179, 235, 184, 0, 33, 10, 0, 0, 0, 0, 0, 64, 214, 222, 152, 122, 119, 123, 134, 153, 171, 181, 189, 194, 196, 196, 197, 201, 205, 206, 206, 205, 201, 253, 196, 42, 109, 93, 33, 0, 0, 0, 0, 167, 256, 203, 170, 172, 180, 183, 186, 192, 196, 197, 199, 202, 205, 206, 209, 215, 220, 218, 211, 207, 208, 258, 207, 74, 153, 157, 100, 0, 0, 0, 17, 238, 244, 199, 192, 201, 206, 205, 202, 201, 201, 202, 205, 211, 216, 219, 222, 225, 223, 216, 211, 218, 228, 274, 215, 91, 186, 193, 152, 68, 0, 0, 82, 250, 228, 204, 204, 205, 205, 206, 205, 203, 202, 204, 211, 218, 227, 232, 231, 224, 216, 211, 221, 243, 259, 286, 204, 93, 200, 221, 189, 133, 27, 0, 120, 227, 215, 208, 209, 209, 209, 208, 206, 203, 201, 204, 213, 224, 232, 235, 230, 218, 205, 212, 242, 270, 282, 280, 192, 99, 210, 240, 224, 180, 134, 90, 157, 205, 199, 203, 210, 215, 220, 221, 218, 211, 204, 205, 217, 232, 238, 237, 227, 210, 200, 218, 267, 294, 292, 272, 183, 120, 220, 260, 246, 221, 192, 175, 194, 207, 204, 206, 209, 212, 216, 217, 211, 208, 208, 211, 220, 235, 244, 240, 230, 214, 207, 225, 269, 297, 288, 260, 178, 89, 179, 207, 203, 193, 177, 166, 168, 172, 166, 164, 162, 163, 160, 154, 142, 132, 135, 149, 170, 188, 191, 178, 157, 139, 140, 180, 225, 243, 232, 210, 143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 31, 53, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 53, 24, 0, 0, 0, 55, 128, 105, 57, 47, 75, 129, 180, 209, 204, 165, 91, 38, 26, 0, 4, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 135, 218, 193, 152, 136, 134, 175, 226, 241, 230, 230, 246, 281, 325, 360, 373, 358, 321, 293, 288, 260, 223, 157, 0, 60, 70, 0, 0, 0, 0, 0, 1, 215, 289, 279, 257, 248, 240, 252, 293, 331, 352, 369, 394, 423, 448, 470, 484, 489, 484, 478, 477, 447, 374, 244, 100, 234, 218, 95, 0, 0, 0, 0, 81, 233, 267, 307, 325, 339, 340, 349, 373, 401, 422, 444, 468, 491, 507, 520, 539, 557, 566, 564, 564, 529, 448, 294, 182, 362, 360, 220, 42, 0, 0, 0, 156, 248, 312, 377, 417, 436, 436, 435, 444, 457, 469, 485, 507, 530, 548, 564, 583, 597, 599, 594, 599, 572, 498, 332, 231, 451, 469, 359, 150, 0, 0, 65, 234, 297, 375, 445, 483, 491, 483, 477, 477, 484, 497, 516, 542, 567, 587, 601, 610, 609, 601, 604, 631, 622, 536, 347, 252, 499, 558, 472, 304, 67, 0, 192, 302, 365, 420, 477, 502, 504, 495, 488, 488, 496, 513, 537, 564, 587, 603, 611, 608, 598, 595, 619, 659, 645, 529, 331, 254, 522, 609, 555, 444, 262, 188, 288, 370, 403, 444, 488, 511, 519, 512, 502, 496, 504, 522, 547, 573, 589, 594, 592, 586, 586, 611, 656, 678, 632, 498, 304, 251, 546, 639, 611, 538, 427, 342, 379, 415, 426, 448, 481, 508, 524, 526, 513, 504, 510, 530, 562, 591, 599, 592, 574, 561, 583, 645, 705, 705, 630, 490, 298, 235, 508, 595, 580, 540, 471, 405, 390, 404, 407, 411, 427, 444, 453, 453, 443, 438, 449, 476, 513, 541, 544, 531, 506, 489, 512, 584, 642, 645, 581, 464, 283, 171, 356, 407, 405, 387, 357, 318, 297, 292, 290, 285, 288, 291, 289, 279, 267, 265, 284, 319, 358, 381, 377, 357, 333, 319, 348, 406, 454, 454, 415, 335, 200, 12, 5, 70, 52, 59, 52, 48, 52, 51, 47, 41, 43, 52, 52, 49, 46, 44, 44, 41, 43, 53, 57, 55, 53, 53, 53, 49, 40, 27, 0, 0, 0, 16, 0, 66, 31, 45, 41, 39, 49, 49, 39, 23, 26, 47, 36, 23, 28, 31, 32, 27, 25, 28, 28, 16, 9, 15, 28, 42, 45, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 28, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 23, 0, 0, 0, 0, 0, 0, 18, 91, 100, 72, 38, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 138, 136, 104, 86, 83, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 157, 151, 80, 50, 61, 35, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 44, 38, 60, 0, 0, 0, 111, 148, 70, 9, 10, 6, 0, 0, 0, 0, 0, 0, 0, 141, 62, 110, 90, 0, 0, 0, 0, 87, 46, 0, 48, 84, 56, 49, 57, 0, 0, 0, 46, 118, 83, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 215, 166, 233, 165, 0, 0, 0, 34, 256, 226, 78, 88, 96, 36, 29, 32, 0, 0, 0, 55, 122, 107, 56, 4, 8, 2, 0, 0, 0, 0, 0, 0, 198, 182, 280, 190, 0, 0, 0, 0, 222, 255, 98, 90, 108, 21, 6, 18, 0, 0, 0, 125, 153, 118, 71, 24, 23, 21, 0, 0, 0, 0, 0, 0, 139, 145, 288, 185, 1, 0, 0, 0, 99, 182, 50, 79, 144, 44, 10, 21, 0, 0, 0, 165, 154, 95, 57, 21, 23, 28, 25, 0, 0, 0, 0, 0, 88, 118, 277, 138, 0, 0, 0, 0, 0, 100, 33, 103, 189, 103, 47, 52, 0, 0, 0, 172, 138, 73, 52, 32, 21, 26, 56, 34, 0, 0, 0, 0, 71, 98, 259, 86, 0, 0, 0, 0, 0, 67, 102, 165, 204, 140, 98, 93, 0, 0, 0, 163, 123, 75, 68, 63, 55, 66, 111, 84, 0, 0, 0, 0, 74, 65, 229, 92, 0, 0, 3, 0, 0, 55, 201, 266, 204, 133, 130, 114, 11, 0, 9, 137, 120, 89, 79, 70, 80, 112, 159, 101, 0, 0, 0, 0, 97, 28, 186, 146, 0, 10, 83, 0, 0, 0, 169, 270, 189, 108, 114, 101, 28, 0, 8, 95, 115, 108, 71, 40, 61, 114, 147, 69, 0, 0, 0, 0, 139, 8, 141, 188, 35, 38, 128, 39, 0, 0, 44, 156, 117, 80, 100, 77, 48, 21, 3, 1, 66, 97, 45, 0, 10, 63, 102, 24, 0, 0, 0, 0, 182, 19, 106, 189, 71, 25, 145, 126, 0, 0, 0, 63, 48, 62, 129, 82, 71, 98, 56, 0, 8, 32, 0, 0, 0, 27, 76, 10, 0, 0, 0, 0, 209, 54, 85, 174, 94, 0, 77, 148, 71, 0, 0, 0, 0, 44, 152, 98, 33, 110, 103, 24, 0, 0, 0, 0, 8, 47, 86, 18, 0, 0, 0, 0, 216, 97, 72, 163, 99, 0, 0, 104, 81, 10, 0, 0, 0, 51, 157, 129, 14, 27, 31, 0, 0, 0, 0, 0, 17, 52, 80, 13, 0, 0, 0, 0, 211, 138, 76, 150, 74, 0, 0, 105, 111, 57, 29, 59, 60, 92, 169, 153, 58, 0, 0, 0, 0, 0, 0, 0, 10, 27, 48, 0, 0, 0, 0, 0, 174, 175, 127, 164, 73, 0, 0, 125, 180, 126, 71, 61, 46, 37, 75, 89, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 59, 142, 176, 222, 126, 0, 5, 125, 133, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 7, 143, 219, 128, 16, 89, 110, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 29, 114, 35, 14, 116, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 10, 117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 55, 38, 44, 47, 46, 35, 31, 39, 43, 36, 33, 42, 60, 59, 44, 35, 32, 27, 17, 19, 33, 48, 54, 47, 35, 24, 16, 11, 0, 0, 0, 165, 183, 172, 184, 185, 185, 174, 166, 176, 171, 130, 100, 116, 169, 192, 179, 171, 171, 153, 113, 84, 98, 135, 166, 182, 178, 161, 137, 116, 65, 0, 0, 172, 213, 208, 219, 217, 219, 217, 214, 228, 221, 151, 70, 83, 180, 235, 238, 243, 230, 166, 70, 0, 0, 27, 84, 135, 177, 202, 188, 154, 90, 10, 0, 170, 228, 236, 238, 218, 214, 218, 222, 240, 253, 208, 97, 65, 154, 224, 240, 240, 215, 132, 9, 0, 0, 0, 0, 0, 79, 166, 207, 175, 92, 4, 0, 169, 237, 280, 278, 217, 203, 216, 222, 237, 272, 273, 180, 84, 99, 139, 145, 144, 148, 107, 0, 0, 0, 0, 0, 0, 0, 94, 202, 210, 109, 6, 0, 115, 170, 247, 281, 207, 195, 219, 220, 212, 239, 270, 210, 75, 0, 10, 25, 31, 61, 90, 18, 0, 0, 0, 0, 0, 0, 26, 163, 232, 146, 15, 0, 13, 30, 107, 166, 136, 168, 223, 206, 145, 130, 164, 131, 23, 0, 0, 0, 0, 19, 117, 96, 0, 0, 0, 0, 0, 0, 0, 95, 218, 193, 38, 0, 0, 0, 0, 2, 25, 122, 231, 195, 66, 0, 0, 22, 0, 0, 0, 0, 0, 14, 138, 148, 10, 0, 0, 0, 0, 0, 0, 15, 159, 208, 82, 0, 0, 0, 0, 0, 0, 76, 240, 246, 105, 0, 0, 0, 0, 0, 0, 0, 0, 20, 122, 140, 4, 0, 0, 0, 0, 0, 0, 0, 76, 172, 112, 12, 12, 0, 0, 0, 0, 36, 235, 345, 271, 34, 0, 0, 0, 0, 0, 0, 0, 14, 103, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 73, 1, 35, 0, 0, 0, 0, 11, 197, 350, 372, 189, 20, 0, 0, 0, 0, 0, 0, 5, 89, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 36, 138, 260, 363, 261, 80, 0, 0, 0, 0, 0, 0, 0, 91, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 84, 101, 168, 284, 243, 75, 0, 0, 0, 0, 0, 0, 0, 93, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 87, 77, 84, 188, 205, 83, 0, 0, 0, 0, 0, 0, 0, 97, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 18, 46, 3, 91, 189, 156, 33, 0, 0, 0, 0, 0, 0, 88, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 16, 0, 0, 146, 217, 145, 9, 0, 0, 0, 0, 0, 49, 75, 29, 0, 0, 0, 30, 70, 50, 8, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 34, 165, 154, 57, 0, 0, 0, 0, 0, 0, 11, 24, 0, 0, 2, 65, 100, 72, 26, 17, 11, 0, 0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 129, 81, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 32, 75, 89, 66, 33, 32, 29, 0, 0, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 44, 58, 53, 41, 46, 42, 0, 0, 148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 181, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 205, 124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 174, 157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 14, 39, 32, 31, 26, 25, 24, 22, 20, 22, 27, 32, 32, 29, 25, 24, 22, 24, 26, 29, 31, 33, 34, 32, 28, 23, 18, 11, 5, 0, 0, 41, 50, 69, 65, 66, 62, 63, 64, 58, 48, 46, 60, 66, 65, 66, 70, 69, 63, 53, 46, 42, 39, 42, 49, 57, 61, 60, 55, 45, 37, 11, 0, 35, 45, 58, 53, 56, 55, 59, 59, 52, 43, 52, 83, 93, 70, 66, 76, 72, 52, 30, 14, 7, 2, 0, 2, 10, 20, 33, 41, 39, 43, 25, 4, 36, 50, 61, 52, 53, 53, 53, 51, 43, 46, 78, 126, 141, 96, 61, 55, 44, 14, 0, 2, 11, 15, 9, 1, 0, 9, 10, 16, 29, 45, 33, 8, 41, 56, 57, 43, 50, 56, 52, 44, 31, 32, 71, 118, 120, 68, 23, 0, 0, 0, 0, 20, 38, 35, 28, 24, 14, 14, 8, 0, 14, 44, 44, 16, 31, 30, 6, 0, 25, 50, 52, 42, 30, 19, 42, 69, 52, 25, 0, 0, 0, 0, 6, 43, 51, 37, 29, 31, 24, 10, 0, 0, 0, 38, 49, 23, 24, 0, 0, 0, 13, 47, 46, 34, 25, 10, 0, 22, 36, 37, 10, 0, 0, 13, 18, 43, 55, 49, 28, 22, 14, 0, 0, 0, 0, 32, 49, 28, 32, 0, 0, 5, 53, 66, 43, 29, 39, 32, 4, 16, 63, 84, 45, 10, 7, 10, 0, 21, 48, 52, 32, 14, 0, 0, 0, 0, 0, 18, 36, 31, 51, 2, 37, 68, 99, 87, 51, 55, 109, 136, 95, 80, 117, 104, 52, 10, 0, 0, 0, 0, 38, 56, 41, 20, 3, 0, 0, 0, 0, 3, 15, 20, 50, 9, 82, 118, 124, 85, 44, 57, 129, 194, 187, 151, 145, 104, 49, 7, 0, 0, 0, 0, 67, 85, 68, 36, 17, 0, 0, 0, 0, 0, 1, 0, 40, 3, 86, 130, 148, 91, 33, 23, 82, 135, 172, 155, 147, 113, 63, 22, 0, 0, 0, 20, 94, 111, 80, 41, 17, 10, 0, 0, 0, 0, 0, 0, 30, 0, 73, 119, 152, 108, 43, 0, 28, 60, 86, 105, 137, 135, 97, 49, 7, 11, 0, 51, 101, 106, 62, 20, 8, 5, 0, 0, 0, 0, 0, 0, 22, 0, 68, 109, 127, 103, 52, 5, 0, 31, 34, 74, 139, 150, 134, 89, 42, 28, 0, 63, 102, 89, 40, 1, 0, 0, 0, 0, 0, 9, 0, 0, 24, 0, 75, 81, 83, 58, 49, 29, 0, 16, 33, 90, 154, 142, 130, 107, 68, 39, 0, 63, 98, 88, 38, 6, 2, 10, 16, 17, 20, 36, 14, 0, 33, 4, 80, 60, 49, 34, 53, 43, 6, 18, 57, 123, 161, 141, 104, 91, 71, 34, 0, 61, 99, 89, 40, 13, 7, 13, 29, 41, 46, 53, 30, 4, 39, 8, 83, 51, 32, 33, 65, 56, 35, 17, 57, 105, 131, 111, 72, 64, 49, 20, 11, 64, 86, 87, 58, 20, 6, 5, 17, 36, 43, 47, 34, 13, 45, 6, 78, 43, 23, 33, 65, 72, 59, 14, 29, 62, 66, 43, 30, 27, 18, 15, 13, 54, 63, 51, 48, 20, 0, 0, 0, 19, 34, 51, 49, 23, 50, 1, 65, 35, 10, 11, 41, 76, 70, 29, 27, 32, 32, 27, 24, 16, 18, 29, 48, 63, 53, 44, 27, 0, 0, 0, 0, 18, 45, 73, 64, 29, 50, 0, 54, 37, 10, 0, 1, 48, 47, 28, 13, 7, 10, 24, 44, 21, 15, 30, 58, 58, 52, 44, 0, 0, 0, 0, 13, 51, 73, 90, 71, 32, 45, 6, 50, 41, 15, 0, 0, 15, 7, 0, 0, 0, 0, 31, 70, 46, 13, 13, 37, 29, 0, 0, 0, 0, 0, 0, 19, 60, 73, 82, 60, 25, 40, 17, 56, 46, 9, 0, 0, 25, 22, 1, 0, 0, 36, 68, 104, 79, 43, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 22, 30, 10, 2, 39, 22, 61, 61, 13, 0, 0, 60, 79, 52, 14, 15, 33, 47, 58, 28, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 26, 55, 32, 20, 36, 109, 101, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 38, 66, 116, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 69, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 67, 60, 15, 0, 0, 0, 0, 0, 0, 0, 0, 98, 93, 76, 57, 35, 26, 23, 17, 0, 0, 0, 0, 0, 74, 87, 108, 142, 150, 133, 117, 145, 214, 289, 323, 294, 211, 106, 20, 0, 0, 0, 0, 42, 14, 0, 0, 0, 0, 8, 6, 0, 0, 0, 0, 0, 91, 212, 273, 264, 139, 0, 0, 0, 0, 0, 51, 165, 216, 168, 58, 0, 0, 0, 0, 151, 160, 101, 33, 0, 11, 27, 44, 79, 105, 107, 74, 103, 228, 343, 347, 241, 51, 0, 0, 0, 0, 0, 0, 0, 103, 189, 142, 16, 0, 0, 23, 270, 335, 274, 150, 49, 11, 6, 24, 115, 288, 392, 305, 139, 79, 93, 69, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 162, 78, 15, 0, 0, 109, 165, 171, 131, 73, 31, 0, 0, 48, 193, 255, 116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 40, 8, 0, 0, 50, 147, 127, 74, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 171, 136, 16, 0, 76, 86, 1, 0, 0, 105, 153, 138, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 147, 156, 108, 0, 0, 0, 0, 0, 0, 0, 22, 152, 212, 147, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 218, 203, 0, 0, 0, 0, 0, 0, 38, 261, 362, 275, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 137, 0, 57, 0, 0, 0, 0, 0, 221, 528, 670, 486, 148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 47, 31, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 132, 82, 0, 48, 288, 480, 393, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 43, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 128, 143, 58, 14, 102, 207, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 103, 183, 109, 18, 0, 0, 48, 117, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 172, 249, 282, 299, 292, 259, 172, 48, 14, 155, 258, 147, 0, 0, 5, 35, 54, 59, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 386, 658, 646, 435, 216, 150, 124, 12, 4, 202, 385, 344, 181, 74, 92, 131, 144, 97, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 187, 456, 441, 183, 0, 0, 0, 0, 0, 0, 171, 316, 321, 217, 104, 54, 17, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 163, 146, 0, 0, 0, 0, 0, 17, 0, 0, 140, 229, 155, 19, 0, 0, 0, 0, 0, 0, 5, 0, 136, 33, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 148, 298, 256, 160, 68, 0, 0, 0, 0, 0, 23, 49, 80, 54, 16, 164, 35, 2, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 184, 24, 0, 0, 0, 0, 0, 65, 124, 105, 91, 58, 40, 192, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 201, 298, 177, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 131, 382, 271, 58, 0, 0, 0, 0, 0, 0, 66, 178, 362, 587, 754, 748, 560, 259, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 132, 492, 552, 386, 135, 0, 0, 0, 236, 552, 544, 378, 293, 322, 362, 349, 264, 124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 209, 439, 556, 438, 99, 0, 44, 412, 561, 378, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 96, 357, 425, 201, 31, 147, 343, 350, 138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 58, 24, 0, 0, 0, 0, 0, 0, 0, 89, 242, 268, 256, 260, 227, 121, 16, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 11, 40, 72, 87, 64, 18, 10, 64, 154, 162, 0, 0, 0, 0, 79, 325, 561, 550, 296, 93, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 12, 49, 93, 118, 99, 32, 0, 0, 63, 206, 304, 255, 0, 0, 0, 0, 0, 232, 584, 693, 431, 180, 100, 97, 76, 34, 0, 0, 0, 0, 0, 0, 9, 52, 94, 101, 44, 0, 0, 0, 52, 167, 220, 181, 0, 10, 34, 29, 0, 50, 267, 397, 299, 152, 120, 158, 179, 175, 147, 98, 43, 0, 0, 0, 0, 32, 65, 49, 0, 0, 0, 0, 49, 102, 110, 95, 98, 228, 273, 267, 216, 175, 197, 224, 203, 164, 166, 214, 268, 310, 328, 321, 300, 271, 240, 221, 222, 231, 232, 223, 215, 229, 267, 312, 327, 293, 238, 154, 272, 476, 528, 500, 474, 430, 390, 358, 324, 295, 283, 296, 315, 331, 347, 375, 424, 489, 545, 571, 553, 505, 465, 473, 555, 684, 775, 758, 648, 520, 398, 231, 0, 63, 44, 35, 23, 20, 24, 23, 19, 19, 22, 23, 19, 18, 23, 27, 26, 25, 25, 28, 28, 26, 30, 38, 41, 37, 28, 21, 19, 26, 29, 19, 0, 56, 30, 29, 14, 10, 19, 19, 15, 15, 18, 11, 0, 0, 10, 30, 31, 23, 15, 11, 5, 0, 0, 3, 20, 31, 34, 35, 35, 46, 71, 22, 0, 70, 60, 61, 46, 38, 47, 51, 50, 57, 72, 67, 21, 0, 24, 61, 60, 48, 47, 57, 47, 15, 0, 0, 0, 18, 42, 63, 73, 83, 117, 37, 0, 90, 80, 83, 72, 60, 63, 64, 64, 70, 97, 112, 46, 0, 12, 49, 55, 59, 79, 103, 83, 34, 3, 0, 0, 0, 13, 51, 88, 106, 135, 43, 0, 69, 50, 74, 88, 77, 69, 63, 51, 32, 44, 83, 39, 0, 0, 24, 46, 52, 65, 92, 62, 14, 0, 0, 0, 0, 0, 13, 70, 111, 146, 45, 0, 41, 0, 28, 82, 88, 77, 68, 54, 21, 21, 66, 61, 21, 8, 18, 29, 32, 34, 54, 16, 0, 0, 0, 0, 0, 0, 0, 31, 101, 153, 52, 0, 29, 0, 0, 47, 68, 71, 68, 61, 32, 10, 45, 92, 72, 16, 0, 8, 8, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 73, 159, 62, 0, 20, 0, 0, 8, 35, 57, 82, 102, 62, 0, 0, 47, 46, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 15, 0, 0, 0, 24, 152, 75, 21, 24, 0, 0, 0, 0, 36, 104, 180, 128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 24, 17, 0, 0, 0, 106, 81, 0, 1, 0, 0, 0, 0, 0, 56, 150, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 59, 0, 0, 0, 0, 22, 37, 0, 0, 0, 49, 72, 0, 0, 0, 0, 0, 0, 0, 0, 19, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 32, 0, 0, 0, 0, 5, 42, 19, 0, 0, 24, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 38, 0, 0, 15, 29, 0, 0, 0, 0, 0, 0, 27, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 12, 0, 12, 11, 0, 0, 0, 0, 0, 0, 29, 41, 0, 10, 41, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 0, 0, 19, 10, 0, 0, 0, 0, 0, 0, 0, 46, 0, 7, 53, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 21, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 88, 30, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 41, 110, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 28, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 18, 33, 49, 116, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 60, 0, 0, 0, 0, 10, 3, 17, 34, 20, 4, 0, 1, 25, 42, 52, 117, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 34, 0, 0, 0, 0, 0, 0, 22, 33, 20, 1, 0, 0, 0, 25, 43, 107, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 30, 34, 38, 17, 0, 0, 0, 0, 14, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 49, 60, 55, 45, 14, 0, 0, 0, 0, 4, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 7, 0, 5, 8, 10, 13, 15, 18, 17, 13, 14, 16, 15, 13, 12, 15, 16, 9, 3, 1, 0, 0, 0, 0, 0, 7, 14, 21, 11, 38, 34, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 66, 35, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 17, 20, 7, 0, 0, 0, 0, 0, 19, 54, 77, 72, 45, 13, 0, 0, 0, 0, 0, 9, 66, 46, 0, 5, 3, 9, 12, 12, 26, 6, 0, 0, 0, 0, 20, 1, 0, 0, 2, 15, 37, 74, 107, 120, 124, 105, 62, 20, 0, 0, 0, 8, 62, 50, 0, 0, 0, 0, 9, 16, 37, 25, 0, 0, 0, 0, 36, 44, 53, 59, 36, 8, 0, 15, 42, 64, 90, 122, 118, 72, 13, 0, 0, 0, 65, 100, 38, 34, 0, 0, 6, 19, 39, 54, 0, 0, 0, 0, 63, 99, 117, 106, 58, 0, 0, 0, 0, 0, 5, 71, 118, 121, 63, 0, 0, 0, 62, 151, 129, 136, 62, 9, 11, 19, 35, 80, 74, 3, 0, 0, 64, 94, 104, 103, 43, 0, 0, 0, 0, 0, 0, 21, 105, 144, 114, 0, 0, 0, 43, 155, 149, 169, 108, 39, 21, 2, 14, 76, 118, 77, 12, 0, 11, 46, 65, 78, 46, 0, 0, 0, 0, 0, 0, 13, 92, 157, 153, 32, 0, 0, 0, 83, 91, 117, 67, 43, 38, 0, 0, 0, 59, 57, 3, 0, 0, 19, 57, 79, 72, 12, 0, 0, 0, 29, 12, 16, 73, 151, 171, 86, 0, 0, 0, 0, 0, 15, 0, 14, 55, 0, 0, 0, 0, 0, 0, 0, 0, 16, 69, 112, 106, 58, 0, 0, 0, 17, 6, 8, 33, 112, 173, 121, 46, 0, 0, 0, 0, 0, 0, 0, 66, 40, 0, 0, 0, 0, 0, 0, 0, 6, 74, 139, 118, 56, 0, 0, 0, 0, 0, 0, 0, 51, 138, 124, 91, 43, 0, 0, 0, 0, 0, 0, 31, 75, 0, 0, 0, 0, 0, 0, 0, 0, 49, 127, 108, 27, 0, 0, 0, 0, 0, 0, 0, 4, 83, 107, 90, 66, 0, 0, 0, 0, 0, 0, 0, 61, 31, 0, 0, 0, 0, 0, 0, 0, 0, 73, 66, 0, 0, 0, 0, 0, 26, 14, 0, 0, 38, 45, 61, 54, 0, 0, 0, 0, 0, 0, 0, 32, 50, 16, 0, 0, 0, 0, 0, 0, 0, 12, 15, 0, 0, 0, 0, 9, 32, 25, 0, 0, 0, 0, 11, 35, 0, 0, 0, 0, 3, 3, 17, 20, 53, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 3, 39, 26, 3, 45, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 42, 11, 0, 5, 57, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 17, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 23, 42, 0, 0, 0, 0, 30, 52, 16, 0, 0, 0, 0, 0, 0, 44, 66, 41, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 75, 49, 9, 0, 0, 45, 101, 48, 0, 0, 0, 0, 0, 47, 93, 101, 64, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 55, 118, 105, 86, 9, 0, 0, 62, 69, 29, 0, 0, 6, 66, 113, 148, 138, 83, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 136, 135, 103, 2, 0, 0, 0, 17, 53, 36, 36, 78, 125, 159, 179, 171, 122, 53, 15, 0, 2, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 45, 10, 0, 0, 0, 0, 0, 39, 102, 125, 143, 157, 171, 178, 178, 150, 109, 88, 73, 85, 74, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 96, 132, 143, 145, 142, 143, 143, 136, 123, 117, 112, 133, 114, 51, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 33, 19, 9, 14, 38, 68, 97, 116, 123, 119, 116, 117, 119, 117, 116, 119, 123, 148, 133, 54, 140, 46, 0, 0, 0, 0, 0, 0, 0, 0, 7, 84, 107, 107, 102, 99, 98, 102, 109, 114, 117, 118, 118, 116, 109, 102, 105, 115, 120, 144, 134, 54, 159, 139, 87, 1, 0, 0, 0, 0, 0, 0, 65, 102, 106, 99, 96, 99, 103, 110, 116, 119, 120, 119, 116, 107, 95, 90, 99, 111, 106, 110, 101, 39, 146, 142, 160, 131, 0, 0, 0, 0, 0, 26, 83, 99, 96, 93, 92, 95, 101, 107, 113, 113, 109, 103, 97, 92, 90, 97, 109, 109, 79, 57, 57, 30, 134, 133, 155, 183, 54, 0, 0, 0, 0, 48, 78, 86, 92, 96, 97, 97, 101, 105, 108, 105, 97, 88, 84, 89, 106, 127, 132, 109, 73, 49, 48, 26, 124, 119, 138, 169, 116, 0, 0, 0, 0, 52, 63, 64, 72, 79, 83, 90, 98, 104, 107, 104, 97, 88, 84, 96, 119, 140, 134, 112, 86, 78, 74, 3, 84, 71, 92, 108, 97, 41, 0, 0, 10, 45, 47, 37, 33, 36, 40, 44, 52, 63, 71, 74, 70, 65, 64, 63, 72, 78, 73, 67, 66, 81, 84, 0, 15, 0, 20, 33, 35, 24, 8, 11, 26, 38, 34, 23, 12, 3, 0, 0, 0, 0, 0, 0, 2, 11, 6, 0, 0, 0, 0, 0, 5, 35, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 15, 12, 1, 4, 4, 2, 3, 2, 0, 0, 3, 9, 12, 9, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 47, 35, 41, 40, 43, 39, 35, 34, 34, 38, 50, 65, 61, 48, 42, 35, 28, 20, 19, 26, 36, 39, 37, 35, 31, 28, 27, 25, 22, 5, 12, 0, 63, 62, 81, 79, 83, 75, 72, 72, 68, 58, 60, 95, 97, 67, 59, 59, 56, 59, 55, 58, 75, 83, 78, 73, 71, 67, 60, 54, 47, 26, 32, 0, 61, 48, 58, 54, 63, 59, 62, 66, 59, 27, 6, 59, 97, 61, 42, 58, 64, 56, 32, 17, 11, 17, 18, 27, 34, 31, 32, 34, 34, 20, 29, 0, 66, 58, 62, 54, 65, 64, 64, 69, 67, 38, 15, 65, 132, 116, 66, 64, 67, 39, 2, 0, 0, 0, 0, 0, 0, 11, 5, 11, 22, 21, 40, 0, 94, 88, 76, 51, 63, 72, 67, 69, 77, 57, 47, 81, 131, 124, 59, 24, 20, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 2, 7, 8, 50, 10, 100, 98, 80, 41, 56, 78, 74, 77, 103, 104, 79, 72, 73, 74, 32, 0, 0, 0, 0, 0, 16, 27, 0, 0, 0, 11, 13, 3, 3, 0, 44, 17, 58, 71, 47, 17, 50, 69, 67, 66, 90, 126, 85, 33, 28, 47, 26, 0, 0, 0, 0, 3, 46, 79, 48, 12, 0, 2, 19, 9, 3, 0, 26, 22, 19, 25, 0, 12, 67, 69, 43, 11, 19, 85, 73, 16, 23, 65, 48, 2, 0, 10, 19, 15, 53, 88, 63, 9, 0, 0, 0, 8, 6, 0, 12, 25, 16, 0, 0, 35, 91, 89, 39, 0, 0, 66, 77, 32, 49, 84, 60, 22, 8, 10, 14, 0, 18, 56, 40, 0, 0, 0, 0, 0, 11, 0, 5, 15, 27, 0, 0, 52, 107, 113, 69, 12, 16, 94, 131, 84, 77, 105, 70, 20, 16, 10, 0, 0, 15, 40, 25, 2, 0, 0, 0, 0, 5, 0, 0, 0, 38, 0, 14, 76, 110, 116, 104, 54, 17, 98, 147, 110, 73, 108, 72, 10, 6, 10, 0, 0, 30, 54, 40, 22, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 7, 83, 105, 101, 117, 79, 25, 59, 112, 83, 69, 92, 69, 13, 0, 13, 0, 0, 41, 64, 40, 18, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 84, 102, 78, 91, 99, 37, 17, 39, 41, 62, 72, 59, 29, 18, 26, 0, 0, 42, 56, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 54, 83, 44, 44, 99, 39, 0, 0, 10, 60, 64, 62, 56, 50, 49, 0, 0, 24, 42, 19, 0, 0, 0, 0, 0, 8, 7, 23, 0, 27, 0, 0, 11, 57, 15, 10, 81, 61, 0, 0, 45, 94, 87, 71, 57, 61, 64, 16, 4, 36, 48, 24, 0, 0, 0, 2, 25, 40, 29, 42, 0, 12, 0, 0, 0, 24, 0, 0, 51, 91, 43, 24, 73, 106, 110, 73, 56, 49, 48, 46, 44, 40, 48, 45, 24, 4, 12, 24, 42, 51, 30, 45, 1, 2, 0, 0, 0, 0, 0, 0, 17, 90, 68, 39, 43, 71, 69, 46, 53, 18, 1, 22, 44, 29, 25, 33, 42, 24, 17, 15, 27, 41, 25, 44, 9, 4, 0, 0, 0, 0, 0, 0, 11, 65, 86, 59, 44, 52, 38, 17, 42, 20, 0, 7, 42, 24, 9, 14, 35, 16, 2, 5, 21, 46, 32, 48, 16, 13, 0, 0, 0, 0, 0, 0, 0, 41, 59, 49, 24, 10, 0, 0, 0, 4, 0, 0, 23, 30, 15, 5, 0, 0, 0, 15, 43, 74, 54, 57, 26, 11, 0, 7, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 41, 8, 6, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 100, 28, 19, 2, 11, 19, 12, 3, 7, 26, 24, 0, 0, 13, 9, 0, 0, 4, 13, 9, 3, 11, 24, 27, 26, 18, 11, 5, 6, 0, 0, 59, 70, 0, 0, 0, 0, 0, 0, 0, 0, 26, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 9, 0, 0, 0, 0, 65, 77, 0, 10, 0, 0, 2, 0, 0, 2, 83, 70, 0, 0, 0, 0, 0, 0, 13, 59, 45, 17, 0, 0, 5, 8, 24, 46, 43, 15, 0, 0, 63, 62, 0, 33, 18, 0, 0, 0, 0, 15, 96, 87, 0, 0, 0, 0, 0, 0, 54, 104, 76, 28, 6, 16, 19, 0, 0, 37, 70, 47, 0, 0, 66, 25, 0, 50, 62, 19, 0, 0, 0, 7, 47, 51, 0, 0, 0, 0, 0, 0, 63, 131, 88, 5, 0, 17, 21, 0, 0, 4, 69, 77, 0, 0, 64, 0, 0, 47, 93, 36, 4, 5, 12, 0, 0, 20, 18, 0, 0, 0, 0, 0, 53, 140, 91, 0, 0, 6, 12, 0, 0, 0, 32, 90, 4, 0, 56, 0, 0, 44, 94, 27, 0, 23, 38, 0, 0, 0, 62, 0, 0, 0, 6, 13, 30, 126, 106, 0, 0, 0, 8, 0, 0, 0, 0, 67, 32, 0, 73, 0, 0, 87, 81, 0, 0, 48, 91, 4, 0, 0, 66, 0, 0, 0, 0, 0, 3, 104, 132, 5, 0, 0, 0, 5, 0, 0, 0, 18, 40, 0, 96, 12, 17, 136, 45, 0, 0, 54, 166, 64, 0, 0, 53, 0, 0, 0, 0, 0, 0, 118, 150, 18, 0, 0, 0, 26, 0, 0, 0, 0, 12, 0, 103, 49, 72, 135, 0, 0, 0, 4, 165, 114, 0, 0, 52, 0, 0, 0, 0, 0, 0, 139, 174, 7, 0, 0, 0, 44, 10, 0, 0, 0, 0, 0, 98, 63, 103, 128, 0, 0, 0, 0, 69, 118, 0, 6, 85, 0, 0, 0, 0, 0, 0, 167, 170, 0, 0, 0, 0, 59, 41, 0, 0, 0, 0, 0, 98, 79, 118, 107, 0, 0, 0, 0, 1, 106, 53, 81, 142, 5, 0, 0, 0, 0, 0, 176, 136, 0, 0, 0, 0, 56, 65, 30, 0, 0, 0, 0, 109, 97, 120, 67, 0, 0, 31, 0, 0, 83, 134, 167, 162, 21, 0, 0, 0, 0, 0, 171, 109, 0, 0, 0, 0, 57, 81, 67, 15, 0, 0, 0, 131, 110, 101, 34, 0, 0, 57, 0, 0, 64, 188, 216, 127, 0, 0, 0, 0, 0, 21, 162, 96, 0, 0, 0, 0, 59, 92, 84, 34, 3, 0, 0, 157, 125, 78, 30, 0, 0, 58, 48, 0, 42, 197, 203, 70, 0, 0, 17, 0, 0, 49, 137, 103, 0, 0, 0, 0, 48, 89, 76, 41, 33, 0, 0, 174, 139, 68, 51, 0, 0, 39, 101, 0, 15, 107, 120, 29, 0, 20, 35, 14, 55, 100, 86, 81, 35, 0, 0, 0, 27, 77, 76, 59, 59, 0, 0, 186, 152, 59, 70, 0, 0, 17, 123, 43, 3, 9, 41, 35, 22, 64, 40, 0, 64, 127, 61, 36, 28, 0, 0, 0, 24, 80, 103, 82, 65, 0, 0, 191, 171, 47, 78, 0, 0, 0, 137, 69, 0, 0, 10, 84, 98, 111, 41, 0, 10, 109, 77, 31, 0, 0, 0, 0, 35, 97, 128, 92, 51, 0, 0, 184, 191, 51, 83, 0, 0, 0, 133, 87, 0, 0, 0, 72, 144, 143, 38, 0, 0, 48, 49, 14, 0, 0, 0, 17, 58, 128, 140, 92, 40, 0, 0, 166, 210, 74, 88, 0, 0, 0, 151, 94, 0, 0, 0, 90, 177, 157, 36, 0, 0, 0, 0, 0, 0, 7, 16, 35, 84, 132, 142, 104, 55, 0, 0, 132, 203, 105, 91, 4, 0, 15, 201, 130, 0, 0, 0, 114, 174, 141, 46, 0, 0, 0, 4, 22, 29, 35, 52, 67, 91, 109, 114, 91, 59, 26, 0, 89, 169, 115, 101, 24, 0, 104, 258, 155, 0, 0, 0, 48, 95, 69, 32, 0, 0, 0, 20, 42, 55, 64, 70, 79, 92, 100, 105, 98, 81, 60, 0, 51, 99, 86, 107, 51, 21, 198, 281, 89, 0, 0, 0, 0, 26, 12, 15, 17, 20, 30, 45, 58, 65, 69, 74, 79, 81, 83, 86, 85, 82, 65, 0, 42, 50, 36, 72, 42, 93, 258, 228, 0, 0, 0, 0, 41, 48, 43, 45, 48, 50, 53, 59, 67, 71, 76, 84, 91, 90, 85, 88, 94, 91, 75, 0, 58, 65, 31, 24, 15, 147, 264, 116, 0, 0, 0, 33, 61, 59, 54, 54, 54, 55, 59, 67, 75, 81, 88, 95, 95, 86, 82, 92, 106, 105, 82, 0, 74, 88, 46, 20, 1, 140, 227, 40, 0, 0, 0, 57, 66, 57, 51, 52, 54, 59, 66, 73, 80, 85, 89, 90, 84, 78, 85, 108, 121, 105, 61, 0, 80, 97, 55, 45, 19, 91, 168, 18, 0, 0, 21, 64, 67, 60, 56, 56, 58, 64, 71, 78, 79, 79, 79, 76, 73, 80, 104, 127, 119, 75, 24, 0, 80, 101, 62, 62, 43, 55, 95, 10, 0, 0, 29, 57, 62, 59, 54, 55, 61, 71, 79, 83, 80, 72, 66, 65, 74, 98, 127, 131, 98, 50, 17, 0, 70, 87, 53, 66, 55, 45, 36, 14, 0, 0, 24, 39, 44, 41, 35, 38, 52, 66, 75, 77, 71, 60, 52, 55, 79, 110, 123, 102, 62, 31, 17, 0, 39, 34, 0, 19, 14, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 26, 25, 12, 3, 1, 6, 35, 64, 58, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 5, 0, 0, 0, 0, 3, 9, 0, 0, 125, 61, 9, 9, 0, 10, 14, 10, 7, 15, 20, 3, 0, 7, 15, 9, 3, 6, 20, 32, 34, 39, 50, 54, 48, 38, 29, 26, 27, 33, 0, 0, 115, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 13, 9, 21, 39, 44, 41, 31, 18, 9, 16, 0, 0, 102, 19, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 26, 40, 21, 5, 6, 24, 42, 47, 53, 51, 31, 23, 0, 0, 99, 17, 0, 5, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 10, 70, 80, 45, 16, 21, 34, 36, 31, 56, 85, 71, 41, 0, 0, 80, 1, 0, 53, 10, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 13, 39, 107, 100, 24, 0, 18, 55, 43, 13, 29, 85, 97, 73, 0, 0, 58, 0, 0, 83, 47, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 21, 57, 51, 107, 119, 17, 0, 0, 66, 57, 14, 6, 50, 103, 104, 0, 0, 66, 0, 0, 95, 56, 0, 0, 0, 0, 0, 0, 21, 35, 0, 0, 24, 70, 51, 89, 127, 38, 0, 0, 51, 73, 38, 9, 15, 76, 124, 14, 0, 110, 0, 0, 73, 17, 0, 0, 31, 0, 0, 0, 0, 32, 0, 0, 4, 52, 29, 62, 119, 60, 0, 0, 4, 79, 72, 27, 0, 30, 119, 56, 0, 134, 0, 0, 58, 0, 0, 0, 60, 56, 0, 0, 0, 0, 0, 0, 0, 18, 5, 49, 122, 58, 0, 0, 0, 72, 96, 51, 3, 0, 82, 78, 0, 128, 0, 0, 21, 0, 0, 0, 25, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 141, 51, 0, 0, 0, 64, 110, 66, 17, 0, 48, 69, 1, 115, 0, 11, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 151, 24, 0, 0, 0, 60, 120, 91, 49, 19, 39, 39, 6, 104, 0, 6, 0, 0, 0, 0, 0, 20, 38, 0, 0, 5, 0, 0, 0, 0, 0, 49, 142, 0, 0, 0, 0, 53, 118, 114, 71, 32, 48, 20, 0, 107, 0, 0, 0, 0, 0, 0, 0, 0, 65, 8, 0, 0, 0, 0, 0, 0, 0, 48, 127, 0, 0, 0, 0, 51, 106, 115, 84, 37, 52, 13, 0, 120, 0, 0, 0, 0, 0, 66, 0, 0, 69, 72, 1, 0, 0, 0, 0, 0, 0, 49, 113, 0, 0, 0, 0, 51, 103, 104, 82, 47, 60, 5, 0, 134, 0, 0, 0, 0, 0, 98, 0, 0, 54, 95, 20, 0, 0, 0, 10, 4, 0, 51, 91, 25, 0, 0, 0, 33, 98, 99, 71, 45, 61, 0, 0, 149, 0, 0, 0, 0, 0, 94, 39, 0, 0, 85, 39, 0, 0, 0, 22, 27, 43, 53, 60, 52, 1, 0, 0, 30, 91, 98, 67, 40, 59, 0, 0, 167, 0, 0, 0, 0, 0, 52, 90, 0, 0, 22, 46, 0, 0, 10, 0, 0, 81, 70, 4, 23, 35, 0, 0, 26, 82, 99, 71, 35, 50, 0, 0, 183, 0, 0, 0, 0, 0, 0, 113, 0, 0, 0, 54, 73, 60, 60, 0, 0, 51, 98, 14, 15, 41, 19, 8, 42, 89, 104, 76, 26, 30, 0, 0, 190, 0, 0, 0, 0, 0, 0, 116, 0, 0, 0, 24, 101, 91, 63, 0, 0, 0, 73, 45, 26, 33, 44, 49, 67, 99, 121, 88, 31, 31, 0, 0, 181, 17, 0, 0, 0, 0, 0, 128, 0, 0, 0, 0, 54, 75, 37, 0, 0, 0, 8, 40, 38, 48, 54, 50, 50, 72, 102, 92, 51, 49, 3, 0, 158, 50, 0, 0, 0, 0, 0, 135, 0, 0, 0, 0, 34, 59, 22, 0, 0, 0, 0, 39, 60, 70, 65, 45, 30, 33, 55, 61, 40, 47, 1, 0, 126, 68, 0, 0, 0, 0, 3, 103, 0, 0, 0, 0, 14, 33, 14, 0, 0, 0, 15, 49, 61, 58, 48, 39, 25, 11, 16, 31, 30, 32, 0, 0, 82, 45, 0, 0, 0, 0, 31, 25, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 21, 36, 40, 35, 27, 21, 13, 1, 0, 1, 3, 7, 0, 0, 66, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 3, 18, 26, 26, 28, 31, 29, 19, 11, 6, 2, 0, 0, 0, 0, 0, 0, 0, 98, 0, 0, 0, 0, 18, 19, 0, 0, 0, 0, 16, 15, 9, 12, 21, 24, 23, 23, 23, 18, 11, 4, 0, 0, 0, 0, 3, 0, 0, 0, 0, 133, 0, 0, 0, 0, 54, 40, 0, 0, 0, 0, 25, 13, 1, 5, 15, 20, 20, 20, 17, 12, 5, 2, 0, 0, 0, 0, 6, 0, 0, 0, 0, 145, 24, 0, 0, 0, 37, 69, 0, 0, 0, 15, 29, 12, 0, 0, 6, 16, 21, 20, 15, 7, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 149, 32, 0, 0, 0, 0, 66, 0, 0, 0, 27, 34, 22, 7, 0, 3, 10, 13, 12, 6, 0, 0, 0, 1, 11, 14, 1, 0, 0, 0, 0, 0, 152, 31, 0, 0, 0, 0, 16, 0, 0, 0, 24, 26, 19, 9, 1, 3, 11, 14, 6, 0, 0, 0, 0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 133, 27, 0, 0, 0, 0, 0, 15, 9, 7, 18, 22, 19, 14, 8, 12, 22, 24, 20, 3, 0, 0, 0, 0, 17, 19, 0, 0, 0, 0, 0, 0, 102, 46, 2, 29, 23, 18, 25, 34, 35, 31, 34, 35, 33, 31, 30, 34, 44, 49, 49, 36, 18, 15, 22, 30, 53, 63, 36, 2, 0, 10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 180, 145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 0, 11, 22, 0, 0, 0, 0, 0, 0, 0, 4, 55, 343, 287, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 77, 0, 0, 0, 40, 46, 25, 49, 87, 49, 0, 0, 0, 0, 0, 0, 0, 67, 405, 354, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 231, 27, 0, 0, 45, 18, 0, 32, 98, 76, 0, 0, 0, 0, 0, 0, 0, 52, 427, 373, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 321, 179, 30, 29, 35, 0, 0, 0, 92, 100, 32, 0, 0, 0, 0, 0, 0, 8, 450, 393, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 290, 287, 152, 35, 0, 0, 0, 0, 82, 134, 37, 0, 65, 71, 0, 0, 0, 0, 452, 415, 0, 167, 0, 0, 0, 0, 0, 0, 8, 27, 0, 0, 130, 293, 214, 16, 0, 0, 0, 0, 79, 217, 67, 0, 96, 164, 4, 0, 0, 0, 408, 439, 0, 215, 0, 0, 0, 0, 0, 0, 33, 187, 48, 0, 0, 264, 253, 25, 0, 0, 0, 0, 40, 285, 149, 0, 54, 163, 74, 0, 0, 0, 305, 443, 0, 230, 0, 0, 0, 0, 0, 0, 0, 308, 209, 0, 0, 249, 275, 61, 0, 0, 0, 0, 0, 296, 223, 29, 0, 95, 120, 0, 0, 0, 177, 401, 0, 170, 0, 0, 21, 0, 0, 0, 0, 278, 317, 0, 0, 286, 289, 93, 35, 0, 0, 0, 0, 274, 280, 80, 0, 21, 149, 94, 0, 0, 77, 304, 0, 62, 0, 0, 130, 47, 0, 0, 0, 109, 314, 0, 0, 349, 312, 117, 94, 0, 0, 0, 0, 294, 308, 101, 0, 0, 137, 162, 14, 0, 36, 192, 0, 0, 0, 0, 143, 20, 0, 0, 0, 0, 198, 0, 0, 375, 355, 134, 141, 3, 0, 0, 0, 361, 333, 106, 0, 0, 74, 157, 73, 0, 61, 123, 0, 0, 0, 0, 117, 0, 18, 0, 0, 0, 29, 0, 0, 321, 355, 144, 170, 28, 0, 0, 105, 421, 323, 90, 0, 0, 0, 79, 83, 1, 144, 134, 0, 0, 0, 141, 153, 0, 0, 119, 0, 0, 0, 0, 0, 228, 248, 125, 190, 42, 0, 0, 166, 430, 307, 88, 0, 0, 0, 0, 48, 15, 227, 204, 0, 0, 0, 259, 247, 0, 0, 139, 0, 0, 0, 0, 115, 214, 131, 69, 173, 26, 0, 0, 136, 390, 309, 97, 0, 0, 0, 0, 14, 0, 287, 281, 0, 0, 0, 277, 335, 0, 0, 87, 0, 0, 0, 0, 218, 238, 67, 31, 95, 0, 0, 0, 42, 292, 343, 143, 0, 0, 0, 0, 0, 0, 326, 345, 0, 10, 0, 212, 404, 0, 0, 0, 100, 0, 0, 0, 180, 196, 52, 43, 3, 0, 0, 0, 0, 146, 318, 166, 0, 0, 0, 0, 0, 0, 361, 395, 0, 56, 0, 120, 424, 87, 0, 0, 138, 0, 0, 0, 23, 78, 48, 108, 0, 0, 0, 31, 0, 82, 256, 131, 0, 0, 0, 0, 0, 0, 401, 430, 0, 74, 0, 48, 401, 202, 0, 0, 130, 149, 0, 0, 0, 0, 1, 203, 81, 0, 0, 57, 94, 130, 178, 48, 0, 0, 0, 0, 0, 0, 429, 436, 0, 47, 53, 7, 348, 267, 0, 0, 103, 223, 67, 0, 0, 0, 0, 271, 229, 0, 0, 51, 135, 143, 80, 0, 0, 0, 0, 0, 0, 30, 406, 386, 0, 0, 80, 3, 294, 260, 0, 0, 87, 343, 169, 0, 0, 0, 0, 266, 355, 97, 0, 43, 86, 67, 0, 0, 0, 0, 0, 0, 9, 39, 303, 267, 0, 0, 42, 7, 252, 183, 0, 0, 90, 479, 302, 0, 0, 0, 0, 188, 335, 191, 70, 25, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 160, 137, 0, 0, 0, 0, 182, 54, 0, 0, 153, 554, 396, 32, 0, 0, 0, 96, 188, 121, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 62, 0, 0, 0, 0, 19, 0, 0, 0, 341, 586, 370, 51, 0, 0, 0, 0, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 52, 0, 0, 0, 0, 0, 0, 0, 97, 544, 509, 228, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 82, 0, 0, 0, 0, 0, 0, 0, 389, 651, 356, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 122, 0, 0, 0, 0, 0, 0, 0, 543, 629, 226, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 131, 0, 0, 0, 0, 0, 0, 0, 489, 498, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 97, 0, 0, 0, 0, 0, 0, 0, 293, 286, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 49, 0, 0, 0, 0, 0, 0, 0, 105, 115, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 22, 44, 40, 0, 17, 2, 0, 0, 0, 0, 15, 38, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 0, 0, 0, 0, 0, 74, 95, 53, 56, 42, 0, 30, 1, 0, 0, 0, 0, 3, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 13, 0, 0, 0, 0, 0, 73, 69, 28, 43, 40, 20, 80, 104, 92, 86, 79, 79, 76, 70, 65, 68, 75, 79, 80, 82, 79, 74, 69, 67, 71, 74, 73, 76, 84, 88, 84, 73, 58, 43, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 65, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 65, 60, 0, 0, 0, 0, 54, 211, 196, 135, 65, 24, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 56, 88, 30, 0, 0, 0, 0, 82, 164, 135, 102, 56, 0, 0, 0, 0, 0, 0, 14, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 51, 17, 0, 0, 0, 0, 0, 11, 46, 79, 90, 41, 0, 0, 0, 0, 0, 44, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 42, 99, 83, 42, 0, 0, 0, 0, 41, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 18, 13, 0, 0, 0, 0, 0, 0, 0, 18, 62, 75, 65, 66, 36, 0, 0, 0, 40, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 46, 38, 0, 0, 0, 0, 0, 0, 0, 87, 129, 85, 28, 23, 8, 0, 0, 0, 42, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 62, 56, 0, 0, 0, 0, 0, 0, 0, 26, 89, 34, 0, 0, 0, 0, 0, 0, 0, 35, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 82, 69, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 106, 75, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 114, 80, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 98, 72, 47, 2, 0, 0, 0, 0, 0, 0, 0, 0, 16, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 88, 72, 36, 0, 0, 24, 91, 51, 0, 0, 0, 26, 107, 130, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 97, 60, 4, 12, 95, 193, 170, 84, 19, 14, 29, 42, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 95, 111, 86, 102, 141, 171, 107, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 87, 105, 130, 140, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 93, 97, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 34, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 20, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 36, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 39, 0, 0, 0, 0, 0, 0, 0, 0, 78, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 60, 77, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 53, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 78, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 21, 5, 0, 0, 0, 0, 10, 21, 26, 28, 26, 19, 14, 7, 0, 11, 20, 0, 83, 129, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 37, 45, 35, 24, 18, 24, 31, 38, 40, 44, 48, 53, 55, 50, 43, 38, 41, 41, 4, 73, 126, 89, 63, 0, 0, 0, 0, 0, 0, 0, 19, 37, 45, 46, 45, 39, 36, 39, 46, 53, 58, 63, 68, 69, 66, 63, 61, 63, 66, 64, 8, 52, 102, 81, 88, 64, 0, 13, 2, 0, 0, 13, 41, 45, 40, 39, 41, 43, 47, 53, 60, 65, 69, 73, 74, 71, 64, 62, 67, 75, 80, 74, 0, 55, 80, 64, 83, 106, 100, 92, 5, 0, 0, 41, 50, 49, 48, 47, 48, 50, 54, 60, 65, 69, 72, 73, 72, 69, 67, 72, 80, 84, 80, 66, 0, 58, 89, 59, 78, 102, 143, 138, 30, 0, 0, 49, 51, 52, 54, 53, 52, 52, 55, 60, 66, 70, 73, 72, 69, 67, 73, 84, 89, 82, 68, 51, 0, 59, 94, 69, 70, 85, 123, 121, 47, 0, 16, 51, 54, 53, 51, 53, 54, 58, 62, 65, 67, 69, 70, 70, 66, 69, 82, 91, 90, 76, 63, 50, 6, 65, 102, 75, 80, 76, 99, 91, 51, 17, 45, 62, 68, 65, 59, 57, 58, 57, 60, 65, 71, 73, 71, 72, 75, 77, 86, 93, 86, 71, 60, 50, 6, 70, 93, 69, 73, 62, 56, 54, 42, 27, 42, 57, 68, 69, 65, 65, 68, 70, 70, 64, 55, 48, 49, 61, 76, 86, 88, 68, 44, 29, 35, 35, 0, 35, 50, 48, 44, 40, 35, 30, 26, 23, 26, 33, 39, 39, 38, 36, 38, 41, 40, 38, 35, 31, 29, 33, 37, 45, 47, 39, 30, 25, 30, 25, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 40, 51, 0, 0, 0, 17, 15, 12, 25, 30, 0, 0, 0, 0, 0, 0, 0, 8, 17, 23, 6, 0, 0, 7, 0, 25, 10, 0, 0, 0, 0, 0, 54, 102, 30, 0, 0, 0, 0, 0, 18, 48, 3, 0, 0, 0, 0, 0, 0, 0, 18, 48, 23, 0, 0, 0, 0, 17, 26, 0, 0, 0, 0, 0, 12, 67, 52, 0, 0, 0, 0, 0, 0, 58, 11, 0, 0, 0, 0, 0, 0, 0, 0, 65, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 48, 0, 0, 0, 0, 0, 0, 65, 39, 0, 0, 0, 0, 0, 0, 0, 0, 56, 80, 0, 9, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 53, 76, 0, 0, 0, 0, 0, 0, 0, 0, 30, 90, 19, 48, 0, 0, 0, 0, 0, 0, 29, 84, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 49, 67, 0, 0, 0, 0, 0, 0, 30, 175, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 49, 60, 0, 0, 10, 0, 0, 0, 0, 179, 220, 50, 0, 28, 0, 0, 0, 0, 0, 0, 32, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 45, 0, 16, 27, 0, 0, 0, 0, 73, 184, 84, 26, 76, 5, 0, 0, 0, 0, 0, 58, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 1, 18, 6, 0, 0, 0, 0, 0, 103, 73, 42, 77, 35, 0, 0, 0, 0, 0, 81, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 17, 29, 0, 0, 0, 11, 0, 0, 37, 76, 73, 67, 16, 0, 0, 0, 0, 0, 90, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 34, 33, 0, 0, 0, 0, 0, 0, 0, 97, 129, 60, 0, 0, 11, 0, 0, 0, 81, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 51, 27, 0, 0, 0, 0, 0, 0, 0, 105, 174, 96, 0, 0, 10, 0, 0, 0, 44, 80, 47, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 102, 68, 16, 0, 0, 0, 0, 15, 0, 0, 33, 126, 103, 26, 0, 0, 0, 0, 0, 0, 40, 75, 8, 0, 0, 0, 0, 0, 0, 0, 2, 0, 117, 88, 8, 11, 0, 0, 0, 23, 0, 0, 0, 23, 55, 23, 0, 0, 0, 0, 7, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 111, 115, 9, 20, 0, 0, 0, 15, 0, 0, 0, 0, 13, 27, 26, 0, 0, 0, 12, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 90, 142, 15, 20, 0, 0, 0, 20, 0, 0, 0, 0, 0, 24, 44, 0, 0, 0, 0, 17, 24, 0, 0, 0, 0, 0, 0, 0, 0, 16, 34, 0, 79, 165, 31, 14, 0, 0, 0, 49, 0, 0, 0, 0, 0, 37, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 15, 0, 72, 186, 70, 31, 0, 0, 0, 67, 20, 0, 0, 0, 0, 85, 117, 78, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 165, 124, 85, 0, 0, 0, 97, 50, 0, 0, 0, 4, 47, 72, 72, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 61, 90, 132, 38, 0, 63, 113, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 59, 54, 67, 135, 109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 125, 201, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 243, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 191, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 2, 0, 0, 1, 1, 2, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 19, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 55, 47, 29, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 43, 62, 64, 69, 68, 49, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 30, 19, 15, 18, 43, 62, 68, 43, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 46, 45, 29, 27, 0, 0, 0, 10, 36, 54, 56, 23, 4, 0, 0, 0, 0, 6, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 51, 60, 28, 6, 0, 0, 0, 0, 31, 60, 74, 42, 4, 0, 0, 0, 0, 0, 0, 23, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 54, 20, 2, 0, 0, 0, 0, 26, 69, 87, 75, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 36, 13, 24, 0, 0, 0, 0, 16, 64, 85, 99, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 21, 0, 0, 0, 0, 0, 49, 69, 91, 82, 29, 18, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 37, 62, 79, 89, 69, 52, 33, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 49, 71, 84, 88, 85, 72, 47, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 63, 84, 92, 80, 67, 59, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 61, 71, 67, 49, 40, 43, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 8, 37, 36, 35, 23, 29, 38, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 33, 22, 0, 0, 0, 0, 0, 0, 14, 14, 22, 26, 28, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 40, 34, 35, 46, 15, 2, 3, 0, 0, 0, 16, 26, 40, 35, 17, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 2, 46, 44, 19, 0, 25, 29, 33, 24, 17, 29, 33, 34, 40, 46, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 33, 43, 13, 0, 0, 0, 10, 25, 36, 52, 65, 61, 59, 58, 46, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 51, 19, 0, 0, 0, 0, 16, 39, 68, 88, 94, 93, 86, 77, 66, 53, 43, 41, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 64, 98, 118, 129, 131, 121, 109, 90, 91, 94, 96, 94, 69, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 86, 118, 128, 125, 118, 106, 96, 93, 98, 107, 116, 111, 81, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 16, 40, 63, 89, 104, 107, 103, 97, 92, 87, 82, 81, 85, 94, 91, 65, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 75, 74, 70, 76, 86, 96, 102, 104, 100, 94, 90, 86, 82, 77, 74, 77, 84, 78, 50, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 89, 91, 89, 87, 90, 94, 97, 99, 98, 94, 91, 85, 78, 70, 67, 69, 74, 75, 57, 27, 0, 14, 26, 7, 0, 0, 0, 0, 0, 0, 1, 76, 91, 87, 86, 88, 90, 91, 92, 92, 90, 86, 80, 72, 66, 63, 67, 75, 75, 64, 31, 2, 0, 14, 51, 47, 0, 0, 0, 0, 0, 0, 35, 83, 85, 79, 82, 86, 88, 88, 87, 86, 84, 79, 73, 67, 64, 68, 78, 85, 77, 54, 28, 8, 0, 12, 50, 64, 39, 0, 0, 0, 0, 0, 56, 78, 71, 68, 72, 76, 79, 80, 80, 80, 80, 80, 76, 72, 71, 76, 81, 80, 70, 62, 58, 39, 17, 4, 28, 47, 53, 8, 0, 0, 4, 34, 59, 65, 53, 48, 48, 52, 55, 55, 55, 58, 60, 64, 66, 66, 62, 58, 46, 38, 43, 58, 70, 52, 28, 0, 0, 4, 23, 10, 0, 0, 24, 47, 43, 34, 20, 15, 11, 6, 0, 0, 0, 0, 8, 21, 28, 25, 8, 0, 0, 0, 0, 28, 47, 44, 19, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 7, 62, 85, 80, 81, 74, 73, 72, 69, 65, 65, 72, 79, 78, 74, 70, 65, 62, 59, 60, 64, 65, 66, 67, 69, 67, 62, 50, 34, 0, 0, 0, 0, 34, 45, 44, 54, 49, 49, 50, 48, 39, 30, 40, 50, 35, 35, 43, 44, 38, 23, 5, 0, 0, 0, 0, 9, 20, 30, 29, 15, 0, 0, 0, 0, 14, 39, 42, 57, 49, 48, 54, 58, 52, 40, 79, 106, 62, 41, 49, 45, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 14, 0, 0, 0, 14, 34, 59, 58, 73, 61, 51, 55, 70, 74, 60, 120, 167, 98, 34, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 34, 45, 30, 59, 61, 49, 49, 67, 63, 16, 42, 93, 36, 0, 0, 0, 0, 0, 0, 13, 39, 31, 15, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 48, 47, 47, 55, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 53, 27, 8, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 38, 29, 21, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 27, 64, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 0, 30, 59, 44, 18, 5, 17, 0, 0, 0, 16, 10, 0, 0, 6, 0, 0, 0, 44, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 88, 76, 119, 103, 74, 46, 62, 151, 171, 79, 26, 42, 13, 0, 0, 0, 0, 0, 0, 36, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 117, 126, 180, 130, 95, 44, 40, 203, 296, 174, 79, 74, 18, 0, 0, 0, 0, 0, 0, 74, 62, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 92, 140, 212, 144, 102, 19, 0, 77, 244, 164, 88, 103, 36, 0, 0, 0, 0, 0, 22, 111, 69, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 56, 138, 220, 126, 89, 35, 0, 0, 170, 131, 80, 136, 89, 0, 0, 19, 7, 0, 40, 104, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 36, 125, 191, 76, 57, 69, 0, 0, 94, 98, 75, 155, 151, 38, 11, 63, 14, 0, 44, 104, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 33, 116, 156, 35, 6, 70, 0, 0, 51, 100, 114, 168, 156, 64, 54, 95, 13, 0, 56, 106, 27, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 67, 31, 117, 152, 28, 0, 70, 45, 7, 35, 116, 186, 189, 131, 47, 50, 91, 25, 0, 55, 101, 36, 0, 0, 0, 0, 17, 48, 0, 0, 0, 0, 79, 47, 106, 159, 49, 0, 65, 92, 21, 0, 33, 130, 134, 58, 11, 31, 60, 29, 0, 21, 52, 41, 17, 0, 0, 0, 6, 39, 0, 0, 0, 0, 100, 83, 79, 148, 58, 0, 56, 118, 31, 0, 0, 19, 49, 0, 0, 9, 31, 25, 0, 0, 0, 3, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 110, 118, 57, 128, 72, 0, 26, 115, 65, 0, 0, 0, 23, 0, 8, 29, 10, 26, 39, 0, 0, 0, 0, 0, 0, 0, 14, 61, 0, 0, 0, 0, 92, 138, 54, 104, 91, 0, 0, 49, 36, 0, 0, 0, 0, 0, 31, 46, 0, 5, 47, 8, 0, 0, 0, 0, 0, 7, 44, 76, 0, 0, 0, 0, 54, 146, 62, 84, 104, 0, 0, 13, 20, 0, 0, 0, 0, 6, 83, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 48, 0, 0, 0, 0, 21, 157, 78, 72, 100, 0, 0, 52, 109, 58, 26, 58, 99, 96, 146, 147, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 164, 112, 104, 140, 37, 17, 127, 195, 119, 59, 54, 47, 20, 34, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 101, 168, 227, 117, 80, 142, 161, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 152, 210, 120, 96, 115, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 118, 82, 82, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 23, 95, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 30, 37, 39, 39, 41, 43, 43, 42, 38, 33, 32, 34, 41, 45, 42, 35, 29, 24, 16, 8, 6, 12, 23, 33, 39, 45, 58, 78, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 47, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 30, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 32, 47, 35, 0, 0, 0, 0, 0, 0, 25, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 4, 33, 48, 42, 11, 0, 0, 0, 0, 16, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 46, 27, 5, 0, 0, 0, 0, 0, 0, 0, 12, 33, 11, 0, 0, 0, 7, 36, 39, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 58, 53, 22, 0, 0, 0, 0, 0, 0, 0, 0, 22, 41, 0, 0, 0, 0, 23, 42, 51, 86, 13, 0, 0, 0, 0, 27, 62, 58, 22, 0, 0, 32, 39, 11, 0, 0, 0, 0, 0, 23, 11, 0, 25, 56, 38, 0, 0, 0, 7, 11, 26, 78, 23, 0, 0, 0, 0, 0, 18, 58, 32, 0, 0, 30, 41, 17, 0, 0, 0, 0, 0, 36, 46, 24, 22, 58, 69, 14, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 10, 0, 1, 36, 58, 50, 25, 4, 0, 0, 0, 23, 45, 27, 11, 31, 74, 61, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 47, 67, 71, 61, 17, 0, 0, 0, 5, 17, 5, 0, 4, 51, 82, 69, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 71, 64, 62, 8, 0, 0, 0, 5, 18, 3, 0, 0, 15, 59, 79, 67, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 31, 34, 0, 0, 0, 0, 21, 36, 25, 0, 0, 0, 17, 48, 68, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 21, 35, 25, 0, 0, 0, 0, 16, 51, 55, 0, 0, 0, 0, 39, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 0, 0, 0, 0, 0, 3, 41, 51, 0, 0, 0, 0, 38, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 36, 49, 0, 0, 0, 0, 3, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 27, 45, 0, 0, 0, 0, 0, 50, 5, 0, 0, 15, 0, 0, 0, 0, 3, 19, 6, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 20, 40, 0, 0, 0, 0, 0, 28, 39, 0, 0, 41, 38, 0, 0, 0, 0, 34, 60, 0, 0, 0, 0, 0, 0, 13, 19, 0, 0, 0, 0, 0, 10, 33, 0, 0, 0, 0, 0, 0, 57, 14, 19, 80, 112, 70, 0, 0, 0, 0, 68, 64, 0, 0, 0, 30, 49, 58, 37, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 39, 13, 19, 91, 132, 84, 0, 0, 0, 0, 0, 64, 46, 19, 30, 58, 82, 74, 46, 10, 0, 0, 0, 0, 3, 25, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 26, 11, 0, 0, 0, 0, 0, 0, 51, 72, 74, 61, 58, 55, 49, 38, 20, 7, 7, 36, 29, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 34, 43, 36, 25, 15, 14, 18, 23, 23, 24, 47, 36, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 15, 0, 0, 0, 0, 1, 12, 11, 7, 3, 1, 0, 0, 0, 0, 0, 0, 17, 8, 28, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 37, 32, 22, 20, 13, 5, 7, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 36, 0, 0, 0, 0, 0, 0, 0, 0, 28, 23, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 20, 0, 0, 0, 0, 0, 0, 32, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 46, 0, 0, 0, 0, 0, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 44, 0, 0, 0, 0, 120, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 10, 0, 0, 0, 0, 0, 0, 14, 0, 0, 29, 69, 14, 0, 0, 0, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 23, 9, 0, 0, 0, 0, 0, 38, 10, 0, 0, 72, 70, 0, 0, 0, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 27, 35, 4, 0, 0, 0, 0, 50, 17, 0, 0, 44, 91, 37, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 22, 46, 22, 0, 0, 0, 0, 63, 22, 0, 0, 3, 69, 58, 0, 7, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 1, 36, 18, 0, 0, 0, 23, 67, 17, 0, 0, 0, 6, 41, 10, 42, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 34, 71, 32, 0, 0, 0, 0, 0, 0, 52, 103, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 61, 32, 0, 0, 0, 0, 0, 0, 36, 117, 0, 0, 0, 17, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 42, 0, 0, 0, 0, 0, 0, 10, 116, 0, 0, 0, 8, 131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 38, 0, 0, 0, 0, 0, 0, 0, 117, 0, 0, 0, 0, 139, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 30, 0, 0, 0, 0, 0, 0, 0, 119, 0, 0, 0, 0, 118, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 35, 0, 0, 0, 0, 0, 0, 0, 120, 0, 0, 0, 0, 87, 130, 0, 0, 0, 28, 2, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 42, 51, 36, 0, 0, 0, 0, 0, 0, 14, 120, 0, 0, 0, 0, 63, 121, 0, 0, 0, 65, 55, 0, 0, 0, 0, 22, 118, 46, 0, 19, 52, 72, 78, 60, 18, 0, 0, 0, 0, 0, 52, 122, 0, 0, 0, 0, 34, 64, 0, 0, 0, 115, 134, 6, 0, 0, 0, 31, 143, 117, 74, 78, 83, 99, 109, 108, 86, 37, 0, 0, 0, 28, 82, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 182, 209, 76, 0, 0, 8, 68, 137, 149, 134, 130, 129, 140, 152, 156, 146, 124, 99, 88, 96, 115, 137, 137, 1, 0, 0, 0, 0, 0, 0, 0, 4, 216, 235, 137, 97, 89, 90, 104, 128, 153, 162, 167, 171, 173, 175, 178, 179, 179, 176, 176, 180, 176, 176, 157, 69, 68, 3, 0, 0, 0, 0, 0, 129, 242, 209, 162, 148, 150, 146, 150, 162, 171, 177, 184, 187, 190, 191, 192, 197, 203, 205, 203, 201, 189, 192, 178, 109, 143, 95, 21, 0, 0, 0, 0, 232, 245, 187, 179, 178, 180, 177, 177, 182, 187, 191, 194, 197, 201, 202, 205, 208, 212, 210, 203, 202, 194, 205, 195, 132, 182, 157, 104, 0, 0, 0, 88, 284, 236, 188, 189, 193, 194, 191, 189, 189, 192, 195, 199, 204, 206, 207, 210, 213, 213, 206, 201, 208, 209, 211, 197, 137, 206, 193, 164, 54, 0, 0, 151, 286, 217, 194, 194, 196, 199, 198, 194, 190, 189, 192, 199, 206, 211, 212, 212, 211, 207, 203, 207, 221, 225, 209, 180, 135, 210, 215, 199, 132, 39, 14, 158, 253, 198, 197, 193, 194, 199, 199, 196, 192, 191, 194, 201, 212, 217, 214, 208, 202, 196, 203, 226, 248, 242, 210, 164, 126, 212, 220, 219, 185, 134, 111, 151, 210, 191, 194, 191, 192, 197, 200, 197, 189, 183, 185, 201, 219, 226, 218, 201, 180, 170, 196, 245, 274, 256, 215, 157, 118, 215, 204, 207, 193, 168, 147, 161, 186, 184, 187, 185, 184, 185, 185, 174, 165, 163, 169, 185, 200, 204, 197, 176, 148, 150, 186, 232, 251, 232, 205, 142, 96, 154, 144, 142, 139, 128, 114, 116, 124, 124, 125, 125, 122, 119, 113, 105, 100, 100, 110, 127, 139, 137, 125, 106, 90, 94, 127, 161, 170, 152, 137, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 28, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 33, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 35, 13, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 53, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 47, 43, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 62, 67, 114, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 81, 75, 160, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 107, 72, 178, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 133, 68, 168, 142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 138, 60, 135, 156, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 129, 44, 96, 143, 31, 0, 0, 49, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 119, 37, 68, 112, 24, 0, 47, 141, 66, 0, 0, 0, 0, 11, 94, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 136, 56, 64, 75, 0, 0, 73, 217, 187, 35, 0, 0, 17, 73, 126, 126, 54, 0, 0, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 2, 0, 44, 184, 123, 93, 64, 0, 0, 74, 228, 255, 172, 81, 75, 100, 113, 116, 101, 72, 37, 17, 14, 21, 42, 68, 83, 80, 70, 63, 51, 53, 57, 1, 74, 205, 175, 130, 71, 0, 10, 126, 208, 203, 142, 92, 77, 100, 106, 99, 80, 59, 55, 60, 74, 86, 97, 110, 123, 129, 127, 123, 118, 128, 121, 34, 94, 202, 182, 158, 85, 36, 85, 194, 198, 141, 89, 74, 77, 77, 79, 79, 77, 76, 78, 86, 99, 112, 121, 129, 138, 146, 147, 149, 149, 170, 167, 57, 109, 172, 149, 156, 124, 98, 168, 236, 167, 90, 79, 90, 94, 91, 90, 89, 90, 92, 96, 104, 115, 127, 139, 148, 155, 156, 159, 166, 174, 200, 199, 80, 112, 177, 128, 137, 137, 177, 246, 255, 136, 64, 85, 106, 111, 106, 99, 98, 101, 104, 111, 120, 131, 143, 156, 164, 164, 159, 160, 173, 188, 209, 204, 98, 117, 182, 148, 126, 150, 202, 278, 252, 144, 82, 98, 115, 124, 116, 105, 102, 106, 114, 122, 131, 140, 148, 157, 162, 161, 159, 163, 179, 194, 196, 172, 79, 120, 187, 156, 152, 144, 188, 239, 201, 125, 92, 99, 119, 131, 128, 117, 111, 114, 122, 131, 138, 141, 142, 143, 147, 157, 171, 184, 193, 185, 168, 135, 54, 128, 198, 161, 162, 156, 152, 178, 142, 87, 80, 98, 120, 132, 133, 127, 120, 121, 131, 145, 150, 143, 135, 132, 134, 157, 196, 224, 210, 173, 147, 117, 45, 102, 191, 162, 151, 151, 137, 123, 101, 77, 76, 86, 105, 114, 116, 113, 115, 120, 131, 146, 157, 146, 128, 118, 117, 147, 196, 229, 218, 172, 141, 110, 45, 61, 143, 137, 120, 120, 112, 96, 81, 69, 68, 71, 79, 83, 82, 81, 82, 89, 101, 115, 126, 125, 114, 106, 109, 126, 154, 177, 175, 145, 114, 82, 41, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 7, 16, 16, 13, 1, 0, 0, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 21, 10, 14, 31, 36, 40, 33, 24, 8, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 18, 14, 30, 56, 50, 40, 42, 30, 14, 0, 0, 0, 38, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 27, 17, 15, 12, 5, 29, 58, 50, 30, 31, 30, 11, 0, 0, 0, 35, 0, 0, 19, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 59, 37, 11, 6, 0, 16, 48, 44, 24, 16, 22, 1, 0, 0, 0, 23, 0, 0, 60, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 57, 35, 8, 5, 0, 0, 13, 34, 26, 3, 0, 3, 0, 0, 0, 1, 0, 29, 78, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 31, 3, 0, 0, 0, 0, 0, 36, 42, 7, 0, 0, 0, 0, 0, 0, 0, 35, 63, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 61, 26, 0, 0, 0, 0, 0, 1, 0, 24, 43, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 73, 53, 13, 0, 0, 0, 0, 9, 0, 12, 11, 0, 2, 0, 0, 0, 0, 0, 32, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 68, 83, 77, 47, 23, 10, 0, 0, 12, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 42, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 63, 92, 93, 76, 56, 38, 0, 0, 11, 0, 0, 0, 0, 0, 19, 0, 0, 0, 1, 21, 5, 0, 6, 35, 26, 0, 11, 0, 0, 0, 0, 9, 57, 88, 97, 97, 88, 53, 0, 0, 7, 0, 0, 0, 0, 0, 35, 12, 0, 0, 0, 0, 0, 6, 54, 79, 72, 50, 51, 31, 11, 0, 0, 11, 48, 67, 83, 99, 103, 56, 0, 0, 0, 0, 0, 0, 0, 0, 35, 50, 15, 0, 0, 0, 0, 35, 75, 86, 82, 85, 86, 59, 28, 18, 1, 13, 38, 52, 80, 101, 94, 35, 0, 0, 0, 0, 0, 0, 0, 0, 27, 63, 19, 18, 14, 14, 33, 55, 69, 38, 40, 73, 104, 76, 53, 31, 6, 9, 30, 51, 79, 90, 69, 3, 0, 0, 0, 0, 0, 0, 0, 0, 12, 45, 9, 0, 0, 24, 50, 51, 36, 0, 0, 31, 87, 67, 53, 36, 10, 7, 17, 47, 78, 80, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 34, 42, 5, 0, 0, 0, 33, 44, 29, 25, 14, 0, 0, 28, 67, 70, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 16, 27, 11, 0, 0, 0, 0, 12, 47, 56, 49, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 26, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 2, 10, 4, 0, 0, 0, 0, 0, 0, 8, 13, 6, 3, 12, 12, 0, 0, 0, 0, 6, 10, 13, 0, 30, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 86, 171, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 6, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 102, 94, 0, 0, 4, 6, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 48, 189, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 143, 186, 49, 0, 20, 0, 0, 0, 0, 35, 73, 36, 8, 23, 0, 0, 0, 0, 46, 199, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 179, 126, 42, 11, 0, 0, 0, 0, 72, 98, 49, 60, 118, 95, 0, 0, 0, 27, 208, 0, 18, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 100, 172, 70, 0, 0, 0, 0, 0, 130, 134, 21, 50, 166, 156, 29, 0, 0, 0, 209, 0, 89, 139, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 26, 197, 115, 19, 25, 0, 0, 0, 141, 184, 37, 18, 114, 151, 92, 0, 0, 0, 188, 0, 83, 136, 0, 0, 27, 0, 0, 0, 0, 141, 0, 0, 32, 235, 139, 46, 85, 0, 0, 0, 74, 212, 110, 2, 29, 113, 130, 44, 0, 0, 138, 0, 11, 61, 0, 34, 137, 1, 0, 0, 0, 234, 32, 0, 86, 274, 165, 85, 128, 5, 0, 0, 21, 240, 203, 23, 0, 72, 148, 112, 0, 0, 63, 0, 0, 0, 0, 166, 207, 62, 0, 0, 0, 218, 105, 0, 121, 306, 180, 123, 178, 0, 0, 0, 64, 284, 255, 42, 0, 39, 146, 145, 0, 0, 15, 0, 0, 0, 0, 247, 205, 87, 0, 0, 0, 93, 14, 0, 89, 334, 196, 134, 222, 0, 0, 0, 177, 350, 265, 46, 0, 0, 92, 137, 37, 6, 26, 0, 0, 0, 0, 310, 145, 40, 91, 0, 0, 0, 0, 0, 31, 334, 209, 133, 252, 0, 0, 0, 280, 371, 231, 42, 0, 0, 3, 95, 65, 65, 86, 0, 0, 0, 0, 399, 90, 0, 129, 0, 0, 0, 0, 0, 26, 261, 184, 149, 260, 0, 0, 0, 302, 350, 217, 58, 0, 0, 0, 54, 66, 97, 145, 0, 0, 0, 42, 498, 113, 0, 79, 55, 0, 0, 0, 0, 134, 186, 101, 142, 218, 0, 0, 0, 252, 303, 217, 69, 0, 0, 0, 44, 39, 82, 173, 0, 0, 0, 24, 523, 235, 0, 0, 117, 0, 0, 0, 8, 245, 133, 23, 95, 115, 0, 0, 0, 125, 259, 246, 82, 0, 0, 0, 21, 0, 37, 187, 0, 0, 0, 0, 478, 366, 0, 0, 132, 0, 0, 0, 27, 210, 72, 0, 52, 0, 0, 0, 0, 0, 211, 268, 93, 0, 0, 0, 0, 0, 6, 211, 0, 0, 0, 0, 385, 460, 0, 0, 109, 87, 0, 0, 0, 48, 0, 0, 87, 0, 0, 0, 0, 0, 146, 219, 77, 0, 0, 0, 0, 0, 8, 237, 0, 0, 14, 0, 275, 494, 35, 0, 15, 195, 133, 0, 0, 0, 0, 0, 198, 0, 0, 19, 37, 18, 113, 123, 26, 0, 0, 0, 0, 0, 30, 244, 0, 0, 40, 0, 179, 488, 110, 0, 0, 224, 254, 3, 0, 0, 0, 0, 302, 113, 0, 13, 81, 86, 73, 23, 0, 0, 0, 0, 0, 0, 43, 232, 0, 0, 18, 0, 123, 449, 71, 0, 0, 230, 325, 39, 0, 0, 0, 0, 365, 278, 40, 2, 23, 21, 0, 0, 0, 0, 0, 0, 0, 0, 26, 192, 0, 0, 0, 0, 100, 365, 0, 0, 0, 294, 441, 142, 0, 0, 0, 3, 286, 319, 164, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 174, 0, 0, 0, 0, 85, 264, 0, 0, 0, 357, 553, 255, 0, 0, 0, 0, 140, 174, 107, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 204, 0, 0, 0, 0, 39, 105, 0, 0, 0, 472, 535, 254, 3, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 251, 0, 0, 0, 0, 0, 0, 0, 0, 259, 551, 376, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 300, 0, 0, 0, 0, 0, 0, 0, 0, 515, 513, 167, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 357, 0, 0, 46, 0, 0, 0, 0, 62, 625, 394, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 382, 0, 0, 37, 30, 0, 0, 0, 121, 573, 277, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 343, 0, 0, 16, 3, 30, 0, 0, 72, 381, 167, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 135, 275, 0, 0, 22, 0, 26, 0, 0, 8, 161, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 104, 139, 240, 0, 0, 72, 17, 40, 53, 1, 20, 71, 45, 0, 0, 0, 0, 16, 9, 0, 0, 0, 0, 34, 56, 43, 0, 0, 0, 0, 75, 171, 155, 155, 220, 0, 0, 74, 29, 35, 48, 36, 33, 42, 38, 17, 6, 8, 13, 14, 0, 0, 0, 0, 0, 55, 69, 43, 0, 0, 0, 0, 109, 161, 124, 119, 145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 33, 58, 89, 102, 86, 46, 0, 0, 0, 0, 0, 0, 83, 77, 26, 32, 14, 9, 6, 0, 0, 0, 0, 0, 0, 0, 38, 40, 44, 65, 70, 48, 14, 17, 69, 139, 181, 182, 149, 84, 17, 0, 0, 0, 59, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 108, 133, 129, 64, 0, 0, 0, 0, 0, 0, 72, 132, 131, 60, 0, 0, 0, 76, 91, 83, 92, 21, 0, 0, 0, 0, 45, 112, 102, 0, 0, 72, 149, 146, 100, 34, 0, 0, 0, 0, 0, 0, 0, 46, 139, 121, 26, 0, 0, 73, 119, 157, 199, 102, 7, 0, 0, 0, 24, 154, 221, 121, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 136, 79, 0, 0, 0, 0, 10, 110, 84, 25, 0, 0, 0, 0, 35, 106, 26, 0, 0, 0, 0, 0, 20, 69, 0, 0, 0, 53, 28, 0, 0, 4, 110, 124, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 183, 108, 0, 0, 26, 65, 0, 0, 0, 56, 137, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 96, 138, 76, 0, 0, 0, 0, 0, 0, 0, 0, 108, 138, 4, 0, 0, 0, 0, 0, 0, 12, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 117, 60, 62, 0, 0, 0, 0, 0, 0, 175, 338, 224, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 26, 68, 13, 3, 0, 0, 0, 0, 74, 326, 413, 221, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 57, 19, 0, 0, 0, 0, 0, 38, 0, 0, 9, 0, 56, 0, 0, 140, 297, 196, 50, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 35, 30, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 80, 62, 0, 22, 154, 70, 0, 0, 0, 0, 0, 0, 0, 0, 68, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 44, 0, 0, 61, 45, 0, 0, 4, 103, 89, 25, 0, 24, 123, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 42, 188, 193, 133, 95, 134, 157, 105, 41, 44, 156, 185, 78, 0, 0, 22, 78, 95, 80, 47, 1, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 244, 393, 328, 179, 82, 56, 47, 31, 29, 117, 233, 209, 84, 11, 55, 107, 125, 85, 14, 0, 0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 245, 232, 63, 0, 0, 0, 0, 0, 0, 52, 171, 173, 94, 46, 51, 47, 7, 0, 0, 0, 0, 116, 1, 0, 0, 0, 0, 0, 25, 0, 0, 0, 64, 106, 0, 0, 0, 0, 0, 62, 0, 0, 51, 97, 44, 0, 0, 0, 0, 0, 0, 0, 0, 162, 84, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 156, 123, 56, 0, 0, 0, 0, 0, 10, 13, 18, 13, 0, 156, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 70, 0, 0, 0, 0, 0, 0, 29, 38, 31, 30, 0, 135, 128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 153, 170, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 146, 226, 126, 31, 0, 0, 0, 0, 0, 0, 0, 52, 209, 314, 393, 389, 291, 129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 123, 256, 289, 236, 76, 0, 0, 0, 56, 170, 197, 154, 139, 145, 160, 165, 138, 78, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 97, 201, 321, 259, 82, 0, 0, 88, 184, 141, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 175, 238, 148, 41, 6, 31, 96, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 34, 20, 0, 0, 0, 0, 23, 0, 0, 35, 128, 188, 182, 59, 0, 7, 1, 0, 2, 3, 11, 16, 13, 4, 0, 0, 0, 1, 13, 25, 38, 47, 40, 20, 9, 31, 57, 0, 49, 5, 0, 0, 41, 179, 353, 248, 58, 11, 3, 14, 2, 0, 0, 0, 12, 13, 9, 9, 16, 31, 51, 64, 55, 22, 0, 0, 32, 90, 124, 30, 50, 19, 0, 0, 0, 109, 320, 369, 197, 79, 58, 66, 48, 19, 0, 0, 0, 0, 0, 0, 8, 26, 47, 55, 31, 0, 0, 0, 2, 54, 75, 1, 52, 20, 0, 0, 0, 0, 113, 204, 142, 71, 65, 89, 101, 95, 74, 48, 23, 0, 0, 0, 0, 0, 13, 13, 0, 0, 0, 0, 0, 6, 10, 0, 132, 143, 122, 123, 95, 69, 87, 118, 106, 84, 92, 117, 145, 166, 178, 185, 184, 170, 148, 123, 107, 107, 115, 129, 147, 155, 146, 142, 132, 122, 86, 7, 187, 274, 271, 258, 243, 221, 203, 196, 181, 165, 160, 168, 175, 183, 193, 209, 239, 274, 302, 310, 292, 263, 247, 260, 308, 380, 417, 394, 324, 259, 189, 83, 83, 43, 74, 51, 54, 50, 42, 41, 40, 39, 39, 42, 51, 55, 52, 46, 40, 39, 42, 42, 47, 57, 64, 65, 60, 51, 40, 30, 17, 0, 0, 0, 56, 3, 62, 42, 56, 54, 45, 45, 44, 36, 15, 3, 21, 37, 39, 44, 45, 41, 31, 13, 1, 5, 17, 33, 48, 59, 57, 45, 25, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 1, 0, 0, 0, 0, 0, 0, 15, 14, 0, 12, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 118, 28, 20, 0, 10, 44, 41, 104, 182, 134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 115, 48, 65, 20, 0, 8, 0, 35, 168, 180, 42, 0, 0, 0, 0, 0, 0, 0, 0, 27, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 21, 81, 56, 0, 0, 0, 0, 31, 103, 27, 9, 13, 0, 0, 0, 50, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 47, 50, 0, 0, 0, 0, 0, 15, 0, 40, 76, 36, 0, 2, 85, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 51, 85, 76, 22, 41, 87, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 29, 75, 88, 68, 42, 26, 51, 72, 0, 0, 35, 0, 0, 0, 0, 6, 13, 16, 9, 0, 0, 6, 0, 76, 1, 10, 20, 0, 0, 0, 9, 0, 18, 69, 85, 23, 0, 0, 11, 19, 0, 0, 24, 11, 0, 13, 0, 0, 0, 0, 0, 0, 0, 17, 0, 113, 36, 21, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 34, 4, 146, 63, 31, 31, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 160, 86, 47, 29, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 139, 88, 52, 41, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 103, 77, 32, 40, 67, 0, 0, 0, 0, 0, 0, 43, 85, 113, 83, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 93, 92, 38, 52, 94, 40, 126, 143, 137, 118, 123, 118, 105, 98, 68, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 82, 111, 109, 143, 157, 88, 147, 148, 130, 68, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 69, 133, 194, 167, 90, 79, 46, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 84, 149, 95, 35, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 99, 31, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 55, 80, 0, 30, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 17, 44, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 20, 22, 21, 21, 18, 13, 5, 3, 13, 29, 44, 54, 57, 35, 0, 0, 0, 11, 11, 64, 46, 43, 40, 35, 14, 0, 0, 0, 0, 0, 5, 18, 34, 50, 66, 77, 76, 70, 62, 61, 81, 110, 127, 129, 110, 80, 38, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 6, 9, 8, 6, 0, 0, 0, 0, 0, 24, 5, 11, 9, 10, 16, 19, 17, 9, 7, 11, 9, 6, 6, 10, 16, 17, 18, 26, 29, 23, 15, 14, 16, 21, 23, 22, 1, 0, 24, 5, 0, 9, 0, 0, 0, 0, 0, 1, 0, 0, 0, 17, 0, 0, 0, 0, 0, 6, 19, 42, 51, 37, 15, 0, 0, 1, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 44, 40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 47, 52, 42, 28, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 93, 95, 79, 81, 89, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 121, 134, 107, 112, 131, 94, 6, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 28, 42, 66, 0, 0, 0, 129, 163, 117, 92, 123, 121, 47, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 80, 94, 111, 113, 12, 0, 0, 103, 166, 121, 76, 89, 116, 79, 0, 0, 0, 0, 0, 0, 79, 31, 77, 47, 0, 0, 0, 0, 4, 0, 0, 17, 95, 108, 126, 127, 28, 0, 0, 53, 133, 110, 72, 63, 94, 94, 36, 0, 0, 0, 0, 0, 100, 50, 123, 91, 0, 0, 0, 0, 13, 0, 0, 17, 88, 80, 98, 106, 24, 0, 0, 18, 104, 110, 77, 52, 79, 90, 64, 0, 0, 0, 0, 0, 61, 12, 126, 99, 0, 0, 0, 0, 7, 20, 0, 0, 78, 46, 53, 82, 0, 0, 0, 22, 102, 126, 99, 59, 70, 80, 81, 12, 0, 0, 0, 0, 0, 0, 126, 73, 0, 0, 0, 0, 0, 7, 0, 0, 69, 28, 23, 72, 0, 0, 0, 42, 117, 138, 116, 79, 72, 81, 95, 50, 0, 0, 0, 0, 0, 0, 149, 44, 0, 0, 0, 0, 0, 0, 0, 0, 61, 27, 29, 83, 0, 0, 0, 59, 123, 134, 123, 99, 90, 86, 120, 80, 12, 21, 0, 0, 0, 0, 175, 41, 0, 8, 0, 0, 0, 0, 0, 0, 77, 47, 52, 102, 0, 0, 0, 63, 114, 127, 121, 102, 98, 96, 131, 96, 18, 33, 0, 0, 0, 0, 176, 58, 0, 38, 17, 0, 0, 0, 0, 54, 105, 75, 87, 116, 0, 0, 0, 64, 122, 138, 124, 94, 91, 105, 144, 107, 8, 37, 0, 0, 0, 0, 151, 92, 0, 49, 107, 0, 0, 0, 0, 101, 119, 100, 124, 131, 22, 0, 0, 22, 104, 142, 117, 68, 62, 96, 140, 80, 0, 34, 0, 0, 0, 0, 103, 131, 0, 15, 151, 50, 0, 0, 0, 113, 120, 124, 159, 128, 68, 22, 0, 1, 83, 128, 82, 35, 31, 68, 115, 35, 0, 21, 0, 0, 0, 0, 38, 158, 16, 0, 131, 108, 0, 0, 0, 89, 77, 113, 171, 107, 50, 87, 57, 31, 69, 93, 58, 27, 31, 57, 90, 0, 0, 9, 0, 0, 0, 0, 0, 158, 35, 0, 77, 139, 84, 5, 0, 41, 0, 48, 165, 101, 45, 91, 76, 45, 54, 63, 40, 34, 37, 48, 72, 0, 0, 2, 0, 0, 32, 0, 0, 142, 31, 0, 0, 103, 111, 42, 0, 0, 0, 0, 120, 108, 78, 97, 87, 47, 45, 36, 30, 55, 45, 42, 65, 0, 0, 7, 0, 0, 31, 0, 0, 132, 16, 0, 0, 0, 40, 15, 0, 0, 0, 0, 48, 87, 55, 53, 31, 7, 0, 0, 0, 25, 34, 39, 68, 3, 0, 28, 0, 0, 0, 0, 0, 121, 0, 0, 0, 0, 20, 18, 0, 0, 0, 0, 0, 63, 32, 7, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 55, 0, 0, 0, 0, 0, 105, 0, 0, 0, 0, 44, 27, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 0, 0, 0, 0, 0, 65, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 13, 0, 28, 8, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 32, 17, 0, 0, 0, 0, 10, 0, 9, 83, 97, 0, 0, 0, 0, 51, 0, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 61, 37, 34, 0, 0, 0, 0, 0, 0, 0, 104, 160, 97, 0, 0, 0, 43, 0, 57, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 71, 32, 52, 0, 0, 0, 0, 14, 0, 0, 79, 162, 168, 46, 0, 0, 29, 0, 48, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 72, 50, 98, 17, 0, 0, 0, 49, 35, 0, 38, 133, 189, 144, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 82, 77, 152, 74, 0, 0, 0, 65, 95, 0, 0, 81, 175, 190, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 76, 94, 195, 76, 0, 0, 0, 66, 115, 2, 0, 18, 143, 184, 59, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 48, 78, 212, 43, 0, 0, 0, 86, 127, 15, 0, 0, 74, 150, 73, 27, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 25, 194, 0, 0, 0, 0, 108, 124, 28, 0, 0, 0, 84, 52, 47, 92, 0, 0, 0, 0, 123, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 149, 0, 0, 0, 0, 112, 129, 50, 0, 0, 0, 0, 0, 14, 100, 0, 0, 0, 0, 244, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 0, 0, 0, 0, 75, 119, 56, 0, 0, 0, 0, 0, 0, 90, 0, 0, 0, 0, 285, 116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 118, 61, 0, 0, 0, 0, 0, 0, 76, 0, 0, 0, 0, 247, 213, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 125, 64, 0, 0, 0, 0, 0, 0, 70, 0, 0, 0, 0, 160, 265, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 126, 72, 0, 0, 0, 0, 0, 0, 69, 0, 0, 0, 0, 57, 284, 0, 0, 0, 31, 44, 0, 0, 0, 0, 0, 130, 0, 0, 0, 0, 0, 52, 134, 93, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 0, 273, 21, 0, 0, 83, 158, 17, 0, 0, 0, 0, 168, 52, 0, 0, 0, 42, 122, 147, 117, 38, 0, 0, 0, 0, 0, 93, 0, 0, 0, 0, 0, 240, 5, 0, 0, 88, 209, 51, 0, 0, 0, 0, 173, 145, 20, 16, 63, 135, 162, 148, 127, 76, 0, 0, 0, 0, 0, 151, 0, 0, 0, 0, 0, 166, 0, 0, 0, 66, 232, 90, 0, 0, 0, 0, 111, 197, 153, 134, 136, 143, 146, 140, 130, 96, 28, 0, 19, 0, 57, 207, 0, 0, 0, 0, 0, 54, 0, 0, 0, 19, 253, 148, 0, 0, 0, 0, 89, 187, 202, 189, 154, 139, 139, 136, 137, 133, 109, 88, 110, 97, 146, 250, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 267, 201, 99, 66, 62, 72, 130, 180, 188, 180, 164, 157, 156, 152, 151, 155, 153, 148, 160, 148, 194, 299, 0, 44, 78, 0, 0, 0, 0, 0, 0, 214, 276, 212, 160, 152, 152, 144, 154, 172, 178, 174, 166, 167, 167, 159, 155, 164, 172, 166, 165, 146, 202, 332, 0, 106, 190, 95, 50, 0, 0, 0, 136, 306, 237, 178, 163, 173, 176, 172, 176, 184, 183, 174, 166, 165, 164, 161, 164, 174, 175, 156, 144, 127, 201, 344, 0, 112, 238, 215, 183, 0, 0, 0, 308, 322, 195, 156, 171, 197, 199, 188, 183, 181, 176, 170, 167, 166, 161, 163, 177, 187, 174, 143, 138, 135, 205, 344, 0, 108, 247, 252, 264, 0, 0, 0, 350, 296, 167, 144, 168, 198, 202, 193, 181, 172, 165, 165, 171, 176, 175, 180, 187, 183, 159, 141, 162, 180, 231, 328, 0, 101, 244, 234, 272, 71, 0, 37, 323, 264, 168, 146, 157, 183, 196, 188, 172, 162, 160, 167, 184, 196, 195, 187, 169, 146, 132, 155, 216, 251, 276, 312, 0, 85, 232, 210, 233, 159, 3, 112, 271, 241, 188, 169, 170, 184, 197, 188, 159, 137, 131, 149, 186, 207, 208, 183, 125, 76, 86, 169, 264, 286, 290, 294, 0, 83, 214, 185, 193, 181, 121, 145, 215, 213, 187, 175, 175, 186, 198, 183, 143, 111, 95, 114, 159, 188, 196, 169, 88, 15, 33, 147, 247, 259, 259, 248, 14, 87, 168, 146, 148, 152, 137, 138, 163, 169, 160, 153, 154, 157, 162, 154, 127, 101, 84, 95, 132, 154, 156, 139, 79, 23, 39, 124, 193, 191, 186, 174, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 44, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 24, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 19, 11, 0, 0, 0, 0, 0, 0, 0, 19, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 17, 3, 0, 0, 0, 0, 0, 0, 0, 11, 15, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 7, 0, 0, 0, 0, 0, 20, 14, 9, 12, 31, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 0, 10, 35, 17, 0, 6, 22, 31, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 7, 16, 2, 0, 0, 6, 24, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 107, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 136, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 138, 96, 19, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 118, 112, 50, 0, 11, 15, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 90, 112, 59, 13, 8, 23, 0, 0, 0, 0, 0, 0, 61, 38, 0, 0, 0, 7, 16, 17, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 93, 34, 0, 8, 69, 68, 34, 25, 23, 29, 67, 119, 117, 86, 62, 42, 28, 33, 50, 64, 55, 25, 12, 11, 13, 16, 23, 0, 0, 0, 0, 37, 67, 6, 0, 0, 128, 185, 179, 147, 128, 91, 92, 124, 129, 111, 103, 93, 95, 108, 124, 136, 136, 125, 109, 107, 112, 108, 86, 11, 20, 4, 40, 32, 26, 0, 0, 11, 152, 225, 185, 126, 89, 61, 56, 81, 104, 116, 123, 135, 146, 157, 165, 167, 167, 163, 161, 163, 165, 161, 120, 20, 69, 29, 35, 19, 0, 0, 0, 49, 161, 198, 151, 113, 98, 90, 93, 105, 119, 133, 142, 151, 160, 165, 166, 170, 177, 184, 189, 193, 192, 184, 135, 25, 119, 78, 57, 18, 0, 0, 0, 76, 153, 149, 128, 132, 140, 147, 147, 149, 153, 156, 157, 161, 167, 173, 179, 187, 197, 203, 207, 208, 206, 201, 162, 51, 159, 150, 107, 36, 0, 0, 0, 97, 142, 135, 133, 159, 172, 168, 161, 160, 162, 165, 169, 175, 182, 190, 200, 209, 212, 208, 203, 208, 215, 221, 196, 82, 175, 183, 158, 85, 0, 0, 43, 141, 153, 149, 152, 178, 181, 172, 163, 160, 163, 170, 178, 186, 193, 198, 205, 211, 209, 202, 200, 211, 222, 222, 187, 70, 176, 196, 188, 146, 64, 37, 95, 164, 164, 158, 170, 184, 188, 185, 176, 168, 165, 170, 179, 189, 193, 195, 194, 194, 195, 200, 214, 227, 222, 201, 147, 40, 171, 196, 205, 187, 131, 87, 98, 142, 150, 141, 159, 171, 181, 187, 185, 178, 175, 180, 190, 197, 198, 194, 185, 178, 184, 205, 237, 251, 234, 201, 135, 35, 151, 188, 214, 212, 187, 152, 136, 144, 149, 141, 145, 150, 159, 166, 165, 161, 161, 170, 189, 207, 216, 209, 188, 173, 177, 204, 253, 280, 269, 230, 165, 67, 107, 162, 184, 187, 177, 162, 149, 142, 142, 136, 134, 131, 131, 128, 122, 115, 114, 124, 146, 170, 182, 177, 164, 152, 150, 175, 211, 228, 217, 190, 150, 78, 0, 46, 101, 86, 89, 79, 79, 84, 83, 77, 71, 73, 81, 82, 83, 88, 89, 87, 81, 77, 75, 68, 60, 61, 68, 75, 76, 73, 70, 72, 85, 82, 0, 0, 68, 52, 60, 51, 53, 62, 62, 51, 40, 49, 66, 47, 40, 59, 74, 72, 58, 42, 32, 19, 0, 0, 8, 24, 38, 53, 60, 76, 115, 115, 0, 0, 41, 27, 36, 26, 28, 39, 36, 23, 15, 53, 104, 53, 9, 36, 54, 38, 8, 0, 3, 1, 0, 0, 0, 0, 0, 0, 29, 67, 128, 130, 0, 0, 46, 27, 41, 35, 31, 37, 30, 12, 12, 81, 155, 96, 10, 11, 13, 0, 0, 0, 43, 52, 28, 0, 0, 0, 0, 0, 0, 53, 136, 138, 0, 0, 20, 0, 13, 39, 36, 33, 24, 0, 0, 31, 100, 79, 0, 0, 0, 0, 0, 0, 67, 76, 50, 23, 12, 0, 0, 0, 0, 25, 136, 149, 0, 0, 0, 0, 0, 29, 43, 34, 23, 0, 0, 0, 34, 61, 39, 0, 0, 0, 0, 0, 54, 65, 26, 13, 34, 29, 0, 0, 0, 0, 124, 161, 0, 30, 0, 0, 0, 17, 37, 26, 24, 30, 0, 0, 16, 93, 104, 37, 0, 0, 0, 0, 12, 58, 24, 0, 2, 31, 4, 0, 0, 0, 96, 164, 0, 94, 0, 0, 0, 31, 19, 6, 35, 93, 74, 0, 18, 115, 119, 36, 0, 0, 0, 0, 0, 52, 50, 0, 0, 19, 22, 0, 0, 0, 59, 146, 0, 91, 16, 0, 21, 52, 0, 0, 50, 183, 207, 62, 29, 107, 98, 29, 0, 0, 0, 0, 0, 66, 84, 31, 0, 18, 44, 20, 0, 0, 18, 100, 0, 47, 0, 0, 51, 62, 0, 0, 3, 140, 204, 87, 36, 113, 100, 39, 4, 0, 0, 0, 1, 111, 112, 59, 0, 16, 55, 51, 0, 0, 0, 57, 0, 5, 0, 0, 55, 60, 0, 0, 0, 0, 76, 37, 21, 123, 131, 60, 30, 31, 0, 0, 36, 127, 97, 38, 0, 0, 48, 59, 29, 0, 0, 35, 0, 0, 0, 0, 40, 29, 14, 0, 0, 0, 0, 0, 2, 123, 163, 90, 48, 68, 0, 0, 26, 104, 69, 9, 0, 0, 14, 42, 41, 18, 32, 49, 0, 0, 0, 0, 26, 0, 0, 45, 0, 0, 0, 0, 9, 100, 138, 103, 66, 76, 0, 0, 17, 95, 63, 8, 0, 0, 0, 24, 41, 48, 64, 71, 0, 0, 0, 0, 32, 0, 0, 65, 0, 0, 0, 0, 36, 71, 57, 62, 60, 62, 0, 0, 19, 95, 71, 24, 0, 0, 0, 18, 35, 49, 74, 90, 0, 0, 2, 25, 70, 0, 0, 45, 32, 0, 0, 0, 54, 62, 0, 0, 22, 24, 0, 0, 8, 83, 86, 33, 0, 0, 0, 0, 7, 29, 79, 108, 0, 1, 16, 41, 100, 0, 0, 18, 55, 0, 0, 0, 9, 23, 0, 0, 0, 0, 0, 0, 0, 40, 80, 51, 0, 0, 0, 0, 0, 15, 90, 132, 0, 8, 18, 34, 93, 18, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 45, 0, 0, 0, 0, 0, 29, 112, 151, 0, 4, 10, 16, 72, 49, 0, 0, 33, 18, 0, 0, 0, 0, 20, 47, 20, 0, 0, 11, 13, 5, 21, 5, 0, 0, 0, 0, 3, 51, 129, 156, 0, 0, 3, 0, 52, 71, 0, 0, 9, 44, 8, 0, 0, 0, 45, 91, 83, 0, 0, 17, 42, 25, 17, 0, 0, 0, 0, 0, 21, 63, 132, 152, 0, 0, 0, 0, 34, 68, 0, 0, 42, 91, 52, 0, 0, 0, 49, 115, 127, 7, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 6, 45, 103, 128, 0, 0, 0, 0, 25, 48, 0, 0, 90, 172, 141, 23, 0, 0, 45, 95, 118, 58, 0, 0, 0, 3, 9, 14, 0, 0, 0, 0, 0, 5, 52, 84, 0, 0, 0, 0, 23, 38, 0, 0, 118, 198, 179, 69, 0, 0, 0, 0, 11, 21, 8, 13, 23, 29, 32, 35, 28, 0, 0, 0, 0, 10, 31, 50, 0, 0, 0, 0, 3, 21, 0, 0, 74, 114, 71, 0, 0, 0, 0, 0, 0, 0, 0, 7, 21, 27, 25, 15, 4, 0, 0, 0, 0, 15, 8, 26, 0, 0, 0, 0, 0, 0, 0, 0, 44, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 74, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 67, 109, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 4, 0, 0, 0, 0, 0, 62, 104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 86, 86, 67, 59, 58, 59, 57, 54, 55, 60, 63, 63, 64, 65, 63, 57, 50, 49, 50, 50, 51, 56, 61, 62, 58, 53, 49, 44, 43, 16, 0, 102, 129, 119, 91, 78, 81, 82, 77, 71, 74, 88, 91, 72, 65, 76, 80, 73, 66, 64, 66, 58, 53, 60, 76, 85, 85, 81, 72, 62, 48, 0, 0, 114, 149, 155, 132, 120, 119, 120, 115, 105, 108, 133, 127, 93, 79, 100, 117, 107, 90, 81, 70, 52, 38, 38, 55, 81, 104, 115, 115, 102, 77, 0, 0, 123, 161, 172, 160, 150, 145, 142, 134, 125, 140, 187, 160, 103, 83, 101, 121, 108, 81, 76, 62, 21, 0, 0, 0, 37, 72, 105, 134, 139, 110, 14, 0, 120, 151, 159, 166, 167, 155, 145, 136, 133, 158, 217, 183, 104, 72, 62, 59, 52, 43, 57, 41, 0, 0, 0, 0, 0, 8, 46, 103, 150, 136, 33, 0, 103, 109, 102, 149, 180, 165, 148, 137, 139, 155, 188, 168, 103, 42, 0, 0, 0, 11, 41, 44, 0, 0, 0, 0, 0, 0, 0, 56, 135, 152, 52, 4, 56, 21, 5, 91, 167, 165, 147, 133, 133, 126, 107, 103, 78, 8, 0, 0, 0, 0, 45, 77, 25, 0, 0, 0, 0, 0, 0, 7, 93, 153, 66, 16, 0, 0, 0, 24, 127, 141, 132, 132, 119, 66, 10, 23, 47, 0, 0, 0, 0, 15, 57, 107, 68, 0, 0, 0, 0, 0, 0, 0, 33, 127, 76, 28, 0, 0, 0, 0, 78, 99, 108, 142, 124, 18, 0, 0, 20, 0, 0, 0, 0, 14, 42, 103, 84, 0, 0, 0, 0, 0, 0, 0, 0, 74, 68, 35, 0, 0, 0, 14, 41, 67, 95, 164, 184, 47, 0, 0, 9, 0, 0, 0, 0, 0, 0, 75, 55, 0, 0, 0, 0, 0, 0, 0, 0, 3, 30, 32, 0, 0, 0, 10, 14, 60, 106, 173, 222, 127, 7, 31, 35, 0, 0, 0, 0, 0, 0, 44, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 65, 120, 150, 206, 185, 91, 96, 73, 0, 0, 0, 0, 0, 0, 48, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 127, 126, 162, 174, 135, 135, 105, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 114, 110, 114, 141, 156, 153, 96, 0, 0, 0, 0, 0, 6, 71, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 93, 88, 123, 177, 161, 71, 5, 0, 12, 0, 12, 62, 105, 26, 0, 0, 0, 0, 4, 38, 42, 26, 35, 0, 0, 0, 0, 0, 0, 0, 0, 20, 70, 76, 123, 200, 174, 62, 17, 37, 54, 35, 60, 111, 135, 86, 4, 0, 0, 0, 34, 72, 80, 75, 88, 29, 0, 0, 0, 0, 0, 0, 0, 0, 42, 58, 109, 159, 151, 70, 30, 52, 41, 26, 79, 132, 127, 117, 60, 0, 0, 0, 41, 85, 106, 116, 126, 41, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 62, 72, 95, 87, 57, 50, 0, 0, 46, 112, 107, 106, 80, 7, 0, 0, 41, 97, 134, 145, 141, 41, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 52, 47, 15, 0, 0, 0, 69, 91, 77, 30, 0, 0, 0, 22, 99, 153, 160, 141, 37, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 5, 0, 0, 0, 0, 0, 58, 123, 130, 104, 10, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 3, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 114, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 298, 118, 3, 40, 33, 36, 16, 0, 23, 30, 0, 0, 0, 58, 92, 25, 1, 20, 31, 17, 18, 78, 171, 224, 222, 175, 111, 45, 0, 0, 0, 0, 316, 154, 46, 76, 57, 66, 64, 59, 94, 93, 0, 0, 0, 0, 145, 126, 133, 167, 128, 7, 0, 0, 32, 149, 226, 267, 266, 183, 70, 0, 0, 0, 301, 175, 111, 127, 53, 39, 63, 76, 120, 143, 3, 0, 0, 0, 177, 248, 272, 278, 156, 0, 0, 0, 0, 0, 0, 124, 262, 286, 161, 0, 0, 0, 272, 226, 276, 290, 124, 42, 58, 79, 111, 174, 152, 0, 0, 0, 138, 244, 257, 246, 124, 0, 0, 0, 0, 0, 0, 0, 178, 336, 263, 16, 0, 0, 180, 196, 350, 404, 201, 76, 71, 72, 58, 127, 224, 175, 0, 0, 0, 49, 85, 111, 93, 0, 0, 0, 0, 0, 0, 0, 85, 315, 351, 117, 0, 0, 23, 0, 169, 275, 114, 68, 105, 55, 0, 0, 89, 139, 0, 0, 0, 0, 0, 49, 144, 34, 0, 0, 0, 0, 0, 0, 0, 235, 382, 236, 0, 0, 0, 0, 0, 0, 0, 0, 151, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 239, 171, 0, 0, 0, 0, 0, 0, 0, 99, 333, 322, 26, 0, 0, 0, 0, 0, 0, 0, 187, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 290, 172, 0, 0, 0, 0, 0, 0, 0, 0, 205, 320, 150, 0, 0, 0, 0, 0, 0, 0, 185, 291, 18, 0, 0, 0, 0, 0, 0, 0, 0, 104, 264, 75, 0, 0, 0, 0, 0, 0, 0, 0, 39, 210, 156, 17, 9, 0, 0, 0, 0, 0, 98, 330, 322, 0, 0, 0, 0, 0, 0, 0, 0, 35, 197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 48, 3, 12, 0, 0, 0, 0, 0, 27, 196, 362, 180, 0, 0, 0, 0, 0, 0, 0, 0, 127, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 44, 67, 258, 243, 0, 0, 0, 0, 0, 0, 0, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 85, 0, 138, 233, 0, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 60, 0, 0, 195, 14, 0, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 103, 188, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 122, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 168, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 147, 189, 124, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 202, 103, 0, 0, 0, 0, 19, 0, 0, 0, 0, 13, 106, 194, 192, 102, 0, 0, 0, 0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167, 121, 0, 0, 0, 0, 0, 35, 0, 0, 0, 65, 133, 172, 162, 83, 0, 0, 0, 0, 0, 160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 41, 33, 36, 46, 57, 74, 56, 0, 0, 0, 0, 0, 215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 257, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 249, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 125, 129, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 96, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 210, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 132, 172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 9, 0, 0, 0, 0, 0, 0, 0, 0, 12, 24, 28, 33, 45, 61, 62, 40, 0, 0, 0, 0, 0, 12, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 53, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 36, 36, 26, 15, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 28, 34, 37, 38, 30, 1, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 35, 47, 50, 4, 0, 0, 0, 0, 0, 19, 41, 49, 36, 0, 0, 0, 40, 0, 12, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 69, 66, 43, 0, 0, 0, 0, 0, 0, 0, 33, 51, 63, 21, 0, 0, 29, 0, 38, 30, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 51, 48, 28, 0, 0, 0, 0, 0, 0, 0, 31, 59, 74, 57, 0, 0, 22, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 32, 22, 18, 0, 0, 0, 0, 16, 15, 28, 64, 74, 87, 7, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 44, 41, 49, 0, 0, 0, 0, 24, 22, 18, 45, 74, 85, 47, 18, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 56, 56, 67, 0, 0, 0, 0, 0, 5, 0, 14, 54, 71, 70, 57, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 53, 55, 0, 0, 0, 0, 0, 2, 0, 0, 27, 62, 67, 87, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 9, 0, 0, 0, 0, 7, 17, 0, 0, 0, 34, 39, 80, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 31, 18, 0, 0, 0, 0, 51, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 5, 0, 0, 0, 0, 22, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 3, 31, 24, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 12, 41, 58, 36, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 40, 0, 0, 0, 0, 0, 9, 0, 0, 0, 23, 64, 84, 77, 43, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 78, 25, 0, 0, 0, 0, 0, 21, 16, 31, 66, 96, 107, 109, 78, 17, 0, 0, 0, 0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 42, 74, 92, 105, 101, 92, 84, 76, 50, 26, 23, 0, 47, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 60, 77, 75, 58, 40, 27, 19, 20, 25, 35, 7, 52, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 26, 25, 14, 0, 0, 0, 0, 0, 0, 0, 9, 70, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 30, 27, 23, 18, 14, 16, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 8, 4, 4, 5, 5, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 199, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 118, 308, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 51, 0, 0, 0, 0, 0, 0, 0, 37, 22, 0, 0, 0, 0, 0, 0, 0, 85, 341, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 239, 234, 0, 0, 8, 0, 0, 0, 0, 50, 104, 62, 0, 0, 0, 0, 0, 0, 64, 344, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 216, 350, 134, 14, 30, 0, 0, 0, 0, 55, 111, 72, 78, 122, 32, 0, 0, 0, 46, 363, 0, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 278, 253, 94, 24, 0, 0, 0, 0, 109, 106, 0, 61, 241, 209, 0, 0, 0, 0, 376, 0, 169, 238, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 116, 295, 129, 1, 1, 0, 0, 0, 185, 178, 0, 0, 226, 283, 116, 0, 0, 0, 361, 0, 265, 327, 0, 0, 0, 0, 0, 0, 110, 194, 0, 0, 37, 330, 174, 12, 58, 0, 0, 0, 177, 284, 29, 0, 104, 249, 225, 0, 0, 0, 301, 0, 201, 249, 0, 0, 101, 0, 0, 0, 32, 415, 0, 0, 90, 375, 216, 74, 134, 0, 0, 0, 86, 348, 187, 0, 0, 168, 277, 172, 0, 0, 191, 0, 68, 53, 0, 160, 282, 59, 0, 0, 0, 433, 120, 0, 189, 431, 248, 157, 222, 22, 0, 0, 47, 382, 304, 0, 0, 73, 275, 280, 0, 0, 79, 0, 0, 0, 0, 284, 355, 193, 0, 0, 0, 287, 104, 0, 221, 498, 267, 214, 310, 1, 0, 0, 137, 436, 352, 1, 0, 0, 204, 283, 53, 0, 40, 0, 0, 0, 0, 344, 265, 204, 57, 0, 0, 55, 0, 0, 132, 543, 300, 220, 373, 0, 0, 0, 301, 506, 361, 14, 0, 0, 61, 203, 88, 53, 99, 0, 0, 0, 0, 466, 110, 54, 239, 0, 0, 0, 0, 0, 12, 461, 274, 216, 413, 0, 0, 0, 410, 516, 326, 39, 0, 0, 0, 91, 62, 129, 192, 0, 0, 0, 97, 682, 70, 0, 233, 0, 0, 0, 0, 0, 32, 298, 165, 203, 409, 0, 0, 0, 402, 470, 296, 52, 0, 0, 0, 15, 12, 142, 266, 0, 0, 0, 179, 850, 196, 0, 131, 137, 0, 0, 0, 0, 197, 167, 12, 141, 312, 0, 0, 0, 274, 409, 299, 59, 0, 0, 0, 0, 0, 92, 307, 0, 0, 0, 108, 876, 416, 0, 0, 240, 0, 0, 0, 0, 300, 116, 0, 55, 124, 0, 0, 0, 40, 315, 346, 91, 0, 0, 0, 0, 0, 22, 341, 0, 0, 0, 0, 782, 616, 0, 0, 265, 65, 0, 0, 0, 184, 38, 0, 47, 0, 0, 0, 0, 0, 199, 343, 119, 0, 0, 0, 0, 0, 0, 383, 0, 0, 0, 0, 617, 732, 0, 0, 174, 236, 0, 0, 0, 0, 0, 42, 206, 0, 0, 0, 0, 0, 129, 264, 93, 0, 0, 0, 0, 0, 7, 418, 0, 0, 0, 0, 419, 759, 90, 0, 42, 354, 273, 0, 0, 0, 0, 98, 448, 16, 0, 0, 17, 21, 142, 142, 15, 0, 0, 0, 0, 0, 34, 419, 0, 0, 0, 0, 251, 726, 144, 0, 0, 457, 491, 87, 0, 0, 0, 91, 606, 302, 0, 0, 46, 92, 96, 43, 0, 0, 0, 0, 0, 0, 32, 368, 0, 0, 0, 0, 174, 664, 65, 0, 0, 550, 669, 191, 0, 0, 0, 16, 565, 473, 160, 56, 32, 27, 0, 0, 0, 0, 0, 0, 0, 0, 35, 321, 0, 0, 0, 0, 143, 556, 0, 0, 0, 564, 772, 301, 0, 0, 0, 0, 349, 406, 233, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 320, 0, 0, 0, 0, 93, 373, 0, 0, 0, 577, 804, 395, 0, 0, 0, 0, 96, 164, 108, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 375, 0, 0, 0, 0, 3, 122, 0, 0, 16, 659, 672, 314, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 456, 0, 0, 0, 0, 0, 0, 0, 0, 454, 709, 429, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 109, 541, 0, 0, 84, 0, 0, 0, 0, 0, 769, 637, 157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 124, 605, 0, 0, 117, 112, 88, 0, 0, 120, 861, 474, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 164, 589, 0, 0, 85, 117, 174, 0, 0, 121, 700, 302, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 202, 501, 0, 0, 47, 54, 153, 0, 0, 36, 405, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 91, 223, 414, 0, 0, 36, 0, 74, 0, 0, 0, 167, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 138, 145, 216, 371, 0, 0, 37, 0, 17, 24, 0, 0, 49, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 3, 0, 0, 0, 0, 48, 173, 141, 186, 311, 0, 0, 45, 0, 10, 30, 15, 12, 30, 30, 4, 0, 0, 7, 18, 0, 0, 0, 0, 0, 26, 48, 35, 0, 0, 0, 0, 63, 133, 93, 114, 185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 3, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 12, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 17, 39, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 3, 16, 27, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 2, 5, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 3, 0, 0, 0, 50, 42, 25, 30, 37, 17, 18, 43, 20, 0, 0, 0, 0, 0, 22, 48, 56, 21, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 5, 0, 0, 23, 84, 81, 47, 40, 29, 0, 0, 0, 3, 0, 0, 13, 46, 70, 86, 95, 96, 84, 60, 45, 43, 38, 54, 4, 38, 12, 0, 0, 16, 3, 0, 22, 47, 31, 0, 0, 0, 0, 0, 0, 4, 27, 43, 63, 84, 98, 104, 106, 103, 101, 99, 98, 95, 85, 89, 3, 66, 48, 7, 0, 0, 0, 0, 16, 0, 0, 0, 0, 23, 44, 54, 63, 71, 79, 80, 89, 100, 103, 101, 104, 108, 112, 112, 112, 110, 100, 97, 0, 84, 96, 56, 15, 0, 0, 0, 2, 0, 0, 1, 43, 77, 93, 89, 90, 91, 91, 95, 99, 104, 109, 114, 120, 123, 121, 116, 116, 120, 116, 111, 5, 95, 110, 93, 61, 17, 0, 0, 4, 0, 6, 45, 77, 96, 95, 89, 89, 91, 94, 101, 108, 115, 119, 123, 126, 122, 114, 109, 115, 129, 124, 113, 0, 102, 106, 110, 99, 61, 27, 4, 14, 17, 33, 68, 95, 98, 96, 94, 92, 93, 98, 104, 111, 117, 119, 118, 114, 111, 109, 117, 131, 139, 110, 83, 0, 104, 115, 116, 119, 93, 59, 29, 23, 28, 40, 73, 92, 97, 100, 101, 99, 98, 100, 106, 111, 115, 114, 110, 105, 105, 117, 136, 148, 138, 86, 59, 0, 105, 116, 125, 115, 111, 77, 60, 38, 33, 40, 69, 80, 85, 89, 94, 96, 100, 107, 114, 117, 118, 114, 106, 101, 109, 132, 152, 153, 130, 91, 67, 0, 103, 106, 121, 114, 105, 92, 91, 75, 60, 67, 81, 81, 77, 73, 73, 75, 83, 93, 106, 115, 116, 113, 106, 104, 114, 132, 144, 135, 117, 88, 71, 4, 81, 64, 52, 56, 47, 41, 42, 41, 30, 34, 46, 47, 42, 36, 32, 30, 32, 36, 42, 46, 44, 46, 49, 54, 58, 59, 53, 41, 36, 25, 22, 0, 31, 9, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 38, 41, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 5, 0, 0, 0, 0, 0, 0, 0, 37, 70, 37, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 28, 0, 0, 0, 0, 0, 0, 0, 24, 78, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 55, 40, 0, 0, 0, 0, 0, 0, 0, 0, 60, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 1, 0, 0, 0, 0, 0, 0, 0, 0, 27, 89, 53, 0, 0, 0, 0, 0, 0, 0, 0, 17, 63, 27, 0, 0, 0, 0, 0, 0, 0, 0, 8, 28, 0, 0, 0, 0, 0, 0, 0, 0, 20, 105, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 0, 0, 0, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 103, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 109, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 98, 17, 0, 0, 0, 0, 0, 0, 0, 0, 11, 46, 0, 0, 0, 0, 0, 6, 32, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 3, 0, 24, 52, 79, 29, 0, 0, 0, 42, 109, 87, 1, 0, 0, 27, 77, 107, 90, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 58, 155, 211, 165, 111, 35, 8, 51, 104, 137, 133, 97, 98, 133, 182, 218, 218, 179, 99, 43, 37, 36, 63, 62, 26, 0, 0, 0, 0, 29, 0, 0, 0, 109, 191, 194, 144, 65, 13, 16, 59, 121, 173, 204, 226, 244, 258, 274, 280, 269, 232, 197, 193, 195, 203, 140, 96, 75, 12, 0, 9, 8, 0, 0, 0, 28, 115, 174, 166, 126, 97, 89, 119, 165, 212, 246, 271, 285, 290, 291, 296, 300, 295, 288, 291, 289, 279, 188, 160, 194, 98, 36, 27, 0, 0, 0, 0, 58, 152, 216, 240, 230, 222, 213, 220, 240, 260, 277, 289, 298, 303, 305, 307, 311, 313, 314, 319, 312, 307, 208, 179, 289, 237, 153, 110, 0, 0, 0, 31, 125, 207, 252, 272, 272, 268, 265, 267, 275, 286, 296, 306, 314, 320, 321, 318, 316, 317, 321, 330, 322, 318, 225, 161, 307, 324, 296, 225, 23, 0, 28, 105, 194, 249, 271, 277, 277, 274, 273, 276, 285, 295, 306, 316, 321, 323, 323, 320, 319, 320, 324, 329, 315, 297, 213, 152, 290, 341, 382, 335, 102, 0, 64, 135, 234, 277, 277, 279, 282, 282, 279, 279, 285, 294, 305, 314, 317, 314, 312, 317, 327, 336, 338, 335, 306, 264, 184, 148, 285, 333, 391, 392, 199, 40, 57, 140, 232, 273, 270, 273, 283, 288, 286, 283, 284, 290, 300, 310, 315, 311, 305, 311, 327, 343, 352, 348, 320, 269, 182, 148, 278, 315, 355, 369, 281, 128, 103, 159, 230, 259, 251, 250, 257, 270, 277, 279, 279, 283, 294, 302, 304, 303, 295, 293, 305, 327, 347, 354, 340, 291, 195, 125, 237, 276, 296, 301, 277, 207, 178, 193, 232, 244, 233, 218, 213, 216, 217, 220, 227, 240, 258, 269, 272, 274, 270, 262, 262, 272, 288, 300, 297, 271, 186, 41, 79, 106, 114, 114, 111, 93, 85, 91, 105, 114, 109, 101, 96, 93, 86, 74, 65, 63, 72, 86, 101, 115, 119, 96, 65, 55, 69, 97, 110, 108, 94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 61, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 156, 169, 139, 94, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 121, 149, 145, 133, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 73, 82, 41, 0, 0, 0, 59, 108, 105, 91, 99, 47, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 138, 137, 48, 0, 0, 0, 0, 67, 71, 67, 90, 91, 0, 0, 0, 0, 0, 0, 42, 158, 92, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 64, 115, 118, 26, 0, 0, 0, 0, 60, 82, 98, 114, 138, 68, 0, 0, 0, 0, 0, 38, 166, 84, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 32, 83, 95, 15, 0, 0, 0, 0, 85, 110, 129, 136, 156, 124, 15, 0, 0, 0, 0, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 63, 91, 22, 0, 0, 0, 0, 65, 96, 117, 122, 141, 148, 95, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 68, 104, 36, 3, 0, 0, 0, 30, 75, 92, 92, 119, 148, 150, 104, 35, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 63, 100, 39, 0, 0, 0, 0, 27, 76, 96, 94, 110, 145, 170, 142, 69, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 52, 13, 0, 0, 0, 0, 52, 113, 130, 124, 125, 137, 153, 122, 44, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 116, 122, 104, 90, 82, 94, 66, 0, 20, 0, 0, 0, 0, 54, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 89, 79, 26, 6, 3, 15, 0, 0, 0, 0, 0, 0, 0, 73, 70, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 18, 0, 0, 0, 0, 0, 32, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 88, 31, 0, 23, 0, 0, 0, 0, 0, 11, 64, 81, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 101, 48, 0, 9, 35, 0, 0, 0, 0, 22, 92, 113, 66, 1, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 69, 0, 0, 49, 29, 11, 0, 25, 18, 74, 131, 79, 10, 0, 4, 10, 27, 46, 66, 54, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 74, 0, 19, 133, 174, 169, 130, 84, 13, 15, 132, 127, 74, 50, 55, 88, 138, 167, 169, 139, 85, 32, 13, 0, 0, 14, 0, 0, 0, 0, 3, 74, 78, 0, 0, 128, 211, 174, 101, 0, 0, 0, 47, 142, 153, 164, 191, 240, 273, 272, 246, 218, 181, 154, 158, 146, 99, 87, 0, 0, 0, 0, 3, 87, 59, 0, 0, 0, 102, 69, 0, 0, 0, 0, 2, 130, 199, 245, 269, 284, 285, 274, 258, 244, 239, 244, 259, 250, 189, 135, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 54, 70, 23, 0, 0, 31, 118, 200, 240, 260, 271, 271, 267, 264, 266, 271, 273, 277, 285, 273, 213, 164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 160, 171, 187, 190, 202, 226, 248, 260, 268, 270, 274, 278, 281, 287, 291, 291, 290, 298, 289, 234, 191, 0, 45, 16, 0, 0, 0, 0, 0, 0, 74, 166, 218, 247, 253, 251, 252, 261, 270, 275, 278, 281, 287, 292, 292, 288, 282, 277, 280, 295, 292, 224, 188, 56, 165, 151, 11, 0, 0, 0, 0, 51, 177, 209, 251, 270, 274, 270, 265, 266, 272, 276, 280, 282, 282, 279, 277, 275, 274, 275, 283, 294, 276, 180, 162, 63, 215, 248, 120, 0, 0, 0, 0, 118, 208, 222, 256, 277, 288, 283, 274, 266, 264, 268, 275, 278, 275, 269, 267, 272, 281, 294, 303, 295, 263, 171, 149, 63, 228, 290, 211, 51, 0, 0, 0, 156, 205, 206, 227, 249, 272, 278, 273, 268, 270, 277, 285, 291, 286, 273, 266, 275, 294, 319, 333, 327, 300, 209, 149, 51, 219, 292, 259, 167, 58, 13, 75, 222, 220, 203, 198, 209, 222, 230, 233, 236, 247, 266, 289, 304, 298, 281, 265, 262, 273, 311, 344, 348, 316, 231, 154, 0, 109, 183, 181, 150, 112, 99, 127, 174, 155, 132, 117, 118, 118, 110, 94, 84, 94, 121, 156, 189, 197, 177, 138, 104, 95, 133, 195, 235, 228, 170, 114, 0, 0, 43, 40, 37, 34, 32, 41, 57, 49, 33, 24, 23, 21, 15, 2, 0, 0, 0, 14, 41, 51, 38, 5, 0, 0, 0, 25, 71, 78, 54, 47, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 9, 9, 8, 4, 0, 0, 0, 1, 5, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 18, 16, 18, 15, 12, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 21, 25, 31, 36, 35, 32, 33, 11, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 15, 13, 4, 0, 10, 26, 41, 51, 50, 50, 35, 5, 0, 0, 0, 12, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 30, 35, 26, 0, 0, 0, 11, 28, 38, 49, 44, 43, 17, 0, 0, 0, 2, 3, 2, 23, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 42, 57, 52, 24, 0, 0, 0, 4, 30, 36, 48, 41, 41, 23, 0, 0, 0, 0, 0, 0, 25, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 58, 57, 21, 0, 0, 0, 0, 33, 42, 51, 47, 36, 30, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 46, 50, 25, 0, 0, 0, 0, 16, 39, 47, 53, 37, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 35, 12, 0, 0, 0, 0, 5, 36, 45, 43, 40, 29, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 0, 0, 0, 0, 0, 4, 37, 50, 42, 37, 36, 33, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 43, 54, 51, 38, 43, 43, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 54, 65, 61, 50, 44, 31, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 54, 65, 61, 49, 41, 22, 5, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 41, 51, 47, 38, 36, 15, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 12, 29, 26, 12, 0, 0, 0, 0, 15, 34, 30, 35, 29, 27, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 10, 21, 39, 47, 29, 12, 6, 0, 3, 14, 26, 31, 40, 27, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 5, 2, 0, 0, 0, 9, 6, 32, 45, 16, 16, 21, 14, 12, 25, 39, 45, 26, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 13, 0, 0, 0, 0, 30, 32, 30, 32, 27, 15, 17, 34, 46, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 10, 29, 23, 31, 24, 8, 4, 14, 27, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 35, 21, 15, 10, 0, 0, 0, 14, 21, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 7, 0, 0, 0, 0, 0, 0, 10, 20, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 77, 0, 9, 0, 0, 0, 0, 0, 0, 0, 3, 2, 7, 9, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 34, 0, 0, 98, 0, 41, 20, 30, 35, 21, 9, 6, 27, 21, 0, 19, 56, 50, 39, 20, 2, 0, 0, 0, 0, 19, 31, 31, 18, 2, 0, 43, 76, 0, 0, 89, 0, 24, 7, 19, 29, 14, 0, 11, 72, 52, 0, 0, 54, 56, 25, 0, 0, 7, 0, 0, 0, 0, 0, 0, 19, 20, 10, 43, 72, 0, 0, 94, 0, 32, 5, 5, 22, 13, 0, 21, 130, 120, 0, 0, 17, 42, 13, 0, 35, 70, 12, 0, 0, 0, 0, 0, 0, 26, 43, 61, 68, 0, 0, 88, 0, 69, 35, 0, 7, 14, 0, 4, 109, 133, 0, 0, 0, 0, 0, 0, 53, 121, 41, 0, 0, 0, 0, 0, 0, 0, 57, 99, 77, 0, 0, 45, 0, 62, 68, 1, 0, 17, 5, 0, 43, 91, 44, 0, 0, 0, 0, 0, 36, 148, 59, 0, 0, 0, 0, 0, 0, 0, 38, 128, 107, 0, 38, 0, 0, 6, 37, 0, 0, 18, 24, 0, 0, 51, 92, 24, 0, 0, 0, 0, 0, 137, 103, 0, 0, 0, 0, 0, 0, 0, 0, 134, 153, 0, 106, 0, 0, 0, 0, 0, 0, 54, 104, 10, 0, 0, 104, 22, 0, 0, 0, 0, 0, 102, 161, 0, 0, 0, 0, 0, 0, 0, 0, 101, 177, 0, 167, 31, 0, 4, 0, 0, 0, 111, 252, 112, 0, 0, 59, 0, 0, 0, 0, 0, 0, 86, 195, 20, 0, 0, 0, 0, 0, 0, 0, 29, 158, 27, 186, 80, 0, 37, 0, 0, 0, 105, 346, 243, 0, 0, 37, 0, 0, 0, 0, 0, 0, 145, 226, 0, 0, 0, 0, 6, 0, 0, 0, 0, 87, 40, 161, 86, 0, 71, 0, 0, 0, 0, 274, 309, 0, 0, 75, 2, 0, 0, 0, 0, 0, 225, 246, 0, 0, 0, 0, 9, 0, 0, 0, 0, 13, 5, 134, 74, 7, 82, 0, 0, 0, 0, 112, 242, 0, 0, 136, 42, 0, 0, 0, 0, 0, 271, 216, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 134, 92, 39, 51, 0, 0, 29, 0, 0, 140, 30, 17, 123, 23, 0, 0, 0, 0, 0, 272, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 151, 128, 54, 28, 0, 0, 72, 0, 0, 74, 127, 121, 51, 0, 0, 0, 0, 0, 0, 233, 131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 182, 160, 44, 47, 0, 0, 69, 0, 0, 13, 191, 206, 0, 0, 0, 0, 0, 0, 0, 161, 105, 0, 0, 0, 0, 0, 3, 0, 0, 0, 39, 0, 222, 189, 3, 80, 0, 0, 35, 3, 0, 0, 164, 208, 2, 0, 0, 0, 0, 0, 0, 43, 66, 30, 0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 263, 222, 0, 90, 0, 0, 0, 67, 0, 0, 15, 97, 22, 0, 0, 0, 0, 0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 13, 86, 0, 278, 264, 0, 74, 0, 0, 0, 111, 0, 0, 0, 0, 32, 0, 41, 6, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 80, 0, 256, 311, 0, 48, 0, 0, 0, 133, 72, 0, 0, 0, 35, 53, 132, 33, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 76, 0, 222, 360, 0, 15, 0, 0, 0, 188, 147, 0, 0, 0, 37, 94, 159, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 0, 211, 408, 0, 0, 0, 0, 0, 291, 233, 0, 0, 0, 28, 101, 130, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 213, 434, 52, 0, 0, 0, 0, 344, 269, 0, 0, 0, 5, 67, 87, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 191, 363, 122, 74, 0, 0, 39, 318, 164, 0, 0, 0, 0, 12, 25, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167, 223, 82, 129, 19, 0, 168, 275, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 186, 123, 0, 71, 45, 90, 310, 193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 15, 0, 0, 223, 116, 0, 0, 21, 219, 418, 114, 0, 0, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 28, 6, 0, 0, 242, 150, 0, 0, 0, 210, 428, 99, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 35, 12, 0, 0, 0, 248, 166, 0, 0, 0, 82, 306, 95, 0, 0, 2, 9, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 23, 45, 27, 0, 0, 0, 0, 249, 169, 0, 0, 0, 0, 109, 49, 0, 0, 0, 10, 8, 0, 0, 0, 0, 9, 14, 5, 0, 0, 0, 0, 28, 77, 70, 0, 0, 0, 0, 0, 246, 179, 0, 0, 0, 0, 0, 8, 0, 0, 0, 20, 23, 12, 5, 16, 45, 61, 56, 25, 0, 0, 0, 8, 80, 128, 81, 0, 0, 0, 0, 0, 163, 138, 0, 8, 5, 0, 0, 3, 0, 0, 7, 20, 20, 17, 14, 25, 53, 72, 75, 52, 7, 0, 0, 18, 77, 120, 88, 4, 0, 0, 0, 0, 37, 27, 13, 21, 23, 25, 25, 25, 26, 27, 27, 27, 28, 28, 26, 24, 26, 28, 27, 24, 21, 21, 21, 21, 19, 20, 22, 22, 24, 21, 16, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 17, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 31, 34, 0, 0, 0, 0, 0, 2, 0, 0, 0, 16, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 19, 38, 39, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 20, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 26, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 6, 7, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 9, 21, 13, 0, 0, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 18, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 14, 10, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 9, 16, 17, 19, 18, 18, 19, 16, 10, 6, 6, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 17, 0, 0, 0, 3, 12, 19, 22, 24, 25, 23, 17, 11, 8, 7, 9, 12, 4, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 24, 14, 8, 12, 16, 17, 20, 24, 25, 24, 21, 17, 10, 3, 3, 9, 15, 13, 0, 0, 0, 28, 26, 0, 0, 0, 0, 0, 0, 0, 0, 28, 20, 13, 10, 13, 19, 22, 24, 24, 22, 18, 15, 13, 10, 9, 13, 18, 15, 0, 0, 0, 0, 24, 32, 2, 8, 0, 0, 0, 0, 0, 2, 26, 20, 14, 10, 11, 15, 20, 23, 22, 18, 16, 14, 14, 17, 24, 28, 23, 6, 0, 0, 0, 5, 23, 28, 1, 19, 0, 0, 0, 0, 0, 7, 27, 23, 15, 11, 12, 15, 20, 20, 17, 13, 10, 12, 18, 26, 34, 33, 16, 0, 0, 0, 0, 10, 24, 24, 0, 15, 5, 0, 0, 0, 0, 5, 24, 18, 11, 8, 11, 14, 16, 15, 11, 4, 0, 1, 11, 19, 25, 19, 0, 0, 0, 0, 0, 7, 7, 14, 7, 20, 19, 9, 0, 0, 5, 15, 22, 18, 14, 13, 17, 20, 20, 17, 10, 4, 2, 8, 20, 29, 24, 9, 0, 0, 0, 9, 7, 17, 0, 0, 23, 28, 27, 27, 23, 17, 20, 22, 23, 20, 18, 19, 21, 17, 14, 10, 8, 10, 17, 26, 28, 23, 13, 2, 1, 15, 30, 32, 31, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 39, 46, 54, 56, 46, 28, 9, 0, 0, 0, 0, 12, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 22, 33, 35, 25, 4, 0, 4, 21, 35, 38, 27, 9, 0, 1, 2, 11, 0, 20, 0, 5, 2, 0, 4, 3, 0, 0, 0, 0, 0, 0, 39, 75, 79, 64, 43, 6, 0, 0, 0, 0, 0, 0, 8, 11, 5, 7, 0, 7, 0, 68, 32, 41, 23, 3, 3, 4, 0, 3, 25, 52, 40, 26, 53, 62, 49, 29, 12, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 17, 1, 3, 0, 97, 48, 54, 35, 11, 3, 13, 14, 25, 52, 72, 49, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 20, 13, 3, 0, 53, 4, 21, 4, 0, 0, 18, 28, 34, 43, 36, 15, 0, 0, 0, 0, 0, 0, 21, 15, 0, 0, 0, 3, 0, 0, 4, 16, 27, 28, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 47, 50, 0, 0, 0, 0, 0, 0, 0, 20, 33, 41, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 34, 23, 0, 0, 0, 0, 0, 0, 0, 7, 48, 55, 55, 0, 28, 0, 0, 0, 0, 0, 12, 39, 13, 0, 0, 0, 0, 0, 0, 0, 3, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 46, 56, 0, 44, 0, 0, 0, 0, 0, 23, 87, 94, 35, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 26, 0, 38, 0, 0, 0, 0, 0, 10, 56, 97, 55, 0, 0, 0, 0, 0, 0, 0, 0, 17, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 5, 19, 59, 10, 0, 0, 0, 0, 0, 0, 0, 0, 24, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 10, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 13, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 53, 75, 65, 29, 9, 17, 5, 0, 0, 10, 34, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 35, 83, 65, 20, 0, 0, 0, 0, 0, 0, 0, 25, 18, 0, 2, 14, 3, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 10, 0, 0, 21, 39, 37, 10, 0, 0, 0, 0, 0, 0, 0, 0, 20, 11, 14, 1, 0, 0, 0, 0, 0, 2, 6, 63, 0, 0, 0, 0, 0, 4, 0, 0, 10, 44, 38, 0, 0, 0, 0, 0, 18, 12, 0, 1, 9, 20, 25, 10, 0, 0, 0, 0, 17, 13, 6, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 32, 3, 0, 0, 0, 0, 7, 8, 14, 22, 30, 26, 4, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 61, 92, 92, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 132, 83, 14, 0, 0, 0, 0, 0, 35, 21, 18, 31, 57, 73, 61, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 88, 105, 95, 41, 0, 0, 0, 15, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 33, 88, 80, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 72, 64, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 95, 120, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 0, 0, 0, 0, 0, 0, 78, 146, 122, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 4, 60, 56, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 43, 0, 3, 0, 0, 15, 11, 0, 0, 3, 19, 28, 31, 31, 29, 24, 20, 12, 0, 0, 0, 0, 11, 21, 25, 11, 0, 0, 0, 0, 0, 75, 105, 76, 66, 58, 46, 42, 35, 27, 26, 29, 37, 42, 45, 48, 57, 73, 87, 95, 93, 78, 62, 62, 74, 99, 129, 133, 107, 65, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 5, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 11, 39, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 37, 18, 4, 0, 0, 0, 0, 0, 0, 0, 0, 17, 8, 0, 0, 0, 0, 42, 0, 10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 45, 10, 0, 0, 0, 29, 0, 43, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 27, 6, 0, 0, 0, 0, 0, 18, 0, 0, 3, 55, 34, 0, 0, 0, 9, 0, 30, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 35, 17, 9, 0, 0, 0, 0, 23, 17, 0, 0, 30, 56, 18, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 40, 35, 23, 14, 0, 0, 0, 6, 37, 0, 0, 0, 54, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 40, 49, 53, 25, 0, 0, 0, 6, 50, 3, 0, 0, 26, 64, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 36, 39, 72, 24, 0, 0, 0, 28, 56, 8, 0, 0, 0, 41, 23, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 20, 71, 8, 0, 0, 0, 46, 61, 17, 0, 0, 0, 7, 11, 20, 34, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 63, 0, 0, 0, 0, 47, 52, 18, 0, 0, 0, 0, 0, 9, 52, 0, 0, 0, 0, 90, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 39, 49, 19, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 104, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 21, 51, 19, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 87, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 36, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 0, 48, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 37, 0, 0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 5, 117, 22, 0, 0, 1, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 24, 15, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 96, 38, 0, 0, 32, 60, 15, 0, 0, 0, 0, 64, 26, 0, 0, 0, 0, 12, 18, 9, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 74, 37, 0, 0, 54, 85, 11, 0, 0, 0, 0, 31, 61, 0, 0, 0, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 63, 6, 0, 0, 0, 78, 14, 0, 0, 0, 0, 0, 52, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 94, 71, 0, 0, 0, 0, 0, 7, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 79, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 85, 63, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 105, 0, 0, 9, 1, 0, 0, 0, 0, 47, 89, 70, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 108, 0, 0, 26, 25, 33, 0, 0, 0, 79, 89, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 113, 0, 0, 28, 39, 45, 0, 0, 0, 66, 73, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 114, 0, 0, 13, 33, 45, 0, 0, 0, 30, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 57, 108, 0, 0, 5, 8, 30, 0, 0, 0, 12, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 34, 61, 101, 0, 0, 8, 9, 19, 21, 0, 0, 13, 23, 8, 1, 2, 6, 11, 8, 0, 0, 0, 0, 0, 9, 14, 1, 0, 0, 0, 0, 35, 55, 69, 105, 0, 0, 49, 47, 48, 53, 43, 33, 32, 36, 31, 29, 31, 33, 36, 32, 23, 13, 9, 15, 31, 44, 52, 50, 30, 8, 4, 29, 61, 65, 65, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 61, 29, 0, 128, 156, 157, 155, 143, 140, 140, 137, 127, 127, 151, 170, 158, 157, 165, 163, 147, 123, 106, 96, 86, 82, 89, 96, 95, 95, 97, 100, 113, 158, 65, 36, 219, 252, 266, 271, 257, 255, 252, 245, 218, 204, 246, 282, 268, 265, 280, 278, 244, 190, 148, 123, 112, 116, 131, 150, 164, 169, 168, 173, 193, 235, 102, 54, 239, 265, 272, 288, 289, 289, 286, 277, 247, 231, 285, 305, 287, 286, 298, 286, 226, 154, 94, 49, 7, 2, 28, 72, 110, 132, 155, 168, 204, 257, 122, 72, 256, 256, 244, 262, 284, 292, 291, 280, 263, 268, 323, 315, 280, 268, 241, 211, 155, 77, 23, 0, 0, 0, 0, 0, 12, 59, 95, 139, 194, 264, 130, 89, 268, 224, 200, 233, 271, 287, 288, 279, 274, 283, 318, 302, 242, 183, 118, 79, 52, 3, 0, 0, 0, 0, 0, 0, 0, 0, 51, 106, 181, 267, 139, 78, 212, 144, 118, 185, 253, 278, 284, 285, 295, 266, 221, 213, 172, 90, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 18, 75, 160, 266, 139, 47, 107, 4, 11, 121, 225, 255, 251, 273, 281, 228, 138, 137, 129, 47, 0, 0, 0, 0, 31, 67, 45, 0, 0, 0, 0, 0, 0, 59, 130, 253, 134, 22, 24, 0, 0, 72, 190, 228, 213, 243, 242, 166, 73, 88, 115, 43, 0, 0, 0, 0, 39, 94, 89, 18, 0, 0, 0, 0, 0, 25, 103, 220, 124, 2, 0, 0, 0, 78, 169, 226, 224, 256, 262, 161, 59, 91, 132, 64, 0, 0, 0, 0, 5, 56, 95, 35, 0, 0, 0, 0, 0, 0, 64, 159, 102, 0, 0, 0, 0, 108, 158, 245, 282, 302, 317, 227, 107, 117, 154, 94, 0, 0, 0, 0, 0, 51, 100, 40, 0, 0, 0, 0, 0, 0, 0, 83, 56, 0, 0, 0, 18, 135, 140, 232, 301, 290, 314, 238, 129, 127, 165, 106, 12, 0, 0, 0, 0, 82, 117, 49, 0, 0, 0, 0, 0, 0, 0, 16, 9, 0, 0, 0, 52, 145, 125, 221, 273, 253, 235, 190, 105, 119, 165, 87, 22, 0, 0, 0, 17, 110, 118, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 121, 97, 180, 228, 201, 155, 101, 61, 98, 147, 75, 26, 0, 19, 0, 43, 120, 107, 20, 0, 0, 0, 0, 0, 0, 0, 18, 7, 0, 0, 0, 45, 69, 43, 102, 170, 148, 106, 68, 76, 103, 115, 61, 37, 8, 22, 0, 59, 111, 88, 16, 0, 0, 0, 0, 0, 0, 0, 78, 42, 0, 0, 0, 20, 29, 0, 14, 95, 100, 94, 110, 148, 151, 97, 41, 24, 1, 0, 1, 77, 102, 87, 16, 0, 0, 0, 0, 0, 0, 20, 141, 81, 0, 0, 0, 0, 0, 0, 0, 28, 54, 101, 138, 187, 166, 83, 20, 1, 0, 0, 0, 82, 90, 89, 43, 0, 0, 0, 0, 0, 9, 72, 202, 114, 0, 0, 0, 0, 0, 0, 0, 0, 17, 41, 98, 111, 110, 35, 0, 0, 0, 0, 0, 32, 59, 90, 52, 0, 0, 0, 0, 0, 48, 128, 251, 135, 0, 6, 0, 0, 0, 0, 0, 0, 21, 19, 35, 27, 19, 0, 0, 0, 0, 0, 0, 15, 12, 29, 17, 0, 0, 0, 0, 18, 92, 171, 268, 139, 0, 37, 0, 0, 0, 0, 0, 0, 0, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 36, 14, 0, 0, 0, 0, 0, 0, 34, 107, 171, 231, 106, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 76, 102, 19, 24, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 74, 0, 0, 0, 0, 0, 0, 27, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 56, 0, 0, 0, 0, 0, 0, 75, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 99, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 29, 41, 48, 49, 53, 55, 55, 55, 55, 56, 54, 53, 53, 54, 56, 59, 57, 54, 47, 40, 35, 32, 32, 34, 39, 44, 50, 56, 72, 84, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 74, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 2, 0, 0, 0, 0, 0, 0, 20, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 32, 34, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 11, 17, 19, 15, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 17, 35, 28, 3, 0, 0, 0, 0, 0, 0, 0, 4, 26, 41, 10, 0, 0, 0, 0, 25, 16, 15, 8, 0, 0, 0, 0, 0, 0, 18, 18, 0, 0, 17, 29, 15, 0, 0, 0, 0, 0, 0, 16, 20, 40, 63, 50, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 42, 40, 7, 0, 0, 0, 0, 21, 21, 17, 28, 54, 68, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 65, 70, 39, 10, 0, 0, 0, 0, 0, 0, 4, 27, 59, 56, 33, 20, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 66, 77, 43, 5, 0, 0, 0, 0, 0, 0, 0, 1, 38, 61, 61, 67, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 45, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 55, 69, 83, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 4, 17, 42, 76, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 3, 60, 67, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 57, 0, 0, 0, 0, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 46, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 36, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 34, 6, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 19, 24, 0, 0, 0, 0, 0, 0, 0, 0, 3, 72, 74, 29, 0, 0, 0, 2, 42, 21, 0, 0, 0, 0, 20, 50, 35, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 5, 24, 116, 138, 75, 17, 0, 0, 0, 0, 0, 0, 0, 19, 67, 96, 94, 70, 29, 0, 0, 0, 0, 18, 42, 0, 0, 0, 0, 0, 0, 0, 7, 0, 45, 65, 18, 0, 0, 0, 0, 0, 0, 2, 43, 85, 109, 119, 108, 84, 44, 16, 0, 0, 26, 65, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 77, 93, 100, 101, 91, 81, 67, 50, 35, 37, 69, 99, 118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 59, 81, 87, 88, 86, 85, 83, 80, 72, 66, 70, 96, 129, 149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 38, 37, 32, 33, 46, 62, 75, 84, 87, 89, 90, 88, 85, 81, 76, 75, 82, 113, 145, 161, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 26, 57, 69, 73, 71, 68, 72, 81, 87, 90, 91, 91, 89, 85, 78, 75, 75, 78, 83, 110, 130, 136, 0, 57, 63, 18, 0, 0, 0, 0, 0, 26, 54, 67, 74, 81, 85, 82, 81, 84, 88, 90, 89, 87, 80, 73, 70, 74, 82, 84, 79, 92, 95, 104, 0, 71, 97, 62, 8, 0, 0, 0, 0, 28, 56, 62, 65, 76, 83, 84, 83, 84, 86, 87, 86, 82, 76, 71, 74, 86, 95, 92, 82, 88, 90, 100, 0, 67, 105, 89, 46, 0, 0, 0, 0, 38, 61, 54, 55, 63, 70, 73, 75, 77, 81, 85, 88, 87, 81, 78, 82, 94, 99, 99, 99, 109, 108, 110, 0, 41, 78, 78, 58, 2, 0, 0, 2, 50, 53, 40, 35, 38, 45, 47, 45, 45, 49, 59, 69, 73, 72, 67, 65, 62, 61, 74, 88, 101, 103, 104, 0, 0, 29, 39, 33, 10, 0, 0, 21, 41, 39, 24, 15, 14, 17, 16, 11, 7, 7, 11, 20, 31, 36, 31, 17, 2, 0, 1, 29, 56, 68, 73, 0, 0, 0, 5, 4, 2, 0, 0, 15, 28, 27, 18, 11, 7, 4, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 15, 32, 35, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 39, 50, 42, 16, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 57, 58, 36, 15, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 0, 0, 0, 0, 3, 34, 42, 27, 24, 10, 0, 0, 0, 0, 0, 8, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 61, 47, 0, 0, 0, 0, 0, 23, 36, 24, 25, 23, 0, 0, 0, 0, 0, 19, 0, 74, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 62, 44, 0, 0, 0, 0, 0, 22, 41, 37, 33, 29, 11, 0, 0, 0, 0, 16, 0, 86, 30, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 19, 56, 36, 0, 0, 0, 0, 0, 25, 53, 55, 31, 29, 18, 2, 0, 0, 0, 6, 0, 58, 9, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 12, 49, 29, 1, 0, 0, 0, 0, 25, 57, 55, 24, 20, 17, 16, 13, 0, 0, 0, 0, 40, 0, 5, 0, 0, 0, 0, 0, 0, 1, 0, 0, 4, 40, 21, 1, 0, 0, 0, 0, 22, 54, 53, 28, 17, 25, 25, 37, 0, 0, 0, 0, 23, 0, 16, 16, 0, 0, 0, 0, 0, 0, 0, 0, 15, 36, 16, 0, 0, 0, 0, 0, 28, 57, 55, 34, 21, 20, 28, 42, 0, 0, 0, 0, 14, 0, 23, 33, 0, 0, 0, 0, 0, 0, 0, 0, 25, 27, 4, 0, 0, 0, 0, 0, 35, 62, 60, 37, 22, 17, 23, 28, 0, 0, 1, 0, 15, 0, 29, 43, 0, 0, 0, 0, 0, 0, 0, 0, 29, 23, 9, 0, 0, 0, 0, 0, 18, 54, 55, 28, 9, 5, 12, 19, 0, 0, 0, 0, 22, 0, 36, 66, 10, 0, 0, 0, 0, 0, 0, 6, 28, 20, 16, 0, 0, 0, 0, 0, 2, 32, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 30, 78, 47, 0, 0, 0, 0, 0, 0, 8, 18, 11, 16, 14, 0, 0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 7, 74, 63, 0, 1, 0, 0, 0, 0, 0, 11, 7, 26, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 60, 78, 25, 17, 22, 0, 0, 0, 0, 6, 3, 36, 45, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 0, 40, 78, 24, 3, 26, 32, 17, 0, 0, 0, 0, 43, 63, 34, 21, 19, 16, 21, 18, 19, 4, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 0, 24, 72, 16, 0, 17, 65, 66, 41, 20, 6, 0, 36, 68, 57, 44, 51, 44, 46, 54, 59, 46, 33, 25, 31, 36, 0, 0, 0, 0, 2, 24, 0, 24, 66, 0, 0, 19, 93, 90, 69, 17, 0, 0, 31, 91, 94, 80, 74, 84, 90, 89, 91, 87, 86, 84, 88, 93, 29, 32, 0, 0, 0, 11, 4, 40, 57, 0, 0, 0, 65, 81, 54, 12, 11, 20, 50, 84, 104, 105, 100, 92, 83, 79, 84, 97, 107, 111, 120, 116, 44, 36, 0, 0, 0, 0, 0, 25, 21, 0, 0, 3, 64, 75, 40, 25, 32, 50, 68, 87, 92, 87, 78, 72, 71, 70, 71, 76, 85, 93, 97, 94, 28, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 84, 79, 74, 73, 78, 80, 81, 82, 77, 72, 68, 67, 68, 67, 67, 69, 76, 79, 77, 76, 7, 17, 32, 0, 23, 0, 0, 0, 0, 0, 6, 91, 83, 82, 75, 76, 76, 71, 68, 68, 68, 66, 66, 67, 68, 68, 70, 72, 74, 70, 64, 67, 7, 27, 43, 21, 46, 0, 0, 0, 0, 0, 44, 104, 74, 65, 63, 65, 64, 62, 62, 63, 64, 64, 65, 66, 66, 66, 69, 71, 69, 62, 57, 62, 10, 30, 39, 28, 71, 17, 0, 0, 0, 0, 73, 100, 68, 61, 61, 66, 67, 65, 62, 60, 60, 61, 62, 62, 61, 62, 66, 68, 65, 62, 62, 64, 12, 22, 37, 27, 78, 45, 0, 0, 0, 9, 83, 84, 52, 46, 51, 60, 65, 65, 61, 58, 59, 61, 63, 63, 62, 61, 58, 55, 60, 66, 69, 67, 22, 22, 28, 17, 71, 58, 32, 24, 39, 47, 84, 67, 44, 36, 37, 40, 42, 44, 44, 48, 55, 60, 64, 66, 61, 51, 44, 43, 57, 69, 76, 71, 28, 25, 0, 0, 11, 7, 5, 7, 18, 21, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 16, 16, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 313, 266, 132, 114, 98, 110, 111, 99, 97, 108, 119, 118, 115, 121, 120, 103, 87, 83, 90, 95, 98, 117, 147, 159, 148, 126, 111, 103, 95, 43, 0, 0, 451, 404, 220, 210, 186, 201, 199, 177, 177, 194, 195, 157, 135, 171, 201, 180, 151, 146, 159, 163, 155, 173, 226, 275, 289, 275, 248, 214, 178, 81, 0, 0, 476, 461, 272, 275, 245, 256, 256, 235, 244, 278, 263, 136, 45, 124, 232, 235, 206, 210, 225, 197, 125, 90, 138, 226, 308, 353, 363, 333, 271, 143, 0, 0, 475, 478, 315, 338, 294, 288, 288, 272, 295, 367, 366, 161, 0, 50, 225, 265, 258, 284, 299, 214, 59, 0, 0, 74, 182, 288, 388, 436, 387, 215, 0, 0, 443, 457, 355, 433, 366, 302, 285, 274, 300, 395, 435, 241, 0, 0, 134, 203, 226, 279, 312, 199, 0, 0, 0, 0, 13, 117, 288, 448, 468, 290, 0, 0, 340, 341, 318, 503, 449, 329, 285, 273, 273, 332, 388, 289, 48, 0, 0, 69, 139, 230, 312, 206, 0, 0, 0, 0, 0, 0, 133, 382, 504, 372, 0, 0, 194, 121, 139, 435, 444, 331, 294, 277, 217, 183, 233, 262, 115, 0, 0, 0, 60, 178, 314, 278, 16, 0, 0, 0, 0, 0, 0, 246, 463, 436, 65, 0, 72, 0, 0, 287, 327, 271, 307, 310, 159, 0, 0, 114, 89, 0, 0, 0, 40, 160, 323, 372, 126, 0, 0, 0, 8, 0, 0, 82, 345, 448, 155, 0, 23, 0, 0, 133, 143, 161, 318, 402, 200, 0, 0, 0, 0, 0, 0, 0, 0, 111, 291, 394, 176, 0, 0, 0, 7, 0, 0, 0, 171, 375, 212, 0, 34, 0, 0, 32, 0, 33, 302, 500, 350, 0, 0, 0, 0, 0, 0, 0, 0, 34, 240, 358, 142, 0, 0, 0, 0, 3, 0, 0, 0, 216, 187, 0, 64, 0, 0, 0, 0, 0, 222, 480, 481, 72, 0, 0, 0, 0, 0, 0, 0, 0, 195, 302, 40, 0, 0, 0, 23, 72, 0, 0, 0, 43, 79, 0, 75, 0, 0, 0, 0, 0, 155, 335, 488, 292, 0, 0, 0, 0, 0, 0, 0, 0, 164, 251, 0, 0, 0, 0, 53, 133, 24, 0, 0, 0, 0, 0, 75, 0, 0, 0, 0, 44, 173, 216, 399, 434, 211, 118, 0, 0, 0, 0, 0, 0, 151, 222, 0, 0, 0, 0, 43, 146, 96, 0, 0, 0, 0, 0, 83, 0, 0, 0, 0, 82, 228, 144, 295, 467, 358, 153, 0, 0, 0, 0, 0, 0, 188, 234, 0, 0, 0, 0, 18, 144, 142, 54, 0, 0, 0, 0, 88, 0, 0, 0, 0, 0, 249, 125, 203, 449, 438, 130, 0, 0, 0, 0, 0, 5, 253, 275, 0, 0, 0, 0, 38, 184, 199, 137, 93, 52, 0, 0, 80, 0, 0, 0, 0, 0, 205, 125, 105, 373, 460, 174, 0, 0, 0, 56, 58, 133, 296, 308, 102, 0, 0, 0, 72, 246, 283, 241, 212, 157, 0, 0, 73, 0, 0, 0, 0, 0, 103, 123, 0, 196, 362, 239, 13, 0, 29, 77, 95, 206, 282, 264, 197, 25, 0, 0, 134, 307, 357, 328, 289, 203, 0, 0, 92, 0, 0, 0, 0, 0, 0, 98, 0, 0, 188, 271, 202, 99, 23, 0, 0, 184, 258, 168, 151, 90, 0, 2, 172, 319, 394, 376, 313, 199, 0, 0, 160, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 190, 278, 183, 0, 0, 0, 44, 223, 130, 65, 65, 27, 52, 170, 310, 404, 384, 297, 171, 0, 0, 241, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 168, 110, 0, 0, 0, 0, 73, 67, 3, 0, 0, 0, 59, 212, 329, 321, 239, 120, 0, 0, 289, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 77, 24, 0, 0, 0, 275, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 154, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 11, 13, 0, 0, 0, 0, 24, 135, 51, 5, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 38, 47, 0, 0, 0, 0, 0, 60, 27, 15, 41, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 72, 61, 0, 0, 0, 0, 0, 1, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 49, 17, 0, 0, 0, 0, 0, 0, 0, 13, 96, 86, 0, 0, 0, 0, 0, 13, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 75, 24, 0, 0, 0, 0, 0, 0, 0, 74, 107, 47, 0, 0, 0, 0, 0, 9, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 93, 106, 60, 0, 0, 0, 0, 0, 0, 0, 77, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 129, 126, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 164, 150, 139, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 175, 161, 151, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 160, 150, 142, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 144, 132, 122, 78, 0, 0, 7, 41, 0, 0, 0, 0, 53, 123, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 145, 145, 132, 79, 0, 4, 141, 207, 85, 0, 0, 25, 75, 112, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 114, 150, 165, 118, 43, 84, 244, 292, 166, 17, 0, 0, 2, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 107, 151, 125, 90, 144, 265, 245, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 46, 93, 74, 94, 176, 231, 135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 23, 2, 22, 22, 92, 209, 203, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 4, 20, 43, 79, 0, 0, 16, 4, 0, 10, 86, 219, 160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 18, 48, 69, 89, 0, 0, 11, 4, 16, 11, 61, 169, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 44, 44, 57, 0, 0, 11, 0, 19, 16, 13, 62, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 22, 0, 10, 0, 0, 40, 28, 38, 46, 21, 9, 1, 0, 0, 0, 0, 1, 6, 5, 4, 11, 21, 27, 27, 21, 13, 13, 25, 56, 88, 101, 79, 29, 0, 0, 0, 0, 43, 30, 37, 40, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 35, 49, 48, 34, 24, 28, 44, 81, 124, 124, 80, 21, 0, 0, 0, 0, 13, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 6, 1, 4, 14, 29, 50, 49, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 31, 0, 0, 0, 0, 0, 80, 99, 81, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 60, 0, 0, 0, 0, 0, 0, 55, 55, 48, 17, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 44, 0, 0, 0, 0, 0, 0, 0, 0, 18, 48, 7, 0, 0, 0, 0, 0, 30, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 41, 6, 0, 0, 0, 0, 39, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 60, 0, 0, 0, 0, 0, 0, 0, 0, 41, 55, 14, 6, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 109, 81, 0, 0, 0, 0, 0, 0, 0, 0, 88, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 136, 111, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 67, 159, 142, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 84, 173, 169, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 158, 169, 109, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 116, 143, 110, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 122, 98, 0, 0, 54, 123, 81, 0, 0, 0, 15, 126, 145, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 134, 114, 6, 11, 132, 252, 233, 114, 44, 37, 47, 78, 77, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 132, 135, 58, 91, 214, 295, 237, 104, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 95, 64, 118, 228, 250, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 24, 40, 48, 43, 32, 28, 32, 0, 0, 0, 0, 0, 0, 1, 116, 217, 138, 0, 0, 0, 0, 8, 8, 3, 0, 0, 0, 0, 0, 10, 22, 33, 46, 56, 58, 53, 47, 58, 74, 12, 0, 7, 22, 0, 0, 0, 137, 220, 63, 0, 0, 0, 14, 17, 11, 6, 2, 0, 3, 10, 19, 30, 43, 57, 62, 56, 45, 45, 63, 101, 116, 33, 0, 18, 48, 7, 0, 0, 134, 189, 33, 0, 0, 9, 20, 17, 9, 4, 3, 6, 13, 23, 33, 42, 52, 59, 55, 40, 32, 46, 79, 112, 103, 14, 0, 15, 57, 32, 0, 0, 63, 93, 1, 0, 0, 21, 32, 34, 27, 16, 8, 9, 16, 27, 36, 42, 44, 42, 36, 32, 44, 69, 85, 77, 45, 0, 0, 20, 61, 48, 29, 17, 6, 0, 0, 0, 0, 10, 25, 36, 39, 34, 28, 28, 33, 39, 43, 43, 37, 28, 27, 48, 84, 104, 90, 46, 16, 0, 8, 53, 82, 77, 70, 73, 50, 0, 0, 0, 0, 6, 15, 24, 31, 39, 50, 65, 81, 92, 88, 75, 62, 56, 75, 125, 166, 165, 116, 65, 32, 0, 0, 38, 62, 61, 58, 62, 57, 12, 0, 0, 1, 4, 4, 1, 1, 3, 12, 32, 58, 75, 72, 57, 44, 43, 67, 114, 148, 128, 79, 45, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 39, 92, 103, 78, 34, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 6, 16, 27, 0, 0, 0, 0, 40, 81, 97, 103, 74, 0, 0, 0, 0, 0, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 110, 110, 94, 10, 0, 0, 0, 0, 0, 9, 70, 109, 75, 0, 0, 0, 0, 100, 73, 97, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 141, 124, 94, 0, 0, 0, 0, 0, 0, 0, 8, 109, 128, 41, 0, 0, 0, 87, 117, 197, 121, 0, 0, 0, 0, 0, 7, 63, 10, 0, 0, 43, 79, 50, 36, 0, 0, 0, 0, 0, 0, 0, 0, 96, 165, 117, 0, 0, 0, 29, 60, 146, 69, 0, 0, 0, 0, 0, 0, 80, 47, 0, 0, 0, 28, 6, 17, 28, 0, 0, 0, 0, 14, 0, 0, 69, 171, 175, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 34, 64, 94, 0, 0, 0, 0, 43, 11, 0, 23, 131, 204, 121, 19, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 47, 71, 115, 132, 0, 0, 0, 0, 24, 0, 0, 0, 62, 184, 165, 101, 0, 0, 0, 0, 0, 0, 0, 48, 51, 0, 0, 0, 0, 0, 0, 0, 50, 77, 137, 137, 0, 0, 0, 0, 7, 0, 0, 0, 0, 103, 150, 120, 49, 0, 0, 0, 0, 0, 0, 0, 94, 13, 0, 0, 0, 0, 0, 0, 20, 48, 121, 113, 0, 0, 0, 0, 38, 26, 0, 0, 0, 20, 72, 96, 61, 0, 0, 0, 0, 0, 0, 0, 48, 71, 0, 0, 0, 0, 0, 0, 0, 0, 70, 70, 0, 0, 0, 0, 54, 41, 0, 0, 0, 0, 0, 41, 48, 0, 0, 0, 0, 0, 43, 0, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 0, 0, 0, 0, 36, 16, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 30, 114, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 129, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 0, 0, 0, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 28, 0, 0, 0, 53, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 37, 81, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 49, 0, 0, 0, 87, 74, 0, 0, 0, 0, 36, 36, 0, 0, 0, 0, 32, 89, 107, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 135, 125, 14, 0, 0, 0, 0, 93, 42, 0, 0, 19, 70, 109, 114, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 78, 0, 0, 0, 0, 0, 5, 70, 64, 56, 58, 70, 88, 85, 62, 11, 0, 0, 0, 0, 15, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 31, 54, 46, 31, 15, 8, 11, 0, 0, 0, 0, 9, 48, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 68, 139, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 37, 25, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 79, 73, 51, 0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 2, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 4, 12, 70, 103, 51, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 6, 104, 156, 0, 0, 0, 0, 40, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 37, 150, 89, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 63, 109, 7, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 51, 0, 0, 0, 0, 0, 27, 15, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 22, 20, 11, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 57, 9, 0, 10, 7, 9, 18, 27, 27, 38, 43, 48, 47, 50, 57, 65, 63, 44, 19, 0, 0, 0, 19, 37, 34, 3, 0, 0, 0, 5, 20, 31, 0, 26, 24, 23, 23, 20, 21, 22, 22, 21, 18, 19, 24, 24, 25, 25, 25, 26, 23, 19, 17, 16, 16, 16, 17, 16, 18, 20, 22, 22, 12, 19, 0, 6, 19, 16, 17, 12, 12, 16, 16, 12, 3, 9, 23, 16, 8, 10, 12, 14, 12, 6, 7, 6, 3, 1, 3, 6, 8, 11, 12, 13, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 59, 21, 26, 17, 18, 21, 19, 16, 17, 20, 21, 20, 20, 21, 19, 14, 9, 10, 13, 13, 14, 20, 25, 25, 24, 19, 15, 12, 8, 0, 0, 34, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 71, 10, 23, 8, 11, 16, 10, 8, 17, 45, 46, 3, 0, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 24, 17, 10, 0, 0, 57, 67, 16, 37, 21, 16, 18, 11, 8, 20, 61, 74, 9, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 0, 0, 3, 11, 28, 36, 27, 0, 0, 51, 53, 1, 42, 38, 20, 16, 10, 1, 3, 42, 54, 0, 0, 0, 0, 0, 0, 4, 29, 11, 0, 0, 0, 7, 1, 1, 17, 42, 47, 0, 0, 38, 21, 0, 23, 48, 30, 18, 12, 0, 0, 18, 19, 0, 0, 0, 0, 0, 0, 23, 61, 33, 0, 0, 0, 0, 0, 0, 3, 31, 61, 3, 0, 45, 8, 0, 9, 45, 28, 22, 18, 0, 0, 0, 1, 0, 0, 0, 0, 0, 14, 28, 70, 51, 0, 0, 0, 0, 0, 0, 0, 9, 57, 21, 0, 59, 12, 0, 22, 48, 24, 24, 37, 33, 0, 0, 0, 18, 0, 0, 0, 0, 5, 21, 60, 56, 0, 0, 0, 0, 0, 0, 0, 0, 33, 36, 0, 71, 15, 0, 62, 42, 8, 16, 62, 108, 48, 0, 0, 40, 0, 0, 0, 0, 0, 12, 42, 58, 0, 0, 0, 0, 0, 0, 0, 0, 9, 26, 0, 82, 15, 0, 86, 24, 0, 0, 48, 132, 85, 0, 0, 56, 0, 0, 0, 0, 0, 0, 49, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 25, 0, 93, 0, 0, 0, 19, 105, 102, 0, 0, 64, 0, 0, 0, 0, 0, 0, 59, 99, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 86, 30, 2, 87, 0, 0, 1, 3, 47, 93, 0, 0, 85, 15, 0, 0, 0, 0, 0, 76, 100, 0, 0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 87, 30, 7, 69, 0, 0, 21, 0, 18, 73, 28, 24, 86, 20, 0, 0, 0, 0, 0, 100, 90, 0, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 90, 39, 16, 49, 0, 0, 27, 0, 0, 49, 53, 69, 82, 11, 0, 0, 0, 0, 11, 107, 78, 0, 0, 0, 0, 0, 18, 26, 1, 0, 0, 0, 96, 52, 16, 27, 0, 0, 35, 0, 0, 26, 69, 94, 66, 0, 0, 0, 0, 0, 19, 103, 69, 0, 0, 0, 0, 6, 32, 33, 10, 6, 0, 0, 104, 64, 9, 15, 0, 0, 23, 17, 0, 8, 71, 84, 17, 0, 0, 0, 0, 0, 28, 69, 47, 0, 0, 0, 0, 0, 25, 25, 4, 16, 6, 0, 116, 72, 1, 30, 0, 0, 2, 45, 0, 0, 27, 46, 0, 0, 0, 0, 0, 0, 34, 22, 2, 0, 0, 0, 0, 0, 21, 27, 14, 31, 11, 0, 129, 79, 0, 50, 0, 0, 0, 49, 0, 0, 3, 22, 20, 0, 0, 0, 0, 0, 54, 22, 0, 0, 0, 0, 0, 6, 25, 38, 30, 41, 11, 0, 133, 91, 0, 52, 0, 0, 0, 45, 0, 0, 0, 0, 11, 16, 23, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 12, 33, 49, 37, 33, 0, 0, 122, 102, 0, 37, 0, 0, 0, 60, 3, 0, 0, 0, 10, 43, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 26, 33, 15, 10, 0, 0, 102, 105, 0, 19, 0, 0, 0, 99, 67, 0, 0, 0, 11, 68, 85, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 100, 0, 20, 5, 0, 0, 138, 112, 0, 0, 0, 7, 50, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 71, 0, 26, 14, 0, 35, 155, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 38, 0, 37, 18, 0, 67, 126, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 30, 0, 22, 28, 9, 78, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 22, 0, 4, 14, 31, 108, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 1, 0, 0, 7, 27, 129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 19, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 60, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 9, 2, 0, 0, 0, 1, 31, 53, 28, 0, 0, 0, 0, 0, 45, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 8, 17, 1, 0, 0, 0, 0, 0, 81, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 137, 80, 0, 6, 0, 0, 3, 0, 0, 0, 9, 0, 0, 0, 17, 2, 0, 0, 0, 0, 0, 0, 3, 29, 35, 28, 12, 0, 0, 0, 0, 0, 167, 99, 0, 19, 0, 9, 11, 0, 0, 19, 44, 0, 0, 0, 23, 15, 0, 0, 0, 0, 0, 0, 0, 0, 29, 45, 48, 33, 4, 0, 0, 0, 161, 104, 12, 58, 24, 22, 27, 12, 10, 55, 108, 28, 0, 0, 22, 31, 12, 12, 32, 19, 0, 0, 0, 0, 0, 20, 56, 83, 61, 27, 0, 0, 147, 86, 21, 104, 54, 17, 19, 12, 3, 53, 134, 64, 0, 0, 0, 2, 0, 9, 57, 59, 0, 0, 0, 0, 0, 0, 14, 88, 106, 65, 0, 0, 120, 37, 0, 142, 95, 21, 16, 17, 0, 27, 102, 74, 0, 0, 0, 0, 0, 9, 89, 100, 0, 0, 0, 0, 0, 0, 0, 53, 130, 114, 0, 0, 99, 0, 0, 126, 109, 23, 25, 32, 2, 0, 15, 52, 0, 0, 0, 0, 0, 0, 88, 138, 18, 0, 0, 0, 0, 0, 0, 11, 108, 154, 0, 0, 108, 0, 0, 92, 65, 0, 38, 70, 32, 0, 0, 1, 35, 0, 0, 0, 0, 0, 69, 159, 66, 0, 0, 0, 0, 0, 0, 0, 48, 156, 45, 0, 134, 0, 0, 67, 0, 0, 40, 130, 108, 0, 0, 0, 32, 0, 0, 0, 0, 0, 40, 164, 90, 0, 0, 0, 0, 0, 0, 0, 0, 108, 83, 0, 156, 0, 0, 62, 0, 0, 18, 173, 213, 6, 0, 0, 18, 0, 0, 0, 0, 0, 25, 176, 107, 0, 0, 0, 0, 0, 0, 0, 0, 39, 60, 0, 172, 0, 0, 66, 0, 0, 0, 141, 294, 126, 0, 0, 24, 0, 0, 0, 0, 0, 29, 200, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 175, 1, 31, 47, 0, 0, 0, 55, 252, 212, 0, 0, 42, 0, 0, 0, 0, 0, 45, 237, 94, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 168, 13, 44, 16, 0, 0, 0, 0, 137, 221, 20, 5, 42, 0, 0, 0, 0, 0, 65, 257, 67, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 175, 27, 35, 0, 0, 0, 46, 0, 37, 183, 111, 62, 19, 0, 0, 0, 0, 0, 72, 242, 38, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 194, 40, 16, 0, 0, 0, 81, 0, 0, 142, 191, 120, 0, 0, 0, 0, 0, 0, 71, 205, 37, 0, 0, 0, 0, 19, 24, 0, 0, 0, 0, 0, 225, 46, 0, 0, 0, 0, 83, 0, 0, 83, 239, 161, 0, 0, 0, 0, 0, 0, 57, 138, 43, 0, 0, 0, 0, 37, 50, 14, 0, 0, 0, 0, 259, 52, 0, 0, 0, 0, 58, 24, 0, 0, 161, 158, 0, 0, 0, 0, 0, 0, 43, 38, 26, 0, 0, 0, 0, 46, 61, 30, 0, 1, 0, 0, 289, 67, 0, 9, 0, 0, 23, 76, 0, 0, 32, 84, 27, 0, 0, 0, 0, 6, 57, 0, 0, 0, 0, 0, 0, 39, 64, 49, 0, 13, 0, 0, 311, 102, 0, 8, 0, 0, 0, 103, 0, 0, 0, 12, 68, 22, 16, 0, 0, 0, 60, 0, 0, 0, 0, 0, 0, 45, 77, 61, 3, 11, 0, 0, 320, 152, 0, 0, 0, 0, 0, 141, 0, 0, 0, 0, 66, 76, 55, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 27, 77, 59, 0, 0, 0, 0, 316, 202, 0, 0, 0, 0, 0, 195, 19, 0, 0, 0, 60, 100, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 27, 0, 0, 0, 0, 297, 238, 0, 0, 0, 0, 17, 217, 41, 0, 0, 0, 75, 114, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 248, 251, 48, 17, 0, 0, 66, 207, 12, 0, 0, 0, 42, 77, 59, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 1, 0, 0, 0, 0, 0, 0, 172, 189, 102, 100, 0, 0, 123, 150, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 6, 7, 9, 10, 4, 0, 0, 0, 8, 0, 0, 104, 88, 64, 141, 81, 66, 178, 55, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 3, 12, 10, 8, 9, 10, 4, 1, 6, 7, 21, 0, 0, 86, 17, 0, 81, 125, 202, 241, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 4, 9, 12, 12, 12, 11, 5, 0, 0, 12, 16, 22, 0, 0, 96, 19, 0, 9, 89, 269, 269, 0, 0, 0, 0, 23, 6, 0, 0, 0, 0, 3, 7, 10, 10, 9, 12, 10, 0, 0, 3, 20, 16, 8, 0, 0, 103, 30, 0, 0, 28, 210, 250, 0, 0, 0, 16, 27, 10, 0, 0, 0, 2, 8, 10, 9, 4, 2, 5, 8, 7, 8, 17, 24, 4, 0, 0, 0, 107, 32, 0, 0, 0, 96, 157, 0, 0, 0, 14, 22, 13, 0, 0, 0, 9, 15, 14, 9, 0, 0, 0, 8, 23, 34, 33, 14, 0, 0, 0, 0, 110, 33, 0, 0, 0, 13, 56, 0, 0, 0, 9, 20, 16, 6, 0, 5, 19, 25, 21, 6, 0, 0, 0, 13, 45, 64, 36, 0, 0, 0, 0, 0, 99, 38, 0, 13, 3, 0, 4, 0, 0, 0, 6, 15, 14, 10, 10, 22, 37, 42, 38, 18, 0, 0, 0, 23, 68, 81, 41, 0, 0, 0, 0, 0, 62, 23, 0, 9, 7, 0, 0, 0, 0, 0, 4, 6, 5, 3, 2, 12, 25, 29, 28, 15, 0, 0, 0, 13, 46, 59, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 30, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 43, 0, 0, 0, 4, 0, 0, 127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 77, 34, 0, 0, 0, 0, 0, 103, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 31, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 103, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 46, 0, 31, 11, 0, 0, 0, 19, 53, 0, 0, 0, 52, 116, 36, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 99, 83, 24, 105, 61, 0, 0, 0, 62, 75, 0, 0, 0, 0, 84, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 95, 105, 34, 152, 97, 0, 0, 0, 82, 71, 0, 0, 0, 0, 14, 36, 10, 15, 0, 0, 0, 0, 35, 0, 0, 10, 0, 0, 0, 0, 0, 0, 35, 70, 14, 149, 78, 0, 0, 0, 81, 46, 0, 0, 0, 0, 0, 0, 7, 50, 0, 0, 0, 0, 144, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 32, 0, 0, 0, 66, 39, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 224, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 26, 46, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 242, 214, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 198, 277, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 9, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 116, 294, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 21, 252, 106, 0, 0, 0, 37, 0, 0, 0, 0, 0, 105, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 187, 100, 0, 0, 85, 174, 34, 0, 0, 0, 0, 160, 150, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 0, 152, 65, 0, 0, 149, 289, 131, 0, 0, 0, 0, 123, 169, 48, 0, 0, 0, 0, 7, 28, 5, 0, 0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 101, 10, 0, 0, 146, 325, 212, 20, 0, 0, 0, 64, 114, 54, 2, 0, 0, 10, 26, 41, 45, 4, 0, 0, 0, 12, 146, 2, 0, 0, 0, 0, 30, 0, 0, 0, 121, 308, 196, 41, 0, 0, 0, 0, 39, 48, 38, 24, 24, 30, 39, 50, 62, 56, 32, 23, 56, 117, 226, 24, 0, 24, 0, 0, 0, 0, 0, 0, 130, 210, 115, 34, 11, 18, 5, 5, 25, 40, 39, 36, 42, 51, 55, 60, 70, 78, 73, 69, 96, 166, 273, 0, 87, 193, 44, 0, 0, 0, 0, 0, 186, 132, 62, 51, 63, 74, 63, 53, 50, 47, 44, 46, 56, 64, 67, 68, 75, 79, 72, 67, 97, 180, 308, 0, 63, 261, 196, 149, 0, 0, 0, 166, 224, 92, 36, 46, 68, 69, 56, 51, 52, 53, 53, 56, 62, 67, 73, 81, 86, 79, 61, 56, 96, 188, 316, 0, 12, 212, 254, 292, 50, 0, 0, 239, 215, 50, 26, 51, 76, 77, 63, 55, 53, 53, 57, 63, 70, 71, 74, 84, 87, 76, 60, 67, 120, 194, 294, 0, 0, 173, 207, 324, 190, 0, 0, 193, 151, 26, 17, 42, 68, 78, 73, 62, 55, 56, 61, 70, 78, 78, 75, 74, 72, 72, 82, 112, 157, 195, 260, 0, 0, 153, 151, 237, 239, 21, 4, 114, 92, 30, 26, 34, 50, 62, 64, 55, 51, 56, 65, 80, 89, 86, 74, 55, 47, 62, 103, 147, 186, 204, 239, 0, 0, 127, 99, 141, 171, 101, 45, 61, 62, 42, 44, 46, 51, 56, 54, 37, 24, 25, 40, 69, 83, 78, 60, 23, 0, 21, 91, 152, 181, 190, 221, 0, 0, 111, 85, 96, 112, 97, 68, 63, 63, 62, 67, 68, 69, 77, 78, 61, 42, 30, 34, 61, 78, 86, 92, 61, 18, 13, 68, 119, 130, 140, 166, 0, 0, 46, 30, 33, 38, 34, 23, 22, 24, 26, 30, 33, 35, 39, 37, 26, 11, 0, 0, 14, 30, 40, 44, 29, 0, 0, 12, 42, 41, 51, 75, 25, 112, 115, 107, 102, 96, 97, 97, 95, 92, 93, 96, 99, 101, 103, 106, 102, 92, 85, 83, 83, 79, 79, 84, 91, 92, 90, 86, 81, 67, 67, 13, 32, 182, 179, 178, 176, 173, 177, 178, 176, 172, 172, 174, 169, 158, 166, 179, 178, 170, 159, 149, 137, 121, 115, 124, 139, 152, 161, 167, 165, 150, 145, 55, 4, 155, 137, 139, 137, 135, 142, 144, 141, 137, 134, 161, 157, 116, 118, 138, 142, 130, 104, 81, 63, 46, 32, 35, 48, 68, 95, 119, 136, 132, 143, 48, 3, 162, 149, 154, 160, 154, 153, 153, 154, 150, 151, 212, 212, 145, 120, 123, 107, 93, 78, 71, 66, 56, 48, 45, 45, 49, 68, 103, 132, 144, 162, 56, 4, 152, 129, 132, 156, 160, 152, 149, 156, 142, 122, 175, 181, 122, 72, 46, 36, 46, 52, 56, 64, 56, 49, 48, 62, 61, 52, 75, 110, 136, 171, 66, 2, 101, 60, 81, 128, 156, 153, 150, 157, 132, 84, 95, 98, 76, 36, 9, 15, 41, 45, 46, 52, 34, 17, 28, 64, 71, 42, 46, 88, 118, 175, 77, 0, 69, 12, 30, 100, 145, 146, 149, 158, 137, 75, 52, 66, 91, 69, 28, 30, 53, 47, 44, 53, 54, 18, 4, 29, 47, 28, 26, 60, 92, 165, 85, 0, 49, 0, 26, 115, 148, 135, 132, 143, 145, 81, 41, 74, 120, 92, 32, 37, 52, 39, 21, 46, 78, 47, 4, 6, 16, 22, 14, 28, 63, 147, 82, 0, 46, 0, 69, 160, 155, 134, 123, 141, 189, 156, 80, 88, 112, 66, 18, 19, 22, 26, 0, 25, 69, 59, 27, 12, 11, 25, 23, 12, 29, 116, 68, 0, 17, 0, 83, 172, 151, 130, 116, 135, 198, 195, 106, 95, 108, 57, 16, 19, 5, 22, 0, 27, 78, 74, 43, 22, 17, 25, 30, 13, 0, 70, 48, 0, 0, 0, 51, 146, 150, 137, 72, 27, 80, 109, 69, 76, 109, 59, 14, 23, 7, 23, 0, 47, 76, 56, 27, 19, 23, 20, 19, 18, 1, 37, 23, 0, 0, 0, 21, 111, 128, 158, 85, 0, 0, 31, 1, 27, 101, 73, 19, 31, 21, 20, 0, 39, 46, 26, 6, 4, 19, 14, 5, 14, 12, 45, 15, 0, 0, 0, 13, 61, 71, 157, 135, 2, 11, 41, 0, 20, 84, 71, 33, 49, 44, 7, 0, 20, 23, 10, 1, 4, 12, 4, 0, 17, 32, 73, 23, 0, 0, 0, 11, 14, 2, 120, 148, 56, 38, 61, 30, 46, 63, 41, 38, 68, 61, 0, 0, 24, 27, 22, 13, 20, 29, 27, 27, 45, 51, 96, 40, 0, 0, 0, 0, 12, 0, 73, 147, 99, 71, 75, 66, 76, 58, 28, 32, 73, 78, 3, 0, 30, 38, 42, 20, 25, 47, 58, 65, 86, 82, 121, 59, 0, 0, 0, 0, 10, 0, 42, 144, 132, 85, 55, 51, 65, 54, 21, 16, 52, 73, 35, 30, 47, 38, 56, 33, 29, 47, 56, 70, 95, 94, 140, 69, 0, 0, 0, 0, 0, 0, 6, 105, 136, 72, 0, 0, 0, 16, 14, 25, 34, 50, 67, 61, 23, 29, 60, 44, 28, 36, 46, 72, 109, 114, 162, 74, 0, 0, 0, 0, 0, 0, 0, 46, 111, 79, 5, 0, 6, 30, 32, 68, 45, 33, 80, 100, 44, 30, 32, 18, 18, 39, 53, 102, 146, 141, 173, 71, 0, 0, 0, 0, 0, 0, 0, 0, 46, 73, 41, 2, 32, 45, 25, 79, 55, 11, 67, 123, 91, 52, 21, 0, 21, 50, 81, 136, 169, 144, 165, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 19, 0, 0, 0, 0, 32, 30, 0, 13, 39, 33, 22, 0, 0, 0, 24, 64, 110, 135, 103, 119, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 21, 0, 29, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 58, 61, 42, 33, 35, 39, 38, 31, 27, 32, 39, 38, 35, 32, 30, 25, 23, 25, 29, 31, 30, 31, 35, 36, 36, 32, 26, 17, 2, 0, 0, 75, 54, 17, 7, 0, 8, 16, 14, 4, 4, 25, 34, 16, 0, 0, 0, 0, 0, 0, 6, 7, 2, 0, 0, 0, 1, 12, 17, 9, 0, 0, 0, 64, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 8, 0, 0, 0, 0, 0, 0, 0, 0, 27, 52, 0, 0, 0, 0, 0, 0, 0, 4, 33, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 63, 96, 66, 41, 43, 44, 13, 0, 0, 0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 90, 98, 42, 26, 50, 49, 21, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 17, 43, 81, 79, 23, 10, 25, 14, 0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 45, 78, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 39, 24, 20, 33, 39, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 73, 0, 5, 149, 136, 17, 0, 0, 38, 27, 6, 56, 82, 4, 0, 0, 19, 0, 0, 15, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 6, 67, 210, 125, 5, 0, 0, 73, 94, 43, 100, 103, 0, 0, 0, 0, 0, 0, 27, 103, 27, 0, 0, 22, 29, 0, 0, 0, 0, 0, 0, 64, 6, 56, 181, 52, 0, 0, 0, 0, 0, 0, 26, 77, 0, 0, 0, 0, 0, 0, 70, 153, 35, 0, 0, 17, 50, 14, 0, 0, 0, 0, 0, 64, 15, 58, 125, 0, 0, 0, 0, 0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 0, 98, 132, 0, 0, 0, 6, 50, 23, 0, 0, 0, 0, 0, 64, 30, 62, 81, 0, 0, 0, 0, 0, 0, 0, 46, 119, 17, 0, 0, 0, 0, 13, 100, 84, 0, 0, 0, 9, 53, 45, 26, 12, 3, 0, 0, 79, 53, 57, 29, 0, 0, 0, 0, 0, 0, 35, 133, 165, 21, 0, 0, 1, 0, 22, 99, 55, 0, 0, 0, 19, 71, 89, 86, 60, 22, 0, 0, 96, 73, 41, 0, 0, 0, 6, 0, 0, 13, 97, 176, 138, 4, 0, 0, 1, 0, 36, 94, 42, 0, 0, 0, 15, 75, 111, 113, 79, 34, 0, 0, 110, 77, 24, 0, 0, 0, 55, 28, 4, 33, 79, 88, 21, 0, 0, 3, 2, 0, 65, 80, 24, 0, 0, 0, 0, 44, 77, 83, 66, 36, 0, 0, 120, 79, 14, 0, 0, 0, 65, 73, 19, 48, 17, 0, 0, 0, 0, 34, 21, 33, 95, 80, 14, 0, 0, 0, 0, 11, 41, 65, 71, 50, 0, 0, 116, 72, 7, 0, 0, 0, 27, 92, 37, 33, 0, 0, 0, 0, 53, 58, 26, 60, 98, 75, 41, 0, 0, 0, 0, 7, 52, 90, 94, 59, 0, 0, 104, 62, 4, 0, 0, 0, 0, 87, 32, 0, 0, 0, 7, 50, 97, 52, 0, 43, 85, 59, 42, 0, 0, 0, 0, 22, 86, 122, 100, 39, 0, 0, 92, 59, 11, 19, 0, 0, 0, 72, 11, 0, 0, 0, 45, 108, 121, 24, 0, 0, 31, 0, 0, 0, 0, 0, 0, 31, 97, 113, 72, 6, 0, 0, 81, 61, 25, 31, 0, 0, 0, 107, 48, 0, 0, 0, 92, 167, 142, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 58, 66, 31, 0, 0, 0, 51, 40, 21, 35, 0, 0, 13, 175, 122, 0, 0, 0, 63, 77, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 225, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 181, 206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 258, 260, 176, 172, 160, 170, 176, 171, 169, 172, 173, 172, 170, 174, 177, 172, 166, 167, 173, 176, 173, 178, 191, 199, 196, 185, 178, 177, 177, 160, 106, 39, 300, 313, 223, 220, 207, 220, 228, 221, 218, 223, 223, 199, 177, 198, 224, 221, 211, 209, 218, 223, 212, 209, 226, 248, 260, 263, 257, 248, 244, 221, 148, 35, 253, 246, 159, 157, 143, 156, 162, 156, 162, 184, 190, 123, 52, 83, 144, 151, 137, 146, 168, 171, 142, 114, 120, 148, 181, 210, 228, 232, 219, 190, 124, 16, 252, 252, 178, 186, 162, 161, 164, 161, 173, 216, 240, 153, 29, 38, 119, 137, 134, 165, 213, 211, 156, 109, 100, 124, 155, 185, 228, 267, 264, 210, 123, 14, 227, 224, 179, 230, 201, 168, 159, 158, 169, 198, 218, 148, 35, 15, 67, 103, 125, 179, 238, 217, 128, 81, 99, 132, 145, 145, 188, 264, 288, 237, 125, 7, 173, 140, 135, 250, 244, 185, 161, 159, 157, 158, 153, 121, 67, 39, 44, 105, 159, 205, 247, 203, 87, 33, 74, 132, 143, 122, 148, 237, 293, 261, 138, 3, 123, 60, 80, 238, 252, 191, 167, 162, 138, 103, 102, 129, 136, 94, 64, 126, 190, 202, 222, 200, 90, 14, 53, 127, 142, 120, 118, 184, 267, 273, 164, 10, 99, 35, 53, 225, 218, 165, 177, 188, 139, 48, 26, 109, 156, 92, 48, 110, 182, 183, 190, 195, 117, 23, 32, 107, 148, 135, 112, 129, 210, 265, 193, 35, 81, 19, 33, 192, 143, 118, 183, 238, 180, 30, 0, 29, 85, 22, 0, 68, 135, 140, 170, 194, 124, 18, 4, 73, 151, 159, 123, 91, 143, 228, 202, 68, 58, 0, 7, 134, 49, 63, 154, 235, 191, 20, 0, 0, 2, 0, 0, 32, 92, 105, 179, 216, 117, 0, 0, 48, 153, 179, 130, 84, 95, 168, 177, 93, 26, 0, 0, 48, 0, 30, 93, 131, 101, 0, 0, 0, 0, 0, 0, 0, 65, 69, 171, 205, 69, 0, 0, 35, 162, 198, 146, 99, 84, 129, 141, 98, 11, 0, 0, 0, 0, 46, 87, 58, 46, 0, 0, 0, 0, 0, 0, 0, 44, 34, 144, 160, 0, 0, 0, 28, 158, 208, 173, 127, 109, 121, 121, 90, 18, 0, 0, 0, 0, 66, 145, 71, 79, 80, 17, 18, 0, 0, 0, 0, 32, 16, 112, 109, 0, 0, 0, 42, 152, 209, 195, 155, 134, 134, 123, 73, 30, 0, 0, 0, 0, 52, 199, 108, 115, 173, 146, 65, 0, 0, 0, 0, 35, 19, 103, 96, 0, 0, 0, 56, 159, 224, 222, 184, 160, 155, 131, 52, 28, 0, 0, 0, 0, 17, 201, 148, 136, 211, 208, 53, 0, 0, 0, 35, 68, 63, 134, 123, 0, 0, 0, 54, 165, 234, 234, 200, 182, 182, 151, 39, 9, 0, 0, 0, 0, 0, 172, 177, 125, 168, 162, 16, 0, 0, 0, 86, 112, 137, 169, 135, 53, 2, 8, 42, 151, 223, 230, 210, 205, 210, 155, 22, 0, 0, 0, 0, 0, 0, 111, 179, 89, 86, 80, 0, 0, 0, 71, 112, 130, 188, 197, 130, 93, 78, 56, 56, 149, 221, 242, 243, 238, 220, 141, 0, 0, 0, 0, 0, 0, 0, 29, 140, 66, 33, 49, 59, 89, 114, 116, 85, 79, 183, 232, 139, 103, 104, 80, 101, 181, 244, 281, 283, 251, 206, 117, 0, 3, 0, 0, 0, 0, 0, 0, 54, 0, 0, 9, 110, 183, 186, 96, 0, 0, 100, 211, 175, 129, 105, 99, 141, 202, 265, 305, 289, 234, 179, 101, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 152, 138, 5, 0, 0, 0, 92, 114, 111, 98, 100, 113, 151, 208, 252, 240, 189, 144, 85, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 30, 0, 0, 0, 0, 0, 38, 50, 53, 44, 33, 38, 66, 97, 102, 82, 56, 22, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
