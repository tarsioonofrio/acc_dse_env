LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias

					-- weights

			118, 367, 0, 
			50, 0, 0, 
			158, 305, 176, 
			

			0, 412, 0, 
			14, 177, 193, 
			0, 74, 169, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 297, 
			0, 0, 0, 
			0, 149, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			42, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 5, 138, 
			67, 0, 20, 
			

			0, 276, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 27, 0, 
			0, 90, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 381, 239, 
			61, 326, 106, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 98, 238, 
			121, 133, 82, 
			

			0, 0, 0, 
			0, 0, 99, 
			0, 5, 144, 
			

			0, 57, 0, 
			0, 0, 0, 
			433, 0, 361, 
			

			198, 0, 344, 
			0, 0, 99, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 60, 
			0, 0, 0, 
			0, 83, 148, 
			

			0, 0, 0, 
			0, 0, 0, 
			499, 0, 23, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 296, 270, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 97, 
			0, 197, 0, 
			

			0, 0, 219, 
			183, 341, 0, 
			194, 0, 216, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 21, 
			

			30, 0, 0, 
			0, 0, 0, 
			0, 0, 80, 
			

			36, 0, 0, 
			0, 94, 0, 
			0, 435, 179, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			187, 264, 262, 
			249, 0, 0, 
			0, 0, 0, 
			

			0, 50, 53, 
			520, 86, 5, 
			0, 0, 0, 
			

			0, 0, 0, 
			16, 0, 92, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			201, 354, 50, 
			252, 107, 0, 
			0, 0, 0, 
			

			24, 0, 0, 
			0, 0, 0, 
			352, 578, 539, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 39, 408, 
			0, 0, 0, 
			194, 421, 355, 
			

			0, 217, 0, 
			418, 130, 13, 
			265, 0, 0, 
			

			0, 0, 27, 
			142, 0, 33, 
			0, 0, 0, 
			

			0, 222, 0, 
			0, 0, 0, 
			559, 505, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			545, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 62, 0, 
			

			0, 98, 199, 
			271, 40, 0, 
			0, 0, 0, 
			

			0, 199, 0, 
			285, 215, 249, 
			0, 0, 0, 
			

			121, 16, 190, 
			0, 184, 47, 
			0, 0, 0, 
			

			22, 0, 0, 
			0, 0, 0, 
			0, 24, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			294, 0, 373, 
			272, 0, 131, 
			126, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			485, 166, 0, 
			190, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 41, 77, 
			

			0, 16, 0, 
			54, 388, 325, 
			50, 329, 411, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			16, 258, 0, 
			0, 0, 247, 
			0, 0, 0, 
			

			0, 53, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 12, 60, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			40, 0, 0, 
			325, 0, 94, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 21, 
			167, 341, 0, 
			149, 0, 0, 
			

			0, 0, 0, 
			5, 89, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 84, 
			0, 192, 31, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			272, 0, 204, 
			523, 0, 116, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 148, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			93, 233, 0, 
			53, 410, 0, 
			0, 0, 0, 
			

			422, 603, 0, 
			20, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 3, 0, 
			0, 0, 81, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 281, 0, 
			

			72, 0, 0, 
			0, 0, 105, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 293, 175, 
			

			0, 78, 0, 
			0, 0, 0, 
			0, 323, 388, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 118, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 499, 0, 
			509, 0, 79, 
			0, 0, 0, 
			

			77, 0, 24, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			244, 0, 0, 
			207, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 150, 
			142, 147, 393, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 123, 227, 
			

			3, 121, 105, 
			0, 59, 146, 
			0, 484, 212, 
			

			0, 102, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			85, 0, 0, 
			237, 286, 0, 
			0, 149, 68, 
			

			0, 0, 0, 
			0, 75, 111, 
			493, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			23, 0, 0, 
			0, 208, 204, 
			172, 0, 0, 
			

			191, 0, 235, 
			338, 0, 0, 
			0, 0, 0, 
			

			0, 187, 0, 
			0, 48, 0, 
			163, 564, 35, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			26, 0, 292, 
			0, 57, 0, 
			0, 0, 0, 
			

			416, 0, 196, 
			0, 38, 188, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 213, 
			0, 18, 0, 
			0, 0, 0, 
			

			39, 96, 53, 
			17, 236, 162, 
			105, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			69, 387, 0, 
			424, 341, 490, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 10, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 72, 0, 
			483, 448, 582, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 462, 
			109, 0, 0, 
			

			0, 0, 239, 
			0, 62, 0, 
			0, 0, 32, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 53, 0, 
			0, 31, 0, 
			0, 0, 0, 
			

			0, 230, 0, 
			107, 0, 0, 
			0, 0, 0, 
			

			240, 322, 0, 
			304, 338, 23, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			101, 0, 31, 
			0, 0, 127, 
			0, 12, 0, 
			

			0, 0, 139, 
			0, 0, 0, 
			0, 0, 0, 
			

			198, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 141, 0, 
			0, 37, 152, 
			215, 148, 95, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			208, 0, 24, 
			182, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			136, 0, 148, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 49, 0, 
			0, 0, 0, 
			0, 166, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			170, 311, 290, 
			220, 330, 414, 
			64, 0, 173, 
			

			0, 81, 0, 
			0, 0, 0, 
			139, 0, 0, 
			

			0, 21, 78, 
			300, 0, 454, 
			181, 235, 164, 
			

			0, 0, 0, 
			0, 36, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 199, 
			0, 0, 139, 
			96, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			156, 0, 0, 
			0, 30, 0, 
			

			0, 0, 0, 
			0, 0, 15, 
			0, 537, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			506, 0, 361, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 276, 0, 
			196, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			15, 0, 18, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			55, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 291, 
			187, 0, 0, 
			0, 112, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			16, 263, 175, 
			146, 65, 0, 
			70, 108, 338, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			91, 264, 150, 
			440, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 486, 130, 
			

			688, 686, 454, 
			437, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 6, 45, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 198, 0, 
			0, 0, 0, 
			

			0, 313, 23, 
			0, 120, 33, 
			0, 0, 0, 
			

			0, 65, 0, 
			0, 0, 0, 
			0, 260, 512, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			153, 0, 266, 
			97, 0, 363, 
			0, 236, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			179, 0, 204, 
			251, 371, 475, 
			352, 705, 218, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			62, 0, 0, 
			249, 0, 0, 
			

			7, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			90, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			39, 0, 57, 
			246, 275, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			260, 0, 0, 
			63, 0, 130, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			107, 0, 0, 
			0, 0, 30, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			7, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			167, 0, 58, 
			0, 34, 0, 
			0, 0, 0, 
			

			250, 0, 187, 
			90, 0, 151, 
			110, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 353, 
			

			0, 70, 0, 
			0, 285, 0, 
			0, 0, 0, 
			

			184, 0, 171, 
			65, 0, 151, 
			0, 6, 179, 
			

			42, 0, 210, 
			0, 334, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			300, 0, 283, 
			140, 30, 181, 
			387, 131, 396, 
			

			0, 61, 198, 
			126, 164, 0, 
			6, 106, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			261, 44, 30, 
			0, 0, 0, 
			

			0, 0, 35, 
			5, 0, 0, 
			0, 556, 109, 
			

			67, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 55, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 12, 222, 
			

			0, 226, 0, 
			0, 0, 0, 
			363, 0, 0, 
			

			265, 65, 16, 
			288, 166, 31, 
			0, 0, 0, 
			

			62, 317, 0, 
			279, 0, 329, 
			0, 0, 449, 
			

			116, 261, 0, 
			89, 0, 46, 
			0, 0, 0, 
			

			344, 649, 333, 
			366, 0, 129, 
			100, 573, 505, 
			

			0, 73, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 38, 
			146, 2, 131, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 53, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			11, 0, 0, 
			86, 290, 133, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			78, 275, 0, 
			0, 0, 102, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 299, 502, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 126, 
			167, 124, 221, 
			0, 69, 0, 
			

			0, 0, 148, 
			503, 0, 151, 
			108, 0, 239, 
			

			0, 0, 0, 
			0, 0, 64, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			
