library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 58, 0, 119, 14, 
    98, 86, 0, 114, 0, 110, 0, 
    76, 34, 0, 71, 43, 68, 0, 
    39, 158, 192, 0, 0, 0, 0, 
    0, 6, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 13, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 
    0, 0, 57, 0, 38, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 
    114, 0, 40, 27, 0, 0, 0, 
    0, 195, 0, 0, 0, 2, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 29, 47, 50, 51, 
    0, 0, 0, 32, 57, 36, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 63, 0, 0, 
    0, 0, 0, 0, 146, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 
    0, 128, 126, 0, 0, 0, 0, 
    0, 111, 0, 0, 0, 80, 44, 
    232, 0, 0, 11, 84, 89, 124, 
    
    -- channel=5
    0, 0, 4, 49, 0, 24, 0, 
    0, 0, 0, 56, 59, 84, 40, 
    111, 132, 0, 62, 50, 56, 0, 
    0, 0, 146, 57, 171, 92, 57, 
    14, 71, 15, 0, 42, 0, 58, 
    0, 148, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 36, 0, 0, 0, 0, 0, 
    0, 0, 0, 61, 0, 0, 236, 
    0, 277, 0, 0, 0, 216, 0, 
    0, 131, 0, 0, 0, 268, 0, 
    0, 0, 90, 0, 0, 70, 0, 
    0, 0, 104, 0, 37, 0, 0, 
    186, 0, 0, 2, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 70, 198, 0, 
    179, 0, 209, 29, 0, 70, 43, 
    0, 0, 0, 0, 0, 0, 0, 
    7, 23, 0, 0, 0, 0, 0, 
    0, 43, 274, 0, 3, 80, 0, 
    0, 0, 0, 151, 26, 0, 42, 
    25, 0, 0, 0, 32, 12, 42, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    45, 62, 0, 0, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 0, 0, 44, 
    2, 0, 0, 0, 0, 0, 0, 
    75, 0, 0, 68, 0, 0, 0, 
    0, 90, 0, 29, 32, 2, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 82, 0, 111, 0, 
    0, 0, 0, 101, 0, 50, 56, 
    0, 0, 0, 78, 0, 0, 53, 
    77, 0, 33, 0, 4, 0, 0, 
    0, 0, 0, 0, 21, 45, 11, 
    0, 0, 0, 21, 39, 18, 0, 
    
    -- channel=11
    80, 65, 51, 44, 45, 31, 47, 
    41, 89, 62, 8, 53, 2, 50, 
    0, 98, 86, 12, 35, 31, 25, 
    0, 52, 26, 0, 32, 48, 68, 
    0, 14, 13, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    0, 0, 0, 106, 18, 0, 71, 
    0, 0, 0, 0, 8, 0, 21, 
    13, 59, 0, 0, 0, 5, 0, 
    0, 0, 99, 68, 13, 3, 0, 
    0, 0, 0, 0, 70, 13, 36, 
    125, 20, 204, 121, 0, 0, 0, 
    13, 167, 0, 0, 0, 8, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    73, 33, 77, 52, 0, 0, 42, 
    0, 0, 0, 0, 31, 0, 3, 
    0, 55, 104, 0, 51, 1, 0, 
    0, 8, 113, 33, 57, 56, 27, 
    0, 0, 0, 0, 0, 2, 21, 
    122, 0, 90, 13, 0, 0, 0, 
    0, 113, 15, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 40, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 88, 145, 265, 281, 
    158, 60, 233, 238, 271, 304, 316, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 35, 0, 0, 
    0, 40, 0, 0, 33, 0, 0, 
    0, 0, 87, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 88, 
    0, 35, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 46, 33, 77, 2, 
    6, 0, 0, 18, 15, 0, 65, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 54, 4, 0, 60, 21, 0, 
    0, 0, 53, 0, 56, 34, 0, 
    39, 0, 0, 31, 0, 0, 0, 
    0, 124, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 
    8, 0, 0, 0, 59, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 
    0, 175, 57, 0, 0, 15, 0, 
    124, 103, 149, 98, 136, 118, 145, 
    186, 145, 123, 68, 59, 95, 70, 
    
    -- channel=24
    7, 31, 11, 63, 12, 55, 28, 
    32, 0, 13, 60, 0, 86, 54, 
    0, 0, 0, 30, 0, 5, 41, 
    0, 0, 0, 40, 0, 62, 41, 
    16, 0, 36, 0, 0, 55, 65, 
    0, 0, 0, 0, 66, 30, 36, 
    14, 0, 88, 80, 82, 57, 60, 
    
    -- channel=25
    109, 79, 96, 107, 39, 46, 89, 
    111, 117, 0, 25, 54, 0, 50, 
    0, 63, 0, 0, 22, 0, 5, 
    0, 35, 13, 0, 0, 5, 53, 
    0, 17, 0, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    193, 199, 182, 234, 140, 121, 128, 
    92, 229, 209, 73, 5, 45, 10, 
    0, 131, 103, 62, 0, 41, 0, 
    0, 43, 56, 29, 24, 10, 0, 
    21, 1, 71, 0, 64, 57, 76, 
    0, 0, 36, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    20, 7, 55, 0, 0, 0, 0, 
    0, 0, 0, 44, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 123, 0, 0, 111, 
    0, 0, 0, 0, 3, 63, 28, 
    0, 0, 32, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    6, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 
    178, 0, 56, 0, 0, 0, 15, 
    109, 0, 14, 0, 0, 0, 77, 
    173, 0, 0, 0, 0, 0, 63, 
    130, 174, 0, 0, 0, 19, 0, 
    0, 175, 0, 4, 0, 0, 12, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 55, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 94, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 39, 139, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    140, 16, 0, 0, 0, 0, 0, 
    48, 0, 234, 0, 141, 0, 39, 
    28, 0, 0, 405, 0, 0, 181, 
    0, 487, 0, 0, 0, 46, 0, 
    0, 165, 42, 0, 31, 0, 117, 
    
    -- channel=35
    0, 0, 0, 27, 140, 132, 3, 
    109, 0, 184, 95, 0, 0, 0, 
    9, 0, 0, 0, 73, 0, 8, 
    0, 55, 0, 0, 0, 0, 0, 
    0, 0, 95, 142, 11, 33, 146, 
    0, 171, 54, 0, 130, 224, 117, 
    0, 0, 0, 0, 37, 0, 22, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    40, 21, 11, 21, 13, 47, 52, 
    16, 57, 7, 45, 51, 18, 2, 
    4, 0, 84, 45, 11, 30, 25, 
    0, 49, 47, 16, 12, 15, 65, 
    2, 4, 0, 0, 23, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    37, 63, 53, 102, 0, 10, 0, 
    0, 44, 53, 44, 0, 0, 0, 
    0, 112, 107, 68, 0, 51, 0, 
    89, 66, 52, 64, 0, 3, 0, 
    70, 0, 0, 0, 65, 0, 0, 
    0, 0, 66, 0, 0, 0, 0, 
    0, 81, 0, 0, 0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 48, 0, 
    0, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 18, 0, 36, 0, 
    0, 0, 245, 0, 0, 144, 0, 
    7, 0, 163, 190, 213, 138, 189, 
    59, 0, 218, 159, 190, 213, 233, 
    
    -- channel=40
    0, 50, 74, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 
    62, 0, 266, 156, 123, 137, 108, 
    206, 10, 151, 82, 96, 117, 72, 
    
    -- channel=43
    52, 189, 1, 0, 0, 0, 0, 
    0, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 69, 
    0, 0, 0, 0, 0, 0, 78, 
    0, 0, 0, 0, 0, 77, 0, 
    0, 0, 0, 0, 12, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 118, 16, 0, 0, 0, 0, 
    0, 68, 21, 0, 0, 29, 0, 
    0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 44, 
    0, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    59, 35, 0, 0, 0, 0, 64, 
    0, 15, 0, 0, 82, 0, 0, 
    0, 113, 0, 0, 7, 0, 0, 
    0, 19, 128, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 42, 
    106, 0, 0, 0, 0, 84, 30, 
    165, 0, 0, 46, 90, 124, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    98, 81, 67, 51, 31, 39, 84, 
    70, 114, 75, 38, 79, 52, 44, 
    121, 79, 102, 79, 65, 49, 31, 
    84, 103, 81, 45, 72, 26, 83, 
    49, 110, 88, 0, 8, 0, 27, 
    9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 40, 0, 19, 
    97, 0, 34, 0, 63, 0, 0, 
    24, 0, 26, 0, 130, 0, 72, 
    152, 201, 0, 0, 0, 0, 17, 
    0, 97, 0, 0, 0, 63, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    54, 0, 0, 1, 0, 21, 133, 
    165, 90, 0, 0, 0, 0, 165, 
    0, 97, 0, 0, 0, 0, 0, 
    0, 147, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 47, 120, 62, 26, 
    55, 141, 0, 0, 112, 38, 6, 
    0, 0, 73, 43, 104, 0, 81, 
    0, 66, 142, 0, 101, 0, 0, 
    0, 100, 64, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    67, 45, 89, 67, 42, 0, 20, 
    8, 38, 24, 0, 0, 0, 32, 
    0, 147, 80, 0, 0, 0, 0, 
    0, 2, 18, 0, 51, 24, 7, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    1, 0, 0, 190, 115, 3, 81, 
    0, 71, 0, 0, 36, 0, 0, 
    5, 26, 155, 0, 0, 59, 0, 
    0, 0, 0, 95, 0, 0, 0, 
    0, 0, 0, 0, 110, 15, 0, 
    93, 0, 412, 126, 48, 52, 19, 
    0, 122, 0, 0, 0, 45, 0, 
    
    -- channel=59
    100, 94, 0, 206, 258, 64, 87, 
    127, 245, 171, 0, 0, 47, 30, 
    0, 0, 82, 5, 0, 191, 38, 
    45, 137, 0, 246, 0, 53, 0, 
    0, 174, 161, 0, 65, 217, 0, 
    0, 0, 245, 86, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 0, 42, 323, 0, 122, 20, 
    3, 64, 81, 207, 57, 186, 11, 
    127, 125, 0, 261, 48, 306, 0, 
    165, 89, 242, 147, 109, 145, 0, 
    0, 109, 118, 20, 402, 0, 0, 
    0, 58, 335, 48, 0, 0, 0, 
    0, 299, 0, 0, 0, 14, 0, 
    
    -- channel=61
    0, 0, 0, 33, 0, 148, 0, 
    151, 0, 52, 182, 0, 191, 184, 
    178, 0, 0, 344, 0, 286, 83, 
    202, 172, 0, 112, 0, 209, 0, 
    63, 106, 202, 89, 60, 30, 0, 
    0, 0, 228, 0, 3, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 42, 
    44, 190, 29, 0, 0, 79, 0, 
    85, 140, 0, 0, 3, 105, 0, 
    0, 0, 104, 58, 40, 32, 0, 
    0, 0, 0, 0, 41, 4, 0, 
    0, 182, 21, 0, 0, 4, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 0, 
    29, 0, 0, 104, 0, 78, 0, 
    52, 0, 0, 63, 0, 113, 0, 
    81, 183, 9, 0, 0, 0, 0, 
    0, 50, 222, 0, 77, 0, 38, 
    0, 0, 149, 55, 35, 66, 75, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 0, 0, 
    32, 0, 0, 0, 97, 0, 10, 
    32, 0, 0, 0, 0, 0, 0, 
    122, 126, 0, 59, 0, 1, 0, 
    231, 134, 0, 106, 112, 134, 151, 
    170, 142, 144, 134, 142, 166, 198, 
    
    -- channel=65
    0, 2, 0, 0, 0, 46, 0, 
    0, 0, 0, 37, 0, 0, 53, 
    0, 0, 13, 134, 0, 106, 149, 
    234, 171, 0, 0, 0, 79, 0, 
    21, 0, 0, 163, 1, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    62, 69, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 
    
    -- channel=67
    240, 315, 71, 167, 0, 0, 136, 
    0, 47, 0, 0, 0, 70, 0, 
    0, 0, 0, 20, 0, 39, 0, 
    0, 0, 0, 66, 0, 14, 0, 
    105, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 55, 
    0, 0, 0, 138, 91, 94, 0, 
    
    -- channel=68
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 36, 0, 
    0, 0, 0, 0, 0, 11, 0, 
    173, 0, 141, 93, 87, 118, 104, 
    71, 110, 155, 133, 128, 173, 137, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 24, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 
    0, 0, 58, 64, 20, 0, 68, 
    0, 94, 80, 0, 69, 81, 44, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    327, 330, 201, 343, 142, 124, 240, 
    184, 252, 108, 0, 0, 0, 32, 
    0, 139, 0, 0, 0, 0, 0, 
    0, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 125, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=72
    0, 0, 12, 0, 30, 119, 0, 
    156, 0, 142, 51, 0, 0, 93, 
    0, 77, 0, 30, 55, 0, 0, 
    14, 35, 0, 0, 83, 47, 0, 
    0, 0, 79, 32, 0, 102, 9, 
    0, 29, 0, 68, 0, 0, 0, 
    40, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 70, 0, 
    0, 0, 0, 72, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 172, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    149, 0, 123, 212, 0, 0, 91, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 169, 
    74, 0, 0, 0, 0, 0, 0, 
    8, 83, 53, 0, 0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 
    150, 26, 0, 0, 60, 0, 0, 
    0, 0, 0, 0, 212, 0, 0, 
    0, 123, 0, 0, 0, 0, 0, 
    0, 368, 82, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=78
    10, 0, 0, 0, 26, 43, 8, 
    53, 41, 0, 32, 82, 0, 78, 
    0, 54, 37, 0, 105, 20, 41, 
    0, 89, 22, 0, 12, 27, 60, 
    0, 68, 27, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 145, 134, 
    124, 0, 0, 142, 162, 166, 105, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 35, 0, 39, 
    67, 0, 2, 0, 38, 0, 0, 
    0, 0, 0, 0, 82, 0, 0, 
    92, 89, 0, 0, 0, 0, 111, 
    137, 242, 138, 84, 95, 130, 129, 
    240, 19, 83, 96, 89, 132, 102, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 0, 203, 0, 0, 
    200, 41, 103, 0, 0, 0, 0, 
    0, 8, 0, 0, 227, 0, 6, 
    0, 61, 0, 0, 0, 0, 0, 
    0, 99, 24, 0, 0, 247, 0, 
    0, 129, 0, 0, 188, 20, 0, 
    132, 0, 33, 0, 43, 0, 117, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 
    46, 0, 0, 0, 0, 10, 24, 
    196, 0, 0, 0, 0, 19, 0, 
    68, 0, 0, 69, 3, 19, 139, 
    90, 9, 0, 0, 0, 0, 0, 
    164, 17, 44, 29, 0, 0, 0, 
    43, 133, 38, 31, 11, 40, 59, 
    
    -- channel=89
    59, 0, 0, 95, 132, 68, 89, 
    108, 25, 0, 0, 2, 0, 44, 
    0, 0, 18, 0, 0, 0, 0, 
    0, 91, 0, 44, 0, 11, 0, 
    0, 0, 0, 0, 0, 98, 0, 
    58, 0, 120, 78, 0, 0, 0, 
    0, 38, 5, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    6, 0, 50, 209, 141, 116, 53, 
    0, 0, 41, 41, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 2, 0, 0, 0, 
    0, 0, 0, 0, 49, 21, 0, 
    0, 0, 174, 157, 11, 0, 0, 
    0, 85, 59, 0, 0, 0, 0, 
    
    -- channel=92
    0, 0, 0, 87, 36, 31, 41, 
    0, 0, 0, 0, 0, 0, 29, 
    0, 48, 0, 0, 0, 15, 0, 
    0, 0, 30, 61, 19, 0, 0, 
    0, 0, 0, 0, 32, 34, 0, 
    20, 0, 138, 134, 0, 0, 0, 
    0, 77, 0, 0, 0, 0, 0, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 61, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 
    0, 232, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 21, 0, 
    0, 0, 0, 109, 0, 33, 277, 
    0, 301, 0, 76, 0, 178, 0, 
    0, 0, 0, 0, 89, 237, 0, 
    0, 0, 216, 0, 0, 23, 0, 
    0, 0, 203, 0, 0, 0, 0, 
    111, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=96
    77, 0, 30, 38, 101, 0, 91, 
    578, 198, 25, 7, 393, 20, 0, 
    394, 89, 0, 19, 850, 0, 0, 
    163, 102, 68, 121, 314, 0, 0, 
    88, 826, 171, 0, 3, 0, 0, 
    0, 430, 252, 0, 16, 0, 0, 
    42, 0, 177, 0, 0, 2, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 51, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 39, 
    4, 0, 0, 58, 51, 79, 0, 
    
    -- channel=98
    0, 0, 117, 0, 0, 2, 0, 
    40, 31, 80, 95, 0, 0, 0, 
    0, 0, 0, 139, 61, 0, 30, 
    0, 0, 0, 0, 0, 39, 0, 
    0, 94, 91, 219, 0, 0, 64, 
    0, 58, 0, 0, 1, 15, 10, 
    0, 0, 2, 25, 26, 0, 73, 
    
    -- channel=99
    116, 61, 148, 99, 131, 66, 102, 
    121, 212, 0, 68, 99, 0, 34, 
    0, 0, 0, 64, 184, 24, 120, 
    0, 161, 0, 0, 0, 10, 8, 
    0, 216, 0, 0, 42, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=100
    0, 0, 0, 137, 0, 39, 0, 
    0, 0, 0, 50, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 
    0, 0, 10, 3, 0, 0, 0, 
    0, 0, 0, 0, 126, 0, 75, 
    0, 0, 176, 87, 48, 95, 131, 
    28, 261, 61, 86, 40, 94, 0, 
    
    -- channel=101
    269, 270, 251, 249, 214, 63, 238, 
    199, 295, 155, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    0, 0, 5, 0, 108, 0, 27, 
    141, 83, 14, 0, 260, 0, 0, 
    88, 0, 0, 0, 420, 0, 0, 
    0, 0, 206, 0, 233, 0, 4, 
    47, 283, 0, 0, 0, 0, 0, 
    2, 261, 0, 0, 0, 0, 0, 
    0, 0, 79, 0, 0, 0, 1, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 
    56, 0, 0, 0, 0, 0, 95, 
    0, 304, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 35, 0, 0, 
    0, 0, 76, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    55, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 42, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 66, 0, 0, 0, 0, 0, 
    0, 3, 26, 0, 0, 116, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    168, 131, 141, 175, 62, 40, 68, 
    0, 151, 51, 19, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    166, 77, 77, 83, 19, 0, 142, 
    22, 132, 0, 0, 116, 0, 0, 
    0, 0, 0, 0, 135, 0, 0, 
    0, 45, 173, 0, 50, 0, 23, 
    62, 81, 0, 0, 0, 0, 42, 
    150, 0, 0, 0, 0, 0, 0, 
    0, 70, 33, 0, 0, 0, 0, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    45, 0, 0, 150, 58, 174, 189, 
    297, 57, 0, 0, 5, 0, 116, 
    144, 0, 0, 0, 19, 0, 45, 
    25, 68, 0, 0, 0, 8, 0, 
    0, 87, 0, 14, 107, 129, 299, 
    157, 24, 70, 160, 189, 105, 148, 
    152, 207, 194, 115, 97, 108, 159, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    1, 83, 65, 65, 0, 42, 4, 
    0, 49, 130, 64, 0, 149, 0, 
    81, 0, 35, 252, 0, 95, 50, 
    33, 0, 0, 75, 0, 29, 0, 
    84, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    146, 0, 205, 103, 0, 0, 82, 
    149, 0, 0, 13, 0, 24, 0, 
    155, 95, 0, 78, 0, 0, 6, 
    57, 45, 203, 71, 139, 41, 59, 
    0, 230, 140, 39, 11, 18, 15, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 
    197, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 325, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 0, 30, 30, 
    0, 212, 0, 0, 85, 0, 0, 
    15, 0, 39, 0, 0, 0, 72, 
    
    -- channel=117
    0, 6, 0, 0, 0, 89, 0, 
    251, 0, 176, 78, 0, 46, 81, 
    0, 66, 0, 67, 143, 0, 0, 
    42, 2, 0, 0, 46, 0, 0, 
    0, 119, 192, 0, 0, 0, 0, 
    0, 64, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    0, 4, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 7, 0, 42, 
    0, 0, 0, 0, 0, 12, 62, 
    35, 82, 0, 0, 0, 0, 26, 
    0, 0, 56, 0, 0, 35, 0, 
    0, 0, 0, 0, 33, 76, 67, 
    75, 0, 0, 56, 79, 54, 3, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 132, 80, 
    0, 0, 6, 26, 88, 88, 77, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 55, 32, 12, 24, 
    41, 0, 0, 3, 0, 59, 0, 
    0, 153, 106, 7, 0, 96, 0, 
    0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 0, 61, 
    0, 0, 0, 0, 0, 193, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 
    
    -- channel=125
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 
    76, 0, 0, 65, 0, 0, 0, 
    0, 0, 0, 0, 0, 162, 0, 
    0, 24, 0, 60, 0, 17, 0, 
    0, 189, 0, 0, 0, 0, 0, 
    0, 0, 229, 0, 42, 0, 0, 
    0, 0, 175, 0, 0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 37, 0, 0, 
    71, 0, 88, 0, 79, 0, 0, 
    0, 5, 70, 22, 75, 0, 0, 
    0, 14, 0, 0, 25, 0, 0, 
    128, 23, 148, 13, 0, 0, 0, 
    71, 205, 59, 0, 0, 18, 0, 
    
    
    others => 0);
end ifmap_package;
