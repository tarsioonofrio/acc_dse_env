library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 2**16) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 38, 42, 42, 47, 47, 36, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 33, 60, 58, 52, 40, 42, 51, 60, 61, 51, 30, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 69, 91, 86, 62, 27, 0, 0, 10, 29, 40, 54, 61, 43, 6, 
    32, 37, 12, 0, 0, 0, 0, 0, 12, 14, 4, 8, 35, 68, 85, 88, 82, 63, 26, 1, 1, 17, 19, 25, 48, 77, 75, 33, 
    66, 78, 38, 0, 0, 0, 0, 0, 17, 50, 32, 23, 11, 21, 38, 52, 72, 70, 40, 8, 6, 32, 40, 45, 52, 81, 94, 62, 
    35, 62, 24, 0, 0, 0, 0, 0, 0, 9, 3, 0, 0, 0, 30, 53, 82, 94, 68, 21, 6, 30, 60, 63, 57, 66, 91, 89, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 40, 66, 106, 132, 96, 38, 1, 17, 47, 57, 53, 46, 71, 97, 
    0, 0, 0, 0, 0, 16, 6, 0, 0, 0, 0, 0, 0, 5, 43, 63, 107, 134, 93, 19, 0, 0, 19, 44, 35, 30, 51, 86, 
    15, 0, 0, 0, 0, 39, 74, 31, 0, 0, 0, 0, 0, 0, 26, 31, 86, 99, 54, 0, 0, 0, 20, 45, 39, 31, 35, 67, 
    44, 15, 0, 0, 0, 52, 145, 130, 48, 7, 0, 0, 0, 0, 2, 4, 66, 79, 49, 0, 0, 11, 46, 62, 53, 44, 30, 31, 
    59, 25, 0, 0, 0, 20, 126, 138, 107, 53, 19, 0, 0, 0, 0, 0, 61, 85, 60, 0, 0, 29, 56, 73, 68, 60, 31, 3, 
    47, 28, 0, 0, 0, 0, 51, 94, 90, 48, 9, 0, 0, 0, 0, 0, 67, 94, 69, 2, 12, 27, 55, 70, 70, 51, 18, 0, 
    33, 26, 0, 3, 9, 0, 16, 62, 80, 40, 2, 0, 0, 12, 10, 16, 70, 91, 63, 1, 0, 8, 38, 57, 57, 34, 7, 0, 
    22, 18, 0, 0, 5, 0, 0, 39, 79, 56, 21, 17, 40, 67, 52, 38, 65, 80, 68, 35, 26, 23, 51, 75, 71, 45, 13, 0, 
    14, 14, 0, 0, 2, 8, 0, 34, 87, 117, 97, 75, 76, 77, 63, 43, 46, 49, 68, 66, 49, 38, 71, 109, 103, 71, 26, 0, 
    13, 17, 0, 0, 18, 23, 0, 24, 83, 147, 150, 101, 76, 52, 28, 31, 39, 65, 73, 83, 77, 84, 107, 114, 93, 43, 3, 0, 
    17, 20, 5, 0, 25, 35, 24, 0, 33, 82, 81, 64, 25, 9, 0, 11, 26, 40, 54, 86, 113, 128, 131, 97, 52, 7, 0, 0, 
    23, 16, 15, 0, 34, 65, 47, 0, 0, 32, 56, 67, 21, 0, 0, 0, 20, 45, 63, 102, 119, 123, 110, 73, 41, 12, 0, 0, 
    29, 9, 14, 0, 35, 73, 48, 0, 0, 16, 46, 46, 25, 6, 0, 9, 56, 106, 145, 154, 145, 134, 108, 100, 79, 64, 48, 48, 
    53, 17, 16, 3, 48, 69, 26, 0, 0, 0, 49, 82, 92, 88, 65, 60, 91, 130, 158, 150, 138, 126, 117, 129, 133, 139, 131, 132, 
    115, 64, 30, 2, 45, 48, 23, 0, 0, 52, 131, 175, 201, 207, 194, 164, 142, 137, 134, 134, 140, 147, 156, 158, 164, 167, 169, 170, 
    184, 142, 66, 23, 44, 50, 33, 31, 100, 192, 246, 272, 283, 278, 258, 223, 192, 172, 169, 167, 172, 179, 185, 183, 182, 182, 184, 183, 
    225, 210, 138, 101, 65, 65, 56, 110, 199, 231, 221, 206, 202, 201, 195, 187, 185, 184, 188, 188, 190, 192, 191, 188, 187, 191, 194, 194, 
    213, 221, 193, 171, 111, 85, 65, 134, 196, 197, 173, 165, 167, 170, 175, 178, 182, 187, 192, 195, 194, 192, 189, 190, 196, 207, 209, 201, 
    201, 203, 200, 211, 175, 120, 81, 136, 190, 183, 175, 171, 171, 173, 177, 179, 182, 188, 193, 195, 198, 200, 199, 204, 214, 223, 217, 198, 
    198, 195, 196, 224, 237, 184, 127, 152, 190, 183, 180, 173, 168, 169, 175, 181, 186, 191, 196, 203, 205, 207, 212, 215, 221, 218, 206, 199, 
    201, 196, 201, 229, 263, 246, 196, 191, 196, 194, 191, 183, 176, 173, 178, 182, 185, 190, 194, 199, 203, 208, 214, 218, 214, 209, 208, 210, 
    204, 202, 202, 223, 257, 260, 236, 220, 204, 200, 197, 194, 192, 186, 185, 185, 187, 187, 185, 187, 194, 201, 207, 210, 208, 202, 195, 194, 
    
    -- channel=1
    195, 192, 198, 205, 208, 205, 204, 201, 203, 209, 213, 216, 207, 194, 174, 147, 134, 122, 117, 111, 111, 117, 125, 140, 154, 164, 165, 160, 
    197, 192, 197, 205, 207, 207, 206, 202, 206, 210, 213, 196, 173, 147, 118, 99, 95, 96, 94, 92, 92, 87, 94, 103, 125, 147, 159, 161, 
    184, 183, 189, 200, 206, 207, 209, 212, 210, 201, 182, 165, 138, 103, 70, 59, 73, 98, 105, 98, 88, 88, 92, 96, 103, 121, 144, 155, 
    154, 172, 190, 199, 203, 205, 207, 212, 188, 149, 131, 123, 88, 50, 41, 51, 81, 107, 109, 90, 75, 73, 73, 76, 74, 96, 126, 148, 
    104, 146, 182, 207, 210, 211, 210, 196, 160, 115, 102, 91, 79, 58, 59, 76, 99, 112, 108, 86, 77, 71, 56, 34, 50, 77, 112, 138, 
    89, 148, 192, 210, 215, 211, 210, 184, 166, 143, 138, 122, 99, 73, 66, 76, 90, 106, 108, 96, 84, 71, 48, 28, 33, 66, 99, 127, 
    107, 182, 222, 220, 207, 202, 199, 187, 169, 160, 159, 129, 87, 69, 57, 58, 78, 102, 109, 103, 95, 75, 51, 38, 31, 52, 79, 108, 
    121, 190, 219, 221, 199, 195, 199, 189, 169, 163, 153, 118, 87, 66, 51, 35, 61, 105, 129, 121, 101, 76, 67, 61, 50, 41, 65, 86, 
    133, 188, 205, 209, 192, 172, 174, 147, 132, 139, 146, 124, 97, 81, 57, 47, 72, 132, 154, 135, 87, 61, 63, 75, 60, 38, 43, 76, 
    136, 178, 195, 194, 171, 136, 116, 94, 104, 140, 163, 148, 120, 97, 70, 66, 97, 155, 157, 112, 55, 40, 56, 69, 61, 47, 43, 69, 
    139, 159, 172, 183, 159, 127, 96, 85, 98, 143, 175, 160, 125, 102, 84, 81, 114, 165, 133, 85, 39, 35, 58, 69, 71, 64, 63, 75, 
    137, 135, 130, 158, 163, 138, 120, 121, 142, 184, 196, 154, 117, 103, 81, 78, 118, 159, 112, 73, 36, 34, 48, 66, 79, 84, 86, 95, 
    133, 106, 108, 148, 165, 140, 124, 135, 165, 192, 164, 103, 71, 83, 72, 72, 116, 147, 112, 78, 56, 52, 55, 76, 95, 101, 97, 118, 
    140, 98, 95, 137, 166, 156, 136, 156, 166, 146, 92, 42, 43, 54, 59, 81, 129, 129, 93, 65, 45, 33, 39, 65, 89, 97, 114, 146, 
    146, 108, 84, 105, 150, 161, 156, 150, 138, 81, 35, 33, 61, 69, 76, 110, 141, 124, 90, 64, 32, 10, 17, 51, 84, 107, 135, 159, 
    143, 114, 73, 77, 118, 143, 151, 127, 90, 37, 22, 47, 77, 90, 100, 127, 144, 113, 75, 42, 5, 0, 15, 54, 89, 128, 163, 187, 
    139, 121, 72, 63, 100, 129, 132, 118, 72, 56, 77, 113, 124, 114, 112, 120, 125, 95, 64, 4, 0, 0, 10, 68, 117, 157, 188, 197, 
    140, 132, 84, 54, 74, 117, 116, 98, 101, 98, 125, 148, 155, 116, 98, 107, 105, 64, 30, 0, 0, 0, 33, 104, 153, 177, 180, 171, 
    145, 140, 93, 59, 78, 129, 132, 98, 77, 96, 129, 147, 149, 94, 49, 57, 39, 0, 0, 0, 0, 0, 32, 90, 133, 145, 130, 115, 
    135, 130, 91, 71, 115, 174, 164, 122, 67, 60, 82, 87, 65, 14, 0, 0, 0, 0, 0, 0, 0, 0, 3, 35, 61, 54, 39, 28, 
    97, 107, 90, 94, 157, 221, 177, 72, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 74, 94, 131, 198, 226, 129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 74, 140, 215, 178, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 132, 203, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 117, 139, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 68, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    420, 425, 421, 422, 425, 428, 424, 415, 396, 403, 417, 433, 439, 434, 416, 384, 334, 292, 260, 248, 246, 262, 284, 305, 332, 356, 367, 362, 
    422, 432, 430, 428, 433, 435, 428, 406, 385, 400, 403, 409, 405, 393, 366, 312, 250, 200, 171, 161, 163, 177, 196, 231, 272, 312, 342, 356, 
    401, 420, 430, 434, 440, 440, 433, 405, 387, 394, 385, 373, 344, 313, 271, 208, 154, 127, 118, 107, 106, 118, 139, 166, 203, 253, 300, 335, 
    334, 367, 404, 431, 442, 442, 436, 410, 392, 372, 334, 298, 256, 207, 162, 116, 99, 100, 99, 89, 83, 92, 104, 122, 152, 187, 247, 304, 
    230, 276, 358, 423, 444, 442, 430, 410, 376, 310, 252, 223, 184, 133, 103, 93, 88, 97, 104, 100, 88, 89, 91, 89, 100, 134, 197, 270, 
    149, 214, 320, 409, 435, 426, 408, 392, 341, 276, 229, 200, 158, 115, 93, 85, 83, 95, 122, 120, 109, 100, 88, 70, 68, 102, 157, 231, 
    121, 196, 305, 390, 409, 377, 361, 350, 298, 231, 204, 182, 136, 99, 79, 77, 79, 87, 118, 127, 126, 109, 82, 66, 63, 84, 127, 186, 
    100, 185, 297, 374, 375, 315, 302, 290, 256, 210, 187, 168, 126, 93, 71, 72, 62, 76, 114, 131, 131, 107, 87, 80, 75, 79, 105, 144, 
    74, 168, 288, 365, 354, 276, 236, 241, 227, 200, 177, 162, 132, 103, 86, 76, 53, 80, 121, 140, 133, 105, 92, 84, 81, 77, 86, 117, 
    44, 156, 273, 359, 359, 276, 189, 185, 168, 170, 170, 172, 156, 122, 100, 85, 54, 83, 126, 143, 125, 90, 80, 79, 77, 72, 76, 105, 
    28, 141, 243, 340, 369, 305, 188, 159, 138, 149, 164, 182, 164, 136, 117, 88, 58, 81, 123, 129, 99, 70, 65, 70, 68, 72, 80, 109, 
    31, 121, 196, 281, 347, 317, 228, 175, 140, 144, 162, 177, 157, 144, 130, 86, 63, 85, 113, 108, 83, 66, 59, 64, 63, 73, 93, 131, 
    46, 92, 140, 202, 294, 295, 244, 170, 134, 151, 163, 152, 132, 131, 130, 89, 75, 95, 113, 106, 87, 72, 60, 62, 75, 98, 130, 168, 
    51, 70, 95, 138, 218, 250, 236, 162, 144, 153, 158, 141, 113, 116, 122, 101, 105, 131, 129, 114, 101, 77, 60, 67, 92, 129, 168, 213, 
    44, 59, 65, 86, 136, 199, 212, 167, 157, 152, 151, 123, 106, 106, 100, 108, 152, 164, 145, 133, 111, 81, 62, 69, 99, 148, 196, 253, 
    33, 50, 44, 49, 71, 142, 173, 162, 150, 116, 106, 91, 100, 101, 89, 111, 171, 179, 145, 125, 108, 88, 68, 79, 117, 179, 243, 303, 
    31, 42, 37, 30, 34, 85, 124, 148, 143, 101, 109, 107, 123, 114, 89, 101, 165, 170, 147, 119, 86, 46, 46, 87, 150, 232, 301, 344, 
    42, 46, 48, 28, 24, 50, 92, 119, 116, 105, 112, 116, 132, 117, 91, 93, 127, 147, 135, 99, 47, 8, 32, 85, 169, 247, 303, 324, 
    53, 58, 61, 30, 19, 45, 81, 106, 87, 87, 73, 76, 96, 100, 78, 74, 83, 73, 43, 1, 0, 0, 0, 35, 108, 174, 213, 215, 
    50, 63, 64, 37, 24, 68, 98, 98, 73, 51, 46, 64, 80, 78, 54, 38, 32, 3, 0, 0, 0, 0, 0, 0, 0, 31, 44, 40, 
    21, 51, 61, 43, 37, 62, 105, 100, 50, 24, 20, 24, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 49, 39, 57, 76, 100, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 20, 55, 91, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 35, 78, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 23, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    25, 26, 29, 28, 29, 29, 28, 22, 21, 32, 44, 44, 32, 28, 29, 20, 0, 0, 0, 2, 3, 2, 0, 0, 0, 3, 11, 19, 
    21, 21, 25, 28, 30, 29, 28, 15, 7, 23, 43, 37, 23, 18, 5, 0, 0, 0, 0, 3, 9, 8, 0, 0, 0, 0, 0, 11, 
    8, 1, 5, 21, 29, 30, 31, 29, 16, 5, 26, 28, 16, 0, 0, 0, 0, 0, 3, 18, 20, 10, 8, 9, 4, 0, 0, 0, 
    0, 0, 0, 17, 28, 30, 33, 45, 32, 5, 3, 11, 9, 0, 0, 0, 0, 0, 10, 29, 23, 7, 3, 10, 7, 0, 0, 0, 
    6, 0, 0, 25, 29, 28, 32, 45, 26, 0, 0, 11, 15, 7, 0, 0, 0, 0, 5, 31, 31, 13, 3, 3, 0, 0, 0, 0, 
    9, 0, 12, 32, 29, 20, 27, 43, 37, 23, 15, 27, 35, 15, 0, 0, 0, 0, 0, 23, 33, 17, 4, 0, 2, 3, 0, 0, 
    15, 0, 29, 43, 22, 0, 15, 39, 59, 43, 27, 41, 47, 27, 12, 5, 0, 0, 0, 21, 40, 28, 9, 0, 3, 11, 6, 0, 
    2, 0, 39, 48, 29, 0, 0, 14, 49, 47, 36, 51, 54, 37, 18, 6, 0, 0, 0, 34, 57, 38, 10, 0, 3, 11, 10, 2, 
    0, 0, 47, 49, 45, 18, 0, 0, 28, 32, 26, 53, 63, 44, 28, 8, 0, 0, 0, 52, 64, 37, 4, 0, 0, 7, 8, 4, 
    9, 15, 49, 41, 46, 38, 0, 0, 18, 10, 19, 56, 69, 57, 36, 19, 0, 0, 10, 64, 61, 34, 1, 0, 0, 0, 2, 4, 
    19, 30, 55, 31, 32, 38, 2, 0, 0, 9, 18, 56, 65, 49, 41, 26, 0, 0, 26, 58, 54, 31, 5, 0, 0, 0, 2, 1, 
    25, 43, 64, 28, 12, 34, 17, 0, 0, 13, 40, 64, 60, 36, 34, 23, 0, 0, 26, 52, 52, 32, 1, 0, 0, 0, 7, 0, 
    32, 53, 67, 37, 5, 19, 17, 0, 0, 4, 59, 66, 46, 25, 16, 14, 0, 0, 20, 49, 46, 32, 7, 0, 0, 0, 4, 0, 
    42, 65, 71, 47, 13, 18, 19, 0, 0, 4, 26, 32, 14, 4, 1, 4, 0, 0, 6, 16, 32, 34, 4, 0, 0, 0, 0, 3, 
    50, 69, 78, 56, 13, 14, 29, 34, 7, 0, 3, 3, 4, 1, 0, 6, 13, 10, 0, 6, 24, 20, 0, 0, 0, 0, 0, 14, 
    51, 68, 87, 67, 26, 4, 23, 45, 17, 0, 0, 0, 0, 13, 17, 10, 7, 13, 11, 5, 12, 1, 0, 0, 0, 0, 11, 23, 
    48, 63, 86, 73, 37, 5, 19, 46, 34, 0, 0, 0, 4, 36, 49, 31, 2, 9, 6, 3, 0, 0, 0, 0, 0, 0, 18, 24, 
    46, 58, 79, 79, 34, 1, 25, 55, 49, 25, 0, 0, 12, 51, 66, 52, 26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 
    44, 60, 73, 75, 26, 0, 35, 83, 87, 40, 15, 7, 17, 57, 66, 45, 37, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    32, 50, 65, 65, 25, 0, 52, 103, 111, 59, 15, 0, 11, 29, 35, 28, 19, 5, 0, 0, 0, 3, 3, 4, 8, 11, 11, 7, 
    14, 27, 49, 53, 16, 5, 80, 126, 97, 50, 18, 13, 15, 17, 19, 23, 24, 19, 13, 12, 15, 16, 18, 21, 22, 25, 30, 31, 
    12, 13, 29, 21, 0, 38, 119, 127, 86, 33, 5, 0, 0, 0, 0, 1, 15, 16, 15, 18, 21, 23, 25, 28, 30, 32, 35, 34, 
    10, 4, 0, 2, 4, 77, 121, 92, 38, 12, 8, 9, 9, 8, 10, 13, 16, 17, 18, 21, 25, 27, 30, 34, 34, 32, 31, 33, 
    18, 2, 0, 0, 10, 94, 110, 76, 28, 19, 24, 27, 25, 22, 20, 19, 19, 19, 21, 24, 27, 30, 34, 38, 35, 29, 31, 40, 
    32, 11, 3, 0, 8, 73, 98, 60, 21, 18, 25, 28, 26, 23, 22, 21, 20, 22, 25, 28, 30, 33, 36, 33, 30, 32, 41, 51, 
    39, 26, 19, 7, 9, 48, 72, 41, 14, 18, 24, 26, 27, 25, 22, 21, 23, 26, 29, 30, 32, 32, 30, 28, 28, 34, 48, 55, 
    42, 33, 28, 13, 7, 22, 41, 23, 13, 15, 21, 24, 23, 23, 22, 22, 24, 28, 33, 34, 30, 26, 24, 23, 29, 43, 56, 50, 
    43, 34, 30, 16, 0, 12, 12, 11, 10, 10, 16, 19, 21, 19, 13, 13, 20, 29, 37, 37, 30, 23, 17, 19, 34, 59, 68, 52, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    136, 141, 141, 147, 151, 149, 144, 139, 143, 150, 148, 142, 143, 143, 132, 109, 90, 81, 77, 70, 72, 83, 103, 122, 133, 127, 112, 97, 
    142, 144, 144, 149, 154, 152, 151, 171, 194, 213, 186, 152, 140, 129, 103, 86, 81, 94, 92, 84, 72, 57, 57, 75, 106, 125, 125, 111, 
    163, 160, 151, 147, 149, 147, 146, 175, 226, 269, 212, 140, 101, 75, 55, 52, 86, 136, 154, 152, 129, 104, 70, 60, 74, 103, 127, 124, 
    128, 160, 169, 155, 146, 141, 137, 132, 151, 171, 145, 98, 48, 21, 25, 50, 107, 168, 191, 189, 176, 149, 109, 68, 49, 70, 115, 137, 
    52, 112, 165, 164, 149, 140, 136, 113, 100, 104, 110, 94, 59, 40, 47, 79, 135, 200, 213, 188, 166, 150, 119, 69, 41, 51, 89, 132, 
    66, 115, 157, 159, 145, 141, 135, 122, 111, 122, 149, 150, 118, 93, 84, 93, 127, 191, 224, 191, 137, 113, 91, 65, 37, 31, 64, 116, 
    155, 202, 207, 173, 150, 172, 195, 201, 168, 176, 207, 192, 140, 100, 82, 72, 90, 144, 207, 201, 144, 100, 75, 65, 43, 18, 29, 78, 
    252, 286, 260, 186, 167, 229, 332, 364, 320, 266, 249, 219, 161, 106, 65, 53, 72, 135, 216, 222, 177, 129, 95, 83, 64, 30, 12, 32, 
    317, 347, 304, 196, 142, 188, 345, 439, 407, 332, 294, 253, 188, 132, 69, 61, 93, 178, 269, 264, 208, 149, 118, 111, 89, 54, 25, 23, 
    335, 379, 338, 227, 118, 95, 190, 326, 364, 344, 337, 294, 228, 165, 98, 91, 121, 231, 313, 277, 200, 135, 120, 117, 108, 86, 63, 46, 
    315, 355, 319, 245, 148, 77, 99, 210, 273, 313, 364, 352, 276, 205, 145, 133, 149, 260, 312, 257, 177, 113, 97, 99, 113, 112, 103, 88, 
    309, 312, 256, 216, 168, 98, 79, 174, 249, 321, 370, 381, 327, 253, 178, 159, 177, 269, 307, 252, 180, 116, 89, 95, 115, 132, 137, 126, 
    329, 297, 239, 198, 168, 123, 86, 164, 276, 362, 370, 334, 295, 257, 200, 162, 177, 260, 295, 245, 183, 138, 114, 120, 147, 162, 156, 141, 
    364, 319, 263, 213, 197, 162, 121, 175, 305, 396, 368, 285, 225, 198, 173, 158, 176, 238, 263, 231, 173, 119, 107, 125, 149, 155, 154, 140, 
    394, 354, 294, 236, 233, 205, 169, 143, 213, 283, 259, 221, 174, 144, 151, 159, 148, 176, 207, 217, 173, 105, 80, 94, 120, 142, 142, 136, 
    410, 383, 309, 253, 244, 253, 209, 130, 122, 140, 158, 163, 143, 132, 154, 165, 154, 124, 100, 124, 114, 65, 48, 72, 105, 137, 145, 147, 
    415, 399, 325, 260, 232, 260, 256, 185, 129, 102, 150, 186, 191, 173, 172, 190, 210, 162, 97, 61, 22, 26, 42, 73, 112, 151, 165, 159, 
    413, 400, 343, 273, 233, 256, 268, 218, 169, 130, 176, 234, 270, 243, 197, 170, 172, 156, 99, 40, 6, 21, 61, 115, 154, 179, 172, 150, 
    408, 389, 338, 286, 274, 307, 324, 273, 204, 179, 211, 281, 352, 329, 249, 167, 86, 33, 25, 22, 24, 24, 67, 120, 162, 177, 158, 131, 
    412, 381, 327, 301, 324, 405, 445, 392, 313, 281, 304, 352, 379, 353, 296, 205, 112, 39, 19, 37, 64, 79, 100, 125, 155, 158, 141, 128, 
    430, 408, 361, 345, 371, 483, 538, 471, 357, 265, 230, 241, 247, 231, 208, 178, 142, 109, 97, 104, 118, 133, 147, 159, 172, 173, 166, 158, 
    380, 420, 409, 407, 443, 513, 494, 382, 252, 176, 147, 125, 122, 124, 126, 131, 130, 132, 138, 144, 155, 169, 183, 192, 196, 199, 198, 198, 
    273, 334, 390, 422, 486, 487, 401, 263, 179, 158, 138, 128, 126, 124, 127, 134, 140, 144, 155, 168, 180, 192, 203, 210, 211, 211, 217, 227, 
    212, 247, 329, 422, 484, 439, 307, 199, 174, 170, 162, 157, 152, 146, 143, 145, 150, 157, 168, 183, 198, 207, 214, 218, 218, 227, 243, 257, 
    199, 207, 281, 409, 480, 407, 262, 178, 173, 171, 169, 164, 159, 153, 151, 154, 161, 169, 181, 197, 211, 215, 212, 208, 223, 244, 263, 278, 
    209, 197, 235, 339, 411, 370, 250, 188, 175, 173, 174, 170, 164, 159, 160, 165, 173, 180, 188, 200, 208, 210, 211, 218, 231, 246, 250, 243, 
    217, 202, 198, 232, 270, 260, 209, 176, 171, 181, 187, 180, 169, 164, 167, 174, 183, 191, 194, 195, 199, 205, 217, 235, 246, 251, 235, 215, 
    218, 206, 194, 178, 168, 148, 139, 141, 136, 153, 170, 180, 184, 181, 177, 183, 194, 198, 197, 193, 193, 206, 231, 256, 266, 262, 239, 209, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 2, 0, 0, 0, 0, 1, 11, 11, 11, 14, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 7, 5, 0, 0, 0, 0, 9, 15, 14, 27, 37, 24, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 11, 3, 0, 0, 0, 6, 18, 18, 29, 43, 46, 21, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 25, 23, 18, 0, 0, 0, 1, 18, 18, 24, 39, 49, 42, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 30, 36, 32, 0, 0, 0, 0, 12, 21, 18, 24, 45, 52, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 28, 41, 34, 0, 0, 0, 0, 8, 29, 18, 15, 34, 52, 45, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 38, 31, 0, 0, 0, 0, 18, 31, 18, 13, 24, 45, 46, 29, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 5, 10, 26, 22, 0, 0, 0, 0, 30, 35, 23, 13, 14, 30, 37, 35, 
    0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 9, 0, 0, 0, 0, 32, 34, 21, 6, 2, 10, 26, 27, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 1, 18, 7, 0, 0, 0, 3, 31, 34, 20, 0, 0, 0, 14, 16, 
    0, 0, 10, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 12, 3, 0, 0, 0, 0, 29, 35, 25, 0, 0, 0, 5, 5, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 44, 31, 7, 0, 0, 0, 0, 
    0, 0, 16, 15, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 4, 38, 56, 35, 8, 0, 0, 0, 0, 
    0, 0, 17, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 42, 50, 31, 4, 0, 0, 0, 0, 
    0, 0, 9, 18, 0, 0, 0, 13, 7, 0, 0, 0, 0, 0, 4, 0, 0, 6, 16, 28, 45, 42, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 0, 0, 19, 20, 0, 0, 0, 0, 0, 13, 19, 8, 33, 42, 43, 55, 37, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 14, 21, 0, 0, 0, 0, 0, 15, 37, 31, 35, 41, 53, 52, 42, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 40, 13, 0, 0, 0, 0, 31, 49, 55, 56, 48, 49, 44, 44, 32, 17, 0, 0, 9, 14, 
    0, 0, 0, 0, 0, 0, 0, 7, 49, 33, 10, 0, 5, 22, 36, 53, 64, 64, 61, 52, 49, 48, 49, 46, 40, 38, 45, 48, 
    0, 0, 0, 0, 0, 0, 0, 25, 52, 60, 50, 36, 36, 41, 48, 55, 62, 58, 57, 57, 59, 58, 58, 60, 62, 62, 64, 67, 
    0, 0, 0, 0, 0, 0, 5, 49, 65, 66, 56, 58, 59, 58, 62, 63, 66, 65, 63, 64, 65, 63, 61, 64, 62, 62, 60, 60, 
    33, 0, 0, 0, 0, 0, 40, 69, 73, 58, 66, 72, 70, 68, 70, 70, 69, 68, 66, 64, 61, 60, 62, 62, 59, 55, 50, 52, 
    72, 30, 0, 0, 0, 0, 67, 75, 62, 57, 68, 75, 75, 71, 68, 66, 65, 65, 64, 63, 59, 60, 65, 70, 64, 50, 52, 57, 
    88, 60, 15, 0, 0, 18, 78, 74, 57, 55, 63, 71, 75, 74, 67, 64, 63, 66, 68, 68, 67, 68, 71, 69, 59, 56, 67, 74, 
    93, 76, 47, 0, 0, 32, 71, 79, 60, 54, 57, 59, 67, 68, 64, 61, 63, 68, 75, 78, 77, 70, 60, 51, 54, 73, 94, 105, 
    94, 82, 70, 46, 31, 50, 67, 79, 65, 58, 60, 63, 67, 62, 55, 49, 51, 62, 78, 85, 79, 63, 40, 29, 46, 80, 110, 112, 
    
    -- channel=9
    6, 10, 10, 7, 5, 5, 4, 0, 0, 0, 0, 0, 11, 30, 48, 53, 46, 24, 7, 0, 0, 13, 25, 35, 34, 24, 12, 2, 
    9, 13, 14, 12, 11, 13, 11, 0, 0, 4, 17, 27, 53, 77, 83, 70, 39, 5, 0, 0, 0, 0, 0, 6, 20, 30, 24, 7, 
    49, 48, 32, 15, 10, 11, 11, 20, 43, 71, 79, 69, 54, 59, 54, 32, 2, 0, 0, 0, 0, 0, 0, 0, 8, 25, 30, 17, 
    46, 50, 36, 18, 11, 11, 11, 22, 39, 51, 46, 37, 11, 4, 5, 0, 0, 0, 0, 0, 0, 2, 2, 8, 7, 17, 27, 26, 
    0, 0, 0, 2, 8, 8, 6, 13, 24, 31, 14, 0, 0, 0, 0, 0, 0, 8, 16, 10, 2, 12, 26, 21, 13, 6, 18, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 26, 26, 21, 0, 0, 7, 11, 0, 0, 6, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 1, 15, 19, 24, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 32, 62, 79, 78, 29, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 16, 5, 1, 0, 0, 0, 0, 
    0, 0, 12, 22, 31, 32, 48, 65, 75, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 31, 28, 14, 8, 8, 0, 0, 0, 
    0, 0, 18, 40, 39, 33, 47, 49, 47, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 20, 24, 9, 0, 0, 0, 0, 0, 0, 
    0, 1, 6, 22, 21, 16, 13, 8, 0, 0, 0, 0, 29, 28, 8, 0, 0, 2, 19, 30, 26, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 45, 51, 56, 44, 17, 0, 7, 25, 27, 18, 7, 1, 0, 0, 5, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 83, 124, 124, 88, 56, 33, 9, 8, 34, 59, 69, 46, 19, 17, 25, 26, 21, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 84, 102, 85, 43, 14, 0, 0, 0, 18, 47, 75, 83, 75, 54, 30, 19, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 47, 61, 34, 0, 0, 0, 0, 0, 10, 7, 37, 73, 70, 34, 2, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 3, 7, 23, 12, 0, 0, 0, 0, 0, 17, 53, 72, 75, 70, 57, 18, 0, 0, 0, 0, 8, 
    0, 0, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 52, 86, 80, 45, 12, 0, 0, 0, 13, 23, 29, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 32, 23, 20, 20, 26, 21, 2, 0, 0, 0, 0, 7, 17, 18, 
    14, 0, 0, 0, 0, 0, 0, 7, 6, 25, 61, 102, 130, 145, 134, 93, 60, 30, 6, 0, 0, 0, 0, 0, 0, 5, 10, 11, 
    72, 50, 15, 0, 0, 0, 4, 64, 111, 114, 102, 113, 131, 142, 126, 84, 44, 19, 2, 0, 3, 8, 11, 11, 13, 19, 25, 23, 
    82, 91, 48, 6, 0, 8, 69, 131, 147, 115, 81, 73, 80, 81, 71, 56, 35, 22, 17, 18, 19, 19, 21, 22, 21, 22, 23, 23, 
    58, 79, 65, 17, 0, 37, 101, 156, 139, 83, 41, 32, 33, 33, 30, 27, 23, 20, 19, 21, 21, 22, 23, 27, 30, 29, 27, 25, 
    45, 50, 50, 26, 26, 62, 105, 115, 80, 39, 23, 22, 21, 22, 21, 20, 20, 20, 21, 23, 25, 28, 33, 38, 36, 34, 32, 30, 
    33, 36, 25, 45, 82, 119, 122, 85, 45, 24, 25, 23, 21, 20, 21, 22, 22, 24, 26, 28, 34, 39, 41, 37, 37, 36, 40, 55, 
    31, 31, 31, 46, 128, 181, 163, 93, 45, 30, 27, 25, 21, 18, 20, 22, 24, 26, 31, 33, 34, 36, 41, 41, 35, 31, 44, 57, 
    36, 30, 33, 48, 97, 158, 148, 85, 50, 48, 47, 44, 35, 26, 21, 21, 22, 26, 29, 31, 34, 35, 32, 29, 28, 35, 48, 57, 
    39, 35, 32, 43, 62, 88, 87, 59, 37, 39, 44, 53, 59, 54, 42, 33, 28, 29, 29, 30, 30, 26, 21, 24, 33, 48, 58, 61, 
    
    -- channel=10
    76, 81, 83, 79, 81, 82, 83, 73, 59, 62, 77, 98, 97, 104, 111, 96, 66, 42, 35, 35, 35, 43, 48, 54, 58, 61, 63, 66, 
    78, 84, 85, 83, 83, 86, 84, 71, 64, 63, 80, 99, 101, 102, 92, 61, 36, 9, 0, 0, 0, 0, 2, 17, 35, 47, 52, 59, 
    80, 81, 77, 83, 86, 88, 87, 80, 84, 82, 97, 95, 83, 70, 53, 34, 5, 0, 0, 0, 0, 0, 0, 0, 1, 9, 31, 45, 
    61, 58, 69, 81, 87, 87, 87, 86, 76, 77, 79, 74, 52, 36, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 29, 
    18, 10, 43, 81, 89, 89, 86, 86, 64, 41, 31, 32, 26, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 3, 68, 89, 78, 79, 77, 68, 47, 23, 17, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 66, 77, 52, 40, 40, 59, 31, 8, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 76, 71, 51, 13, 26, 37, 25, 5, 10, 12, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 75, 79, 52, 6, 19, 44, 38, 12, 2, 15, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 75, 80, 40, 4, 0, 31, 21, 3, 7, 17, 8, 0, 0, 0, 0, 0, 13, 24, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 69, 83, 61, 9, 0, 0, 0, 0, 23, 25, 1, 0, 0, 0, 0, 0, 5, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 37, 72, 76, 33, 0, 0, 0, 0, 29, 37, 13, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 52, 46, 0, 0, 0, 0, 30, 28, 23, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 30, 0, 0, 0, 16, 18, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 17, 0, 0, 28, 19, 9, 0, 0, 0, 0, 0, 0, 17, 15, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 21, 26, 3, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 14, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 26, 24, 0, 0, 0, 0, 0, 0, 0, 38, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 
    0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 54, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 29, 53, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 36, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    49, 36, 34, 36, 38, 38, 39, 37, 25, 14, 14, 29, 38, 37, 45, 62, 82, 99, 112, 119, 123, 127, 125, 119, 105, 86, 69, 63, 
    47, 36, 34, 35, 38, 38, 39, 33, 21, 6, 8, 28, 53, 65, 87, 105, 117, 117, 114, 114, 120, 125, 129, 133, 135, 121, 95, 75, 
    72, 68, 53, 43, 39, 40, 43, 41, 46, 40, 40, 62, 94, 119, 138, 148, 140, 121, 108, 106, 114, 121, 131, 136, 151, 149, 128, 94, 
    126, 130, 98, 59, 40, 35, 41, 61, 79, 84, 97, 117, 120, 137, 151, 155, 145, 129, 115, 117, 129, 142, 144, 151, 160, 173, 155, 118, 
    150, 159, 116, 70, 42, 32, 32, 60, 85, 103, 107, 98, 99, 121, 143, 150, 166, 155, 136, 128, 147, 166, 171, 178, 186, 187, 170, 139, 
    124, 133, 97, 64, 47, 28, 16, 19, 42, 63, 68, 68, 85, 120, 155, 178, 197, 184, 155, 136, 147, 165, 181, 190, 194, 183, 180, 161, 
    105, 91, 68, 57, 51, 27, 4, 0, 0, 13, 41, 59, 92, 145, 176, 204, 217, 202, 156, 123, 125, 142, 164, 177, 178, 178, 175, 174, 
    108, 77, 49, 57, 52, 47, 17, 0, 0, 0, 22, 52, 93, 142, 175, 192, 206, 188, 128, 89, 93, 123, 147, 161, 163, 166, 168, 173, 
    122, 93, 61, 67, 59, 86, 78, 48, 15, 28, 33, 47, 75, 111, 155, 162, 176, 152, 97, 67, 87, 129, 158, 167, 164, 160, 160, 162, 
    145, 105, 82, 77, 74, 106, 134, 123, 113, 89, 57, 43, 53, 88, 126, 136, 156, 133, 90, 79, 115, 162, 185, 184, 175, 167, 154, 147, 
    158, 109, 98, 101, 90, 95, 138, 142, 133, 108, 60, 45, 48, 80, 108, 120, 154, 132, 105, 104, 146, 180, 195, 191, 184, 171, 153, 138, 
    141, 100, 107, 128, 106, 87, 114, 124, 124, 92, 53, 48, 77, 100, 106, 126, 164, 145, 117, 118, 148, 169, 181, 183, 178, 160, 147, 137, 
    111, 94, 108, 135, 111, 96, 108, 114, 112, 81, 58, 72, 117, 147, 136, 154, 176, 154, 121, 122, 147, 164, 178, 178, 172, 156, 149, 142, 
    88, 88, 101, 122, 106, 103, 102, 126, 131, 120, 107, 136, 166, 177, 165, 177, 185, 163, 144, 138, 152, 166, 190, 195, 182, 171, 158, 140, 
    81, 85, 100, 115, 113, 114, 102, 136, 166, 177, 186, 200, 204, 182, 168, 171, 168, 159, 172, 181, 181, 193, 211, 219, 202, 178, 145, 104, 
    84, 86, 113, 123, 133, 119, 117, 140, 175, 200, 219, 194, 165, 146, 135, 154, 153, 148, 168, 192, 207, 223, 229, 220, 190, 146, 103, 76, 
    100, 98, 120, 132, 146, 124, 122, 126, 138, 173, 169, 143, 111, 102, 104, 143, 146, 151, 162, 189, 219, 238, 221, 187, 152, 109, 79, 69, 
    114, 106, 119, 132, 145, 128, 107, 95, 109, 148, 126, 105, 80, 69, 90, 134, 155, 185, 202, 218, 234, 229, 191, 166, 143, 118, 98, 95, 
    118, 107, 115, 128, 148, 127, 72, 48, 72, 93, 104, 92, 79, 78, 98, 138, 179, 215, 245, 255, 239, 219, 188, 175, 159, 155, 147, 151, 
    124, 109, 104, 119, 145, 100, 45, 29, 67, 92, 117, 116, 119, 131, 151, 171, 196, 222, 235, 233, 220, 212, 205, 201, 193, 192, 197, 202, 
    151, 131, 108, 113, 131, 66, 41, 61, 113, 169, 210, 238, 254, 265, 264, 253, 244, 236, 233, 230, 227, 222, 225, 231, 236, 238, 243, 244, 
    224, 185, 138, 128, 112, 72, 85, 145, 234, 289, 305, 297, 302, 302, 297, 287, 277, 263, 254, 248, 248, 247, 248, 250, 254, 254, 254, 251, 
    272, 248, 186, 166, 121, 105, 139, 217, 287, 304, 281, 263, 265, 269, 272, 273, 275, 273, 270, 265, 261, 260, 257, 256, 256, 253, 248, 246, 
    286, 264, 231, 198, 153, 132, 170, 255, 294, 277, 254, 249, 253, 259, 265, 269, 272, 273, 270, 265, 262, 261, 259, 261, 258, 255, 251, 248, 
    281, 267, 246, 224, 180, 155, 198, 273, 282, 259, 254, 256, 260, 263, 265, 264, 264, 265, 266, 266, 266, 265, 264, 266, 273, 273, 267, 261, 
    276, 268, 264, 256, 236, 220, 250, 284, 274, 256, 254, 256, 257, 257, 259, 259, 259, 261, 265, 272, 276, 276, 275, 274, 276, 272, 269, 272, 
    274, 266, 274, 282, 282, 291, 317, 312, 290, 277, 267, 258, 253, 251, 253, 252, 252, 257, 264, 274, 280, 280, 275, 269, 261, 255, 257, 280, 
    274, 268, 273, 286, 290, 309, 333, 325, 303, 299, 294, 286, 276, 265, 257, 249, 247, 250, 258, 268, 275, 277, 268, 256, 244, 244, 254, 281, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 1, 22, 23, 19, 20, 29, 26, 20, 4, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 27, 9, 0, 0, 0, 0, 0, 25, 50, 54, 49, 35, 26, 14, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 41, 75, 75, 58, 41, 46, 47, 28, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 37, 66, 98, 88, 57, 28, 27, 30, 20, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 25, 14, 14, 23, 39, 60, 74, 64, 39, 12, 0, 0, 0, 0, 0, 0, 0, 
    41, 12, 0, 0, 0, 2, 56, 65, 38, 28, 47, 29, 11, 4, 11, 8, 24, 35, 41, 32, 17, 4, 0, 1, 0, 0, 0, 0, 
    116, 64, 0, 0, 0, 56, 192, 213, 169, 103, 70, 31, 4, 0, 0, 0, 3, 39, 74, 65, 51, 36, 25, 25, 9, 0, 0, 0, 
    146, 101, 9, 0, 0, 28, 154, 202, 182, 129, 88, 46, 7, 0, 0, 0, 12, 82, 122, 96, 72, 53, 46, 41, 31, 12, 0, 0, 
    140, 124, 43, 0, 0, 0, 66, 121, 118, 103, 103, 83, 47, 12, 0, 7, 42, 113, 137, 98, 60, 37, 37, 32, 31, 21, 0, 0, 
    137, 128, 33, 0, 0, 0, 18, 58, 68, 91, 126, 129, 105, 77, 37, 42, 72, 126, 130, 88, 52, 27, 22, 15, 17, 19, 4, 0, 
    130, 114, 27, 0, 0, 0, 0, 31, 75, 137, 163, 156, 131, 123, 78, 58, 78, 117, 119, 84, 60, 38, 31, 34, 39, 37, 12, 0, 
    133, 113, 58, 8, 0, 0, 0, 44, 137, 221, 221, 180, 141, 114, 74, 44, 58, 98, 122, 108, 75, 43, 44, 65, 72, 46, 0, 0, 
    152, 133, 101, 47, 20, 0, 0, 45, 155, 222, 200, 151, 98, 62, 37, 21, 28, 73, 103, 122, 102, 72, 72, 74, 59, 8, 0, 0, 
    177, 152, 123, 84, 61, 46, 25, 31, 79, 100, 79, 60, 29, 24, 18, 15, 10, 17, 33, 83, 97, 82, 61, 28, 0, 0, 0, 0, 
    194, 161, 128, 104, 85, 85, 67, 46, 27, 26, 36, 33, 21, 31, 31, 30, 31, 35, 56, 75, 61, 52, 29, 0, 0, 0, 0, 0, 
    199, 165, 139, 117, 97, 91, 79, 51, 24, 16, 35, 48, 57, 54, 43, 35, 62, 96, 119, 95, 50, 42, 32, 13, 0, 0, 0, 0, 
    192, 164, 147, 122, 103, 92, 90, 37, 12, 12, 41, 98, 141, 133, 110, 72, 59, 70, 80, 67, 51, 43, 54, 55, 59, 60, 57, 57, 
    210, 174, 138, 100, 109, 129, 137, 114, 90, 114, 170, 236, 272, 261, 229, 160, 92, 54, 41, 46, 62, 71, 86, 97, 109, 109, 108, 106, 
    265, 225, 150, 107, 129, 205, 244, 261, 259, 245, 258, 288, 296, 277, 244, 186, 125, 89, 82, 87, 99, 115, 127, 135, 137, 134, 132, 130, 
    278, 279, 210, 180, 184, 261, 304, 307, 279, 241, 207, 194, 190, 179, 163, 144, 125, 120, 121, 126, 133, 140, 147, 150, 153, 154, 153, 152, 
    227, 261, 247, 227, 236, 289, 302, 260, 211, 174, 141, 127, 125, 124, 123, 125, 125, 126, 134, 140, 143, 148, 153, 159, 161, 163, 164, 162, 
    196, 203, 224, 252, 283, 295, 256, 195, 172, 152, 133, 127, 122, 120, 120, 120, 122, 129, 137, 144, 151, 160, 169, 176, 178, 180, 179, 180, 
    176, 178, 195, 274, 325, 295, 215, 163, 155, 143, 136, 130, 124, 122, 122, 124, 130, 138, 148, 159, 170, 179, 183, 179, 180, 188, 202, 220, 
    164, 169, 199, 261, 332, 305, 235, 181, 159, 141, 137, 130, 124, 124, 129, 135, 142, 149, 159, 168, 176, 179, 177, 171, 176, 197, 220, 223, 
    164, 166, 196, 236, 264, 272, 236, 193, 163, 157, 155, 148, 138, 129, 129, 137, 146, 152, 156, 162, 165, 164, 164, 170, 187, 204, 203, 180, 
    166, 165, 174, 196, 185, 175, 176, 163, 143, 154, 163, 164, 162, 152, 147, 148, 150, 151, 151, 150, 149, 150, 160, 183, 201, 202, 180, 158, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 37, 41, 39, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 35, 39, 19, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    191, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 55, 45, 12, 0, 0, 0, 0, 2, 5, 0, 0, 
    223, 82, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 51, 91, 78, 34, 4, 0, 2, 1, 6, 15, 9, 0, 
    233, 86, 0, 0, 0, 0, 0, 0, 0, 0, 18, 18, 0, 0, 0, 0, 81, 112, 89, 31, 7, 0, 5, 0, 1, 14, 10, 0, 
    226, 94, 0, 0, 0, 0, 0, 0, 0, 22, 32, 29, 13, 12, 0, 6, 88, 103, 77, 22, 20, 15, 17, 9, 9, 8, 0, 0, 
    227, 127, 12, 0, 0, 0, 0, 0, 0, 69, 56, 22, 7, 2, 0, 0, 48, 58, 44, 23, 33, 26, 28, 31, 23, 0, 0, 0, 
    239, 170, 102, 29, 0, 0, 0, 0, 8, 53, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 17, 22, 5, 0, 0, 0, 
    270, 217, 164, 128, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    296, 254, 209, 178, 128, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    286, 265, 222, 192, 179, 108, 46, 0, 0, 0, 0, 0, 0, 10, 21, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    246, 244, 212, 190, 194, 155, 103, 49, 0, 0, 0, 18, 51, 64, 62, 55, 0, 0, 0, 0, 0, 29, 58, 31, 0, 0, 0, 0, 
    220, 219, 193, 181, 201, 201, 144, 83, 64, 57, 74, 119, 145, 155, 136, 108, 17, 0, 0, 38, 95, 139, 153, 132, 66, 0, 0, 0, 
    242, 230, 188, 164, 212, 227, 217, 193, 194, 178, 184, 184, 189, 185, 177, 170, 128, 92, 126, 178, 222, 252, 268, 271, 230, 174, 137, 132, 
    274, 261, 217, 185, 244, 257, 262, 243, 251, 251, 240, 221, 203, 195, 215, 243, 254, 260, 282, 304, 327, 351, 374, 386, 379, 360, 349, 354, 
    301, 283, 246, 231, 281, 274, 266, 247, 256, 271, 251, 220, 209, 220, 250, 291, 325, 345, 366, 382, 397, 413, 428, 440, 446, 448, 447, 451, 
    334, 292, 262, 278, 312, 267, 225, 207, 257, 307, 327, 318, 318, 324, 338, 357, 373, 383, 401, 416, 430, 444, 454, 462, 466, 472, 478, 485, 
    401, 321, 286, 331, 337, 277, 219, 268, 343, 387, 396, 390, 385, 377, 376, 380, 388, 402, 421, 439, 454, 468, 475, 479, 482, 492, 508, 516, 
    464, 389, 347, 366, 339, 281, 248, 334, 389, 405, 406, 401, 394, 384, 383, 390, 403, 419, 440, 462, 476, 485, 489, 490, 497, 514, 527, 527, 
    498, 449, 407, 379, 307, 258, 281, 369, 396, 403, 408, 406, 402, 393, 394, 403, 418, 437, 455, 474, 485, 487, 484, 488, 508, 535, 542, 526, 
    515, 484, 440, 385, 284, 237, 285, 368, 380, 392, 398, 401, 404, 400, 403, 411, 428, 446, 460, 469, 472, 468, 473, 491, 524, 555, 548, 504, 
    515, 492, 459, 400, 313, 257, 294, 353, 367, 379, 386, 387, 385, 385, 394, 411, 433, 450, 459, 461, 456, 453, 464, 493, 534, 560, 547, 500, 
    
    -- channel=14
    234, 226, 224, 226, 230, 230, 229, 230, 233, 234, 230, 222, 222, 210, 193, 185, 187, 191, 191, 186, 186, 182, 183, 187, 199, 209, 214, 211, 
    233, 228, 226, 225, 229, 227, 227, 225, 216, 204, 195, 189, 191, 174, 162, 159, 166, 176, 177, 165, 164, 174, 189, 196, 200, 208, 214, 212, 
    211, 223, 232, 232, 230, 230, 229, 221, 203, 177, 163, 156, 162, 157, 153, 157, 165, 170, 150, 116, 111, 129, 152, 165, 182, 203, 215, 217, 
    190, 217, 236, 239, 235, 234, 233, 234, 223, 203, 185, 166, 170, 165, 165, 171, 176, 178, 153, 108, 96, 105, 119, 126, 152, 187, 214, 219, 
    188, 239, 260, 245, 235, 231, 228, 227, 218, 210, 199, 183, 153, 137, 148, 162, 170, 174, 158, 124, 100, 109, 107, 106, 122, 160, 207, 223, 
    155, 228, 266, 251, 237, 235, 230, 217, 198, 185, 176, 146, 112, 104, 122, 143, 162, 180, 170, 142, 115, 120, 122, 110, 115, 144, 186, 215, 
    100, 182, 222, 224, 232, 226, 216, 180, 137, 131, 142, 120, 96, 92, 109, 135, 168, 197, 197, 162, 120, 118, 131, 128, 120, 128, 157, 196, 
    89, 163, 194, 200, 207, 192, 168, 123, 81, 81, 116, 107, 85, 92, 109, 128, 164, 200, 207, 153, 94, 91, 113, 137, 123, 115, 134, 176, 
    99, 170, 178, 192, 196, 190, 163, 124, 80, 75, 108, 110, 78, 89, 104, 117, 158, 189, 186, 113, 65, 71, 99, 137, 130, 108, 117, 151, 
    109, 171, 157, 174, 203, 209, 192, 164, 130, 110, 131, 122, 77, 77, 100, 108, 150, 190, 172, 91, 43, 69, 100, 138, 138, 115, 113, 133, 
    108, 151, 136, 157, 196, 195, 198, 199, 209, 169, 158, 117, 79, 71, 85, 106, 144, 189, 168, 88, 47, 80, 113, 149, 153, 138, 125, 133, 
    102, 135, 119, 157, 201, 196, 186, 201, 223, 193, 156, 90, 66, 69, 80, 112, 146, 184, 162, 87, 56, 83, 122, 156, 168, 159, 141, 149, 
    88, 107, 83, 138, 212, 212, 186, 197, 217, 182, 127, 70, 64, 77, 88, 126, 161, 193, 160, 92, 57, 70, 99, 140, 162, 157, 162, 176, 
    75, 80, 49, 85, 180, 208, 184, 181, 180, 146, 89, 64, 85, 116, 120, 152, 176, 183, 155, 119, 88, 77, 96, 136, 165, 173, 185, 194, 
    64, 66, 35, 42, 129, 190, 178, 182, 177, 149, 104, 104, 115, 149, 152, 175, 198, 183, 150, 104, 74, 62, 97, 147, 187, 203, 210, 216, 
    65, 64, 35, 21, 84, 158, 163, 169, 173, 184, 164, 176, 169, 160, 144, 172, 210, 208, 179, 128, 87, 73, 111, 169, 207, 220, 225, 219, 
    77, 70, 42, 23, 62, 135, 151, 119, 128, 156, 176, 191, 164, 129, 103, 125, 155, 150, 135, 118, 103, 97, 133, 188, 213, 222, 221, 214, 
    101, 81, 49, 30, 58, 133, 146, 83, 77, 119, 171, 192, 151, 101, 70, 76, 116, 103, 74, 79, 80, 98, 128, 172, 197, 200, 199, 194, 
    125, 89, 55, 34, 64, 132, 144, 62, 43, 81, 123, 148, 108, 53, 26, 39, 97, 116, 85, 77, 81, 94, 105, 134, 160, 163, 150, 139, 
    137, 96, 71, 61, 92, 146, 112, 3, 0, 0, 44, 72, 48, 0, 0, 0, 33, 69, 76, 65, 58, 50, 49, 72, 97, 110, 100, 90, 
    120, 88, 78, 81, 116, 158, 73, 0, 0, 0, 12, 43, 33, 0, 0, 0, 0, 13, 23, 25, 25, 21, 18, 19, 30, 40, 37, 28, 
    87, 79, 79, 111, 144, 139, 30, 0, 0, 0, 29, 70, 68, 47, 31, 15, 13, 17, 17, 14, 10, 7, 4, 0, 0, 0, 0, 0, 
    80, 91, 115, 149, 169, 110, 0, 0, 0, 0, 17, 27, 26, 23, 20, 16, 15, 14, 11, 6, 1, 0, 0, 0, 0, 0, 0, 0, 
    44, 83, 127, 171, 171, 74, 0, 0, 0, 0, 0, 0, 0, 4, 7, 6, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 100, 158, 148, 33, 0, 0, 0, 7, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 59, 113, 98, 0, 0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 35, 77, 72, 4, 0, 0, 3, 7, 3, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 56, 36, 0, 0, 18, 18, 8, 0, 0, 0, 5, 8, 3, 0, 0, 0, 0, 0, 7, 12, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 21, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 27, 35, 3, 0, 0, 0, 0, 0, 0, 
    47, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 22, 0, 0, 0, 0, 0, 0, 49, 43, 5, 0, 0, 0, 0, 0, 0, 
    54, 41, 14, 0, 0, 0, 0, 0, 0, 0, 0, 28, 36, 0, 0, 0, 0, 0, 0, 41, 32, 1, 0, 0, 0, 0, 0, 0, 
    63, 63, 49, 0, 0, 0, 0, 0, 0, 0, 18, 47, 37, 0, 0, 0, 0, 0, 0, 30, 26, 2, 0, 0, 0, 0, 0, 0, 
    76, 78, 91, 0, 0, 0, 0, 0, 0, 0, 20, 36, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    99, 92, 121, 57, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    122, 111, 133, 103, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    120, 115, 129, 126, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    100, 101, 111, 128, 67, 7, 20, 39, 9, 0, 0, 0, 0, 12, 42, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    87, 91, 103, 122, 72, 10, 23, 58, 50, 0, 0, 0, 14, 50, 85, 46, 4, 0, 0, 1, 0, 4, 2, 0, 0, 0, 0, 0, 
    94, 94, 100, 106, 58, 25, 57, 110, 131, 85, 40, 41, 68, 97, 121, 99, 55, 31, 31, 41, 51, 63, 76, 67, 57, 54, 62, 65, 
    100, 101, 96, 94, 50, 40, 99, 199, 217, 166, 116, 103, 111, 126, 140, 133, 112, 93, 87, 89, 99, 112, 125, 130, 127, 127, 134, 138, 
    114, 100, 102, 87, 53, 74, 166, 249, 244, 176, 124, 107, 111, 117, 126, 127, 123, 119, 117, 125, 133, 138, 143, 150, 153, 154, 157, 159, 
    130, 101, 95, 80, 68, 119, 220, 254, 207, 158, 129, 122, 120, 119, 121, 122, 122, 123, 126, 135, 143, 148, 154, 162, 167, 167, 165, 166, 
    150, 112, 89, 65, 83, 158, 254, 245, 183, 144, 136, 136, 130, 123, 120, 119, 121, 127, 134, 143, 153, 162, 171, 178, 179, 173, 175, 186, 
    176, 137, 100, 68, 90, 188, 260, 221, 157, 134, 137, 140, 134, 126, 123, 123, 128, 136, 147, 159, 166, 174, 183, 183, 180, 177, 189, 206, 
    190, 165, 128, 83, 84, 175, 233, 188, 136, 128, 134, 139, 137, 132, 128, 130, 137, 146, 157, 166, 172, 176, 175, 175, 178, 189, 208, 223, 
    196, 178, 160, 116, 103, 150, 195, 162, 126, 121, 128, 136, 138, 134, 131, 132, 140, 151, 161, 168, 167, 162, 155, 159, 175, 204, 224, 230, 
    195, 179, 170, 143, 120, 136, 156, 139, 120, 119, 125, 129, 129, 127, 124, 127, 138, 152, 165, 167, 158, 146, 138, 149, 182, 221, 239, 223, 
    
    -- channel=16
    102, 99, 101, 105, 110, 112, 113, 115, 117, 111, 113, 112, 111, 105, 98, 98, 100, 98, 98, 92, 88, 82, 83, 85, 88, 95, 99, 102, 
    104, 101, 102, 105, 108, 110, 111, 117, 117, 107, 104, 92, 89, 85, 82, 86, 88, 87, 80, 66, 62, 60, 62, 69, 77, 86, 94, 102, 
    97, 97, 101, 107, 110, 112, 112, 110, 98, 94, 103, 92, 96, 89, 84, 78, 75, 69, 64, 55, 55, 56, 61, 59, 65, 71, 82, 91, 
    99, 98, 105, 108, 110, 110, 111, 103, 97, 104, 105, 98, 90, 76, 64, 64, 62, 58, 50, 44, 44, 44, 46, 46, 53, 60, 64, 78, 
    84, 85, 96, 111, 115, 116, 117, 110, 103, 100, 95, 78, 75, 73, 66, 59, 57, 49, 44, 39, 41, 40, 39, 36, 42, 47, 50, 66, 
    61, 74, 90, 103, 120, 124, 121, 113, 114, 106, 99, 79, 70, 66, 57, 47, 46, 44, 48, 51, 53, 49, 48, 43, 38, 35, 44, 57, 
    61, 71, 89, 100, 119, 126, 115, 96, 87, 77, 72, 63, 56, 55, 48, 44, 42, 46, 49, 56, 51, 53, 51, 45, 36, 36, 36, 47, 
    53, 66, 83, 98, 111, 104, 85, 63, 56, 60, 49, 50, 51, 47, 40, 40, 41, 36, 48, 50, 40, 51, 57, 53, 46, 38, 37, 45, 
    43, 58, 81, 91, 92, 76, 49, 41, 34, 39, 40, 45, 51, 47, 44, 43, 50, 42, 44, 41, 36, 46, 53, 56, 52, 40, 35, 37, 
    31, 43, 70, 77, 78, 65, 39, 25, 44, 42, 58, 55, 55, 57, 45, 48, 49, 47, 34, 36, 33, 42, 46, 53, 53, 46, 40, 42, 
    20, 31, 62, 72, 88, 73, 44, 31, 38, 44, 54, 50, 52, 55, 49, 51, 54, 41, 30, 39, 38, 43, 47, 59, 60, 50, 47, 53, 
    16, 17, 56, 71, 95, 97, 77, 64, 68, 57, 59, 46, 50, 43, 42, 51, 48, 39, 31, 36, 23, 33, 36, 50, 57, 48, 51, 62, 
    21, 7, 42, 68, 89, 106, 95, 80, 70, 41, 31, 22, 31, 32, 39, 50, 40, 39, 38, 42, 34, 43, 53, 53, 52, 47, 54, 64, 
    22, 6, 24, 53, 86, 106, 100, 77, 43, 24, 1, 11, 21, 30, 48, 59, 45, 30, 35, 26, 22, 27, 33, 37, 41, 52, 62, 73, 
    23, 11, 13, 38, 69, 88, 93, 72, 34, 37, 32, 41, 51, 49, 62, 63, 53, 57, 58, 40, 23, 18, 22, 31, 42, 52, 65, 72, 
    21, 15, 8, 22, 46, 60, 75, 65, 47, 32, 35, 36, 33, 45, 57, 63, 65, 64, 59, 30, 27, 25, 29, 32, 41, 53, 69, 82, 
    22, 18, 8, 12, 31, 49, 60, 49, 43, 41, 40, 61, 56, 45, 49, 54, 50, 48, 33, 17, 6, 13, 24, 33, 49, 63, 79, 92, 
    28, 21, 8, 9, 18, 21, 29, 36, 45, 63, 58, 59, 60, 34, 29, 46, 44, 52, 43, 30, 34, 28, 34, 59, 64, 75, 88, 99, 
    38, 27, 12, 21, 22, 26, 7, 0, 8, 22, 45, 34, 23, 2, 0, 4, 25, 26, 25, 20, 13, 12, 17, 37, 53, 75, 90, 99, 
    27, 23, 17, 23, 19, 24, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 6, 21, 30, 29, 
    0, 0, 8, 24, 28, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 31, 40, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    81, 89, 95, 99, 106, 108, 104, 94, 101, 134, 145, 129, 98, 79, 64, 34, 3, 0, 0, 0, 0, 0, 0, 13, 35, 48, 53, 53, 
    88, 91, 94, 99, 106, 107, 102, 98, 130, 186, 191, 137, 75, 39, 1, 0, 0, 0, 25, 48, 46, 17, 0, 0, 3, 24, 41, 54, 
    74, 72, 76, 89, 100, 101, 96, 89, 115, 168, 178, 105, 24, 0, 0, 0, 0, 25, 97, 136, 132, 98, 64, 26, 5, 0, 16, 44, 
    20, 27, 57, 84, 96, 97, 91, 63, 50, 66, 75, 37, 0, 0, 0, 0, 0, 60, 141, 180, 171, 133, 97, 65, 15, 0, 0, 35, 
    0, 0, 59, 102, 103, 98, 93, 61, 17, 0, 11, 47, 45, 17, 2, 0, 19, 70, 150, 178, 158, 108, 79, 53, 16, 0, 0, 13, 
    43, 45, 101, 126, 105, 89, 97, 90, 66, 52, 90, 136, 134, 88, 46, 22, 10, 36, 122, 166, 139, 83, 44, 26, 17, 0, 0, 0, 
    172, 174, 201, 166, 103, 85, 141, 195, 193, 162, 169, 192, 168, 103, 47, 16, 0, 0, 80, 162, 161, 100, 39, 24, 29, 20, 0, 0, 
    245, 266, 288, 212, 101, 83, 177, 301, 328, 278, 237, 236, 201, 120, 53, 10, 0, 0, 94, 200, 219, 149, 77, 46, 55, 44, 4, 0, 
    279, 326, 348, 240, 90, 33, 104, 289, 366, 325, 276, 279, 244, 164, 89, 37, 0, 44, 166, 265, 258, 168, 84, 50, 62, 62, 33, 0, 
    276, 335, 371, 253, 85, 0, 0, 137, 263, 275, 288, 328, 299, 218, 133, 83, 36, 88, 220, 302, 250, 138, 61, 36, 46, 62, 63, 45, 
    271, 320, 356, 243, 99, 0, 0, 26, 146, 213, 286, 366, 344, 256, 183, 126, 68, 111, 235, 292, 219, 114, 49, 22, 33, 60, 90, 95, 
    286, 313, 321, 206, 106, 35, 0, 20, 118, 216, 306, 371, 353, 263, 199, 139, 82, 123, 228, 273, 211, 121, 53, 21, 33, 72, 112, 124, 
    318, 329, 318, 210, 117, 63, 18, 27, 124, 255, 332, 332, 279, 210, 169, 118, 74, 118, 216, 256, 211, 140, 75, 42, 54, 93, 120, 122, 
    355, 361, 354, 259, 162, 120, 78, 48, 112, 221, 290, 244, 163, 120, 114, 90, 73, 100, 155, 187, 175, 122, 52, 19, 36, 78, 100, 104, 
    391, 393, 386, 298, 208, 168, 135, 73, 58, 114, 156, 133, 96, 72, 83, 95, 82, 66, 81, 111, 118, 72, 0, 0, 1, 50, 83, 100, 
    410, 413, 402, 320, 230, 194, 190, 109, 33, 1, 20, 49, 73, 93, 117, 127, 100, 56, 20, 23, 43, 2, 0, 0, 0, 65, 110, 127, 
    405, 415, 403, 333, 235, 197, 220, 197, 103, 22, 26, 74, 135, 175, 185, 164, 126, 87, 23, 0, 0, 0, 0, 0, 35, 96, 130, 127, 
    383, 404, 398, 344, 235, 188, 229, 265, 197, 90, 69, 119, 209, 268, 262, 202, 121, 70, 18, 0, 0, 0, 0, 32, 84, 111, 116, 94, 
    364, 392, 380, 337, 240, 228, 304, 354, 297, 188, 148, 176, 267, 333, 313, 226, 94, 0, 0, 0, 0, 0, 3, 51, 85, 101, 88, 61, 
    348, 377, 363, 323, 261, 298, 428, 495, 424, 284, 198, 189, 235, 266, 257, 206, 103, 0, 0, 0, 18, 38, 60, 77, 93, 92, 77, 60, 
    294, 345, 365, 338, 297, 358, 508, 553, 442, 277, 154, 118, 113, 112, 121, 125, 109, 75, 63, 71, 88, 104, 119, 129, 131, 129, 126, 121, 
    204, 272, 341, 345, 344, 418, 500, 464, 317, 151, 53, 12, 0, 4, 25, 55, 81, 95, 106, 117, 128, 138, 151, 164, 170, 175, 177, 177, 
    125, 166, 245, 296, 362, 438, 449, 323, 157, 83, 73, 72, 70, 69, 79, 94, 105, 109, 118, 133, 147, 158, 171, 184, 188, 187, 189, 198, 
    132, 113, 150, 221, 347, 431, 402, 252, 136, 123, 142, 143, 135, 126, 118, 116, 118, 122, 131, 147, 163, 177, 189, 199, 197, 194, 208, 227, 
    177, 129, 118, 172, 291, 396, 349, 217, 134, 139, 151, 151, 141, 129, 123, 122, 126, 136, 148, 163, 178, 191, 199, 195, 190, 198, 221, 243, 
    205, 163, 129, 133, 199, 290, 270, 189, 132, 139, 149, 153, 149, 137, 130, 132, 141, 152, 163, 174, 183, 188, 185, 181, 187, 207, 236, 247, 
    218, 189, 154, 110, 109, 145, 159, 134, 113, 124, 142, 151, 149, 142, 138, 140, 150, 164, 176, 177, 173, 169, 170, 182, 205, 241, 257, 229, 
    219, 195, 172, 123, 72, 63, 70, 82, 84, 95, 113, 130, 137, 135, 131, 136, 156, 176, 187, 185, 171, 158, 161, 187, 234, 275, 275, 229, 
    
    -- channel=18
    311, 313, 314, 314, 317, 318, 318, 312, 297, 300, 308, 317, 313, 301, 278, 247, 218, 191, 170, 162, 162, 170, 179, 195, 216, 242, 263, 272, 
    305, 310, 313, 315, 318, 320, 318, 307, 283, 264, 267, 266, 255, 234, 208, 184, 158, 128, 106, 90, 94, 106, 130, 152, 178, 208, 237, 260, 
    256, 272, 295, 314, 323, 325, 323, 306, 263, 229, 224, 219, 202, 178, 153, 133, 110, 82, 54, 38, 43, 56, 77, 99, 129, 163, 201, 237, 
    206, 230, 273, 310, 326, 328, 324, 301, 261, 222, 206, 184, 162, 133, 113, 98, 76, 47, 22, 16, 20, 28, 37, 55, 80, 114, 164, 209, 
    154, 197, 263, 312, 327, 328, 319, 293, 257, 214, 181, 157, 134, 101, 81, 73, 47, 26, 12, 20, 28, 26, 26, 32, 46, 77, 129, 180, 
    102, 160, 245, 304, 322, 312, 297, 275, 249, 203, 161, 119, 96, 67, 45, 43, 31, 28, 28, 38, 44, 46, 42, 34, 36, 61, 98, 147, 
    38, 113, 217, 278, 300, 269, 225, 192, 179, 146, 111, 76, 63, 48, 30, 35, 31, 30, 42, 53, 56, 54, 50, 45, 39, 48, 75, 118, 
    0, 69, 185, 261, 270, 216, 128, 74, 80, 75, 62, 55, 53, 42, 28, 37, 34, 33, 36, 43, 46, 49, 48, 46, 42, 41, 61, 87, 
    0, 33, 155, 247, 255, 182, 71, 0, 5, 21, 37, 43, 54, 51, 34, 45, 34, 24, 16, 17, 17, 34, 36, 41, 41, 31, 45, 71, 
    0, 6, 121, 224, 241, 183, 69, 8, 12, 33, 34, 37, 57, 54, 39, 54, 25, 8, 0, 0, 0, 20, 27, 37, 39, 30, 36, 66, 
    0, 0, 94, 197, 235, 207, 108, 40, 40, 42, 31, 12, 40, 40, 36, 53, 5, 0, 0, 0, 0, 22, 31, 39, 42, 36, 40, 69, 
    0, 0, 65, 161, 230, 224, 158, 88, 57, 42, 18, 0, 15, 12, 24, 43, 0, 0, 0, 0, 0, 14, 26, 34, 39, 42, 58, 91, 
    0, 0, 28, 105, 196, 213, 182, 106, 47, 0, 0, 0, 0, 8, 20, 41, 15, 7, 0, 5, 5, 18, 24, 29, 35, 45, 75, 120, 
    0, 0, 0, 46, 124, 174, 171, 107, 27, 0, 0, 0, 0, 19, 45, 59, 45, 27, 9, 2, 0, 12, 19, 18, 33, 62, 111, 160, 
    0, 0, 0, 0, 48, 106, 137, 97, 25, 0, 0, 17, 25, 39, 58, 74, 89, 75, 54, 18, 3, 2, 7, 21, 52, 96, 151, 200, 
    0, 0, 0, 0, 0, 38, 77, 73, 43, 22, 26, 57, 57, 42, 59, 62, 88, 93, 73, 37, 20, 12, 17, 41, 86, 141, 194, 229, 
    0, 0, 0, 0, 0, 0, 19, 30, 47, 42, 62, 69, 49, 22, 41, 32, 63, 65, 41, 11, 8, 10, 25, 63, 120, 175, 217, 242, 
    0, 0, 0, 0, 0, 0, 0, 13, 42, 40, 51, 43, 12, 0, 4, 9, 40, 34, 11, 0, 0, 0, 17, 45, 93, 137, 174, 192, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 53, 76, 82, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    277, 267, 267, 278, 287, 288, 284, 275, 274, 272, 284, 280, 272, 259, 237, 215, 209, 205, 196, 185, 185, 188, 199, 214, 235, 243, 242, 233, 
    276, 272, 273, 281, 288, 289, 286, 284, 292, 299, 299, 274, 244, 218, 191, 172, 170, 173, 176, 169, 157, 151, 160, 181, 206, 230, 245, 245, 
    267, 277, 288, 289, 287, 286, 287, 293, 310, 313, 294, 255, 214, 175, 138, 120, 145, 189, 211, 197, 177, 163, 159, 163, 179, 206, 234, 246, 
    231, 270, 297, 299, 288, 283, 286, 298, 296, 280, 256, 216, 159, 108, 96, 123, 175, 229, 250, 230, 201, 185, 167, 148, 140, 164, 215, 240, 
    160, 227, 291, 304, 292, 282, 281, 277, 257, 232, 216, 199, 158, 123, 132, 166, 207, 262, 285, 265, 224, 203, 173, 133, 111, 130, 183, 230, 
    126, 210, 291, 309, 288, 274, 258, 237, 215, 212, 228, 223, 185, 150, 150, 175, 206, 264, 289, 274, 229, 192, 160, 120, 102, 107, 148, 206, 
    154, 242, 312, 318, 284, 273, 261, 247, 214, 220, 248, 245, 206, 165, 149, 159, 182, 229, 262, 270, 231, 176, 145, 130, 110, 98, 112, 164, 
    231, 303, 349, 330, 282, 270, 310, 317, 291, 267, 282, 261, 214, 171, 140, 127, 144, 198, 259, 278, 237, 182, 159, 159, 132, 102, 89, 118, 
    306, 380, 394, 338, 284, 263, 323, 351, 354, 321, 317, 290, 230, 184, 145, 113, 141, 217, 292, 293, 235, 187, 168, 179, 158, 111, 86, 93, 
    336, 415, 409, 342, 294, 245, 277, 330, 367, 359, 359, 333, 266, 202, 161, 139, 162, 251, 330, 308, 222, 179, 167, 183, 176, 138, 108, 107, 
    330, 404, 382, 331, 294, 234, 227, 278, 338, 359, 383, 366, 311, 243, 191, 180, 198, 292, 353, 305, 208, 169, 163, 177, 184, 170, 148, 149, 
    324, 364, 317, 293, 286, 247, 224, 259, 324, 376, 408, 377, 332, 284, 220, 213, 236, 322, 350, 296, 205, 163, 159, 175, 193, 209, 209, 207, 
    321, 329, 271, 255, 280, 268, 232, 256, 331, 400, 400, 352, 315, 287, 240, 236, 262, 329, 342, 298, 224, 179, 161, 187, 222, 241, 251, 253, 
    333, 325, 270, 230, 268, 291, 266, 280, 338, 389, 373, 315, 272, 259, 233, 254, 284, 314, 308, 287, 224, 163, 145, 181, 229, 254, 274, 270, 
    356, 343, 291, 222, 253, 304, 293, 288, 314, 333, 304, 277, 248, 230, 225, 267, 299, 303, 281, 257, 203, 143, 132, 166, 224, 251, 265, 268, 
    385, 364, 308, 236, 238, 303, 307, 283, 256, 241, 224, 239, 233, 217, 225, 264, 295, 269, 222, 195, 153, 100, 100, 140, 200, 242, 269, 274, 
    420, 388, 327, 259, 230, 282, 307, 269, 212, 194, 229, 262, 263, 233, 222, 237, 267, 243, 202, 143, 76, 44, 85, 156, 222, 266, 284, 282, 
    446, 409, 342, 270, 226, 261, 288, 238, 199, 178, 214, 263, 281, 250, 229, 206, 228, 199, 141, 82, 26, 24, 85, 170, 243, 275, 278, 269, 
    456, 419, 349, 277, 252, 288, 310, 232, 160, 157, 210, 286, 319, 281, 237, 179, 152, 108, 41, 4, 0, 12, 53, 134, 205, 238, 233, 211, 
    447, 417, 348, 291, 288, 351, 368, 302, 188, 156, 205, 269, 288, 243, 188, 139, 93, 40, 0, 0, 13, 24, 43, 81, 123, 147, 139, 119, 
    397, 402, 359, 344, 355, 437, 441, 340, 205, 150, 164, 185, 167, 116, 75, 45, 27, 22, 16, 15, 16, 18, 23, 38, 59, 69, 64, 52, 
    286, 349, 369, 407, 438, 500, 450, 290, 129, 50, 36, 34, 19, 0, 0, 0, 6, 13, 14, 16, 18, 21, 27, 34, 42, 43, 39, 30, 
    172, 253, 337, 425, 497, 510, 353, 128, 0, 0, 8, 11, 10, 6, 8, 14, 15, 16, 19, 21, 22, 26, 35, 42, 44, 39, 37, 35, 
    100, 158, 265, 411, 514, 452, 230, 25, 0, 17, 23, 19, 18, 19, 18, 16, 15, 16, 17, 21, 29, 36, 41, 39, 36, 37, 45, 55, 
    48, 85, 191, 352, 462, 353, 149, 16, 17, 34, 30, 21, 17, 19, 19, 17, 17, 17, 18, 23, 33, 38, 34, 26, 23, 37, 55, 61, 
    11, 44, 135, 264, 335, 242, 95, 28, 38, 41, 38, 30, 19, 17, 17, 17, 19, 18, 20, 25, 29, 31, 26, 18, 24, 41, 51, 37, 
    0, 17, 91, 163, 176, 120, 44, 7, 32, 42, 42, 37, 27, 23, 23, 25, 26, 23, 20, 22, 22, 25, 30, 40, 47, 42, 18, 0, 
    0, 5, 40, 86, 63, 20, 0, 0, 16, 35, 38, 32, 28, 30, 37, 45, 47, 41, 28, 19, 20, 33, 57, 82, 81, 48, 0, 0, 
    
    -- channel=21
    165, 177, 181, 181, 182, 185, 182, 184, 204, 229, 228, 210, 181, 170, 147, 107, 71, 49, 38, 32, 23, 20, 26, 51, 81, 107, 120, 117, 
    170, 183, 185, 183, 183, 185, 181, 182, 216, 262, 270, 216, 145, 106, 72, 40, 27, 37, 57, 73, 61, 32, 6, 1, 19, 53, 92, 113, 
    131, 153, 170, 179, 182, 183, 176, 157, 164, 203, 206, 152, 74, 22, 0, 0, 0, 44, 100, 120, 104, 77, 40, 9, 0, 0, 45, 95, 
    44, 77, 131, 172, 185, 184, 176, 140, 98, 98, 114, 96, 38, 0, 0, 0, 0, 59, 125, 140, 109, 75, 44, 12, 0, 0, 0, 65, 
    0, 16, 98, 169, 187, 186, 179, 153, 103, 78, 83, 94, 77, 25, 0, 0, 0, 51, 122, 135, 93, 45, 16, 0, 0, 0, 0, 21, 
    74, 72, 134, 183, 181, 191, 211, 212, 186, 150, 148, 162, 130, 56, 0, 0, 0, 0, 88, 130, 97, 29, 0, 0, 0, 0, 0, 0, 
    178, 185, 226, 217, 175, 197, 282, 349, 343, 272, 237, 214, 150, 57, 0, 0, 0, 0, 65, 150, 144, 66, 3, 0, 0, 0, 0, 0, 
    235, 259, 288, 242, 165, 165, 282, 424, 454, 379, 296, 259, 183, 83, 0, 0, 0, 0, 109, 207, 199, 114, 35, 0, 0, 0, 0, 0, 
    237, 287, 323, 270, 158, 83, 161, 318, 411, 385, 334, 297, 233, 130, 43, 0, 0, 54, 182, 268, 217, 114, 34, 0, 3, 6, 0, 0, 
    212, 282, 325, 283, 179, 58, 38, 146, 260, 305, 322, 340, 300, 194, 98, 55, 27, 93, 222, 270, 196, 78, 4, 0, 0, 8, 11, 12, 
    205, 263, 283, 241, 189, 103, 22, 55, 157, 237, 307, 375, 339, 248, 151, 93, 55, 105, 219, 248, 169, 54, 0, 0, 0, 9, 36, 49, 
    235, 261, 247, 179, 154, 121, 51, 56, 149, 253, 324, 369, 328, 250, 171, 102, 61, 105, 212, 235, 161, 64, 2, 0, 0, 30, 63, 69, 
    285, 290, 259, 163, 131, 128, 79, 62, 153, 283, 347, 325, 240, 182, 138, 80, 51, 94, 184, 207, 151, 69, 8, 0, 14, 50, 67, 73, 
    332, 329, 285, 195, 141, 147, 114, 76, 116, 221, 278, 230, 134, 79, 69, 62, 51, 73, 127, 155, 124, 53, 0, 0, 0, 26, 59, 84, 
    363, 358, 309, 226, 152, 162, 153, 83, 44, 76, 120, 104, 72, 33, 42, 56, 53, 45, 50, 72, 72, 20, 0, 0, 0, 21, 72, 107, 
    373, 366, 322, 240, 158, 162, 182, 129, 47, 1, 22, 48, 79, 77, 81, 76, 89, 69, 12, 0, 0, 0, 0, 0, 0, 54, 112, 143, 
    362, 357, 329, 250, 165, 141, 192, 182, 109, 26, 21, 86, 154, 176, 155, 102, 95, 92, 40, 0, 0, 0, 0, 0, 30, 98, 141, 150, 
    342, 348, 328, 261, 191, 174, 222, 240, 170, 88, 77, 157, 250, 295, 241, 133, 47, 9, 0, 0, 0, 0, 0, 0, 47, 100, 120, 116, 
    332, 345, 315, 265, 216, 254, 342, 392, 296, 201, 178, 225, 304, 341, 284, 176, 34, 0, 0, 0, 0, 0, 0, 0, 16, 44, 57, 46, 
    319, 348, 323, 290, 255, 342, 472, 504, 412, 289, 216, 215, 236, 247, 221, 150, 54, 0, 0, 0, 0, 0, 0, 5, 16, 24, 27, 19, 
    257, 326, 340, 323, 320, 395, 515, 505, 378, 208, 88, 51, 49, 45, 37, 29, 11, 0, 0, 0, 1, 15, 25, 26, 31, 33, 33, 28, 
    132, 222, 299, 322, 358, 420, 457, 376, 217, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 21, 34, 45, 50, 53, 54, 56, 
    27, 88, 177, 267, 346, 417, 398, 255, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 37, 53, 67, 69, 69, 76, 86, 
    13, 17, 75, 187, 316, 392, 321, 157, 31, 7, 17, 16, 4, 0, 0, 0, 0, 0, 8, 26, 44, 59, 69, 68, 64, 72, 90, 117, 
    36, 17, 35, 122, 262, 345, 265, 105, 16, 13, 23, 16, 4, 0, 0, 0, 5, 14, 26, 38, 50, 58, 57, 52, 53, 69, 104, 126, 
    54, 35, 32, 59, 150, 224, 179, 68, 7, 15, 25, 26, 18, 10, 6, 9, 19, 27, 32, 33, 35, 38, 43, 48, 58, 85, 105, 83, 
    64, 50, 31, 13, 17, 46, 39, 0, 0, 0, 14, 23, 25, 21, 17, 25, 36, 43, 41, 31, 23, 22, 35, 65, 102, 126, 111, 61, 
    63, 51, 40, 6, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 13, 30, 49, 59, 59, 41, 23, 21, 48, 97, 145, 159, 124, 57, 
    
    -- channel=22
    22, 28, 26, 13, 8, 9, 7, 0, 0, 0, 0, 1, 39, 71, 120, 154, 148, 105, 77, 79, 99, 125, 140, 128, 92, 50, 21, 7, 
    13, 22, 26, 24, 24, 28, 24, 0, 0, 0, 0, 57, 131, 203, 249, 222, 123, 9, 0, 0, 0, 16, 63, 96, 111, 88, 45, 12, 
    106, 87, 51, 30, 30, 36, 36, 49, 73, 125, 173, 186, 210, 256, 241, 163, 35, 0, 0, 0, 0, 0, 0, 25, 95, 109, 72, 26, 
    201, 141, 64, 29, 26, 29, 33, 88, 170, 258, 233, 161, 133, 135, 101, 40, 0, 0, 0, 0, 0, 0, 0, 26, 78, 98, 80, 44, 
    132, 67, 19, 14, 19, 11, 15, 61, 119, 152, 90, 23, 0, 0, 0, 0, 0, 0, 0, 31, 62, 73, 72, 68, 68, 77, 76, 60, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 74, 92, 62, 42, 57, 86, 94, 55, 31, 41, 63, 77, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 38, 86, 107, 80, 24, 0, 0, 18, 29, 1, 0, 0, 46, 87, 
    0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 58, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 53, 
    0, 0, 0, 0, 67, 146, 187, 184, 144, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 65, 22, 0, 0, 0, 0, 0, 
    1, 0, 40, 45, 88, 180, 312, 353, 315, 142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 145, 133, 83, 44, 3, 0, 0, 0, 
    5, 62, 157, 122, 86, 120, 221, 270, 243, 81, 0, 0, 0, 0, 0, 0, 0, 0, 26, 127, 146, 102, 70, 44, 6, 0, 0, 0, 
    0, 76, 165, 127, 70, 73, 98, 87, 28, 0, 0, 83, 99, 46, 2, 4, 0, 0, 71, 118, 106, 53, 25, 0, 0, 0, 0, 0, 
    0, 20, 67, 51, 4, 13, 15, 0, 0, 0, 73, 242, 256, 198, 113, 67, 22, 27, 102, 111, 90, 54, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 69, 202, 345, 395, 346, 269, 160, 65, 42, 115, 208, 178, 125, 108, 102, 82, 73, 69, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 58, 229, 433, 481, 372, 246, 156, 87, 23, 35, 162, 272, 258, 231, 218, 189, 146, 103, 49, 0, 0, 
    0, 0, 3, 6, 0, 0, 0, 24, 186, 343, 321, 191, 60, 0, 0, 0, 0, 80, 181, 285, 334, 275, 162, 67, 10, 0, 0, 0, 
    31, 12, 19, 24, 15, 0, 0, 0, 82, 139, 82, 0, 0, 0, 0, 0, 26, 91, 166, 283, 322, 228, 82, 0, 0, 0, 0, 0, 
    60, 37, 47, 46, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 19, 147, 263, 292, 264, 182, 102, 4, 0, 0, 0, 35, 83, 
    57, 50, 75, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 53, 152, 255, 260, 158, 44, 0, 0, 0, 0, 36, 93, 117, 
    77, 49, 46, 14, 0, 0, 0, 0, 0, 2, 76, 181, 303, 358, 306, 202, 117, 73, 46, 0, 0, 0, 0, 0, 0, 42, 71, 73, 
    197, 114, 22, 0, 0, 0, 0, 196, 326, 356, 375, 443, 522, 524, 435, 271, 105, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 8, 
    316, 248, 110, 0, 0, 0, 293, 547, 557, 418, 324, 335, 361, 343, 276, 178, 84, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    308, 333, 220, 60, 0, 146, 467, 593, 444, 228, 108, 75, 78, 75, 62, 39, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    174, 265, 225, 84, 40, 258, 475, 435, 223, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 17, 0, 0, 0, 
    55, 129, 166, 145, 187, 347, 405, 262, 92, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 25, 37, 18, 0, 0, 40, 
    3, 39, 124, 237, 385, 479, 411, 202, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 34, 30, 2, 0, 0, 42, 129, 
    0, 3, 82, 240, 437, 525, 410, 209, 84, 48, 32, 12, 0, 0, 0, 0, 0, 0, 0, 7, 27, 28, 0, 0, 0, 0, 43, 107, 
    4, 3, 32, 136, 270, 350, 283, 166, 93, 88, 94, 88, 73, 42, 10, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 26, 52, 
    
    -- channel=23
    158, 157, 157, 155, 152, 152, 150, 135, 122, 119, 141, 153, 157, 160, 163, 166, 159, 144, 129, 129, 138, 144, 152, 150, 150, 146, 143, 139, 
    151, 155, 157, 157, 157, 159, 157, 138, 101, 89, 122, 152, 158, 173, 187, 181, 138, 90, 56, 58, 69, 91, 110, 129, 136, 138, 141, 138, 
    159, 166, 168, 164, 163, 166, 165, 159, 137, 134, 161, 180, 185, 193, 192, 152, 89, 43, 21, 18, 19, 25, 44, 82, 109, 127, 133, 134, 
    178, 177, 167, 162, 162, 164, 164, 171, 186, 197, 187, 169, 158, 143, 119, 89, 46, 28, 28, 43, 36, 29, 30, 54, 91, 103, 120, 125, 
    147, 146, 151, 153, 158, 155, 154, 159, 170, 160, 124, 95, 81, 61, 48, 54, 33, 31, 38, 70, 68, 59, 57, 67, 74, 84, 100, 119, 
    56, 76, 119, 144, 146, 136, 127, 136, 132, 107, 68, 50, 60, 48, 35, 55, 63, 66, 56, 74, 81, 78, 75, 66, 64, 73, 85, 109, 
    0, 24, 89, 134, 128, 97, 54, 52, 74, 66, 58, 55, 73, 59, 53, 68, 79, 76, 63, 62, 67, 65, 55, 45, 43, 55, 82, 99, 
    0, 17, 81, 131, 133, 88, 32, 26, 66, 60, 64, 66, 64, 56, 51, 72, 55, 36, 31, 41, 50, 53, 34, 30, 29, 39, 62, 91, 
    2, 28, 90, 131, 153, 143, 121, 109, 132, 98, 67, 61, 60, 45, 43, 58, 23, 5, 16, 45, 66, 75, 46, 29, 29, 26, 42, 61, 
    17, 46, 102, 139, 160, 174, 177, 168, 179, 124, 64, 47, 62, 36, 24, 45, 9, 11, 28, 82, 96, 97, 65, 44, 38, 25, 26, 41, 
    12, 74, 128, 156, 160, 155, 152, 140, 148, 107, 54, 39, 70, 43, 15, 45, 6, 19, 52, 105, 101, 86, 67, 54, 44, 30, 24, 36, 
    2, 78, 133, 140, 148, 145, 127, 94, 73, 62, 65, 82, 90, 73, 46, 68, 24, 30, 60, 91, 78, 59, 44, 36, 27, 26, 35, 45, 
    0, 51, 96, 85, 112, 126, 104, 65, 26, 35, 86, 138, 135, 110, 84, 89, 55, 50, 69, 90, 74, 60, 41, 26, 29, 38, 61, 69, 
    0, 23, 63, 38, 52, 84, 92, 72, 57, 81, 132, 183, 157, 136, 110, 91, 68, 77, 89, 94, 89, 82, 64, 50, 63, 78, 91, 88, 
    4, 10, 50, 35, 9, 46, 77, 103, 130, 191, 214, 204, 143, 107, 84, 67, 84, 128, 136, 117, 105, 100, 96, 83, 87, 89, 90, 96, 
    19, 11, 42, 55, 10, 19, 52, 93, 136, 170, 158, 129, 80, 55, 58, 34, 59, 111, 136, 138, 149, 145, 111, 86, 78, 73, 84, 99, 
    40, 19, 31, 63, 25, 25, 39, 58, 98, 85, 76, 47, 19, 20, 60, 34, 45, 61, 91, 132, 140, 122, 69, 49, 59, 76, 94, 118, 
    61, 31, 31, 63, 28, 7, 43, 63, 73, 59, 41, 31, 11, 10, 55, 58, 93, 122, 124, 127, 102, 69, 41, 21, 39, 72, 102, 122, 
    65, 43, 47, 75, 19, 0, 0, 37, 31, 12, 0, 3, 5, 11, 44, 47, 89, 129, 126, 86, 42, 14, 4, 6, 26, 54, 85, 96, 
    62, 47, 53, 67, 8, 0, 0, 0, 15, 6, 13, 55, 91, 106, 108, 73, 48, 35, 21, 0, 0, 0, 0, 0, 0, 23, 40, 43, 
    75, 54, 34, 39, 0, 8, 21, 86, 119, 131, 138, 164, 192, 184, 158, 105, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    96, 80, 59, 44, 6, 23, 110, 190, 206, 163, 123, 128, 137, 125, 96, 58, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 92, 96, 57, 26, 59, 174, 202, 152, 75, 28, 15, 16, 15, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 73, 72, 43, 24, 94, 186, 150, 65, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 32, 48, 28, 47, 108, 160, 77, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 58, 84, 144, 146, 49, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 24, 80, 119, 165, 156, 62, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 28, 
    0, 0, 0, 44, 82, 106, 109, 54, 22, 16, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    272, 263, 258, 263, 269, 269, 267, 266, 268, 261, 256, 257, 261, 248, 225, 208, 201, 207, 210, 203, 204, 210, 217, 221, 232, 241, 245, 245, 
    264, 258, 257, 262, 268, 268, 267, 262, 259, 237, 215, 213, 216, 202, 180, 171, 182, 188, 178, 161, 157, 167, 183, 204, 220, 237, 246, 250, 
    237, 244, 258, 269, 271, 272, 272, 267, 259, 223, 199, 191, 198, 184, 166, 165, 187, 181, 167, 145, 143, 145, 159, 171, 195, 222, 243, 247, 
    223, 255, 277, 277, 271, 270, 271, 272, 259, 223, 202, 196, 176, 157, 154, 170, 185, 182, 160, 133, 127, 134, 142, 136, 153, 199, 235, 244, 
    198, 262, 294, 288, 275, 273, 270, 255, 227, 207, 207, 186, 149, 148, 165, 170, 178, 177, 162, 132, 127, 145, 136, 117, 124, 173, 219, 241, 
    160, 235, 272, 280, 278, 275, 267, 241, 208, 204, 200, 177, 144, 138, 151, 150, 168, 182, 175, 145, 138, 149, 148, 131, 126, 148, 197, 228, 
    141, 207, 241, 260, 263, 260, 240, 185, 153, 163, 170, 156, 131, 130, 145, 146, 162, 189, 191, 166, 135, 131, 148, 149, 136, 133, 165, 212, 
    141, 199, 233, 248, 246, 225, 197, 145, 114, 129, 142, 129, 119, 124, 132, 132, 158, 192, 185, 158, 126, 118, 144, 159, 146, 131, 136, 184, 
    143, 194, 219, 239, 236, 217, 179, 128, 76, 103, 124, 124, 116, 126, 132, 120, 164, 190, 171, 134, 110, 103, 137, 161, 152, 132, 123, 149, 
    141, 182, 200, 222, 225, 199, 165, 133, 114, 127, 158, 139, 112, 125, 137, 116, 160, 190, 161, 112, 84, 99, 132, 162, 157, 142, 129, 141, 
    134, 159, 179, 220, 227, 185, 159, 146, 143, 160, 161, 137, 104, 120, 140, 116, 164, 184, 153, 97, 88, 111, 141, 168, 173, 162, 142, 152, 
    128, 120, 137, 215, 242, 214, 192, 176, 189, 184, 161, 124, 103, 113, 127, 116, 167, 178, 141, 96, 86, 104, 129, 157, 176, 175, 165, 177, 
    122, 94, 92, 188, 239, 227, 203, 197, 201, 168, 119, 75, 101, 118, 125, 129, 171, 184, 148, 117, 106, 115, 132, 156, 172, 176, 182, 195, 
    109, 96, 66, 138, 220, 227, 210, 200, 184, 140, 69, 46, 88, 127, 140, 164, 185, 169, 137, 114, 98, 96, 116, 149, 170, 185, 200, 229, 
    96, 103, 59, 91, 181, 222, 207, 202, 181, 133, 98, 101, 129, 146, 160, 195, 213, 190, 159, 134, 96, 78, 104, 149, 184, 201, 226, 245, 
    86, 104, 67, 55, 136, 186, 181, 182, 148, 124, 128, 143, 161, 150, 146, 199, 213, 177, 161, 146, 111, 83, 116, 168, 204, 227, 245, 248, 
    89, 101, 79, 46, 105, 163, 165, 146, 114, 135, 169, 188, 183, 149, 116, 166, 174, 147, 125, 96, 77, 83, 131, 180, 219, 241, 245, 240, 
    104, 105, 87, 46, 82, 136, 146, 115, 112, 155, 177, 178, 162, 126, 86, 122, 157, 150, 107, 74, 85, 105, 139, 181, 214, 221, 218, 215, 
    122, 116, 95, 57, 92, 145, 124, 63, 55, 94, 127, 141, 121, 80, 38, 51, 98, 104, 89, 81, 81, 87, 98, 138, 171, 187, 179, 177, 
    112, 114, 101, 72, 105, 143, 115, 35, 0, 17, 55, 52, 27, 0, 0, 0, 28, 46, 51, 60, 54, 53, 46, 63, 85, 99, 98, 93, 
    75, 81, 87, 83, 127, 141, 87, 0, 0, 0, 17, 27, 9, 0, 0, 0, 16, 37, 37, 34, 32, 21, 13, 11, 15, 26, 28, 22, 
    56, 72, 77, 103, 154, 129, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 17, 12, 8, 3, 0, 0, 0, 0, 0, 0, 
    27, 63, 79, 128, 160, 108, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 8, 10, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 34, 69, 137, 148, 61, 0, 0, 0, 0, 0, 0, 2, 7, 10, 9, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 52, 114, 112, 0, 0, 0, 0, 1, 0, 0, 0, 4, 6, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 73, 64, 0, 0, 0, 0, 4, 2, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 38, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 15, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 
    
    -- channel=25
    546, 559, 557, 548, 542, 540, 536, 527, 515, 509, 518, 532, 542, 539, 518, 474, 413, 358, 319, 306, 308, 320, 340, 359, 386, 420, 453, 462, 
    529, 553, 561, 556, 550, 548, 542, 515, 486, 478, 478, 485, 480, 467, 437, 380, 317, 258, 220, 204, 215, 244, 273, 300, 326, 362, 402, 432, 
    463, 494, 532, 554, 561, 561, 557, 532, 497, 446, 415, 410, 399, 378, 348, 303, 245, 184, 135, 110, 106, 124, 160, 201, 245, 290, 344, 396, 
    376, 406, 470, 536, 567, 571, 566, 557, 524, 464, 410, 374, 351, 322, 280, 226, 173, 137, 118, 104, 84, 81, 93, 118, 165, 222, 291, 355, 
    322, 355, 426, 505, 552, 560, 548, 541, 513, 455, 381, 317, 262, 208, 158, 129, 114, 115, 124, 130, 117, 103, 84, 81, 109, 165, 239, 317, 
    231, 284, 380, 476, 528, 531, 511, 493, 453, 383, 310, 238, 180, 131, 94, 93, 102, 116, 131, 146, 158, 144, 113, 85, 89, 132, 196, 272, 
    146, 204, 317, 431, 484, 463, 439, 430, 405, 347, 274, 215, 171, 125, 92, 95, 113, 140, 155, 164, 172, 165, 136, 98, 80, 109, 167, 233, 
    107, 166, 284, 400, 445, 398, 354, 332, 331, 300, 259, 217, 182, 143, 112, 110, 119, 146, 176, 179, 166, 139, 114, 88, 70, 85, 137, 201, 
    77, 137, 266, 390, 458, 417, 324, 275, 280, 276, 255, 229, 196, 151, 118, 110, 111, 139, 163, 174, 158, 122, 99, 77, 64, 64, 102, 167, 
    62, 124, 247, 372, 474, 472, 386, 319, 279, 260, 237, 225, 209, 170, 124, 108, 109, 134, 154, 173, 152, 122, 99, 78, 60, 51, 73, 129, 
    78, 137, 235, 344, 446, 478, 418, 339, 294, 264, 239, 218, 200, 174, 131, 104, 105, 123, 149, 168, 148, 126, 105, 87, 68, 60, 72, 114, 
    91, 137, 221, 311, 392, 437, 392, 298, 249, 244, 239, 203, 170, 157, 136, 116, 110, 127, 146, 154, 133, 109, 95, 89, 85, 83, 93, 125, 
    96, 113, 174, 241, 316, 369, 355, 269, 214, 222, 240, 231, 190, 154, 133, 130, 138, 154, 159, 147, 119, 86, 62, 63, 78, 100, 129, 168, 
    100, 92, 115, 155, 214, 272, 289, 240, 210, 196, 200, 203, 192, 173, 148, 146, 168, 191, 181, 158, 132, 109, 84, 75, 95, 130, 177, 231, 
    101, 81, 81, 96, 122, 177, 227, 246, 242, 223, 214, 207, 189, 177, 152, 155, 201, 232, 208, 163, 126, 106, 100, 99, 132, 184, 244, 315, 
    94, 72, 62, 75, 79, 116, 166, 232, 262, 262, 255, 225, 196, 170, 138, 134, 184, 252, 267, 217, 151, 119, 122, 145, 186, 241, 306, 373, 
    91, 70, 56, 68, 74, 82, 110, 166, 204, 213, 197, 164, 158, 146, 134, 122, 141, 182, 212, 191, 160, 124, 117, 146, 201, 280, 354, 404, 
    99, 82, 64, 63, 69, 88, 127, 150, 161, 160, 148, 154, 160, 147, 146, 143, 144, 139, 121, 103, 88, 67, 56, 74, 144, 235, 306, 336, 
    106, 104, 86, 67, 59, 86, 139, 174, 184, 164, 135, 132, 123, 106, 99, 105, 138, 147, 108, 56, 28, 20, 11, 23, 71, 123, 166, 182, 
    84, 103, 101, 91, 92, 119, 135, 146, 131, 108, 95, 112, 112, 91, 58, 34, 35, 44, 35, 0, 0, 0, 0, 0, 0, 33, 54, 58, 
    49, 66, 77, 95, 117, 138, 144, 137, 106, 84, 87, 105, 119, 105, 63, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 46, 44, 67, 110, 152, 170, 131, 77, 67, 89, 122, 137, 118, 72, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    87, 75, 45, 52, 97, 160, 175, 124, 77, 31, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 64, 50, 42, 80, 137, 129, 61, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 35, 39, 63, 90, 63, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 59, 77, 53, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 69, 105, 72, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 71, 62, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 32, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 51, 47, 27, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 26, 2, 8, 35, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 17, 0, 0, 29, 42, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 29, 6, 0, 0, 0, 0, 0, 24, 13, 0, 11, 45, 23, 0, 0, 
    62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 47, 46, 30, 8, 0, 0, 0, 7, 54, 42, 1, 0, 32, 52, 0, 0, 
    78, 0, 0, 0, 0, 0, 0, 0, 10, 16, 0, 37, 63, 46, 44, 30, 0, 0, 0, 39, 79, 53, 5, 0, 16, 60, 40, 0, 
    71, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 71, 52, 53, 33, 0, 0, 0, 69, 100, 56, 2, 0, 0, 37, 48, 0, 
    87, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 80, 64, 58, 26, 0, 0, 17, 91, 114, 69, 12, 0, 0, 5, 33, 8, 
    111, 85, 24, 0, 0, 0, 0, 0, 0, 0, 0, 32, 57, 57, 60, 21, 0, 0, 22, 92, 120, 84, 28, 0, 0, 0, 1, 0, 
    122, 143, 115, 0, 0, 0, 0, 0, 0, 0, 34, 59, 40, 19, 19, 0, 0, 0, 0, 72, 104, 67, 22, 0, 0, 0, 0, 0, 
    127, 173, 189, 66, 0, 0, 0, 0, 0, 0, 11, 42, 19, 0, 0, 0, 0, 0, 0, 23, 77, 73, 18, 0, 0, 0, 0, 0, 
    144, 180, 229, 153, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 46, 0, 0, 0, 0, 0, 0, 
    166, 182, 250, 208, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 
    163, 173, 238, 233, 124, 7, 6, 17, 0, 0, 0, 0, 0, 49, 59, 0, 0, 0, 0, 0, 6, 17, 0, 0, 0, 0, 0, 0, 
    130, 149, 208, 231, 148, 43, 58, 102, 56, 0, 0, 0, 0, 106, 134, 69, 0, 0, 0, 14, 49, 36, 0, 0, 0, 0, 0, 0, 
    104, 130, 182, 203, 122, 40, 113, 187, 172, 75, 0, 0, 37, 138, 205, 167, 76, 30, 47, 89, 112, 112, 84, 31, 0, 0, 0, 0, 
    101, 140, 177, 168, 85, 19, 142, 257, 285, 185, 72, 33, 61, 136, 201, 213, 170, 143, 159, 174, 187, 199, 201, 176, 131, 108, 114, 121, 
    89, 135, 170, 140, 72, 33, 158, 305, 348, 254, 155, 102, 115, 168, 223, 253, 253, 238, 242, 250, 265, 283, 303, 306, 291, 282, 290, 303, 
    98, 109, 135, 97, 52, 73, 218, 336, 371, 327, 251, 216, 219, 240, 270, 293, 298, 294, 302, 316, 327, 334, 345, 360, 366, 366, 372, 377, 
    167, 117, 89, 64, 48, 143, 286, 383, 393, 350, 314, 300, 296, 298, 307, 315, 320, 322, 332, 343, 354, 360, 368, 379, 384, 388, 387, 387, 
    281, 171, 84, 42, 68, 228, 374, 435, 393, 346, 339, 337, 329, 321, 320, 324, 330, 337, 348, 361, 370, 381, 390, 394, 394, 390, 391, 408, 
    386, 271, 137, 41, 79, 281, 427, 444, 365, 334, 345, 350, 340, 329, 326, 329, 336, 349, 366, 377, 385, 398, 412, 414, 399, 396, 415, 426, 
    442, 365, 223, 86, 78, 268, 412, 407, 335, 326, 340, 351, 351, 339, 332, 335, 347, 365, 382, 393, 399, 403, 409, 407, 408, 430, 457, 448, 
    459, 416, 325, 185, 140, 239, 355, 369, 309, 309, 321, 339, 349, 342, 334, 338, 353, 372, 394, 406, 401, 387, 376, 382, 418, 470, 506, 485, 
    462, 428, 387, 303, 249, 270, 332, 346, 308, 300, 303, 314, 323, 321, 318, 321, 341, 373, 402, 407, 389, 359, 334, 351, 419, 499, 531, 495, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    48, 48, 49, 50, 55, 57, 55, 46, 44, 53, 60, 55, 58, 64, 71, 69, 56, 42, 40, 44, 46, 46, 48, 55, 60, 62, 59, 53, 
    64, 64, 58, 53, 55, 57, 55, 49, 61, 88, 99, 83, 79, 80, 70, 43, 28, 37, 57, 58, 57, 50, 48, 54, 64, 68, 67, 62, 
    85, 86, 75, 57, 51, 52, 51, 47, 51, 71, 90, 71, 50, 32, 18, 16, 26, 47, 54, 55, 57, 56, 53, 48, 57, 62, 66, 66, 
    60, 62, 69, 64, 56, 54, 53, 51, 37, 44, 44, 31, 22, 19, 27, 38, 40, 46, 55, 50, 48, 53, 53, 49, 42, 50, 59, 68, 
    35, 52, 71, 70, 58, 51, 50, 48, 34, 28, 40, 59, 51, 42, 47, 47, 44, 46, 62, 61, 48, 39, 43, 39, 30, 32, 49, 64, 
    53, 74, 92, 78, 56, 44, 45, 44, 38, 38, 59, 63, 57, 46, 41, 47, 39, 39, 48, 61, 46, 30, 25, 21, 28, 25, 35, 51, 
    70, 86, 99, 82, 60, 50, 72, 97, 80, 63, 58, 60, 54, 39, 28, 35, 24, 15, 32, 60, 50, 36, 27, 31, 31, 31, 25, 38, 
    69, 97, 115, 85, 52, 46, 71, 113, 110, 76, 58, 52, 48, 36, 28, 20, 23, 20, 52, 68, 64, 52, 42, 38, 36, 34, 24, 25, 
    59, 106, 127, 94, 54, 18, 15, 71, 107, 74, 55, 61, 50, 40, 31, 20, 29, 33, 66, 73, 66, 60, 41, 40, 41, 35, 34, 25, 
    46, 106, 134, 111, 70, 11, 0, 18, 68, 52, 46, 71, 61, 46, 38, 38, 33, 31, 73, 74, 59, 51, 35, 39, 40, 37, 37, 41, 
    43, 88, 118, 103, 74, 31, 0, 1, 57, 56, 61, 82, 92, 66, 46, 50, 36, 32, 72, 67, 47, 41, 28, 28, 31, 35, 43, 52, 
    42, 71, 91, 90, 75, 52, 6, 0, 46, 61, 73, 71, 91, 79, 58, 58, 30, 35, 60, 72, 57, 51, 43, 37, 43, 46, 55, 61, 
    45, 68, 76, 80, 83, 74, 35, 19, 55, 82, 88, 84, 80, 66, 56, 59, 28, 32, 53, 67, 55, 41, 36, 44, 53, 60, 70, 66, 
    49, 68, 85, 68, 77, 98, 64, 35, 40, 83, 97, 79, 60, 51, 48, 59, 43, 44, 55, 70, 63, 49, 38, 39, 51, 62, 62, 51, 
    53, 66, 87, 59, 68, 90, 82, 53, 26, 34, 42, 38, 26, 29, 40, 64, 57, 39, 30, 40, 57, 55, 40, 27, 31, 40, 50, 54, 
    56, 61, 82, 62, 53, 76, 97, 65, 24, 16, 20, 54, 49, 47, 51, 62, 63, 54, 35, 29, 38, 25, 9, 10, 26, 46, 57, 56, 
    60, 55, 72, 69, 40, 49, 81, 72, 51, 48, 38, 65, 61, 61, 54, 54, 72, 86, 68, 49, 36, 10, 23, 46, 62, 68, 69, 66, 
    68, 58, 66, 71, 46, 44, 74, 67, 45, 26, 35, 57, 60, 68, 70, 44, 54, 47, 39, 18, 0, 11, 19, 48, 74, 83, 87, 82, 
    81, 65, 58, 60, 49, 50, 84, 73, 69, 50, 56, 72, 83, 91, 101, 68, 47, 23, 0, 0, 15, 30, 27, 38, 53, 73, 73, 68, 
    101, 80, 59, 66, 52, 49, 87, 100, 83, 78, 77, 79, 86, 76, 71, 62, 37, 25, 23, 29, 26, 20, 21, 21, 29, 43, 48, 48, 
    86, 88, 82, 95, 66, 61, 93, 105, 88, 50, 20, 1, 0, 0, 0, 0, 7, 9, 11, 9, 3, 0, 3, 7, 10, 13, 20, 21, 
    41, 60, 77, 96, 65, 83, 81, 58, 26, 0, 0, 0, 0, 0, 0, 3, 4, 2, 0, 0, 0, 0, 0, 2, 5, 4, 5, 4, 
    19, 32, 55, 79, 71, 91, 49, 21, 0, 1, 8, 5, 4, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 6, 
    10, 13, 45, 61, 88, 73, 44, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 
    1, 6, 26, 46, 73, 70, 51, 14, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 1, 17, 19, 37, 47, 49, 13, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 5, 0, 0, 8, 17, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 1, 8, 9, 5, 0, 0, 
    
    -- channel=29
    133, 123, 122, 126, 131, 135, 136, 129, 120, 114, 121, 125, 123, 121, 122, 125, 128, 131, 133, 133, 131, 128, 127, 131, 139, 143, 145, 150, 
    131, 124, 124, 127, 131, 134, 135, 124, 103, 90, 110, 118, 119, 117, 121, 128, 131, 123, 120, 127, 130, 129, 128, 129, 136, 141, 145, 151, 
    131, 132, 133, 133, 131, 134, 135, 121, 101, 100, 128, 127, 129, 136, 138, 131, 121, 109, 119, 131, 144, 142, 140, 143, 142, 143, 146, 147, 
    136, 142, 148, 144, 134, 131, 134, 136, 126, 111, 129, 148, 147, 139, 137, 139, 125, 114, 116, 140, 154, 150, 160, 172, 164, 141, 139, 141, 
    139, 136, 149, 148, 135, 127, 129, 138, 128, 117, 130, 147, 150, 147, 154, 160, 130, 114, 117, 143, 152, 161, 174, 194, 192, 164, 139, 136, 
    136, 120, 135, 145, 132, 117, 107, 110, 112, 106, 97, 120, 155, 163, 167, 173, 146, 121, 121, 140, 153, 159, 176, 199, 206, 186, 149, 135, 
    116, 98, 127, 145, 126, 96, 64, 55, 64, 61, 68, 102, 149, 167, 175, 188, 167, 124, 107, 133, 153, 152, 165, 186, 206, 198, 162, 133, 
    89, 83, 123, 147, 124, 66, 6, 0, 33, 40, 49, 91, 133, 162, 176, 190, 164, 109, 75, 106, 138, 158, 154, 171, 191, 199, 182, 141, 
    71, 69, 117, 151, 130, 78, 21, 3, 25, 28, 33, 76, 126, 151, 176, 179, 142, 83, 58, 89, 131, 166, 158, 163, 183, 195, 191, 157, 
    67, 66, 107, 147, 157, 120, 50, 19, 45, 45, 42, 68, 119, 133, 162, 171, 121, 58, 52, 99, 139, 173, 164, 164, 179, 187, 187, 176, 
    54, 61, 104, 137, 168, 143, 90, 49, 72, 54, 32, 53, 106, 121, 146, 168, 116, 57, 59, 113, 149, 179, 176, 170, 173, 181, 182, 180, 
    52, 69, 108, 124, 153, 157, 133, 76, 68, 44, 22, 56, 107, 116, 134, 160, 119, 62, 70, 123, 159, 179, 175, 160, 153, 162, 178, 183, 
    42, 75, 122, 114, 130, 164, 153, 92, 55, 31, 27, 50, 95, 126, 142, 164, 132, 80, 80, 126, 161, 184, 179, 155, 145, 153, 176, 177, 
    22, 70, 135, 119, 103, 144, 156, 114, 62, 46, 69, 103, 113, 135, 148, 169, 149, 105, 105, 131, 162, 180, 176, 155, 148, 153, 165, 170, 
    8, 55, 130, 133, 84, 122, 150, 136, 94, 86, 102, 144, 145, 139, 154, 162, 153, 125, 129, 148, 179, 192, 184, 169, 165, 162, 162, 157, 
    16, 44, 123, 144, 85, 92, 124, 148, 126, 109, 120, 147, 145, 133, 148, 145, 152, 137, 121, 149, 194, 202, 185, 166, 163, 151, 146, 141, 
    40, 46, 112, 149, 101, 71, 110, 142, 135, 110, 115, 118, 108, 119, 148, 132, 135, 139, 143, 162, 184, 198, 175, 152, 147, 137, 137, 138, 
    63, 53, 100, 150, 115, 50, 75, 123, 138, 129, 95, 74, 56, 89, 140, 124, 119, 161, 181, 182, 185, 184, 162, 132, 120, 120, 127, 132, 
    69, 53, 89, 143, 106, 43, 45, 99, 111, 95, 49, 27, 19, 60, 120, 135, 130, 157, 183, 200, 190, 169, 145, 123, 108, 111, 123, 133, 
    55, 47, 80, 129, 72, 2, 2, 56, 95, 85, 54, 34, 27, 59, 116, 148, 161, 165, 176, 187, 184, 167, 147, 136, 117, 118, 128, 141, 
    50, 45, 69, 95, 39, 0, 0, 51, 117, 112, 93, 78, 74, 94, 136, 165, 175, 186, 182, 178, 173, 165, 155, 147, 141, 143, 156, 164, 
    60, 53, 67, 66, 19, 0, 0, 101, 156, 148, 123, 115, 116, 127, 152, 172, 186, 192, 185, 176, 168, 161, 157, 156, 157, 157, 160, 162, 
    78, 71, 71, 50, 0, 0, 67, 129, 159, 172, 166, 158, 159, 165, 177, 190, 190, 187, 182, 176, 170, 162, 158, 158, 158, 154, 152, 149, 
    116, 89, 67, 36, 0, 31, 121, 170, 180, 186, 175, 173, 175, 177, 183, 186, 186, 184, 178, 172, 165, 160, 159, 160, 157, 150, 141, 137, 
    160, 111, 78, 34, 9, 64, 163, 190, 189, 176, 171, 175, 176, 178, 179, 179, 178, 174, 172, 168, 165, 163, 161, 159, 154, 144, 142, 149, 
    174, 148, 105, 48, 30, 103, 199, 206, 192, 172, 171, 174, 175, 176, 174, 171, 167, 167, 168, 169, 167, 167, 167, 161, 149, 144, 151, 160, 
    175, 164, 138, 80, 51, 134, 222, 213, 199, 183, 180, 181, 177, 173, 166, 162, 160, 162, 167, 173, 175, 173, 167, 154, 142, 145, 157, 163, 
    172, 168, 164, 130, 96, 144, 219, 216, 201, 193, 190, 191, 191, 182, 170, 161, 155, 156, 167, 178, 181, 172, 153, 136, 132, 146, 168, 182, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    73, 14, 0, 0, 0, 0, 0, 0, 27, 20, 13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    87, 19, 0, 0, 0, 0, 0, 0, 0, 0, 2, 20, 0, 0, 0, 0, 0, 0, 7, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    98, 37, 0, 0, 0, 0, 0, 0, 0, 0, 5, 27, 18, 0, 0, 0, 0, 0, 14, 28, 0, 0, 0, 0, 0, 0, 0, 0, 
    111, 63, 0, 0, 0, 0, 0, 0, 0, 0, 33, 40, 19, 0, 0, 0, 0, 0, 8, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    122, 90, 24, 0, 0, 0, 0, 0, 0, 20, 55, 54, 12, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    137, 111, 81, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    162, 136, 127, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    183, 159, 147, 86, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    174, 163, 145, 112, 53, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    141, 149, 132, 111, 67, 53, 44, 27, 0, 0, 0, 0, 1, 34, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    122, 138, 123, 101, 85, 79, 105, 97, 63, 1, 0, 17, 65, 77, 74, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    119, 142, 126, 107, 103, 108, 149, 168, 141, 99, 60, 63, 73, 71, 65, 36, 0, 0, 0, 0, 0, 21, 44, 43, 35, 17, 4, 0, 
    102, 120, 122, 121, 129, 153, 190, 220, 188, 125, 78, 62, 56, 57, 59, 50, 35, 26, 37, 51, 66, 83, 99, 111, 110, 102, 99, 98, 
    103, 101, 99, 123, 148, 189, 219, 216, 155, 99, 70, 59, 59, 59, 64, 70, 69, 71, 79, 93, 104, 116, 128, 140, 144, 145, 144, 147, 
    117, 92, 84, 109, 164, 205, 212, 168, 120, 98, 89, 83, 79, 76, 77, 80, 81, 87, 97, 111, 124, 136, 145, 153, 155, 158, 164, 174, 
    142, 97, 79, 102, 177, 207, 200, 155, 123, 112, 109, 105, 99, 90, 85, 87, 92, 101, 112, 127, 141, 153, 160, 160, 159, 166, 184, 196, 
    160, 125, 94, 114, 156, 183, 171, 149, 118, 111, 117, 113, 106, 96, 92, 95, 103, 115, 128, 141, 153, 160, 164, 165, 169, 179, 195, 196, 
    176, 150, 129, 109, 116, 125, 125, 122, 94, 102, 113, 118, 114, 105, 103, 110, 120, 129, 141, 149, 154, 155, 157, 166, 182, 200, 212, 201, 
    184, 165, 151, 123, 93, 84, 80, 84, 74, 83, 95, 104, 108, 109, 112, 118, 131, 142, 149, 150, 147, 142, 148, 170, 201, 226, 225, 201, 
    183, 168, 154, 134, 95, 74, 68, 68, 67, 71, 77, 84, 83, 86, 96, 111, 133, 149, 154, 150, 138, 132, 143, 175, 215, 234, 223, 192, 
    
    
    others => 0);
end ifmap_package;
