library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    126, 150, 122, 103, 56, 70, 114, 
    158, 134, 108, 77, 57, 74, 95, 
    77, 97, 0, 73, 76, 63, 61, 
    0, 94, 19, 45, 86, 63, 70, 
    0, 66, 47, 0, 28, 27, 40, 
    0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    106, 134, 136, 112, 115, 103, 92, 
    192, 174, 186, 132, 111, 134, 117, 
    153, 180, 115, 177, 162, 149, 108, 
    135, 180, 88, 138, 150, 119, 93, 
    96, 217, 167, 88, 87, 82, 46, 
    0, 179, 86, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 14, 0, 132, 0, 88, 62, 
    32, 0, 0, 123, 0, 112, 62, 
    102, 0, 0, 139, 0, 173, 23, 
    95, 37, 0, 111, 0, 140, 0, 
    0, 0, 0, 0, 118, 42, 0, 
    0, 0, 215, 79, 69, 0, 0, 
    0, 52, 61, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    73, 69, 87, 85, 69, 59, 86, 
    144, 100, 74, 64, 129, 72, 89, 
    160, 174, 105, 110, 221, 94, 39, 
    118, 142, 141, 91, 192, 87, 61, 
    132, 226, 105, 66, 72, 0, 48, 
    39, 209, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 76, 29, 0, 
    83, 0, 50, 18, 117, 54, 0, 
    144, 18, 112, 78, 101, 33, 20, 
    236, 105, 47, 80, 51, 12, 32, 
    269, 239, 155, 240, 190, 248, 286, 
    337, 306, 272, 289, 323, 358, 384, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    41, 77, 18, 7, 29, 35, 27, 
    0, 48, 2, 16, 45, 40, 0, 
    105, 0, 70, 31, 0, 46, 3, 
    152, 14, 42, 92, 34, 21, 53, 
    182, 71, 22, 91, 40, 11, 67, 
    180, 48, 81, 173, 165, 198, 240, 
    225, 169, 192, 220, 235, 259, 249, 
    
    -- channel=10
    18, 0, 0, 30, 5, 11, 23, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 66, 49, 0, 0, 0, 0, 
    13, 0, 59, 19, 6, 2, 0, 
    11, 0, 0, 0, 33, 28, 23, 
    116, 27, 86, 103, 10, 12, 32, 
    122, 130, 75, 46, 44, 66, 65, 
    
    -- channel=11
    123, 132, 116, 72, 64, 68, 103, 
    99, 128, 96, 65, 74, 73, 81, 
    85, 121, 114, 86, 70, 84, 61, 
    27, 98, 64, 56, 75, 66, 87, 
    5, 38, 68, 48, 28, 0, 58, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    152, 153, 129, 111, 105, 107, 155, 
    144, 122, 54, 110, 112, 115, 118, 
    204, 141, 133, 127, 142, 171, 80, 
    179, 186, 139, 153, 121, 144, 126, 
    144, 180, 88, 103, 112, 22, 86, 
    149, 62, 94, 54, 36, 0, 26, 
    47, 83, 20, 9, 0, 0, 0, 
    
    -- channel=13
    71, 30, 53, 123, 58, 47, 76, 
    80, 39, 60, 0, 18, 21, 72, 
    5, 117, 20, 0, 12, 15, 0, 
    0, 16, 73, 54, 70, 53, 0, 
    0, 0, 38, 0, 83, 89, 32, 
    59, 41, 138, 99, 0, 0, 0, 
    71, 168, 48, 0, 0, 0, 16, 
    
    -- channel=14
    48, 100, 15, 0, 18, 0, 0, 
    0, 82, 47, 0, 23, 0, 0, 
    0, 0, 38, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 40, 
    16, 0, 0, 21, 0, 0, 21, 
    8, 0, 0, 44, 73, 189, 181, 
    143, 0, 75, 173, 217, 228, 234, 
    
    -- channel=15
    0, 0, 20, 21, 8, 69, 0, 
    50, 0, 37, 123, 0, 139, 81, 
    184, 0, 72, 284, 3, 207, 128, 
    253, 131, 0, 145, 0, 163, 0, 
    229, 217, 63, 135, 72, 65, 0, 
    8, 144, 188, 13, 77, 0, 0, 
    0, 42, 55, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    35, 0, 12, 120, 62, 36, 58, 
    8, 52, 37, 0, 0, 0, 16, 
    0, 14, 43, 0, 0, 0, 0, 
    0, 0, 52, 14, 0, 1, 0, 
    0, 0, 19, 0, 108, 71, 41, 
    72, 0, 158, 94, 0, 0, 0, 
    9, 144, 0, 0, 0, 1, 0, 
    
    -- channel=20
    258, 292, 250, 151, 122, 133, 175, 
    98, 230, 175, 78, 101, 84, 92, 
    44, 131, 129, 85, 47, 42, 89, 
    53, 117, 143, 61, 85, 57, 157, 
    61, 0, 20, 104, 38, 0, 122, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    132, 106, 134, 93, 96, 51, 89, 
    111, 125, 102, 15, 96, 21, 49, 
    100, 206, 221, 23, 137, 36, 56, 
    52, 90, 104, 49, 85, 37, 65, 
    60, 100, 67, 55, 43, 57, 72, 
    127, 208, 134, 25, 0, 25, 0, 
    30, 39, 0, 0, 0, 1, 9, 
    
    -- channel=22
    97, 144, 53, 62, 51, 46, 69, 
    0, 70, 33, 27, 15, 27, 0, 
    3, 0, 0, 0, 0, 3, 0, 
    82, 18, 74, 82, 51, 5, 41, 
    106, 0, 0, 16, 11, 2, 28, 
    64, 0, 0, 117, 56, 12, 92, 
    94, 110, 121, 98, 103, 92, 81, 
    
    -- channel=23
    10, 0, 15, 4, 0, 18, 0, 
    26, 0, 38, 30, 0, 9, 0, 
    55, 10, 49, 32, 0, 14, 35, 
    84, 19, 0, 0, 0, 28, 0, 
    53, 40, 89, 60, 38, 67, 20, 
    122, 104, 237, 148, 173, 228, 211, 
    216, 165, 216, 216, 232, 258, 275, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    274, 275, 224, 175, 202, 129, 212, 
    250, 308, 193, 0, 89, 0, 51, 
    0, 147, 0, 0, 186, 0, 0, 
    0, 75, 33, 0, 36, 0, 23, 
    0, 65, 69, 25, 0, 29, 173, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    85, 1, 23, 25, 0, 0, 0, 
    0, 0, 0, 7, 0, 5, 0, 
    0, 8, 0, 0, 0, 0, 0, 
    0, 32, 136, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 34, 0, 56, 0, 
    80, 0, 0, 109, 0, 116, 141, 
    163, 3, 0, 196, 0, 216, 58, 
    164, 128, 0, 97, 0, 168, 0, 
    63, 104, 130, 16, 88, 45, 0, 
    0, 0, 225, 0, 70, 0, 4, 
    104, 0, 78, 23, 2, 10, 33, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    196, 209, 160, 160, 85, 56, 132, 
    45, 114, 51, 28, 4, 0, 38, 
    0, 113, 35, 0, 3, 0, 0, 
    0, 38, 15, 11, 22, 4, 25, 
    0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    48, 46, 49, 52, 26, 17, 41, 
    60, 28, 11, 17, 0, 0, 75, 
    0, 0, 0, 0, 23, 0, 28, 
    0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    6, 14, 16, 14, 15, 17, 1, 
    0, 0, 0, 22, 7, 49, 22, 
    41, 12, 29, 14, 0, 61, 39, 
    70, 0, 14, 35, 18, 66, 34, 
    112, 0, 53, 62, 95, 106, 91, 
    245, 121, 331, 332, 328, 418, 423, 
    474, 369, 382, 429, 468, 516, 541, 
    
    
    others => 0);
end ifmap_package;
