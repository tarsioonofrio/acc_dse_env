library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 13, 0, 62, 0, 0, 
    13, 29, 27, 0, 152, 0, 0, 
    0, 0, 48, 0, 244, 0, 0, 
    0, 0, 182, 0, 101, 0, 33, 
    53, 103, 0, 76, 0, 0, 78, 
    0, 271, 0, 0, 0, 48, 13, 
    0, 0, 0, 0, 22, 0, 26, 
    
    -- channel=1
    30, 57, 43, 42, 54, 58, 46, 
    105, 106, 89, 75, 77, 82, 78, 
    69, 147, 42, 89, 127, 112, 53, 
    61, 101, 43, 60, 104, 68, 57, 
    7, 145, 132, 41, 28, 2, 16, 
    0, 55, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 66, 0, 0, 
    82, 48, 0, 27, 88, 0, 37, 
    0, 152, 0, 0, 224, 10, 0, 
    0, 113, 0, 0, 51, 0, 0, 
    0, 144, 43, 0, 0, 89, 6, 
    0, 20, 35, 0, 107, 78, 21, 
    66, 0, 96, 9, 50, 20, 5, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 3, 0, 
    25, 0, 0, 25, 34, 30, 39, 
    8, 0, 0, 29, 62, 15, 84, 
    42, 0, 2, 0, 17, 34, 52, 
    50, 62, 5, 62, 51, 73, 64, 
    144, 123, 95, 180, 238, 274, 279, 
    300, 224, 277, 272, 293, 310, 350, 
    
    -- channel=5
    156, 172, 149, 145, 113, 114, 154, 
    192, 182, 149, 125, 85, 115, 145, 
    101, 145, 46, 118, 120, 127, 96, 
    22, 129, 73, 93, 96, 93, 94, 
    0, 75, 111, 43, 89, 61, 71, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 11, 0, 30, 26, 
    32, 0, 10, 87, 89, 160, 151, 
    102, 44, 129, 169, 176, 187, 170, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    74, 84, 108, 0, 33, 45, 25, 
    107, 96, 194, 74, 0, 16, 3, 
    43, 25, 55, 42, 0, 0, 71, 
    49, 31, 9, 0, 0, 0, 49, 
    0, 7, 180, 130, 0, 113, 73, 
    0, 0, 0, 15, 17, 61, 34, 
    11, 0, 37, 26, 37, 3, 30, 
    
    -- channel=9
    0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    225, 240, 215, 173, 109, 84, 142, 
    125, 224, 145, 78, 75, 64, 62, 
    52, 169, 76, 111, 117, 72, 40, 
    56, 109, 96, 65, 73, 65, 70, 
    41, 84, 43, 42, 12, 0, 1, 
    0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    73, 31, 53, 131, 48, 45, 80, 
    79, 59, 86, 0, 14, 10, 34, 
    0, 137, 54, 0, 11, 12, 0, 
    0, 30, 107, 59, 19, 15, 0, 
    0, 0, 99, 0, 114, 62, 28, 
    121, 16, 169, 108, 0, 0, 0, 
    1, 164, 0, 0, 0, 0, 0, 
    
    -- channel=14
    36, 34, 75, 83, 17, 50, 36, 
    144, 59, 81, 144, 100, 151, 72, 
    166, 113, 83, 266, 249, 213, 84, 
    186, 160, 126, 164, 157, 189, 37, 
    239, 261, 129, 105, 142, 33, 9, 
    75, 294, 126, 0, 10, 0, 0, 
    0, 144, 46, 0, 0, 1, 53, 
    
    -- channel=15
    42, 76, 51, 34, 37, 36, 42, 
    73, 68, 35, 39, 69, 78, 58, 
    117, 76, 41, 97, 98, 73, 53, 
    57, 45, 19, 80, 124, 46, 71, 
    93, 110, 39, 0, 0, 0, 10, 
    0, 97, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    84, 128, 75, 67, 32, 34, 64, 
    39, 139, 28, 43, 25, 56, 5, 
    86, 0, 15, 73, 6, 65, 31, 
    21, 41, 0, 37, 16, 0, 39, 
    33, 87, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    31, 0, 34, 106, 60, 58, 58, 
    109, 66, 85, 18, 30, 37, 58, 
    29, 82, 89, 2, 10, 39, 9, 
    18, 55, 115, 110, 15, 47, 12, 
    0, 57, 133, 2, 135, 131, 23, 
    121, 16, 241, 138, 0, 0, 0, 
    31, 216, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    39, 17, 49, 99, 71, 41, 46, 
    112, 82, 61, 67, 87, 52, 45, 
    72, 115, 40, 93, 165, 82, 32, 
    10, 58, 103, 83, 137, 85, 24, 
    6, 152, 34, 4, 72, 12, 0, 
    0, 125, 129, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 
    95, 0, 152, 57, 4, 39, 0, 
    141, 0, 5, 53, 7, 0, 0, 
    159, 103, 70, 73, 0, 5, 0, 
    87, 203, 292, 165, 135, 164, 160, 
    138, 121, 151, 139, 162, 185, 201, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    42, 38, 26, 14, 19, 27, 9, 
    0, 40, 43, 0, 25, 0, 0, 
    44, 0, 14, 0, 0, 0, 14, 
    86, 28, 16, 16, 2, 0, 25, 
    86, 8, 47, 24, 14, 0, 30, 
    53, 17, 53, 56, 85, 134, 138, 
    174, 9, 102, 149, 151, 157, 145, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 4, 98, 0, 44, 
    0, 102, 0, 4, 257, 22, 0, 
    0, 33, 0, 0, 139, 42, 0, 
    0, 115, 0, 0, 0, 27, 0, 
    0, 123, 60, 0, 32, 7, 0, 
    117, 0, 114, 15, 28, 39, 34, 
    
    -- channel=29
    79, 67, 59, 92, 71, 58, 83, 
    97, 110, 108, 67, 32, 24, 29, 
    0, 117, 21, 21, 77, 34, 0, 
    0, 68, 7, 6, 14, 21, 13, 
    0, 46, 104, 0, 18, 25, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    101, 157, 112, 106, 63, 58, 61, 
    30, 133, 131, 84, 7, 92, 12, 
    18, 60, 45, 104, 0, 56, 34, 
    21, 32, 34, 101, 29, 31, 53, 
    50, 0, 52, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    39, 17, 47, 84, 42, 35, 44, 
    65, 54, 51, 63, 32, 42, 0, 
    158, 124, 158, 67, 64, 89, 0, 
    106, 68, 75, 91, 33, 53, 0, 
    90, 166, 105, 38, 87, 17, 20, 
    100, 141, 301, 84, 79, 53, 51, 
    34, 39, 55, 7, 3, 28, 10, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 43, 0, 59, 0, 
    56, 0, 0, 148, 0, 136, 51, 
    193, 0, 0, 249, 0, 270, 58, 
    227, 108, 0, 169, 0, 215, 0, 
    122, 59, 66, 19, 65, 37, 0, 
    0, 0, 210, 0, 70, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 
    
    -- channel=34
    21, 64, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 10, 43, 51, 
    53, 0, 39, 91, 104, 100, 39, 
    
    -- channel=35
    67, 38, 57, 77, 30, 0, 52, 
    12, 28, 28, 0, 30, 5, 8, 
    26, 99, 100, 0, 7, 11, 0, 
    0, 12, 95, 57, 50, 24, 17, 
    0, 0, 0, 0, 44, 0, 0, 
    54, 54, 141, 34, 0, 0, 0, 
    0, 98, 0, 0, 0, 0, 0, 
    
    -- channel=36
    13, 28, 0, 0, 0, 0, 0, 
    0, 10, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 28, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 16, 0, 
    0, 0, 0, 124, 0, 11, 27, 
    77, 0, 0, 0, 0, 22, 0, 
    0, 61, 61, 76, 0, 0, 0, 
    0, 0, 96, 0, 67, 61, 49, 
    29, 0, 107, 70, 88, 65, 120, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 16, 61, 40, 
    81, 0, 148, 162, 195, 246, 238, 
    229, 126, 210, 235, 256, 275, 278, 
    
    -- channel=39
    259, 271, 203, 201, 100, 62, 146, 
    45, 193, 64, 1, 0, 0, 0, 
    0, 98, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 80, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    0, 0, 37, 40, 17, 68, 27, 
    118, 26, 95, 103, 3, 75, 92, 
    118, 104, 45, 156, 53, 104, 80, 
    89, 88, 7, 42, 50, 96, 0, 
    42, 143, 158, 98, 96, 92, 51, 
    29, 182, 220, 45, 89, 54, 30, 
    29, 59, 44, 0, 0, 0, 21, 
    
    -- channel=41
    60, 36, 71, 53, 60, 32, 35, 
    8, 47, 41, 24, 22, 0, 8, 
    18, 85, 117, 0, 17, 21, 2, 
    15, 65, 76, 0, 15, 38, 11, 
    0, 0, 19, 50, 27, 20, 26, 
    0, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 
    51, 59, 105, 0, 34, 0, 0, 
    0, 0, 30, 0, 82, 0, 24, 
    0, 0, 0, 0, 0, 0, 27, 
    0, 68, 168, 123, 0, 0, 75, 
    0, 66, 0, 0, 32, 171, 94, 
    0, 0, 0, 15, 84, 38, 106, 
    
    -- channel=43
    123, 150, 80, 0, 29, 0, 55, 
    39, 114, 0, 0, 52, 0, 0, 
    0, 8, 0, 0, 113, 0, 0, 
    0, 13, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 68, 
    0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 
    0, 0, 71, 0, 0, 0, 2, 
    62, 0, 53, 0, 0, 0, 0, 
    218, 0, 0, 32, 0, 0, 0, 
    154, 87, 0, 103, 57, 131, 132, 
    8, 220, 0, 102, 152, 164, 204, 
    
    -- channel=45
    35, 10, 19, 18, 16, 0, 27, 
    0, 0, 4, 0, 8, 0, 2, 
    0, 54, 44, 0, 0, 0, 0, 
    0, 0, 51, 1, 13, 0, 7, 
    0, 0, 0, 0, 0, 50, 11, 
    63, 0, 0, 49, 0, 0, 0, 
    9, 93, 0, 0, 0, 0, 0, 
    
    -- channel=46
    172, 142, 87, 146, 127, 107, 142, 
    67, 160, 58, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 0, 31, 64, 181, 
    0, 0, 0, 17, 40, 86, 103, 
    34, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    1, 0, 0, 18, 7, 13, 42, 
    151, 7, 26, 44, 109, 23, 109, 
    0, 211, 0, 17, 272, 76, 0, 
    0, 83, 86, 0, 186, 64, 0, 
    0, 117, 110, 0, 46, 42, 13, 
    43, 129, 31, 0, 0, 0, 0, 
    97, 56, 51, 0, 15, 14, 40, 
    
    -- channel=49
    42, 43, 3, 0, 14, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 7, 
    38, 0, 0, 47, 0, 20, 65, 
    14, 57, 23, 75, 77, 77, 58, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 6, 0, 0, 0, 33, 21, 
    95, 39, 0, 23, 11, 0, 84, 
    0, 0, 0, 0, 67, 0, 17, 
    0, 64, 0, 0, 0, 0, 0, 
    0, 46, 73, 0, 0, 10, 26, 
    0, 0, 0, 0, 23, 49, 0, 
    20, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 0, 0, 36, 0, 
    56, 0, 1, 0, 0, 0, 41, 
    11, 0, 0, 0, 0, 0, 7, 
    2, 0, 0, 0, 0, 0, 0, 
    0, 0, 128, 0, 37, 101, 56, 
    101, 0, 155, 192, 162, 213, 208, 
    253, 94, 147, 162, 175, 201, 190, 
    
    -- channel=54
    83, 109, 20, 33, 1, 0, 52, 
    0, 39, 0, 0, 6, 0, 0, 
    0, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 79, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 
    103, 0, 0, 0, 6, 0, 0, 
    101, 0, 0, 41, 34, 65, 95, 
    190, 107, 61, 125, 143, 156, 166, 
    
    -- channel=57
    33, 69, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 50, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 40, 22, 
    0, 0, 0, 52, 69, 60, 9, 
    
    -- channel=58
    147, 142, 137, 151, 117, 110, 150, 
    177, 178, 127, 80, 107, 83, 116, 
    106, 179, 104, 75, 129, 90, 71, 
    39, 112, 97, 83, 102, 62, 90, 
    0, 93, 110, 47, 93, 35, 101, 
    14, 19, 23, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 47, 0, 
    0, 2, 0, 0, 0, 66, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 106, 0, 0, 0, 0, 0, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 81, 0, 
    113, 0, 15, 42, 0, 0, 81, 
    0, 0, 0, 43, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 96, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
