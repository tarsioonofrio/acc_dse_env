library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    28389, 4094, 2684, -7314, 2181, 899, 12211, 6059, 16087, -2835, -7048, -29240, -13051, -55056, -157, -12551,

    -- weights
    -- filter=0 channel=0
    25, 60, -18, 43, -28, -45, 15, -1, -50,
    -- filter=0 channel=1
    9, 9, -52, -6, -56, -75, -22, -9, -77,
    -- filter=0 channel=2
    14, -22, 4, 69, -6, 6, 18, 4, 5,
    -- filter=1 channel=0
    0, 2, -58, -72, -79, -93, -52, -43, -60,
    -- filter=1 channel=1
    95, 43, 4, 35, 82, 27, 46, 2, 40,
    -- filter=1 channel=2
    90, 64, 21, 12, -9, 62, 63, 8, 27,
    -- filter=2 channel=0
    -15, -76, 5, -49, -59, -43, -62, -76, -29,
    -- filter=2 channel=1
    51, 12, -28, 36, -30, 30, 54, 20, -23,
    -- filter=2 channel=2
    39, 78, 47, 70, -4, 12, 16, 1, 77,
    -- filter=3 channel=0
    -4, -33, -13, -6, 24, -10, 5, 32, -34,
    -- filter=3 channel=1
    -29, 7, -10, -35, -27, 48, 40, -24, 20,
    -- filter=3 channel=2
    -2, -37, 16, 41, -22, -17, -8, -47, -21,
    -- filter=4 channel=0
    45, 70, -20, 35, 37, 0, -15, 6, 36,
    -- filter=4 channel=1
    -11, 56, 24, 58, 46, -27, 15, -12, -15,
    -- filter=4 channel=2
    -25, 17, -53, -22, 18, 17, -72, -74, 9,
    -- filter=5 channel=0
    37, 50, -41, -35, -48, 47, 43, 8, -16,
    -- filter=5 channel=1
    33, 5, -55, 30, -45, 36, -51, -32, 31,
    -- filter=5 channel=2
    28, 0, -18, 44, -9, 22, -33, -26, -12,
    -- filter=6 channel=0
    21, -7, 9, 50, -6, -12, -46, 45, -6,
    -- filter=6 channel=1
    4, 41, -23, 27, 30, 9, -27, -40, -2,
    -- filter=6 channel=2
    -22, -41, 45, -47, 36, -38, -56, -47, -22,
    -- filter=7 channel=0
    13, -45, -5, -43, -22, -4, -18, -26, -8,
    -- filter=7 channel=1
    59, 54, 40, 74, 0, 76, 80, 2, 79,
    -- filter=7 channel=2
    -48, -47, -12, -58, -34, -29, -19, 16, 27,
    -- filter=8 channel=0
    67, 58, 89, 62, 31, 40, 40, 60, 75,
    -- filter=8 channel=1
    59, 107, 74, 14, 17, 111, 59, 74, 34,
    -- filter=8 channel=2
    -132, -67, -109, -150, -60, -69, -144, -110, -145,
    -- filter=9 channel=0
    -45, 19, -33, -42, 21, -14, -44, 23, -22,
    -- filter=9 channel=1
    11, 36, -34, -9, 16, 18, 13, -21, 42,
    -- filter=9 channel=2
    10, 4, -47, 39, -22, -10, 0, 50, 45,
    -- filter=10 channel=0
    -33, 0, -3, -4, 36, 16, -47, -41, -42,
    -- filter=10 channel=1
    -31, -10, -44, -6, 30, 28, 29, -17, -8,
    -- filter=10 channel=2
    -45, 24, 1, 34, 3, -34, -49, 30, -13,
    -- filter=11 channel=0
    3, 29, 16, -43, 23, -8, -27, 26, -44,
    -- filter=11 channel=1
    66, 61, 92, 66, 24, 86, 43, 59, 28,
    -- filter=11 channel=2
    -26, -18, 51, -20, 19, 47, 53, 3, -11,
    -- filter=12 channel=0
    33, 16, -13, -20, -35, -43, 20, 32, -42,
    -- filter=12 channel=1
    -16, 26, 18, -25, 18, -21, -11, 5, -12,
    -- filter=12 channel=2
    3, -6, 37, 45, -12, 65, 12, 39, 42,
    -- filter=13 channel=0
    7, 2, 9, 54, 39, 55, 27, 47, 64,
    -- filter=13 channel=1
    -63, -40, -40, 12, 8, -50, 27, 2, 29,
    -- filter=13 channel=2
    67, 0, 84, 61, 69, 47, 109, 71, 92,
    -- filter=14 channel=0
    -38, 50, 51, -36, -15, 25, 0, 4, -37,
    -- filter=14 channel=1
    23, -36, 52, -58, -56, 29, -38, -48, -41,
    -- filter=14 channel=2
    7, 76, 87, -15, 44, 64, -42, -27, 69,
    -- filter=15 channel=0
    18, -43, -5, -1, 13, 23, 9, -33, 34,
    -- filter=15 channel=1
    20, 11, -30, 4, -24, -32, 4, 8, -41,
    -- filter=15 channel=2
    -1, -17, -36, -32, 5, 48, 39, 14, 25,

    others => 0);
end iwght_package;
