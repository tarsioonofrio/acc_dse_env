library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    -11774, -1473, -5599, 14140, 15406, -18950, 18901, -4627, -455, -5733,

    -- weights
    -- filter=0 channel=0
    0, 16, -9, -13, -9, 9, 7, -5, -20, 19, 0, -12, 26, 1, 17, -19, -28, 13, 6, -5, -25, -10, -2, 7, 23, 7, -19, 24, 11, -8, -5, 7, 14, -1, -13, 12, -16, 11, -6, -14, 13, -6, -15, 2, 1, 1, 4, -2, -7, 5, 10, 4, -5, 6, 0, 0, -5, 0, 0, 1, 17, 18, 0, -24, -26, 7, 2, 27, -25, 20, -18, -2, 9, -5, 6, -3, 2, 2, 19, -9, 17, -9, 10, -12, -2, -14, -4, -22, 22, -2, 4, 8, -12, 0, 28, 11, -50, 39, -18, -20, -2, -16, 1, 10, 8, -24, -20, 17, 16, 9, -12, -14, 9, 5, -4, 12, 20, 3, -8, -14, 2, 13, 8, 0, -33, -16, 7, 16, 14, -20, 4, -25, 38, -17, -12, 11, -2, 0, -1, 0, -2, -13, -27, -8, 18, 18, 33, 5, -5, -14, 5, -3, 2, -4, -3, -3, 1, 3, 0, -4, 8, -19, 4, -17, 3, 14, 19, -15, 22, -17, 2, -2, -13, 7, 6, -4, 2, -7, 0, 8, -16, 7, 13, 3, -13, 16, 21, -24, -6, -12, -3, -12, 27, -10, 10, -1, -11, -12, -4, 15, -8, -3, -3, -7, 0, 13, 5, 3, -3, 16, -3, 4, -24, 27, 11, 3, 20, -10, -12, -3, -5, -1, 1, -3, 4, -8, 0, -6, 0, 14, -8, -3, -24, 19, 15, 24, 9, -6, 7, -20, -1, -21, 6, -11, -5, -4, 33, -13, 9, 8, 12, -16, 8, 11, -7, -18, 6, 4, 14, -11, 6, -2, -8, -19, -11, 14, 4, 7, -7, 17, 2, 1, -6, -16, 22, -27, 25, -7, -17, 7, -1, -11, 7, 29, -3, -38, 30, -10, -25, 15, 2, 5, 10, -12, -16, 12, -4, 5, -16, 17, -27, -18, -14, 20, -10, -9, -9, 16, 17, 21, -8, 9, 6, -3, -7, -3, 0, 8, -7, 8, -14, -1, 12, 9, -6, -15, 20, -3, 17, -14, 17, 11, 0, 10, 0, 7, -13, -6, -32, 21, -10, 0, -9, 4, 21, 1, 16, -17, -21, -10, 0, 15, -1, 7, 2, 13, -16, 3, -16, 1, -15, 13, 33, 11, 10, -12, -16, -4, 0, -12, 26, -7, 51, 29, -1, -32, -17, -37, 23, -34, -19, 9, 11, 6, -11, 15, 32, -23, -7, -17, 0, 5, 3, 13, 1, -3, -5, 1, 13, -15, 0, -10, -12, 17, 9, -16, -6, -11, 21, 13, 17, 5, -3, -17, 4, -5, -3, -18, 28, -3, 1, -3, -4, -3, 0, -4, 3, -1, -3, 0, 2, 6, -29, -1, 20, -8, -2, 21, 13, -4, -1, 0, 9, 0, -4, -4, 4, 2, -4, -2, 8, -20, 15, 7, -22, -24, 13, 22, 10, -17, 6, -6, -22, -11, -10, 33, 12, 7, 13, -20, 10, 21, -5, -5, 8, -11, 0, -10, -20, -5, -13, 0, 5, 3, -27, 12, 6, -3, 15, -4, -1, -15, 3, 17, 0, 16, -22, -15, 34, -28, 10, 2, -17, 11, 4, -25, 13, 4, -8, -12, 40, 1, -12, 13, -9, -7, 6, -3, -20, -10, -8, 1, 3, -12, 0, 18, -10, 10, -19, 5, 8, 2, 0, -19, -26, -7, 10, 5, -9, 29, -18, -9, -9, 1, 14, -11, 15, 20, -20, 19, -13, 17, 3, 17, -19, 10, 16, -14, 0, -13, 23, -26, -9, 21, -1, -8, 7, -25, 36, -19, -18, 42, -6, -3, -9, -12, -5, -14, 12, 16, -10, 1, -2, -4, -2, -3, 0, -10, 31, 8, -11, 8, -1, 13, 2, -12, -2, -2, 3, -4, -17, 14, -10, -7, 11, 11, 21, -15, 4, -2, -1, 6, -9, -7, -4, 9, 4, -4, 5, 13, 0, 3, 2, -5, 2, 0, -12, 0, -5, 14, 33, 34, -17, 15, -19, -43, -2, 3, -28, 29, -2, 3, 2, 3, 3, 4, -3, -4, -1, 2, -4, 0, -4, 8, -1, -4, -18, 22, -10, 4, -5, -6, 0, 4, -1, -1, 0, -2, -1, 11, -5, -1, -7, 5, 3, 5, -24, -7, 7, 6, -11, 1, 11, -3, -7, 0, 7, 7, 3, 0, -20, -12, -10, 14, 4, -14, 16, 19, 17, -10, 19, -22, 31, -8, 39, -14, -22, -29, 29, -26, -6, 8, -4, 0, 0, 3, 8, -1, 10, -3, -24, 28, 17, 1, 1, -31, 1, -15, -3, 35, -10, -13, -23, 3, 21, 14, -14, 8, 6, 4, 19, -5, 21, -11, 0, 19, -11, -31, -1, 16, 14, -7, 2, -16, 13, 29, -3, -20, -4, -19, -2, 0, -15, 8, -2, 9, 5, -11, 1, 4, 5, 4, 3, -18, -1, -10, 18, 1, -11, -5, -11, 8, 3, -6, 17, -14, -10, 5, 0, 0, -6, -1, -27, 15, 19, 0, 0, 0, 9, -11, 37, 22, -36, -21, -28, -24, 1, 30, 6, 7, -1, -17, 3, -10, -14, -14, 1, 22, 14, 19, 4, -3, -7, -9, 10, 8, -3, -1, -6, -5, 8, 1, -14, 9, -9, 5, 11, 3, -16, 8, -6, -5, 7, 40, -7, -32, 13, -11, 1, -8, -31, -15, -29, 29, 6, 21, -10, 9, 18, -16, 11, 18, 14, -12, -12, 1, -3, -16, 5, -4, 5, 21, -16, 6, -5, -22, 34, -11, -2, -6, -13, 29, 6, 3, -7, -21, -2, 0, -6, 9, 16, -10, 1, 15, -12, 11, -9, 9, -11, -11, -9, 0, 17, 13, -6, -11, 5, -12, 1, 5, 0, 0, -10, 6, 10, -4, -2, -3, 1, 17, -20, -12, -8, 47, -12, 2, -3, -9, 13, -1, -21, -4, 34, -9, 21, -12, -4, -3, 3, -2, -22, -5, 37, 8, -4, -13, 8, -25, 3, 3, 2, 26, 8, 5, -18, 0, 4, 1, -14, -5, 5, -4, -25, 25, 7, -10, 16, 7, -1, -13, -1, -22, -35, 7, 13, -22, -2, 14, 22, 23, -3, 11, 1, 5, 2, 0, -7, -5, 0, -5, 0, 0, -5, -1, -2, 6, 6, 0, 0, 0, 0, -4, -14, -12, 2, -11, 12, 21, -8, 0, 1, 0, -2, -6, -4, 7, 4, 1, -5, 0, 6, -8, -10, -14, 7, 11, 13, 1, 2, -7, 24, -10, -14, -3, 14, -22, -5, -9, 7, 0, 5, 34, -1, -26, 22, -2, 6, -16, 2, -17, 3, 3, -10, -7, 10, -1, -6, 15, -6, 1, -4, 19, 9, 5, -6, 9, -15, -5, -12, 6, -3, -1, 25, -6, -15, 12, -3, -2, 0, -6, -1, 8, 3, 0, 14, 7, -18, -7, -9, 12, -22, -16, -2, 26, -20, 20, 0, 4, 19, 4, 0, 5, -3, 3, -5, 0, -2, -2, 2, -5, -11, 23, -16, -17, 31, 6, 8, -31, 9, 0, -4, 0, 15, -6, 18, -2, -19, 8, -9, -7, 6, 0, 1, -25, 6, 34, 9, 2, -17, -11, 0, -2, -5, 0, -1, -4, -2, -3, -5, -6, 1, -30, 9, 1, -8, 19, -9, -3, -13, 16, 36, 8, -14, -13, 9, -44, 13, -7, -21, 26, 2, 11, -17, 5, 1, -27, -27, -13, 22, 27, 1, -5, 6, -10, 5, 0, -1, -7, 5, 7, -10, -9, 0, 11, -17, 13, 8, 14, -12, 17, -20, 3, -5, 31, -7, -13, -5, -6, 3, 18, 7, -5, 22, -15, -33, -8, 2, 38, 0, -2, 3, 3, -9, -10, 28, -16, 9, -8, 3, -3, 6, -2, 6, 7, 0, -2, -9, -5, 1, -1, -11, -1, 3, 23, -1, -8, -12, -11, -3, 4, -10, -5, 2, 2, -4, 1, 3, 3, 18, -1, -8, 10, 0, -3, -12, 10, 13, -10, -12, 7, 2, -2, 1, 2, 3, 0, 2, -2, -1, 4, -20, -1, 1, 14, 31, -10, 41, -9, -22, -12, 22, -31, 12, -26, 37, -31, 8, 26, -6, -14, -8, 0, 21, -4, 12, 0, -13, 30, -7, -35, -3, 37, -14, 9, -16, 1, 25, -33, 20, -15, 1, 5, 0, -27, -22, 1, -1, 34, -3, 16, 10, 13, -4, -1, 6, 3, 23, 0, -21, -29, -15, -12, 7, -4, -18, 21, 22, -6, 0, 1, -38, 12, 9, 8, -7, 22, 28, 2, -18, -18, 23, -7, 7, 21, -17, -19, 3, -10, 0, -6, -11, 24, 27, -14, -41, -7, 6, -9, 12, 8, -9, -25, -31, 21, -5, 35, -9, 37, 3, -25, -25, 21, -27, -5, -12, -14, 12, -11, 16, 33, -23, -6, 1, 10, 27, 6, 19, -20, -12, -20, 6, -4, 3, 24, 2, 16, -8, -18, -8, -2, -2, 0, -14, -7, 5, 5, 9, -4, 3, -3, 17, -1, 4, -23, 10, 16, -12, 24, 5, -23, -29, -7, 0, 32, -24, -23, 16, 0, 43, 7, -18, 0, -25, 41, -8, 14, 27, -28, 4, -19, -1, -14, -4, 1, -28, -7, 47, -7, -9, 9, 1, -8, 7, -8, 4, 2, 3, -2, 6, 6, 12, -6, 2, -17, -12, 10, 8, 0, -7, 8, -6, 0, 13, 5, 0, -8, -4, 9, -3, 7, -4, 9, 21, 0, 14, -30, 1, -1, -11, 0, 3, 0, -6, -20, 17, 14, 19, -16, -6, -1, 14, -3, -4, -10, -27, 12, 19, -5, 27, -27, 0, 3, 7, 8, 1, -13, -3, -2, 0, -3, -27, 9, -7, 17, 23, 19, -16, 21, -11, -21, -17, -10, -28, 13, 13, 5, 14, 12, -23, 8, 0, 0, -1, -5, -3, -3, -4, 3, 3, 1, 8, 2, -1, -4, -9, 1, -3, 7, -2, -8, 3, 5, -16, -1, -24, 26, -9, -18, 23, 3, 14, -7, 3, -20, 2, 12, -2, -1, 9, -6, -31, 6, 32, 18, 14, -20, 5, -29, -5, 4, 14, 4, 12, -38, 10, 11, 22, -15, 2, -9, 8, 4, -8, 3, 0, 4, 3, -10, -4, -4, -2, 4, -9, 1, 10, 10, -25, 19, 9, -18, 12, -30, 32, 2, 13, 20, -8, 10, -4, -38, 0, 4, -1, 8, 1, 0, 7, -14, 5, -3, 9, -1, 8, 0, -3, -2, -2, 4, -8, 2, 13, -9, 3, -9, -2, 11, 0, -9, 9, -10, 20, 5, 6, -5, -5, -4, -10, -18, 19, 7, -5, -5, 4, -1, 0, 6, -2, 0, 0, 0, 20, -20, 27, 8, 7, -12, -8, -14, 11, -28, -2, -5, 1, -4, 15, -3, -9, 0, 0, 3, -6, -2, 8, 7, -13, 15, 14, -13, -11, 8, 37, -4, -14, 19, 16, 0, 20, -17, -38, -17, -10, -6, 8, 19, -3, 5, -16, -3, -13, 1, 18, -18, -9, -29, 25, -29, 20, 11, -10, 10, 3, 1, 15, 16, -5, -9, -1, -1, 3, 0, -30, -12, -13, 11, 37, -28, 18, 17, 6, -16, 16, 24, -11, -11, -12, -10, 1, 6, -6, 1, 9, -4, 25, -27, 8, 18, 5, -9, -8, -10, -16, 13, 18, 0, -5, 11, -15, 10, -14, -10, 1, 0, -2, 6, 4, -6, -5, 5, 2, 3, -6, -2, 7, -5, 7, 10, 0, -6, -9, 20, 20, -14, -32, 7, -5, 24, -12, 6, 13, -3, 9, 28, -1, 12, 0, -22, -12, -9, 16, -4, 4, -21, 12, 22, -10, 36, 17, -27, -11, -25, -11, -2, -2, -7, 0, 0, 5, 0, 13, 3, 1, -2, 3, 3, -3, -3, 2, 4, 3, -3, 31, -58, 6, 0, 33, 1, -12, -11, 21, -25, -3, 24, 0, -4, -3, -11, -5, -9, 15, 17, 6, 28, 30, -7, -30, 22, -4, -24, -18, -5, -7, 6, -25, 25, -3, 6, -6, -11, 2, 0, -29, 24, 48, -14, -7, 4, -24, -7, 1, 22, -20, -9, 8, 7, 0, -36, 4, 1, 11, 45, -5, -23, 11, 9, 2, 22, 7, 23, -12, -33, 8, 4, -15, -13, -8, -4, -13, 26, -2, 21, 4, 15, 24, 5, 28, -20, -28, -17, -8, -20, -14, -15, 3, 16, -17, -2, 19, -13, 47, -20, 4, -27, -1, 23, -10, -4, -5, 6, 0, 6, -35, 0, 18, 12, 5, -17, -26, -6, 18, 23, -17, 4, 30, 22, -3, -38, 22, -33, 15, -4, 17, 9, -20, 0, 19, 0, -12, -11, 22, -17, 20, -16, -8, 0, 1, 1, 4, -13, 25, -14, 1, -4, -8, -6, 15, 27, 19, -12, -7, -11, 6, 1, -10, -20, 6, 33, -24, 14, -6, -10, 34, -5, -12, -20, -3, -17, 10, -16, 49, -16, -3, -8, 0, -8, 6, 22, -16, 2, 0, 10, -6, 6, -4, -13, 5, 6, -12, 6, -3, 11, -9, 17, 0, -23, 14, 11, 25, -22, -8, -1, 0, -22, 8, -3, 0, 32, 7, -19, 2, 7, 26, 2, 42, 10, -12, -23, -16, 6, -23, -17, -11, -13, 23, 29, 15, -6, -8, -3, -3, -15, -27, 9, 9, -18, 24, 20, -8, 13, 9, -14, -17, -1, 2, 9, 4, 8, -13, 5, 12, -5, -9, -1, -6, -2, 9, 2, -12, 10, 6, 12, 2, 5, -6, 9, -6, 3, 0, 3, -1, -1, 11, 4, -5, 18, -14, -16, 1, 22, -14, 3, -13, -4, 16, -23, 7, 5, 9, 6, 2, -6, 0, -3, 0, -14, -11, -7, 7, 22, 8, -5, 0, 6, -1, -2, -2, 3, -3, -6, -4, 4, -5, 3, -12, -2, 17, 2, 7, 1, -37, 28, 4, 13, 4, -9, -15, -10, -3, 12, 8, -7, -3, -3, 0, -11, 15, -5, 2, -4, 0, 8, -10, 1, -6, 12, 2, 0, 0, 8, 2, -5, -12, -11, -1, 17, -13, 6, 14, -4, 6, -13, 8, -4, 5, 2, -7, 11, 0, 6, -8, -7, 28, -1, -20, 0, -9, -31, -2, 9, 9, 10, -14, 4, 5, -11, -16, 17, 4, -6, 21, 1, -3, -3, 14, -2, -24, -9, 16, 11, -16, 5, -9, 10, -13, -5, -2, -9, 0, 33, 0, -6, -2, 0, 2, -3,
    -- filter=0 channel=1
    0, -4, 6, -1, 8, -4, -2, -1, -2, 0, 0, 2, -5, 4, 1, 4, 43, -16, 20, -26, -14, -4, 2, -19, 24, -11, -25, -15, -6, 26, -3, 6, -13, 10, 2, 13, 46, 4, 0, 1, -6, 2, 0, 4, -34, -4, -34, -16, 15, 24, 26, -2, -16, 19, 8, -29, 0, -10, 9, 15, 14, -3, 7, -26, -3, -4, -16, -10, 6, -19, 33, -14, 19, 6, -7, -17, -14, 30, 4, -15, -21, 2, -10, 9, -19, 34, 24, 13, -1, 0, 1, -43, 4, 22, -5, -8, -11, -2, 15, 2, -19, 6, -1, 14, -6, 9, 5, 17, 0, -3, 23, -31, -17, -10, 23, -3, -2, 0, 11, -7, 1, 4, 3, -5, 0, -2, 5, -17, 11, -5, -21, 1, 26, -9, -6, 6, 17, -38, 28, -4, -18, -5, 15, -4, 0, 19, -8, 1, 0, 5, 0, -1, 0, 1, 2, -4, -3, 9, -10, -8, -3, -19, 5, 2, 17, 1, -13, 20, -17, 18, -14, 3, 15, -31, -4, 9, 5, -5, -18, -29, 26, 6, 17, 6, -21, 7, 6, -22, -1, 22, -41, -6, 24, 8, 6, 8, 8, 5, -10, 5, 8, -7, 4, 1, -7, 4, -17, -1, -14, 5, 5, 12, -16, 20, -2, 6, 3, 2, 7, -10, 0, 19, 10, -3, -19, 0, -19, 30, 7, -25, -10, -9, 31, -8, 5, 8, -4, 1, 0, -6, 8, -9, -10, 0, 18, 7, 3, 6, -3, -11, -14, 6, 7, 2, -10, 5, 7, 35, 0, -7, -1, 3, 1, -7, -12, -10, 0, 1, 9, -14, -2, 16, 11, 0, -1, -13, 7, 13, -21, 20, -10, 14, -9, -20, 9, 0, 20, 24, -15, 0, -34, 14, -7, 17, 2, -19, 6, 6, -16, 0, 10, 2, -3, 8, -2, -4, 9, 0, -2, 1, -2, -4, -1, -8, 25, -14, 1, -24, 9, -2, 1, 8, -4, -14, 5, 12, 6, 23, 9, -2, 4, -19, -6, -2, -14, 0, 2, 1, 15, -1, 2, -3, -3, -10, 1, -2, -9, 11, -22, -1, -6, -3, -15, -2, 24, 20, 2, -5, -4, -14, 0, -5, -7, 18, -21, 16, -10, -17, -7, 5, 0, 0, -7, 9, 12, 21, 20, -19, 27, -10, 28, 0, -3, -24, 4, -9, -17, -1, -24, 2, -14, -4, 8, 25, 11, 10, -15, -1, -2, 0, 10, 8, -1, -12, 18, 0, 16, 2, -11, -10, -10, 16, 12, 2, -13, -2, -7, 13, -3, 0, -14, -3, -13, -10, 20, 16, 16, -11, -2, -14, 5, 22, 1, -13, 20, -13, 22, -12, -15, -4, -23, -11, -6, 7, 16, 40, 31, -25, -15, -9, 11, 0, -9, 24, -32, 25, 5, 12, 7, -4, 16, 9, -31, -12, -20, 13, 0, 2, -1, -7, 4, 5, -9, 0, 2, 4, -8, -2, 30, 28, -28, 10, 20, -11, -16, -31, -3, -13, -7, 12, 0, 7, 0, -10, -11, 29, -12, -3, 12, 14, -26, 15, -14, -3, -5, 14, 31, -12, 3, -8, 2, 9, -19, 34, -28, -5, 10, -7, 0, 6, 0, -9, 5, -4, 4, -7, -4, -14, 10, 12, 9, 16, -41, 44, -5, -26, 5, -2, -9, 3, 14, -21, 10, 3, 7, 1, 1, 7, -11, 14, -3, -18, -5, 11, 0, 3, 0, 25, -12, 11, -10, -11, -24, 6, 15, -10, 6, -5, 8, 10, 3, -22, 5, -1, -12, 3, -11, -20, -6, 38, 20, 17, -20, 9, -1, -28, -4, 0, -1, -1, 9, 0, 1, -7, -2, 8, -14, -4, 7, 9, -10, -2, 0, 8, 15, -5, -20, 5, 1, -15, 0, 0, -7, 9, 1, 15, 2, 3, -3, -2, -2, 4, -1, -4, 1, -3, 7, 3, 11, 7, 28, -16, -42, 26, 2, -21, 25, -9, 0, -9, -5, 5, 10, 0, -5, -7, -25, 30, 0, 12, -22, -5, -3, -12, -8, 20, -12, -7, -4, -10, 0, 7, -2, -3, 11, 1, 11, 1, -13, -3, 4, 6, -7, -8, 4, -1, -2, 2, 4, 1, 5, -3, 0, 0, -4, -3, -6, 0, -5, -4, -3, 13, 3, 2, 11, 0, 14, -8, -8, -10, 7, 5, -6, 8, -1, 4, -9, -12, 5, -32, 34, -23, 27, 27, -20, 2, -8, -19, -11, 19, 14, 11, 5, 18, -4, -6, 22, 4, -19, -18, -14, -10, -2, 2, -5, 22, 3, -6, 48, 6, -18, 23, -7, -36, -16, -6, 24, -22, -1, -21, 15, -8, -42, 24, 30, 1, -14, 6, -4, -14, -9, -1, 12, 6, 18, 5, -13, 0, 14, -4, 20, -9, 12, -5, -12, -11, -23, 29, -7, -7, -12, -14, -27, 3, 20, 37, 0, -5, -10, -2, -2, 11, -9, 10, -4, -1, 17, 5, -13, 16, -24, 2, 24, -15, -9, 0, -1, -3, 5, 4, 14, -26, 8, -9, 23, -17, -23, -3, 5, 7, -3, 1, -21, 21, 22, 5, 9, -12, -8, -14, -4, 26, -31, 18, 7, 7, 1, -15, 11, 16, 31, -19, -29, 18, 4, -17, -7, 7, -11, 19, -19, 10, 7, -17, -7, 8, -1, 4, 0, -3, 4, 2, 4, 3, 0, -4, -39, -33, -29, 42, 19, 15, -6, -4, 12, 26, -1, 3, 13, -20, 2, 8, 6, -9, 3, -1, -10, -8, 3, 10, -1, -12, -1, -6, 9, -5, -3, -8, -6, -5, 16, 0, -7, 0, 5, 2, -32, -23, 23, 22, 29, 9, 14, -11, -29, -1, 9, 23, 10, -6, -8, 22, -5, 5, -22, -13, 28, 17, 14, -13, -15, 9, -30, -22, 32, -6, -15, -11, -2, 20, 0, -2, -4, -5, -7, 24, 8, 6, 7, -15, -31, 1, 9, 21, -2, -9, 3, -3, 4, -4, 3, 2, -3, -3, 3, 2, -14, -7, 3, 23, -5, -25, 2, 0, 5, 0, 14, -6, -7, -21, 15, 5, -21, 7, 4, 15, -13, 26, -17, -28, 6, -21, 10, -15, 29, 29, 16, -12, -13, -18, 25, 4, 5, 6, -26, 9, 26, -18, 10, 27, 6, 11, 0, 0, -34, -17, 4, -4, 0, 2, -3, 9, -5, 1, 0, -7, -7, 34, 1, -5, 13, 11, -9, -13, 2, -14, -4, -16, 2, -14, -10, 24, -9, 24, -17, 18, 13, 15, 9, -2, -4, -13, 2, -13, -23, 7, 0, 11, -1, 0, 28, -29, 26, -22, 8, -12, -2, 24, -3, 13, 17, -25, 3, -14, 15, -26, -23, -2, -25, -13, -14, 29, 13, 11, -6, 24, -10, 5, -2, -6, 11, 0, 1, 5, -8, 2, -1, 4, 2, 4, 3, 3, -5, 4, 1, 6, 33, -1, 17, -13, 3, -10, -3, -18, -7, -2, 5, 22, -5, 8, -1, 2, -12, -11, 0, -10, 2, -27, 21, -28, 1, 6, 14, 27, -12, 0, -8, 15, -17, -7, -2, 12, 10, 12, 6, -14, 14, -7, 13, -13, -8, 2, 3, 9, -4, -2, -4, 0, -2, 7, -5, 1, -5, -4, -2, 4, 6, 6, 19, 2, 0, 2, -7, -17, -26, 15, -4, -1, 0, -2, -1, 1, -3, 0, -1, 3, 10, -15, 26, 24, -5, -11, -23, 12, -17, -2, 6, -8, -2, -28, 2, 11, -21, 31, -7, 17, 17, -1, -11, 7, 5, -4, -8, -7, -7, -10, -17, -3, -4, -20, -4, 13, 4, 0, 13, 14, -1, 0, -5, 16, -15, 21, -18, -9, 4, 7, 32, -18, 22, -20, -2, -5, 8, -36, 18, -2, -4, -20, -15, 9, 15, 4, -20, 15, 23, -3, 0, 3, -11, -10, 0, 9, -4, 7, -3, -6, 17, 3, -9, -3, 5, -18, 8, -5, 13, -15, 19, -5, 11, -8, 14, 10, -6, -6, 1, -19, -11, 30, -1, 13, -11, -14, 18, -6, -25, 12, -32, 14, -18, 10, 27, -7, -22, 23, 12, -15, -9, -5, 10, -6, 17, -2, 19, 7, -10, -5, 7, 2, 0, 4, 0, -4, 0, -5, -6, 0, -10, -10, -3, -19, -8, 28, 11, 21, -14, -10, 4, -43, 33, 20, -17, -1, -20, -12, 16, 8, -35, 34, -54, 5, -2, 14, 20, -20, 39, 0, -5, -26, 8, -7, 6, 7, 0, -2, 16, -3, 27, 4, -20, 0, -5, 20, -2, 0, -8, -7, 25, 3, -12, 26, 9, -11, 0, -5, -22, -8, -8, -2, -5, -19, -7, 29, 15, 0, -10, 11, 11, -10, 0, -26, -7, -5, 25, -11, 3, 17, 4, 3, -17, 20, 9, 12, -2, -18, 4, -10, -20, -4, 7, -1, -6, 0, 18, -4, 2, 7, -3, -9, -8, 0, -17, -19, 12, -13, 10, 29, 24, -11, 0, -13, 29, -6, -11, 0, -19, 8, 9, 29, -24, 1, -8, -41, -1, -1, 18, 9, 17, 3, 0, 2, -2, -24, -3, 12, -14, 6, -46, -4, -4, 9, 6, 10, 6, 8, 34, -21, 20, -4, -9, -14, 6, 7, 15, 3, -11, -10, -2, -17, -8, 16, 3, -11, -26, 28, -9, 27, -4, -5, 13, 7, -20, 12, -4, -4, 16, 1, -1, 35, 8, 0, -21, -18, -1, 12, -13, 7, 15, 0, 1, -10, 18, -5, -31, 18, -25, 10, 16, -10, 3, -18, -2, -22, -6, -7, 20, 24, 19, 18, -22, -6, 2, -2, -15, 2, -12, 12, -16, -8, -10, 10, 16, 15, 15, 5, 0, -11, 1, -7, 1, -4, 10, -6, 2, 0, 3, 0, 9, 2, -12, -11, 17, 11, -4, -9, -6, 12, -2, -2, 6, 11, -3, -9, -2, 1, 7, 1, -1, 1, -8, 28, -17, 3, 14, -8, -3, -10, 19, -9, -13, 16, 0, 26, 7, -5, -27, -15, 1, 2, -28, -15, 13, 16, -14, 34, -1, -14, 15, -5, 20, -21, 19, 23, -18, 14, -27, -28, 21, -10, 13, -10, 22, -15, -4, -16, -8, -14, -5, -2, -3, 18, -12, 6, 3, 0, -19, 14, 17, -4, -6, -9, -8, -13, -14, 17, 21, -13, 7, -7, -8, 14, 0, -12, 9, -4, -5, -14, -12, 2, 2, 4, 2, -1, 2, -1, 4, -4, -4, -13, -32, 21, 15, 35, -12, 18, -5, -21, -5, 1, 0, 0, 0, 8, 0, 4, 4, 3, 12, -5, -15, -4, 7, -22, 27, 3, -13, 25, -12, -7, 10, 3, 17, -14, 9, 10, -17, -13, 17, -12, 6, -7, 15, 17, -13, 13, -19, -21, -2, 0, -29, -7, 3, 0, -10, 22, 2, 8, -5, 0, 0, -6, 1, 0, -4, -4, 13, -15, 1, -5, -4, 12, 10, -16, 0, 0, 4, 1, -21, -4, 19, 14, -10, -15, -5, 21, -3, 2, -6, -2, -32, -17, -12, 45, -1, 8, 8, 4, 1, 2, -1, -3, 0, -7, 3, 4, -5, 4, 21, -27, 10, 2, 6, -1, -19, 4, -21, 18, -19, -1, 4, 12, -5, 0, 0, 5, 7, 1, 11, 5, 18, 1, 5, -21, -1, 3, 4, -9, -10, 17, -14, 27, -23, 17, -15, 17, -10, -7, -5, 2, -11, -13, -13, 6, 30, 8, -15, 12, 21, -2, -6, -4, -15, -14, -3, 1, 6, 7, -1, 2, 20, 19, -9, 36, -25, -31, 5, -11, -5, -1, -17, -3, 21, 11, -18, 18, -9, 0, 10, -6, 0, 4, 0, -2, 5, 0, -12, 9, 11, -4, 4, -14, -1, 2, -18, 8, 8, 4, 0, 5, 6, 0, 4, 6, -6, 0, 2, 4, 7, -1, 5, -1, 9, -1, 0, 4, -2, -4, -5, -3, -10, -6, 5, -3, -5, 0, 5, 14, -10, 11, -7, 0, -8, -2, -18, 0, 18, 10, -7, 17, -11, 6, 0, 4, 21, -7, 0, -10, -9, -11, -7, -1, -4, 20, -33, 38, 9, -2, -10, -3, -12, 0, -12, 17, 1, 1, 6, 7, 3, -5, -7, 14, -17, 5, 6, 0, 4, -11, -7, -19, -3, 23, -21, 31, -11, 9, 10, -8, -3, 5, -6, -1, 1, 10, 1, 0, 5, 2, -3, -7, 8, -25, 17, 0, -7, 10, -1, 1, -3, -4, -10, -4, -2, 19, 5, -2, 5, -2, -7, -16, -24, 7, -12, 27, 16, -14, -3, 20, 24, 20, -2, 27, -19, -6, 2, -4, -31, -26, -13, -4, 2, 6, -25, 20, 10, 6, -4, 14, -2, -6, -14, 19, -3, 34, 1, -18, -2, -7, -30, 9, 1, 5, -13, -2, 0, 1, 25, 12, -18, -3, 10, 29, 11, 1, -12, 4, -11, -18, -15, 15, 2, 24, -4, -14, 14, -26, 15, -9, -9, 15, 15, -37, 27, 14, 8, -7, -18, -17, -14, -20, -16, 10, 4, 0, 8, 3, 31, -3, -13, 0, -16, -2, -6, 27, -20, 22, 5, -9, -20, 10, -9, -13, 9, 15, 9, 13, -9, -6, 11, 2, 17, 4, 0, -10, -6, -4, 1, -13, -5, 3, 22, 8, 0, -20, -5, 0, 4, 0, 31, -10, -6, -9, 3, 15, -36, 12, 21, -23, -3, -5, 2, 11, 0, -9, 6, 2, 2, -2, -36, -13, -2, 13, 32, 22, 5, 15, -13, -29, 3, -1, -1, 11, 2, 3, -7, -7, 0, -3, 8, -7, -6, 17, 4, -1, -7, -3, -6, -7, 16, -11, 29, -1, 17, 14, 19, -44, -30, -2, -9, 14, -2, 10, -4, -29, 27, -28, 21, 1, -13, -13, 3, -3, 9, 3, -5, 3, 7, 6, 16, -9, 27, -29, 10, -7, -16, 19, -11, -20, 26, 10, 12, -3, 1, -19, -1, -19, 25, -19, -4, -10, 3, -3, 4, 16, -5, 0, 0, 0, 2, 3, 4, -1, -5, -14, 8, 0, -11, -2, -19, 8, 5, -19, 1, 23, -17, 33, 11, -13, -11, -6, 11, 23, 6, 6, -8, -18, -11, 22, 0, -4, -8, -11, -9, 20, 4, -6, -9, 7, 14, -15, 1, 8, -5, -14, -16, -18, 21, 0, 0, 15, 28, -23, -26, 9, -13, 16,
    -- filter=0 channel=2
    -3, -3, 33, 4, -9, 6, -7, -18, 2, 7, -16, -1, 4, -32, 17, 20, -17, 3, 33, -20, 3, 0, 1, -1, 7, 5, 2, -16, -14, 22, -8, -10, -10, -8, 14, 7, -1, 11, -8, -3, -5, -1, 5, -1, 3, -1, 0, 0, -6, -7, 1, 2, 7, 1, 11, -8, 5, -11, -13, 3, 11, -5, 13, 0, 4, -15, -6, -7, -15, 14, -2, 19, -9, 33, 0, -38, 25, 25, -11, 14, -21, -7, -17, 8, -14, 13, 5, 2, 20, -25, -9, -2, -8, 13, 1, -5, -8, -9, -6, 9, 7, 5, 21, 17, 17, 8, -13, -4, -23, 17, -17, -23, 15, -20, 1, -1, -8, -6, 7, -14, 18, 3, -3, -2, -1, -3, -9, 1, -4, 8, -1, -5, -15, 3, -16, 34, -13, 45, 20, -20, -35, -13, -52, -22, 3, 12, 23, 12, 11, 36, 11, -10, 0, 8, -15, 2, 1, 14, 3, -3, -6, 0, -24, -10, -3, -2, -14, -6, 21, 23, 13, 5, -21, 26, 24, -5, 21, 0, -1, -20, -10, -4, 8, -30, 16, 9, 6, 20, 6, 3, -19, -10, -6, -2, 19, 4, -13, -9, 8, -6, -3, -1, 0, -3, -1, -4, 6, -6, -5, 5, -7, 14, -19, -3, 18, -16, 20, 13, -7, -35, 12, 22, -3, -7, 0, -6, 7, 9, -2, 0, 5, -3, -9, 3, -5, 7, 13, -9, -3, -8, 2, 3, 14, 2, -6, 1, -11, 12, -16, 19, -23, 18, 0, -1, 6, -2, 14, -21, 34, -11, -3, -12, 16, -13, -24, -10, -5, -8, 5, 19, -7, 29, 6, 17, 14, 8, 4, -14, -10, -27, -6, 3, -1, -4, 4, 4, 0, 0, -3, -3, -3, 0, -13, 3, -2, 0, 18, 0, -7, 5, 8, -8, 4, 4, 9, -47, 36, 19, -22, 20, 0, -12, -18, -4, 16, -14, 23, -11, 23, 14, -19, -12, 1, -13, 15, 12, -9, 3, 5, -14, 0, 5, 23, 26, -16, -27, 19, -17, -29, -28, 31, 29, -10, -12, 18, 14, -24, 9, -7, 2, -5, 11, -14, 3, 12, 0, 3, -1, -24, -14, 26, 2, 8, 22, -5, 5, -22, 19, -25, 1, 9, -11, 0, -1, 11, 6, -18, 2, -27, -5, 16, 24, 24, -23, 9, 9, 11, -7, -35, 22, -37, 27, 2, 3, 2, 0, -5, -9, -3, 8, -2, 1, 15, 0, 5, -9, 9, -5, 8, 21, -16, -4, 22, -17, 17, 0, 30, -5, 7, -18, -30, -18, 15, -31, -9, 17, -17, -14, 30, 10, -13, 20, -1, -9, -3, 0, 7, 3, -1, 0, -4, 5, 6, 4, 4, -15, 6, 0, 6, -6, 0, 6, -4, -3, 8, -5, -1, 5, -5, -3, 1, 3, -3, 11, -28, -6, 3, -20, -12, 7, 21, 39, 5, 3, -5, 0, -5, 0, 2, 6, 0, -5, -4, 22, -11, 0, -16, 28, -28, 6, -2, 7, 7, -9, 13, 6, -5, -11, -3, -5, 3, 2, 22, 27, -23, 10, 7, -24, -11, 4, 2, -10, 3, -2, 38, -19, 0, 0, -33, 24, 4, -17, 18, -15, 19, 6, 10, 8, 7, -15, -15, -13, 1, -20, -12, 25, 1, 14, 17, -21, 0, 2, 20, 21, -12, -8, -4, 22, -4, -19, 23, -26, -31, -5, 54, -6, 51, -14, 21, -8, -33, -31, 0, 24, 15, 0, -25, 1, -23, -18, 15, 7, -4, -1, -2, 4, 1, -5, -1, 0, -3, 2, 1, 6, -4, 2, -2, -16, -4, -3, 17, 10, 1, 13, -14, 3, 2, -12, 12, 14, 8, -8, -4, -15, -17, 16, -4, 16, 10, -3, 2, 9, -3, -5, 3, 11, 2, -6, -8, 2, -10, 21, 13, 10, 7, -2, 9, 17, -10, -26, -11, 2, 5, -7, 9, 11, -2, -23, 28, -14, -4, 0, 28, 12, 5, 3, -16, -16, 0, -36, -5, 18, -6, -27, 10, -3, -21, 29, 6, -7, 2, 22, -15, -14, -9, 9, 11, 27, -11, 8, 3, -9, 10, -5, -3, -5, 8, -12, 3, -7, 22, -13, -5, 0, 14, -29, 14, -25, 21, -4, 9, -2, 14, 2, 11, -3, -4, -12, 0, 4, -6, 1, -1, 5, -19, 14, 13, -2, 0, 1, -7, 1, 44, -14, 1, -15, 11, -19, -4, -28, 31, -19, -14, 9, -17, 0, -16, 17, 24, 14, -24, 20, 7, -26, -4, 36, -27, 57, -3, 12, -19, -24, 34, 9, -26, 1, 0, -12, -2, -28, 27, 1, -18, 1, 7, -6, 20, 0, 10, -8, 4, -15, 2, 5, 0, 8, -5, 26, -11, -9, -20, 2, -31, -15, -26, 10, -1, 21, -12, 29, 23, -6, -5, -1, -9, 3, 0, 5, -2, 5, 6, -5, -7, 5, -22, 24, 1, -3, 17, -18, 16, 7, 18, 3, -6, -8, -3, -14, 3, 0, 6, 1, -3, 24, -6, -16, -10, -16, -27, 0, 23, 11, -2, 3, -2, 10, 14, -7, -6, 2, 0, -6, 21, -1, 12, 6, -6, 19, -17, 0, -14, -17, 12, 2, -3, 9, 6, -8, -5, 13, -5, -12, -11, -4, -10, 7, 13, -6, 2, 18, 2, -6, -1, 1, -7, -7, 0, 8, 0, 2, 5, -4, 2, 21, -4, -7, -5, -4, 3, -18, 8, -6, -9, -5, 0, 3, 8, 0, 10, -20, 3, -3, 3, -5, 4, 13, -1, -9, -6, -5, 1, -1, 25, -7, -6, -12, 11, -13, 7, -16, 25, -9, 4, -1, -3, -5, 3, 12, -2, -5, 4, -4, 1, 4, 33, 1, -11, -9, -13, -10, -6, 3, -8, 5, -2, 0, 0, -12, 0, 2, 5, 9, -17, 5, 16, 9, 29, -5, -4, -5, -25, -7, -5, 10, 13, 9, -18, -2, -11, 14, -25, 11, 0, -15, -36, 0, -1, 32, -8, 12, 11, -2, 0, 0, 0, 0, 0, -1, 5, 0, 4, -5, 33, -9, -7, -22, 4, -6, 1, -10, 32, -7, 12, -6, 0, -13, 12, 7, -12, -8, 29, -22, -11, -26, -2, -8, 28, 23, 0, 8, -29, 7, 4, -9, 16, -10, -12, 0, 13, -21, 22, 9, 0, 2, -4, 0, 5, -5, -1, 4, 0, 3, -1, 2, 1, -3, -5, 0, 5, -3, 0, 2, 5, -1, -36, 19, -1, 4, -31, 36, 5, 0, -8, 21, 13, -9, -3, -23, 15, -10, 12, -23, 2, -10, -6, 19, 12, -3, -6, 0, -11, 7, 10, -23, 25, 29, -1, -9, -9, -10, -14, 13, -24, -26, 16, 11, 23, -8, 7, -25, -1, 32, 12, 0, 20, -7, -22, 22, 2, 13, -18, -7, 15, -16, -24, 0, -2, -4, 6, 19, 31, -25, 6, -3, 20, 4, -9, -15, -4, 3, 4, 0, 6, -7, 3, 1, -5, -2, -2, -6, -5, 12, 2, -6, 7, -14, 0, 16, 3, -5, -1, 9, -3, -8, -18, 10, -3, 29, -5, 10, -35, 25, -4, -7, 11, 18, -30, -24, 49, -9, -10, 8, 27, 0, -7, 5, -7, 9, -18, -20, 15, 0, 4, 4, 4, -4, -1, 0, -1, 0, -3, 0, 30, -2, 9, 27, -10, 12, 13, -11, -40, -22, -13, 4, 19, -12, 23, -20, -26, 41, -13, -8, -8, 2, 24, 18, -42, -4, 23, 4, -12, -1, -3, -11, 0, -7, -8, 10, 2, -6, -8, 20, 5, -24, -11, -7, -26, 30, 0, -6, 26, 4, -22, 15, 21, 1, -14, 31, -16, -13, -20, 24, 6, -1, 14, 10, -24, 5, 17, -11, -24, 15, -7, -20, 18, -1, 5, 0, 0, -1, -7, 0, 23, 9, -10, -21, 5, -1, -5, -21, 14, 25, 5, -13, -9, -8, 21, 4, 2, 13, -29, 11, 2, 33, -7, -5, -3, -20, -11, -6, 2, 20, -1, 1, 6, 0, 1, -8, -3, -1, 9, -2, -12, -34, -20, 10, -12, 24, -3, 5, 11, 20, 13, 19, -17, -9, 12, -2, 19, -15, 0, -5, -20, 16, 0, -20, 9, 52, 1, -3, -28, 0, -6, 33, -7, -16, -16, 25, 21, -24, -8, -3, 6, -6, -9, 0, -3, 1, 8, -3, 3, 1, 1, 3, -2, -7, 2, 0, -7, -5, 7, 10, 0, -20, 7, 14, 10, 30, -17, -22, -3, -14, 18, 0, 11, -14, -26, 19, 11, -15, -11, 6, 27, -12, 6, 21, -25, 29, 3, -28, -3, -16, -12, -14, 11, 2, 19, 10, 16, -4, -9, -1, 1, -1, -8, 14, 0, -2, -5, 3, 4, -7, 16, 3, 5, -3, -7, -22, 8, 3, 0, 0, -20, 9, 12, 4, -23, -18, 19, -4, 2, 0, -2, 1, 0, -6, -2, 3, -3, -3, 4, 0, -8, 8, -15, 0, -12, 0, 28, 14, -41, 29, -13, 18, -2, -4, 9, 4, 26, -4, -19, -7, 2, 0, -9, 26, -14, -2, 19, -13, -9, -12, 4, -5, 1, -18, -16, 16, -13, 26, 0, -8, 4, 6, 3, -1, 8, -6, -11, -8, -7, 10, -4, 7, -18, 10, 6, 2, 21, -3, -29, 10, 30, 1, 7, -16, -14, 6, 0, 10, -22, 2, -15, 4, 13, 18, -3, -13, 37, -25, -4, -18, -14, -29, 24, -19, -1, 17, 14, 7, 3, -22, -11, -1, -19, 3, 13, -10, 22, 19, -7, -9, 11, 8, 21, 1, 3, -10, -4, -10, -12, 6, 0, -9, -2, 6, 28, -10, -23, 13, -9, 1, -1, 5, -6, -22, -6, 0, 2, 14, 0, 19, -13, -1, 6, -4, 43, -31, 25, 1, -2, -8, 31, 1, -20, -19, -24, 5, 24, 9, -19, 12, 0, 0, 2, -1, -4, 3, 3, -5, -3, 0, 9, -8, 9, 7, -21, 12, 11, -7, 5, -7, 37, 0, 4, 4, -20, -8, 9, -10, -24, -7, 5, 16, 17, 9, 6, 0, -5, -35, 4, 3, -6, 14, 4, 0, 0, -23, 15, -9, -15, 10, -21, -13, -9, 0, -12, 26, -2, -13, 32, 15, -14, -24, 8, 7, 5, 23, 22, -29, 17, -29, 5, 11, 12, -2, 11, -29, 16, -21, 0, -5, 12, -9, 25, -18, -1, -11, 6, 10, 0, -11, 2, -5, 39, 4, -3, -7, -18, 2, -6, -5, 8, 1, 11, 0, 3, -6, -8, -6, 0, 9, -5, -13, -5, 0, 27, -31, 6, 11, 7, -9, 27, 0, 27, -2, -2, 9, -18, 0, -23, -14, -9, 8, -3, 8, 6, -10, 0, -3, 3, -2, 15, -21, 33, 11, 10, 2, -20, -15, 20, -26, 18, 5, -6, 15, -22, 22, 12, -1, -12, -27, 0, -26, -5, 26, 24, 33, 12, -3, -23, -34, 2, -9, -2, 0, -4, 1, 1, 1, 4, 1, 2, 3, -2, -9, -2, 7, 9, 3, 4, 0, 6, -2, -16, 0, 1, 5, 0, 3, -2, -2, 4, 11, 3, -1, -1, -7, -9, 0, -9, 0, 14, -10, 1, -8, -9, 0, -2, -8, 28, -18, -5, -8, 5, 17, -13, -10, 13, 14, 1, -12, -25, 34, -10, 34, -11, -7, 18, -18, 2, -21, -1, 8, 8, 4, -7, -11, -5, -6, 8, 1, 11, -11, 16, -31, -3, -9, 34, -21, 3, 15, -21, 6, -16, 12, 14, 3, -4, 2, 11, -1, 8, -3, 12, -16, 5, -9, -5, 6, -2, 0, 11, 13, 21, 8, -8, -1, 2, -30, 23, -28, -1, -6, 11, 8, -1, -1, -7, 0, -5, 0, -11, -3, -4, -22, -19, 26, -28, 26, 5, 22, 16, 8, -10, 4, -22, -6, 8, 28, -12, 0, -10, -18, -25, 2, 11, 20, 44, 16, -29, -20, 3, 12, -15, 6, -1, 0, -20, -9, 6, 15, -12, -6, -4, 14, -6, -20, -13, 32, 10, -7, -14, 3, 8, -12, -9, -8, 0, -6, 42, -11, -4, -17, 15, -17, 17, 3, -28, 22, 0, 3, 13, 12, 2, 19, 17, -13, -31, -44, 13, -3, 32, -19, 7, -22, -4, 0, -12, 7, 37, -24, -5, -12, -2, 17, 10, 24, 8, -25, 8, -14, -12, 0, 4, -5, 25, 6, 36, 4, -32, -20, -10, 0, 41, -18, -3, 10, -38, 1, 8, 14, 4, 0, 11, 27, -5, -27, 3, -4, -13, 0, -5, -5, -3, -1, -6, -6, 3, 8, 0, 8, 27, -43, 20, -17, 24, -40, -4, 40, -30, 26, 5, 4, -3, -7, -4, -1, -10, -7, -12, 10, -8, 9, -3, 15, -9, 29, -14, 4, -8, -2, -9, -2, 6, -5, -1, 0, -6, 5, -2, 3, -4, -21, 0, 16, -3, -23, 22, 23, -18, 15, 13, -22, -2, -7, -12, 19, -13, -3, 24, 0, 2, 1, 10, 15, 7, 12, -34, 28, -19, -25, 2, -1, -2, -2, 3, -6, 4, 0, 1, 10, 0, -4, 30, 11, 4, -23, -28, 33, -12, -21, -7, -11, 1, 11, -14, 22, -23, 32, -32, 24, -8, 14, -5, 5, -19, 4, 19, -9, 2, -2, -10, 10, -15, -23, 7, 2, 22, 17, -5, 3, 1, 7, -13, 8, -33, -5, 10, 23, 8, 17, -3, 6, 5, 0, -11, -20, -9, 7, -2, 14, 18, -24, 22, -18, -17, 7, -11, 7, 12, -23, 25, -9, 5, -28, -17, -2, 1, -10, 7, 33, 15, 2, -6, -5, -18, 13, -2, -14, 37, -7, -6, 7, 3, -9, -1, -4, 0, -1, 9, -8, -16, 23, -11, -7, -20, 17, -7, 8, 8, 3, -28, -19, -6, 34, 5, 18, 4, 9, 6, -17, -12, 5, 12, 7, -6, 3, 2, -10, 7, 0, -4, -9, 21, -4, 0, -15, 19, -12, -2, -5, 51, -2, -11, 8, -6, -21, 0, -19, 17, -23, -17, -5, 19, 16, -13, -15, 2, 14, 8, -10, 16, 18, -18, -3, 0, -40, -21, -2, 27, 21, 18, 3, 8, -10, -13, 11, -2, -10, -8, -3, -5, 22, 9, 5, -30, 6, 19, -5, -20, 0, 8, -22,
    -- filter=0 channel=3
    12, -1, 11, 0, 11, 25, -22, -27, 3, 4, -5, 0, 6, 0, -6, 3, -3, 7, 0, 0, -24, 18, 26, -18, -14, -13, -7, 11, -13, 21, -14, -13, 14, 1, -19, -6, 12, 3, 0, 7, 0, 2, 9, 8, -13, -23, 14, 7, -7, 0, 8, -3, 6, -10, 0, -1, 2, 0, 25, 24, -20, -4, 32, -33, 6, 8, -17, -23, 0, 4, -4, 3, -6, 0, 0, 6, -1, -6, -14, -8, 3, 12, 17, -11, -14, -4, 7, 3, -26, -12, -11, 9, 19, 0, 29, 2, -6, -18, 1, 4, -2, -7, 6, -6, 6, 5, -9, 4, -10, -7, -36, 17, 2, -19, 7, 20, 19, 6, -25, -19, -7, 1, -18, 19, 16, 20, 4, 10, -4, -3, 0, -13, 9, 0, 3, -14, -5, 1, 1, 13, 0, -8, 3, -12, -27, -16, 25, 19, 5, -10, -5, -24, -10, -12, 43, -5, -4, 4, 34, -4, 11, -16, -5, -2, 0, -20, -4, 9, -1, -14, -18, 2, 2, 8, 13, -13, 12, 13, 13, -23, 1, 7, -4, 23, -28, -10, 8, 3, -10, -19, 31, -21, 3, 13, 24, 9, -7, -36, -2, -5, 7, 10, -1, -8, 10, 0, -1, -2, -16, -12, -1, 28, 10, -4, -22, 5, 6, 2, -20, 38, 25, -3, -35, -8, 26, -13, -24, 6, 9, -15, -10, 11, -7, 27, -15, -9, -9, 17, 20, -31, 33, 20, 19, -18, -22, 1, 11, -27, -7, 2, -5, -2, -2, 7, -31, 0, 16, 25, -6, 6, 16, -5, -3, 8, -5, 18, -30, 11, 12, 16, -5, -9, -17, 21, 2, -17, -32, 33, -17, 6, -4, -3, 2, -6, -6, 8, 19, -8, 2, -7, 14, 21, -6, 23, -29, -20, 7, -8, 1, 5, -25, 14, 27, -13, -5, -4, -6, 0, -1, 0, -1, 2, -12, -3, 11, 10, 0, 0, 17, 7, -5, -18, 16, -22, 0, 17, 11, -12, -4, -5, 2, 3, -5, -6, 2, 6, 10, 1, 17, 13, 26, -24, -50, 7, -23, 31, -18, 16, -16, 0, -7, 0, 9, 24, -19, 17, -7, -20, -7, -23, -9, 27, -19, 1, -4, 0, 11, 29, 18, 25, -6, -23, 4, -4, -11, -24, -3, 28, 15, -6, 34, 33, -22, 27, -8, -27, -12, -34, -11, -15, 6, 17, -11, 6, -12, 2, 9, 2, 14, -3, 0, 17, -1, -8, -3, 9, -21, 13, -14, 0, 31, 16, -9, 21, 20, -29, -19, -19, 1, 10, -4, 20, 0, -5, -11, -2, -5, -7, 24, -30, 14, -9, 15, -4, 7, -24, 6, 2, -2, -9, 5, -8, 8, -11, -7, -2, 24, 0, 19, -25, 24, 22, 7, -9, -28, 32, -29, -9, 4, 1, 0, -5, 1, 8, -5, -4, -3, 2, 4, 5, 8, 5, -4, -4, -1, 0, 3, -6, -2, 2, -5, -2, -3, 0, 1, 3, 4, 3, -2, -15, 30, 20, -27, 11, -14, -6, 10, 13, -7, -16, 24, -22, 18, -7, 13, 27, -11, -24, -7, -5, 6, 1, -18, -13, -13, 38, 12, -3, 6, 0, -17, 10, -12, -9, 2, 16, -19, 13, 2, -1, 0, -3, -5, -3, 6, -3, -3, -3, -8, -11, -3, -16, 0, 13, 21, 5, -21, 8, -11, 12, 26, 7, 2, -31, 20, -20, -5, 11, 1, -1, 1, 0, 0, -8, 8, -3, -4, 0, 34, -7, 16, -1, -15, -11, -11, -19, 27, -14, -2, -32, 8, 23, 8, 23, -13, 17, -13, -11, -8, 1, -4, 23, -7, -23, -3, -4, 0, 23, 3, 6, 0, -4, 4, 8, -3, -10, 8, -5, 5, 11, -19, 9, -3, -5, 15, -2, 4, -14, 17, -51, 25, 15, 4, 17, 13, 11, 3, -36, 16, -9, 10, -14, -13, -10, -3, -13, 30, 11, -6, 7, -9, -11, -15, 18, -9, 23, 2, 4, -21, 15, 48, -47, -11, 5, 22, 2, -3, -18, 9, 10, 2, -18, -3, -24, 0, -12, -5, 34, 20, -8, -1, 4, 2, -9, -8, -2, -17, -2, 14, 10, -5, 16, 15, 20, -36, -19, 8, -14, -16, 0, 3, -10, -8, 9, 2, -3, 4, 15, 0, -1, -3, -2, -5, 5, 0, -1, 8, 5, 21, 0, -42, 0, -1, -20, 1, -6, 18, 23, 21, -3, 12, -2, 0, -20, -10, 3, 10, -12, 2, 27, 14, -3, -15, 2, -8, -5, -39, 17, 6, 7, 0, -4, 0, -4, -2, 2, -1, -1, 17, 0, 14, -23, -9, 1, 10, -19, 1, 4, 12, -1, 3, -12, -3, 2, 4, -17, 13, -2, -9, 5, 10, -5, 1, -2, -2, 5, 6, 0, -9, -5, -14, -16, 11, 13, 33, -2, -2, -7, -20, 9, -9, -6, 8, -20, 32, -18, 8, -9, -3, 8, -2, 9, -3, 11, -11, 1, 0, -1, 13, -20, 4, -1, 10, -10, 37, -21, -4, 10, 13, -9, -14, -3, 0, 1, -7, 11, -7, -9, 8, 0, 8, 11, -1, -18, 8, -7, -16, 2, -9, 5, -4, 9, 2, -3, -9, -2, 0, -11, -11, 14, -14, -5, 12, 8, 3, -26, 8, 6, 1, -3, 0, -2, 2, -1, 3, -6, 19, -5, 0, 25, 8, -9, -29, -12, 6, 11, 8, -9, 3, -6, 4, -25, 0, 3, 2, 2, 10, 4, -4, -17, -12, 12, -3, 19, -7, -4, -4, 8, 18, -14, 12, -7, -11, -10, 7, -8, 20, 4, 24, -4, -12, 0, 7, -9, -14, 12, -8, 0, -8, -4, 4, -4, -5, 0, -1, -1, 8, 1, -25, -1, -6, 8, 5, 29, 10, 15, -14, -26, 2, 7, -1, -3, -3, 0, 3, 0, 2, -6, 2, -27, 1, 18, 0, -11, 4, -7, 25, -10, 12, -11, 2, -14, 5, 2, 13, 1, 13, -16, 27, -2, 9, 2, -7, -12, 3, 0, -27, -5, 3, -18, 15, 3, -25, 6, 2, -8, 28, -3, 26, 25, -10, 9, -2, -19, -9, 15, -17, -8, -16, 19, -6, 10, 26, -12, 14, -22, 11, -12, 18, 16, 11, 16, -21, 2, -13, -11, 2, -21, -6, -14, -12, 32, 0, 21, 38, -29, -27, -12, 3, 12, -16, -4, 13, 5, 5, 5, 6, -19, -10, 11, 12, -19, 0, 19, -1, -8, -8, 2, -9, 30, -5, 3, -14, 19, -11, -24, 18, 3, 14, -3, 0, 15, 0, -9, -28, 9, 28, -17, -6, 2, 14, -1, -10, 0, 3, -5, 7, 0, -5, -20, 18, -31, 26, 0, 18, 14, -12, -15, 3, -3, -2, 0, -5, 9, 0, -2, 1, -5, 14, -11, 6, -13, 2, -5, -2, 0, 13, -4, 5, 15, -1, -25, -2, -16, 0, -8, 16, 25, -9, 12, 0, -2, -7, -17, 0, -7, 22, 16, 9, 12, -12, -10, 1, -11, -1, -7, 11, 15, -4, -1, -5, 4, 8, -10, 2, 1, 9, -3, -7, -4, 12, 0, -23, 0, -9, 14, 14, 4, 0, -4, -17, -21, 5, 17, 1, 5, 10, -7, 5, 7, 1, -12, 6, 13, 1, 9, 2, -23, 4, 11, -2, 3, -1, 2, 0, 0, -7, -8, -20, -4, -20, 0, 15, 0, 17, 28, -3, -19, 2, 5, 9, -1, -3, 0, 10, -16, -2, 8, -14, -12, -9, 0, 6, 30, -21, 10, 3, 0, -11, 19, -4, 15, -18, -33, -22, 14, -8, 42, 0, 0, 0, 2, 3, -3, -13, 3, 0, 0, 2, 3, 17, -2, -3, -13, 0, 4, -4, -1, -14, -9, 31, -4, 17, -17, 30, 4, 0, -28, 4, 1, 0, -2, -1, 3, -1, 1, 5, 2, -8, 9, 6, -14, -23, 18, -18, 30, -13, 4, -3, 13, 0, 12, -12, 6, -20, 16, -7, 6, 26, 0, 3, -1, -13, -9, -6, 18, 20, -29, -11, -13, -25, 0, 8, 15, -4, 29, -6, -9, 16, 2, -6, 0, -1, 4, -5, -2, -13, 12, -9, -2, -4, 10, 4, 11, -8, -11, -5, -1, -13, -26, 22, 18, -10, 8, -29, 5, 15, 9, -1, -4, 1, 3, 3, 2, 0, -4, 0, 1, -25, -14, 24, -9, 15, -9, 38, -29, 8, 7, -16, -12, 17, -4, 12, -5, 6, -26, 38, -12, 19, -1, 4, -11, -15, -2, -5, -18, 37, -11, 13, 2, 24, -14, 11, 6, -8, -29, 7, -10, 1, 26, -10, -14, -28, -12, 13, 3, 15, 5, 17, -16, 18, 0, -11, -12, 0, 26, -18, 2, -7, 5, -3, 22, -8, 6, -1, -9, 15, -12, 0, 0, -15, 9, 7, -2, -28, -8, 13, 27, -3, -10, 19, 7, -4, -23, 35, -13, -8, -2, 4, 5, 8, 0, 11, 0, 5, -17, 3, 8, 1, -23, 14, -15, 24, -21, 0, -10, 8, 7, -6, -2, -1, -24, 18, 5, 21, 18, -2, -18, -10, -6, -7, 15, 7, 28, -8, -7, 4, -6, -40, 25, -6, 0, 17, 27, 9, 3, -4, -28, 1, 4, -9, 6, 6, 3, 5, 2, -1, -4, 0, 0, -13, -6, 4, 4, -20, 32, 2, 0, -4, 0, 5, 24, -23, -12, 11, -21, 15, -1, 22, 20, -11, -3, -27, 3, -12, -17, 21, -17, 5, -5, -9, -5, 26, -13, 20, 0, -13, -9, 33, 5, -24, -11, 6, -5, -14, -27, 20, 8, 2, 2, 8, -7, -2, 4, -6, -1, -10, 7, 13, 26, 14, -17, -14, -12, 3, -7, 7, -9, -14, -27, 15, 15, -8, 17, -15, 9, 0, 15, -1, 34, -9, -21, -12, 0, -14, -7, 20, -5, -7, 0, 1, -4, -5, 13, 0, -11, 4, -6, -7, 2, -8, -14, 2, 26, -4, 0, -7, 6, -5, -10, -22, 10, 2, 31, -40, 36, -8, -6, -3, 0, -32, 14, 21, 2, -16, 13, -22, 16, 37, -1, -5, 14, -3, -10, 2, 0, -29, -5, 13, 17, -8, -1, -8, 4, 4, -7, -14, 0, 3, 6, -4, 1, -2, 0, 5, -6, 7, -6, -13, -6, -20, 18, -15, 23, -8, -25, 25, 16, 0, 22, -4, -8, -4, 10, 5, 15, -19, -13, -4, 9, 6, -4, 5, 0, 7, -1, 2, -1, 13, 4, 6, -11, 2, 7, -1, -8, -4, -3, 19, -3, -1, -2, 1, 10, -4, 1, -20, 0, -1, -4, 0, 25, -3, 13, -11, 11, -1, -21, 4, 1, 2, 2, 2, 2, 1, 2, 3, 6, 0, -9, 6, -2, -4, -8, -4, 6, 0, 0, -4, 0, -14, 3, 12, -3, -6, 1, 4, 12, -6, -12, 0, -8, -6, 10, -2, -17, 15, -2, -17, -4, 22, 3, 8, 6, -10, -13, 5, 0, -13, 13, 1, -4, -3, 3, 9, 6, -13, -11, 19, -4, -3, -9, -4, 5, 9, -4, -2, -7, 14, 2, -16, 11, 8, -14, 0, 19, -21, 14, 29, 36, -27, -23, 3, -27, -31, -19, 20, 36, 3, 26, -20, 3, -14, -14, -22, -16, 28, 30, -3, 23, -7, -9, 8, -23, -12, 0, 0, 18, 1, -5, 3, 0, -2, 2, 1, 2, -5, -5, 12, 7, 9, -3, 10, 9, -4, -15, -10, -13, -9, -18, 21, 5, -27, -13, -2, -2, -2, 33, 8, -13, -18, 16, 2, 4, -19, 6, 16, -5, -14, 26, 0, 27, -19, -8, 7, -3, -26, 2, 1, 6, -5, 7, -18, -4, -13, 6, -7, 30, 4, 2, 2, 19, 33, -20, -28, 5, -13, -12, 16, 16, -6, -28, -22, 28, -2, 3, 16, -24, 0, 10, -1, 6, 0, -4, -6, -2, -3, -10, -9, -10, 40, 9, 0, 24, -13, -27, 0, -11, 3, 2, -5, 2, -6, 0, 3, 0, 2, -2, -9, 7, -11, -2, 8, 7, -10, 9, -12, 7, 1, -3, 0, 13, -22, 0, 19, -3, -21, 12, 2, -16, 35, -14, -22, 27, -6, -6, -16, 19, -19, 16, -19, -5, -16, 0, -10, 4, 27, 24, 2, -35, 20, 10, -5, 0, -24, 22, 0, 8, 22, -27, -24, 22, 4, 24, -37, -14, 17, 21, 23, 17, -16, 2, -11, -20, -13, -6, 29, -8, -32, 11, -12, 17, 2, -1, -21, 10, 24, 12, -14, -8, -4, 6, 0, -13, -3, 0, 33, -9, 6, -6, -6, -6, -3, -2, 15, 8, -12, -10, -2, 0, -7, 6, 3, 3, 1, 4, -12, 5, 34, 1, -12, 14, 11, -15, -6, -9, -30, 16, 7, 5, 12, -2, -8, -11, 3, 0, 7, 0, 0, -32, 42, -8, 2, 12, 18, 4, -24, -36, -2, 10, -2, 12, 16, -15, 11, -9, -3, 7, -3, 3, 3, 1, -2, -2, -3, -2, 2, 0, -1, -29, 17, -11, 30, -27, 3, 21, -8, -8, -19, 13, -25, 0, -4, 0, 17, 20, 10, -21, -3, -11, -5, -13, 2, -10, 43, 14, -11, -4, -6, 35, -14, -13, 4, -13, 18, -9, 13, -29, 11, 4, -4, 6, 3, 5, 4, -15, -2, -4, 8, 0, 5, -18, -14, 1, 28, -1, -3, 12, -17, -23, 29, -14, 21, 25, 17, -4, -13, -24, -10, -8, 1, 0, -25, 16, 11, -9, 23, 11, 8, -4, 3, -29, 29, -14, 14, -25, 7, -3, -7, -12, 8, -14, 7, -3, -21, 3, 13, 24, 3, -13, -7, -14, 1, 2, 0, 0, 22, 8, 8, -7, 9, -7, -11, -5, 19, -5, 2, -3, 0, 3, -4, -6, 13, 10, 0, 0, -2, -3, 1, -19, 11, 21, -8, 19, -22, -10, 5, 3, -3, 0, -15, -1, 8, 5, 5, -2, 3, -8, 0, 11, 9, 4, -9, -28, 14, 8, -6, 8, -6, -1, 7, 3, -4, -5, -3, 1, 1, -1, 18, 17, -2, -4, -1, -9, -37, -18, 20, 13, -13, 8, -10, -8, -24, 23, 27, -21, 9, 5, 9, 6, -10, -7, -2, 2, 11, -7, -6, -10, 2, 6, 3, 10, -38, 8,
    -- filter=0 channel=4
    -9, 23, -47, 31, 25, 2, -7, 7, -11, -14, -2, -3, 17, 1, -8, -1, -1, -4, -15, 16, 4, -1, -3, 15, 10, -5, 3, 0, -4, 6, -25, 19, -2, -4, 21, -16, -13, 25, -16, 26, 8, -17, 14, -28, -6, 1, 16, -7, -8, -14, 9, 3, 8, 1, 2, -1, 3, 4, 0, -5, -2, 0, 0, -1, -12, 29, -6, 0, -24, 3, 23, -20, 22, -10, -6, 23, -13, 4, -5, 18, 17, -21, 0, -2, -14, 8, 14, 11, -4, -15, 2, -15, -1, 14, -12, -17, -6, 29, 0, 19, -4, -12, 10, -9, 12, 24, -14, 9, -5, -34, 2, -10, 10, 7, 13, 4, 0, 2, -3, 0, 3, -4, -9, 1, 4, -9, 1, -6, -12, -6, -5, 13, 22, 2, -36, 9, -11, 21, 4, 14, 20, -5, -27, 14, 25, 18, -9, -20, -5, -20, 2, -13, 12, 10, 1, -11, -19, 0, -9, 25, 6, 2, -7, 6, 11, -6, -15, -32, 13, 3, -17, 40, -5, 12, 21, -1, -16, -26, 0, 13, -18, 29, -18, 8, -27, 3, 6, -13, -7, 7, 14, 10, 11, -4, 20, 9, 1, -10, -30, -25, 3, 21, 23, -11, 11, -15, -3, 5, 14, 6, -28, 17, 1, -16, 1, 8, 10, -11, -12, 2, 14, -1, -6, -3, -18, -3, -10, 7, 16, -5, -16, 22, 6, -2, 1, -7, -3, -1, -7, -1, -5, 26, -7, -3, 11, -13, 8, 3, -9, -16, 12, 2, -2, 0, -23, 37, 25, 8, -20, 20, -17, -5, 1, -10, -8, 6, 9, -7, 6, 2, 1, 3, 9, -10, 9, -2, -2, 1, 1, 4, 4, -6, 0, -8, 0, -1, -4, -8, 10, 15, 6, -4, -16, 16, -5, -17, 26, 6, -3, -17, -5, 2, -3, -4, 9, 8, 3, 9, 5, 6, 2, -19, -10, 10, 6, 11, -7, -5, 7, -5, 6, 11, 0, -21, 2, -7, 6, -10, 19, -3, -4, -4, 4, 5, 0, 1, 5, 15, -6, -10, 0, 9, -5, -6, 4, -16, 5, -3, -4, 20, -36, -4, 18, 1, 16, 8, -6, -2, -34, 4, 10, 13, -26, 11, 0, -1, -8, 7, -8, -9, 15, -6, 23, -11, 23, -13, 7, 12, -9, -26, 5, 23, -18, -8, -7, -8, 18, 21, -23, 11, -16, 0, -4, 16, 18, -13, -3, 0, -2, -9, -6, -11, 26, -3, -4, 6, 6, 27, -4, -15, -7, 13, -6, -21, -3, 10, 0, -12, 6, -6, 19, -7, 0, 7, 18, -8, 8, -13, 8, -17, -16, 18, 7, 5, -7, -31, -19, 21, -9, 14, 5, 2, -9, 24, -3, -2, -10, -19, -16, -11, 23, 17, 4, 24, 5, -13, 6, 14, -22, -11, 22, -2, 3, 0, -22, -22, -4, 18, -13, 23, 43, -10, -4, -6, 6, 9, -4, 19, -13, -29, -14, 9, 12, 2, 6, -17, 13, -23, -14, 27, -6, 13, 3, 0, 37, -8, 17, 1, -12, 37, 12, -39, -21, -23, -3, -7, -3, 1, 3, -3, 2, 1, 2, 0, -6, 5, 3, 1, -10, 25, -8, 4, -27, 14, 6, -8, 0, 7, -3, 1, -31, -4, 9, 15, -1, -2, -1, 0, 3, 0, -3, 0, 2, 0, 12, 8, -7, 3, 22, 10, 2, -20, -10, -15, 12, 9, -14, 1, 1, -19, 14, -30, 19, -2, 3, 6, 0, -5, 3, -4, 3, 5, 0, -7, -4, 16, 8, -10, 16, 11, -32, -20, -12, 29, -5, 2, -11, -12, -15, 25, 54, -23, -22, 7, 2, -19, 17, 20, 14, 0, 0, -7, 0, -29, -3, -13, -11, -14, 8, 8, 5, 18, 0, -7, 0, 20, -21, -12, -4, -7, 19, 6, 19, -12, 14, -17, -15, 4, 8, -22, 9, 0, 8, 9, -26, -10, -5, 3, 13, 8, 29, 7, -23, 13, -30, 5, 3, 21, -15, 3, 6, -6, 21, 1, -30, 0, 11, -3, 30, -9, 14, -8, -32, 11, 10, -17, -5, -11, 33, 3, -12, 24, -30, -5, 32, 2, 13, 0, -3, -25, -5, 11, 5, -31, -11, -20, 7, -6, 2, 14, -24, 32, -4, 10, -4, -6, -10, -2, 1, 6, 9, -13, 4, 16, -6, -9, 14, -18, -7, 0, 34, -1, -13, -4, 10, -19, -3, 5, -24, -19, 16, 26, 10, 10, 0, 12, -4, 8, -11, 1, 2, -9, 14, -18, -11, 17, 1, 1, -14, -13, -4, 9, 0, 11, -8, -11, -14, 7, 10, -18, -15, -3, 18, 38, -6, -4, 6, 3, 1, 3, -5, -1, 4, -7, -8, 7, 6, -16, 0, -7, 25, -12, 3, -4, 4, -11, 8, 8, -4, 26, -23, -9, 10, -1, 6, -2, 2, -4, 0, -3, 2, -5, 12, 6, -4, 0, 0, 15, -21, -1, -29, 6, 5, 28, -16, -11, 29, 29, 38, -33, 10, -28, -5, -14, -1, -14, -6, 5, -12, -2, 13, 25, -22, 22, 0, -14, 29, -14, -7, -1, -11, 39, 4, -29, 10, -4, -1, -1, 9, 21, -17, -1, 9, -17, -1, 8, -14, 14, 13, -6, -12, 4, -9, 8, 6, -6, -22, 8, 3, 7, -32, 33, -2, 8, -5, -4, 32, 2, 0, -4, -9, 5, 0, -1, -3, 13, 0, 1, -3, -6, -1, 4, 5, -14, 2, 18, -9, -3, 32, 0, 1, -35, -3, 21, 41, -32, 1, -21, -4, 16, 0, -15, 19, -19, -10, 13, -7, 10, -25, 27, 1, -23, -13, 26, 0, -16, -1, 3, 4, 10, 6, -20, -4, 12, 0, 0, 6, -6, 6, 6, 0, -6, -5, 0, -10, -7, 0, 16, -3, -18, -2, 5, 17, -6, -17, -12, 22, 3, 0, 8, -4, -15, 0, -1, -1, -4, -8, -20, 17, -1, 22, 4, 9, -1, -14, -4, -11, -5, -9, 11, 3, -20, 0, 35, 6, -25, 23, -10, -8, 0, 8, 0, -9, 8, -15, -28, -12, 3, 33, -33, 58, 10, -15, 8, 2, 7, 5, -14, 12, 0, 0, 0, 4, -15, -8, 9, 4, 6, 0, -6, -6, 2, 6, -11, 25, -18, 23, -16, 0, -1, -1, -26, 2, 19, 7, -2, -5, 0, 7, 1, 0, 5, 0, 2, 4, 5, 12, 25, -21, 10, -17, -23, 6, 3, -1, -3, 7, -10, 1, -1, 12, 4, -3, -11, -7, 0, -4, -9, 8, 10, 0, 1, 11, 4, -1, -11, 11, 2, 10, -10, 34, -11, -13, -21, 16, -8, 0, 31, -19, 34, -24, -20, -9, -11, 21, -30, 30, 0, 13, -5, -4, -9, 8, -8, 9, 13, -19, -21, 3, 17, -20, -2, 14, 12, -5, -16, 40, 19, 31, -16, 0, -14, -23, -27, 5, 4, 0, -5, 11, 3, 3, 0, 4, 0, 7, 13, -15, -8, 2, 0, 0, 0, 4, 2, -7, 23, 24, -21, -7, -8, 6, -12, -1, -5, -7, -17, 3, 20, 2, -22, -9, 23, -8, 17, 0, -8, 6, 0, 2, -21, -10, 22, 18, -22, -10, -16, 6, -5, 1, -8, 26, 12, -11, 11, 3, -22, 14, 6, 5, 14, 24, 6, -29, -34, 34, -2, -10, 5, -18, -4, -6, -15, 20, -4, 15, 1, -14, 2, -8, -16, -10, -17, 26, 16, 0, -2, -8, 11, 1, 1, -7, -2, 4, 6, -8, -37, -1, 6, -30, 14, -9, 4, 30, 38, -22, -5, 12, 0, 1, 13, -23, 15, -1, -3, 23, -10, 12, -23, -13, 1, 4, -25, 47, -17, 0, 9, 2, 6, -15, -15, 17, -5, 2, 2, -1, 4, -4, -8, 1, 7, 4, 4, 1, -4, 7, -5, -3, -11, -10, 22, -2, 13, -14, 0, -14, -4, -1, -15, -13, -14, 0, 12, 6, 24, 0, 7, 1, -14, -2, 0, -21, 4, 6, -4, 0, -20, 35, -21, -1, 16, 16, -33, -2, 1, -6, -1, 19, -16, -18, 29, -1, -28, 4, 5, -12, -2, 17, 1, 0, -7, -4, -5, 2, -1, -14, -2, -6, 13, 29, 3, 8, -5, -6, -17, -4, -2, -14, 7, 12, 11, -3, -1, -8, 0, -5, 1, -20, 4, -4, 2, 15, 7, 2, -14, -9, -11, 26, 0, 20, 2, -31, 3, 3, -9, 3, -11, -14, -5, -2, 19, -7, -1, 22, 1, -13, -11, 6, 8, -5, -1, 4, 13, 2, 3, -10, -14, -18, 3, 11, -15, -14, 26, 29, -3, 7, -1, 9, -5, 37, -20, -5, -22, 24, -28, -14, 29, 18, 10, -15, -14, -11, -1, -12, 0, -17, -5, 29, 8, -3, -27, 13, 11, -17, 3, -11, -4, -1, -7, 14, 9, 8, -2, -9, 0, 4, -1, 3, -4, 1, 11, -6, 1, 3, 0, -36, -3, 14, 13, 30, 0, -9, 8, -6, -9, 29, -20, 24, -7, 11, -10, -13, 18, 5, -23, -10, 20, -15, -23, -8, 32, 12, 2, 0, -4, 3, -10, 14, 5, 4, -9, -14, 0, 15, -9, 14, -3, -2, -21, 0, -9, 0, -13, 6, 29, -7, -22, 28, 22, -16, 14, -11, 18, -23, 7, 40, 11, -9, 1, 0, -10, -4, -22, 6, 0, -7, 4, -9, 13, 7, -1, -10, -8, 12, -12, -4, -18, -15, -2, 18, 6, 32, 10, -17, -7, -19, -13, -6, 23, 11, -8, 8, 7, 11, -13, 43, 14, -23, -10, 4, 23, -21, -29, 5, -1, -3, 1, 6, -6, 1, 3, -3, -4, 0, 0, -14, 5, 0, 2, 15, -25, 29, -9, 3, -13, -19, -1, 18, 29, -12, -34, -15, -19, 22, 15, -2, 6, -4, 7, 0, -2, -4, -8, -2, 0, 17, 3, 45, -8, 18, -15, -5, 4, -37, -22, 4, -4, 1, -6, 5, -3, 4, -1, -7, 1, 2, -12, 11, 0, 1, 0, 5, -1, 6, 8, -2, 13, 9, 18, -3, -3, 13, -19, -15, -12, 20, -9, -13, -9, 0, 6, 5, -5, 15, -7, 7, 0, -13, 8, 8, 0, -11, -9, -1, 0, 2, 35, 17, 2, -32, 1, 5, 0, -11, -18, -3, -10, 13, 0, 10, -21, -10, 18, 9, -6, 11, 31, -18, -11, -8, -13, -22, -9, 12, 16, -16, -12, -18, -5, 14, -3, 0, 18, 9, -11, 20, 6, 20, -10, -3, 31, -18, -13, -15, -6, -8, -2, -11, 36, 12, 13, -1, -19, -21, -12, -13, -20, -6, 10, 6, 1, 13, -4, 7, -12, 3, -19, -24, 0, -34, -7, 27, 24, 13, 10, 10, 2, -10, 5, -18, -9, -21, 16, 13, 2, 8, 0, -18, 4, 9, -29, -11, 6, 17, 8, 12, -12, 3, -15, 21, 2, -3, -3, -30, 15, -11, 5, 9, 2, -11, 4, 11, 13, -20, 17, 11, 14, 20, -6, 16, 1, -23, -33, -13, 8, 21, 1, 0, -14, -1, 24, -12, 9, -27, -6, 10, -15, 12, -21, 12, -32, 1, 25, -24, 12, -5, 2, 3, 6, 4, 3, -4, 0, 3, -2, 0, 2, -11, -4, -8, -2, 18, 6, -4, 6, 7, 23, 8, -21, -13, 0, 9, 10, -5, -13, -6, 8, -10, -11, -2, -9, -5, 3, 25, 11, -12, 17, -24, 23, -7, -24, 13, -3, -19, 38, 19, -25, -1, -2, 2, 6, 7, -5, 18, 4, 7, -6, 9, -8, 10, -3, -20, 14, -15, -11, -3, 0, 3, 1, -6, 0, 4, -6, 7, 3, -4, -5, -3, 2, -10, 5, -2, -7, -1, 13, 2, -5, -2, -5, -12, -8, -5, 11, 10, 11, 2, -2, -2, -9, -1, 8, 6, -1, 0, 7, -2, 9, -33, 12, 15, -28, 23, 11, 17, -16, 15, -3, 39, -17, 1, 12, -6, -30, -6, -7, -1, -15, 1, -4, 8, 3, 24, 14, -22, 1, 0, 1, 5, -4, 0, -9, 0, 8, -2, -5, -41, 5, 10, 9, 30, 16, 20, 17, -17, -40, -7, 10, -9, 27, 1, 8, 8, -48, 4, 12, 4, 2, 0, 0, -6, 3, -2, 1, -5, -2, 1, 7, -1, -1, -3, -1, -7, 3, 0, -1, -5, -7, 0, -1, 2, 0, -5, -7, -6, 2, 1, 0, -16, 17, 8, -10, 22, 2, -12, -10, -11, 7, -12, 14, -26, -2, 16, 6, 9, -4, 47, -20, -34, 37, 1, 24, 23, -14, -37, -31, -1, -1, -20, -13, -4, 1, 10, 17, -9, 18, -7, -11, 0, 43, -21, -9, 51, -30, -29, -3, 22, -3, 15, -9, 16, 32, -28, -7, -12, -8, -5, 7, 17, 0, -4, -3, 10, -7, 0, -3, 7, -7, 5, -2, -2, -22, -1, -8, 28, 9, 9, -8, -12, -6, -14, -15, 6, -20, 43, 6, 2, 8, -11, 0, 3, -13, -1, -7, 10, 4, -18, 13, 9, 8, 14, -20, 9, -13, 15, -17, -14, 15, -5, -2, -1, -9, -8, 12, 6, -10, 19, 0, 0, -35, 28, 10, 25, 5, -19, -26, 3, -2, -3, -12, 24, -34, 18, 9, 13, -4, -13, -21, -31, 22, 4, 14, 37, -7, -4, 0, 4, -21, 22, 0, -3, -10, -18, 5, 7, 3, 15, 0, 0, -4, -3, -4, 6, 2, -4, -2, -1, 7, 1, 2, -11, -7, 8, 7, 0, -8, 0, 2, -6, -4, -1, 9, -2, 1, -2, -4, 1, 17, 18, -21, 8, -4, -17, 6, -12, 1, 16, 1, -11, -15, -10, -28, 0, 0, 21, 25, -4, 1, -3, 3, -1, 3, 5, 2, 2, -5, 49, 0, 7, -5, -16, -13, 0, -39, 7, 10, -15, 40, 7, 15, -14, -31, 37, -16, -8, -15, 0, 14, 7, 17, -17, -9, -7, 0, -5, -8, -10, 15, 2, 7, -10, -11, -9, 4, 7, -11, -5, 18, 5, 22, 11, -17, -13, 9, -19, 0, 12, -1, 2, 4, -9, -6, -24, -15, 19, 18, -5, -4, 9, 2, 2, -3, -6, 1, -7, -4, 7, 2, -8, 13, -2, -3, 2, -2, -11, 0,
    -- filter=0 channel=5
    -7, 30, 4, 14, -11, -22, -13, 8, -16, 21, -4, -15, 3, 18, 27, 0, -19, -9, -10, 7, -20, 1, 22, 7, 12, 11, 23, -36, -3, -4, -10, -1, 17, 3, 17, -7, 4, -11, 2, 0, 20, 27, -18, -9, -9, -26, -16, -3, 28, 19, 6, -32, 39, -12, -9, 0, -9, 19, 0, 3, 7, 16, -17, -7, -9, -5, 0, 35, -13, 3, 6, -7, 6, 10, 6, 0, -5, -4, -4, 0, -19, -13, -5, 11, 13, 11, -8, 24, 10, -16, -4, -14, -12, 27, 19, 5, -19, 9, 11, -15, -3, 2, -1, 10, 3, -4, -8, 1, 5, 0, -24, -29, -25, -11, 14, 24, 15, 17, 19, -8, -17, -9, -35, -4, 17, 10, 10, 27, -3, 0, -5, -3, 2, -4, -10, -8, -3, 2, 12, -7, 10, -18, 13, -11, 18, -37, 14, 6, -3, 1, -19, 24, 9, 3, 3, -6, 0, -8, -16, 3, -13, 9, -2, -7, -28, -7, 16, 29, 13, -4, 4, 5, 7, 29, -14, 16, -13, -4, 4, -20, -5, -2, 18, 17, -6, -14, -6, 5, -7, -5, -10, -3, 10, -3, -1, -1, 7, 1, -5, 2, 19, -17, -10, 4, -7, -5, -3, -23, 35, -17, -4, 8, -24, 10, 34, 2, -29, 4, -5, -2, 11, 21, -16, 2, 6, -1, -22, -21, 2, 31, -1, 3, 2, 1, 3, 0, 2, 1, 3, -7, -14, 13, -5, 3, -2, 11, -19, -9, -1, 12, -8, 23, 27, 9, -9, 7, -24, -1, -12, -13, 8, -7, 11, 15, 17, -51, 20, -17, 6, -3, -1, 19, 5, -22, 24, -15, 7, -6, 14, -20, 19, 7, 0, 14, 8, -11, -11, 12, -18, 0, 0, 6, -2, 4, -8, -3, 12, -11, -14, 9, 1, 13, -4, 32, 0, 29, -3, -27, -30, -23, -27, 2, -18, 10, 14, -5, -6, 6, 12, 20, -4, -12, -21, -17, -4, 22, 20, 16, -11, 16, 19, 6, -21, -6, 1, -17, -16, 3, 5, 26, 0, -7, 1, 2, 6, -4, -9, 5, -9, 10, -6, 19, -9, -21, -5, -1, 17, -19, 8, 13, 4, 3, -4, -25, 6, 9, 19, -1, 4, -11, -10, 6, -30, 1, 0, -24, 35, 0, 36, -18, -13, 25, -15, -9, -2, -10, -18, 6, 6, 27, 5, -2, 24, 0, -15, -11, -2, 6, -3, -8, -4, -19, 29, 26, -31, -33, -9, 4, 18, 18, 11, 7, -22, 0, -12, -22, 19, -5, 11, 20, 33, -19, -5, -8, 23, -24, -34, 45, -27, 15, -15, -17, 9, -5, 30, -11, 39, -5, -19, 2, -16, -23, -5, 25, 28, 30, 16, -27, -28, -5, 0, 0, 3, 13, 3, -12, -3, 1, -1, 3, 29, -16, 5, 41, 0, 31, 7, -34, -48, -22, 7, 12, -9, 6, -17, -22, 19, 19, 5, -14, 5, -6, -3, 6, -17, -3, -7, 4, 17, -4, -10, -1, 11, -29, 8, -13, 23, 20, -3, -6, 6, -12, -8, -12, 14, -27, 7, 40, -14, 0, -6, -20, 13, 0, 2, -13, 21, -15, 2, 19, 2, -14, 21, -5, 8, -5, 15, 3, -12, -18, -16, 12, -7, 37, -15, 7, -4, -9, -6, -2, -17, -17, -3, 8, 33, 20, 15, -9, -19, -21, -3, -3, 5, 0, -13, 3, 11, -1, 4, 0, -12, -4, 12, 0, -15, 22, -19, -3, -14, 25, -10, 0, -11, -8, -5, 0, -3, 22, -1, 4, -11, 6, 9, -2, -14, 7, -2, 6, -12, 7, -1, 0, 7, -5, -20, 28, -9, 6, 2, 0, 2, 4, -1, 3, -6, -1, 2, 2, 2, 3, 18, -1, -12, 0, -6, -15, -18, 18, 1, 20, 3, -31, 14, 8, 10, -19, -18, 30, 22, -2, -4, -10, 7, -2, 12, 11, -11, -1, 8, 5, -2, 24, 5, -5, 10, -23, 9, 18, -29, 8, 2, 1, 11, 10, 1, -12, -3, 2, -1, -2, 4, -17, 32, 11, 0, -18, 3, -11, 23, -30, -1, -2, -3, 0, 6, 1, -4, 3, -4, 3, 11, 3, 5, 12, -8, -10, 2, 9, -3, -3, -12, -7, -3, -20, 18, 12, -5, -6, 8, 0, 4, -5, 0, 2, 8, 2, -4, -2, -4, 7, -7, -5, -5, -28, 33, 9, -6, 16, -11, 0, 16, -8, 4, 4, -3, -14, 14, -14, 3, 4, 0, -2, 1, 2, -7, -8, 8, -3, -2, -5, -3, -9, 5, 12, 4, 10, -14, -9, -11, 10, 0, 19, -14, 2, 8, -8, -2, 8, -8, -10, -15, 0, 3, 26, 18, -2, 52, -51, -17, -18, -4, -22, 31, -33, 3, 8, 6, -11, -1, 22, 31, -10, -8, 10, 8, 0, -2, -5, 18, -28, 6, 8, 2, -5, 3, 7, 0, -11, -2, 0, 29, 16, -18, -7, 2, -30, 4, -29, 19, 14, -8, -2, -1, 7, 8, 13, -14, -9, -8, 7, -3, -20, 23, 19, -6, 4, -13, -22, 21, -2, 17, 3, -21, 0, 30, -3, -34, 25, -8, 0, 31, 12, -5, -29, 7, 2, -1, 0, -10, -12, -1, 0, 3, -4, 0, 5, 1, 2, -4, -1, -6, -7, 19, -17, 6, 25, -4, -14, 2, -11, -17, 4, -6, -1, -1, -9, -7, 3, 33, -4, -4, -8, -1, -10, 20, -8, 18, -1, 22, -18, 1, -4, -10, -10, 7, 0, 7, -2, 6, 12, 12, 14, -7, -4, 17, -22, -17, -2, 21, -8, -4, 3, -4, 5, 16, -6, -9, -18, 10, 19, 13, 1, 6, 1, -12, 0, 7, -11, -12, 1, 5, -3, 1, 1, 1, 0, 4, 0, 6, -6, -31, -18, 5, 21, 44, 32, 14, -6, -24, -42, 0, -1, 0, 4, 2, -4, -5, 4, 3, 3, -9, 22, -8, 18, -34, -17, 3, 28, -9, -3, -6, -8, -4, -9, 15, 7, 6, -7, 5, -2, 11, 45, 3, 2, 9, -2, -15, -15, -15, -16, -22, -31, -13, 20, -22, 17, 3, 21, 18, 7, -7, 3, -2, 14, -29, 3, 18, -6, 13, 6, -6, -6, -2, -3, -3, 3, -3, 10, 6, 4, 19, 3, 3, 0, -4, -7, -12, -9, -8, 7, -21, 37, 15, -10, -19, -12, 14, -4, -5, 2, 17, 28, 17, 4, -8, -25, -30, 16, -29, 7, 14, -12, -11, 15, 5, -3, -6, 0, 0, 18, -5, 0, -3, -11, 8, 8, -5, 10, 0, -4, -2, 12, 23, 7, 5, -9, -4, -14, -23, 12, 0, -8, -4, 2, -1, 6, 1, 0, -3, 1, 1, 2, -8, 7, -4, 5, 1, -6, -2, 2, 11, -17, 3, 9, 14, -16, -18, 5, 11, -20, 26, -24, 7, 18, -41, 10, 6, -16, 1, 9, -20, 22, -11, 20, 22, -20, 16, -21, 3, -10, -14, 25, 0, 17, -4, -13, -21, -6, -14, 14, -5, -1, -3, 3, -1, 1, -5, 6, 1, 3, -28, 33, 9, -35, -15, -7, 14, 11, -6, 30, -8, -8, -3, -10, 1, 0, 5, 0, 2, 9, -19, -10, 10, 11, 0, 16, 9, -7, 5, -11, 1, -2, -3, 0, 6, -5, -8, -6, -6, 1, 21, -11, 14, 2, 1, -29, -7, 3, 2, 2, -25, 6, 0, -6, 4, 0, -19, -1, 22, 5, 12, 21, -2, -18, -13, -4, 0, -11, -11, 27, -8, 22, 0, -23, -5, 25, 1, -16, -14, 15, -4, 7, -8, -4, -5, 4, 1, 11, 5, -7, 25, -2, 2, -24, 16, 7, -5, 25, -18, -18, 0, -7, 27, 5, -6, 12, 20, -6, -34, 9, 20, -11, 15, 11, -14, 20, 9, 3, -17, -29, -6, -6, -9, 6, 0, 17, -16, -17, 14, 20, 6, -20, 2, 0, -4, 28, 2, -21, -15, 14, 28, -27, -5, -13, -8, -5, 4, -14, 36, 6, -17, 16, 5, 16, -22, 10, 33, -22, -17, -5, -25, 10, -2, 0, 2, -7, -7, 5, 31, 6, 18, -29, 30, 10, 1, -15, -31, 13, -5, 0, 29, -8, -9, 0, 6, -13, -7, 1, -13, 3, -1, 29, 2, 1, -1, 0, -1, 1, -6, -14, -16, -12, 7, -22, 33, -13, 42, -16, 0, -6, -1, -3, -1, -7, -5, 2, 4, 1, -3, 7, 43, -11, -14, -13, -7, 7, -7, -15, 29, -9, -17, -3, -39, 9, -9, -21, 0, 36, 15, 29, 2, -12, 1, -6, -8, 3, 9, 3, 3, -3, 27, 0, 1, 5, -1, -16, -4, 0, -7, -3, -11, -2, -26, 10, 43, 5, -4, -23, 19, -13, -8, -12, -29, 31, -21, 38, 26, 0, -7, -15, -12, -8, 6, 14, -9, 1, -16, 12, 9, -10, 6, -2, 18, 6, -1, 21, -24, 29, -16, -33, 9, 29, 1, -11, -18, -5, 0, 1, 18, -24, 0, 5, 1, 1, 1, 1, 0, -2, -2, -6, -4, -2, -9, 9, 19, -13, -1, -5, 7, -8, -8, -17, 11, 10, 4, -23, 7, 16, 4, -6, 7, -10, -10, 24, -35, 14, 30, 0, -11, -10, 3, 0, 25, -21, 18, -9, 19, -18, -11, 2, -12, 4, -13, 11, -32, 27, 23, -11, 16, -20, 20, -4, 27, -8, -10, 11, -14, 6, -4, -17, 33, 12, -16, -3, -16, -8, 17, 1, -21, -6, -14, -16, -9, 0, 20, 21, -5, -2, 19, -6, -37, 23, -3, 15, 3, 23, 5, 7, -11, -24, -4, -6, 2, -4, 12, 4, 0, 0, 1, 2, -3, 4, 5, -1, 3, 10, 2, -4, 4, -2, 3, 0, -3, -5, 3, 1, 10, 2, -8, -5, 18, 4, -17, 13, 2, -16, -6, -8, 4, 0, 10, 3, -9, 9, 0, 14, -9, -7, -4, 9, -21, -15, -13, 18, -11, 24, -2, 7, 9, 8, -1, 1, -17, -14, -24, 10, 21, 22, -11, 10, 2, -6, -21, -11, 1, 18, -1, 36, -2, -8, 5, 2, -3, -7, -4, 0, -1, 2, 0, 5, 0, -1, -19, -15, 30, 17, -20, 26, -18, -6, -14, -13, 16, 18, 17, 27, -7, -20, -10, -8, -18, 12, -10, -6, -4, -19, 15, 15, 9, 5, 19, -9, 17, 39, 20, 16, 16, -27, -45, -35, -5, -13, 17, -5, 17, -8, 14, -16, 7, -9, -16, 5, 1, -8, 10, 14, 24, -18, -25, 26, -2, -2, 2, 4, 3, -4, 3, 2, -4, -1, -3, 0, 9, 17, 0, -5, -9, 2, 0, 0, -3, -4, -6, 2, 6, -9, 0, 3, 4, -7, -2, 1, 22, -7, -23, -11, 0, 16, 0, 5, 25, -19, 18, -13, -10, -5, 0, 16, 10, -21, 10, -38, 35, 3, 13, 2, 35, -14, -10, -37, 4, -3, 0, -13, 0, 4, 5, -14, -3, 14, 3, -1, -1, 0, 25, 0, -2, -18, 3, -2, 12, -1, 6, 1, -7, -3, -9, 17, -7, 3, 9, 17, -7, 9, -7, 0, -21, 27, 7, -16, 6, 22, -31, -28, -9, 12, 21, -12, 0, 18, 0, 0, 2, 14, 0, -2, 5, -11, 0, -3, 23, -8, -10, 0, -21, 7, 19, 18, -16, 2, -31, -8, 23, -20, -8, 26, 21, 14, -8, -19, -3, -13, 29, -4, -18, -2, -2, 19, -7, -6, -6, -6, 8, 24, 26, 13, -20, -7, -8, -27, -7, -1, -1, -10, 2, 2, 33, -3, -15, 12, -13, -32, -14, -5, 11, 8, 50, 10, -36, 19, 1, 6, 6, -8, -4, 6, -2, 0, -2, -3, 13, 2, 10, -10, 25, 11, -15, -22, -3, 6, 9, 7, 4, 4, -2, -11, 13, -19, -13, 20, 13, -31, 26, 10, -8, -17, -1, 0, 11, 6, 18, 2, 12, -8, 0, -26, 1, -19, 21, -10, 5, 2, 13, -1, -4, -1, -1, -4, -8, 5, 12, -43, 30, -17, 11, -14, 5, 26, -15, 5, -3, -4, -5, -1, 2, -5, -1, 0, 12, -6, -12, 1, 0, -3, 14, -9, -5, 21, 4, -3, 0, -18, 5, 6, -25, 10, 3, 26, 7, -18, 0, -4, 0, 4, -2, 1, 0, 7, -4, -9, 1, 7, -5, 16, 6, -6, -5, -7, -4, -4, -5, -1, -6, -6, -1, -7, -2, 2, 19, 7, -2, 3, 9, 4, 4, 0, 0, 2, 6, 0, 0, -3, -8, 3, 13, 19, -5, -2, -7, 1, 10, -9, 9, 6, -15, -7, 0, 22, -28, 8, 3, 19, -12, 15, 4, 1, -13, 9, -23, 11, -14, 3, 1, 0, 9, 29, 4, -24, 11, -20, -29, 11, 18, -15, 3, 8, 12, -26, -8, 25, -10, -9, -7, 22, -3, -1, 17, 8, 0, -14, 14, 6, 2, -11, -44, -14, 35, 23, -1, -16, 16, 17, -12, -2, 4, -9, 0, -11, 0, -15, -2, 11, 4, 14, -14, 10, 9, -42, 8, 3, -5, -7, 8, 12, -27, 21, 16, 4, -1, -16, -14, 4, 7, 10, -15, 25, -4, -1, -4, -2, 10, 26, -9, 0, 30, -20, -12, -7, -18, 0, 3, 5, -5, 14, -1, -4, -13, 1, 0, -4, 5, -5, 7, -25, 17, -5, -18, 39, -23, 8, -9, 23, -10, -1, -9, -13, -25, -3, 10, 29, -2, 0, -1, 2, -13, 5, 0, 2, -5, 1, 15, 14, 6, 0, -25, 20, -26, 18, -19, 9, -18, 3, 17, 9, 0, -18, -1, 0, 3, 15, 1, 8, 31, -22, 8, -17, -5, -6, -13, 11, 4, 10, -12, -25, 6, 1, 0, -6, -1, 23, -1, -3, 33, -3, -9, 7, -7, 4, -20, 18, 9, -10, -10, 3, 20, -11, -18, -17, 23, 6, -10, 9, -9, 0, -3, -20, -4, -6, 16, 21, -8, 8, -1, 13, -16, -6, 5, -5, -7, -1, -3, -36, 25, -17, 16, 38, 8, 29, -14, -39, 7, -6, 4, 8, 8, -14, -3, -12, -6, -5, 16, -9, 1, -6, 2, 10, -3, -4, -12, 6, 11, -11, -1, -20,
    -- filter=0 channel=6
    -26, 1, 0, 40, -20, 21, 1, -25, -18, 18, -4, 14, 8, -15, 12, 17, -8, 6, 23, -9, -2, 3, -5, -7, 10, -12, 5, 4, 9, -2, -9, 7, 2, 0, -7, -4, 7, 6, 15, 29, -6, -36, -13, 26, -20, 2, -16, 5, 12, 17, -9, -21, 3, 8, -27, 33, -8, 25, 1, -5, -13, -15, -22, -7, 4, 34, 11, 1, 28, -18, 33, -7, -26, -3, 10, -18, -6, -3, -15, 12, -1, -1, 16, -15, -2, 12, -4, 18, 2, -7, 10, -5, 0, -16, 0, 4, 5, 25, 11, -28, 10, -25, 5, -7, -17, 18, 7, 26, -23, -11, 12, -30, -26, 0, 7, 40, -8, -12, -10, 16, 12, 25, -4, 15, -37, 14, -2, -7, -4, 6, -35, 14, 14, -4, -2, 10, 19, -4, -1, -1, 12, -12, -29, 24, -8, -2, -5, 1, -1, 8, 5, -3, -4, 0, -2, -6, 4, 3, 7, -5, -8, 9, 12, 1, 9, -15, -17, -13, 7, -21, 29, 18, 0, -1, -9, 0, -19, 18, 2, 5, -6, -10, -11, -4, 0, 12, 19, 3, -13, 7, -12, -3, 12, 5, 0, -12, 6, 30, -9, -14, 9, -9, 16, -3, -13, -16, 0, 5, 4, 7, 2, -1, 2, -4, 4, -6, 30, -24, 13, -15, -26, 33, 13, -15, 17, -12, 3, -1, 2, -5, 7, -4, 0, 0, 0, 6, -1, -3, 1, 11, -3, -4, 0, 1, -5, 5, 6, -7, 5, -7, -14, -1, 23, 3, 5, -3, -28, -3, 23, -12, 6, -8, 24, -21, 22, 8, 1, -14, 0, 6, 0, -6, 21, -15, -6, 13, 2, 1, 6, -15, -18, -8, 13, 4, -12, 12, -25, -6, 18, 0, 0, 2, -10, -10, 10, 17, -1, -18, 0, -5, -2, 5, 3, 32, -20, 0, 1, 16, -4, 0, -18, 6, -22, 12, 4, 3, -3, -2, -6, -2, -3, 0, -1, 12, 0, 7, 4, 8, 0, 3, 2, -11, -7, 12, -11, 6, -17, -6, 6, -6, 1, -5, 0, 12, 10, 4, 34, -14, 1, -12, 0, 17, 8, -37, -15, -1, 10, 5, -23, -3, 6, 7, -16, 29, 0, -6, 3, 6, -4, 0, -6, 1, 2, -2, -1, -1, -12, 25, -6, -5, -4, -7, 6, -15, -4, 14, 3, -1, 7, -4, -10, 8, -4, 0, 7, -3, -8, -12, -22, 0, 28, -4, 0, 9, 7, 5, 4, -2, 3, -9, -1, 7, 6, 1, -3, 1, 8, 37, 15, -9, -33, -4, -6, 7, -14, -2, 5, -8, -9, 3, 14, -1, -5, 5, 1, 0, -8, 2, 15, -1, -11, 8, -1, -6, -2, 5, 22, 13, -18, 7, 0, -18, 3, -1, -2, -6, 3, 14, 16, -7, 5, -18, -5, -5, 2, -12, -7, -12, 6, -11, 36, 13, -19, -5, 18, -13, -11, -7, 11, 7, 0, -5, -3, -4, -4, 3, -2, -9, -6, 5, 0, 2, -7, 9, -3, 12, -6, 36, 16, -8, -27, -12, 5, -8, -1, 7, 26, -13, 1, -20, 8, 10, -18, 16, -17, 0, 1, 0, 7, 9, -4, -6, -3, 1, 5, -4, -21, 11, 14, 8, 6, -16, -2, 8, 6, 2, -28, 3, 0, -7, -11, 6, -15, 7, 6, 32, -6, -11, -4, -16, 25, 12, -12, 0, -6, 9, -17, 15, -6, 2, 5, -8, -18, -1, 12, 33, 12, -14, -11, 16, 17, -13, -18, 5, -20, 12, 0, 0, 6, -3, 7, 2, 1, 5, -3, -1, 13, 8, -27, -12, 13, -28, -7, -7, 7, 27, -14, 3, -11, 11, 17, 16, -31, 8, -3, 0, 19, 14, -16, 0, 53, -41, -31, -11, -1, 15, 18, 0, 8, 16, -23, 4, 2, -11, 1, -21, -5, -7, -12, 5, 0, 3, 8, -2, 3, 0, 10, 21, 7, 22, 9, 8, -18, -28, -16, 1, -10, 1, 30, 12, 8, -31, 21, -23, -14, -5, 3, 2, -19, 2, 19, 1, -8, 0, 5, -9, 1, -9, -14, 22, 9, -1, -10, -5, 15, -5, -15, -6, -19, 23, -17, -3, 12, 12, 12, -8, -17, 4, -6, 37, -2, 8, -24, -4, -3, 13, 2, 3, -14, 3, 7, -6, 0, 0, 13, -17, -11, -7, 12, 0, -4, -17, 2, 0, 5, 14, -5, 30, 2, -11, 12, -29, 17, -24, -1, 11, -3, -4, -2, 8, -15, -26, 50, -19, 0, -3, -1, 0, -1, -3, -1, -1, -1, -3, -4, -3, 1, 2, -3, 2, -1, -6, -6, 0, 1, -2, 9, 11, -18, 5, 25, 8, -19, -3, -4, -16, -3, 21, -5, -32, 22, 2, 8, 0, -13, -12, -13, -1, 29, 0, 9, -7, -10, -21, 4, 1, 5, 0, -14, -4, 7, 0, 7, 6, -9, 2, 17, 3, -3, -12, 3, -10, -18, 2, 14, 5, -25, 26, 9, 21, 1, -11, -2, -25, -21, 7, -1, 0, 2, -2, -2, 7, -4, 0, 2, -4, -18, -15, -25, 20, 3, 26, 21, 10, -16, -13, 8, 11, -11, -24, 2, 18, 15, 2, -12, -18, -7, 18, -8, -18, 3, -14, 7, 4, 0, 30, 9, -14, 46, -1, 15, 6, -11, -6, -3, -38, 34, 16, 2, -17, -23, -21, -6, -19, 58, -35, 5, 13, -13, -14, -13, 33, 4, -21, 6, -9, 9, 31, -22, -3, 11, -23, -10, -16, 5, 19, 22, -19, -9, -18, 25, -24, 1, 20, -29, 32, -11, -8, 2, 15, 23, -12, -8, 3, 6, -16, -12, -4, -7, 0, -7, 0, -15, 16, 8, 9, -8, 11, -10, -16, -14, -14, -8, 20, 4, 45, 2, -2, -4, 4, 0, -1, 4, -5, 0, 1, -7, 27, -20, 12, -4, -36, -29, 22, -3, 24, 4, -26, 21, -2, 14, -9, -35, 20, 26, -1, -20, 15, -2, -14, -11, -5, -6, -3, 10, 26, 0, 4, 2, 0, 1, 2, -3, -2, 1, -4, -7, 10, -4, -4, -1, -16, 2, 1, 26, 10, -12, 19, -11, -1, 10, -6, 2, -14, 0, -6, -3, 8, 0, -38, 6, -6, 19, 24, -13, -5, -13, -10, -7, 0, -17, 15, 3, 12, 14, 3, -3, 1, 1, 0, -5, 1, 15, -2, 2, -9, 8, 2, 8, 0, -24, 10, 12, 8, -4, -2, -8, -10, -6, 6, 6, -2, -3, -1, 9, -4, -3, 5, 12, 6, 11, -8, -4, -13, 6, 3, 5, 3, -15, 8, 7, -13, 10, 14, -8, -4, 0, 7, -11, -2, 43, -15, 4, -3, -6, -4, -1, -2, -3, 2, 7, -12, -7, 12, -8, 0, 10, -1, 0, -2, 10, -3, -19, 15, -18, 1, 11, -7, 43, 0, 1, -5, -8, -48, 12, 1, 5, 18, 22, 6, -12, 12, -15, -18, -22, 13, -6, 0, -11, 4, 5, -1, -2, 8, 2, -8, -15, 14, 2, 19, -15, -13, 28, -18, -9, -4, 3, 29, -8, -12, -15, -3, 7, 3, -22, 12, -18, -1, 0, -11, -1, 12, 0, 7, 3, -6, 0, -23, -12, 42, -24, 19, 5, -17, 20, -13, -15, 17, -7, 19, 0, 18, -25, -14, 4, -17, 23, 9, -20, 7, -2, -7, -16, 3, -2, -2, -1, -50, 28, 1, 6, 25, -1, 0, -23, 5, 18, 20, 1, -7, 12, -7, -40, -13, 1, 22, -6, -6, -1, 3, 4, -3, 0, 5, -3, 9, -12, -14, -15, 8, -3, 23, 8, 11, 11, -12, 10, 10, -15, 11, -3, -8, -22, 8, 19, -12, -15, 0, -20, 13, -1, 12, 11, -6, 7, -4, -6, -9, 5, -5, -39, 3, -4, 24, 15, 12, -7, 3, 8, -5, -5, 6, -3, -4, 3, 4, -6, 0, -1, 0, -1, 3, 5, -4, -4, 0, 0, 7, -4, 0, -5, -4, 13, -7, 0, -8, 30, 16, -14, -18, -12, -8, 3, -7, 3, 13, 2, -12, -14, -7, 15, 13, 24, -2, -6, -4, 1, -17, 1, 14, -15, -6, 4, 1, 12, -11, -8, -22, 33, -23, 10, -7, 0, 10, 7, -3, 8, -15, -17, 3, 22, -5, 7, 9, -4, -7, 0, 0, 0, 5, -6, -8, 11, 2, -2, -2, -4, -14, 2, -24, 0, -2, 27, 17, 7, -11, 0, 6, -16, 10, 27, -8, -42, 42, -19, -2, -2, 2, -9, 8, 15, -19, 16, 3, -9, -1, -15, 23, -3, 18, -16, 1, -26, 5, 12, -10, 18, -3, 23, -4, -34, 1, 16, -22, 35, -24, -15, -3, -7, 19, -4, -19, 15, -13, 21, -4, 11, 0, 3, 10, 4, -7, -5, -3, 0, 2, -4, -3, 1, 1, 4, -5, -7, 5, 14, -5, -6, 27, 8, -27, 6, 10, 20, -17, -4, -19, -15, -11, 0, 13, -15, -21, -10, 16, 20, 19, 11, -28, 18, 14, 11, 11, -7, -17, 9, -23, 0, -8, -5, -1, 1, -6, 1, 6, 2, 8, -4, -6, 24, 19, 13, -27, 7, -17, -2, -6, 20, 18, -12, -1, 6, -21, -12, -15, 17, -17, -11, 1, -3, 0, 3, 15, -13, 1, 4, -10, 21, -18, 0, -12, 25, -13, -35, 22, -13, 5, -21, 3, -13, 15, -17, 30, 19, -21, 0, 0, 0, 23, -7, -19, 9, 11, 2, -29, 14, -5, 25, -9, 5, -10, 12, -8, 7, -1, -18, 1, 1, -1, 4, 5, 1, -7, -3, -5, -4, 0, -8, -5, -16, 18, 0, 37, 4, -3, -2, -23, 27, 13, 37, 9, -8, 6, -28, -16, -11, -26, -1, 5, 17, -12, -2, -3, -3, -2, -7, -2, 19, -6, 9, -3, -23, 21, 6, 0, 7, -15, 14, -1, -23, -22, -9, 22, 4, -11, 13, 17, 13, 4, 8, 11, -5, 4, -24, -1, 16, -22, -8, 1, 0, 10, 3, -3, -3, -5, 3, -5, 14, -3, 0, -7, -5, 8, 11, -9, -2, -17, 22, 24, 9, 9, -36, -6, 14, -7, -29, 12, 12, 16, -29, -3, -16, 0, -38, 19, 12, 30, -3, -17, -7, -26, 30, 11, 14, 11, -12, -11, 11, -13, 15, -13, 1, -12, 5, 14, -3, -11, 2, 3, -5, 8, -10, 0, 7, 2, -2, -6, 27, -9, -1, 3, 13, -36, -5, -3, 29, -4, 7, 2, 5, 4, -4, -2, -4, 0, 3, -8, -2, -25, -12, 3, 30, 9, 14, 15, -18, -13, 6, 10, 24, -15, 21, -7, -1, -9, 6, -14, 0, 1, 7, -6, 6, -6, -4, 0, 0, -4, 10, 19, 21, -16, -17, -2, -15, -22, 29, 5, 12, -32, 12, 4, 7, -1, 21, -16, -14, 16, 1, -11, 0, -15, 20, -2, -26, 4, 8, 14, -10, 6, 2, 19, 7, 6, -23, -2, 7, -9, 7, 1, -6, 9, 0, -8, 7, -8, -4, -3, 19, -24, -3, 5, -17, 1, -6, 4, 15, 8, -20, -10, 14, -22, 17, 2, -2, -20, 9, 21, 15, 0, 15, 1, -6, -7, 4, 7, -16, 1, 0, -4, -7, 3, 0, -3, 1, 2, -2, 6, -17, -18, 3, -14, 11, -12, -14, -4, 40, 15, 10, 9, -14, -26, -19, -9, -2, -4, 37, 22, 11, 0, -7, 40, -24, 16, -20, 11, -22, 4, 7, 4, -20, 4, -11, 15, 7, -6, 6, -11, 3, 0, 5, -4, -3, 14, -2, 1, -2, -6, 1, 24, 0, 6, -1, -12, 0, -2, 20, -23, 2, 14, 15, 7, -11, -5, -13, -8, 0, -6, -5, 1, -3, 0, 2, 0, 0, 2, 4, 3, -3, -8, -15, 1, -18, -4, 0, 28, -9, 24, -11, 0, -13, 10, 15, -10, -9, 4, 10, 6, 4, 22, 13, -5, 4, -14, 12, -5, 2, -17, 13, 9, 0, 14, 1, -27, -2, -9, 14, 4, -6, -6, -6, -2, 4, 16, 1, -10, 7, 0, 1, 4, -15, 8, 0, -15, -7, 11, 3, 16, 1, 0, 12, 13, -8, 4, -12, -4, 3, -6, 15, 25, -12, -5, -17, -17, -20, 21, -2, 9, 27, -28, -15, -15, 24, -4, -6, 21, -3, 9, 5, 7, -21, 43, -7, 24, -19, -6, -21, -14, 5, -6, 18, 5, 7, -3, -1, -8, 3, 0, 0, 4, 13, -1, 3, 10, 19, -17, -7, -4, 13, -4, 0, -22, 21, 25, -4, -6, -22, -4, 2, 20, 0, -13, -22, -15, 8, 9, -13, 14, 3, 15, -20, 3, -5, -3, -7, 5, 11, 7, -11, -7, 17, 12, -13, -8, -9, 12, -5, 6, -5, 1, 11, -1, -1, 10, 1, -9, 1, 0, 3, 1, -1, -2, 1, 0, -3, 3, -2, 3, -7, 56, 0, -4, -19, -13, -20, -27, 9, 33, 0, 5, 3, -4, 1, 0, 2, -1, -3, -1, 5, -18, 2, -14, 5, 0, -20, 33, -22, 31, 1, -2, -14, -10, 0, -2, -19, -2, 15, 14, -13, -17, 23, 6, 20, 0, -15, 1, 6, -2, -2, 8, 2, -2, 2, -14, -4, 12, -6, -1, -16, -6, 0, 15, -3, 19, -31, 17, 8, -14, 14, -18, 0, 19, -13, 13, 4, -7, -11, -3, -5, -2, -4, -3, -3, 0, 5, 12, -7, 0, -7, 21, 13, 1, -18, -7, 25, -6, -27, -11, -5, 6, -2, -20, -14, 22, 0, 5, 19, -4, -33, -12, -17, -1, 15, 23, -4, 27, 5, 10, -5, -4, -6, -1, 16, -2, 6, 8, 5, -12, -2, -3, -2, -4, 0, 0, 3, 4, -5, 1, -21, -17, 2, 18, 15, 21, 14, -3, -21, 1, -8, -5, -7, 21, 0, 0, 7, -7, -12, 13, -14, 2, -1, -4, -4, -6, -18, -8, 32, 16, 10, 4, 7, 26, -14, -15, 0, -1, -24, 0, 27, 2, -4, 4, -5, 10, -7, 11, -15, -11, 5, 3, -12, 15, 22, -19, -17, 4, -6, -1, 5, -21, 15, 0, 2, 30, -9, -6, 10, -17, 8, -15, -10, 37, 0, -19, -13, 7,
    -- filter=0 channel=7
    2, 0, 3, 20, 30, -19, -11, -3, -5, 7, -30, 9, -1, -9, 1, -4, -8, -9, -8, 13, 28, -16, -10, -15, 24, -14, -6, 8, 9, -20, 0, 25, -8, -5, 4, 5, -10, 25, -27, -14, -1, 23, 0, 0, 1, -7, 0, 6, 3, 8, 0, -2, 23, -27, -6, -3, -6, 6, 14, -8, 12, 2, 42, -11, 1, -16, -8, -11, -10, -28, 30, 6, 2, -12, -12, 4, 4, 16, -13, 4, 3, 18, 24, -1, 10, 0, 24, -5, -10, 5, -9, -13, -4, 10, 4, 1, -7, 1, -14, 25, -11, -5, -1, -9, 12, -2, 0, -10, 26, -11, 1, -1, 21, 20, 30, -4, -13, 17, -12, -8, -29, -17, 0, 14, 22, -34, -14, 31, -9, 12, -12, -17, -11, 18, -32, -10, 22, -2, -6, 12, 7, -6, 16, -27, 32, -14, 9, 20, -21, -9, 2, -22, 1, -1, 0, 0, -3, 2, 2, 4, 4, 3, 0, 0, 0, -3, 5, -5, -3, 1, 0, -2, -14, 8, 18, -10, 2, 16, 0, -29, 14, -8, -11, -8, 4, 2, 8, -5, 0, 6, 9, -3, 0, 25, -23, 11, -6, -27, 0, 2, 35, -23, -34, 35, 33, -14, -12, -28, 40, -29, -2, 15, 3, -6, -10, 6, -2, -18, 16, 15, 2, 0, 6, -6, -6, -5, 1, 7, -14, 21, 6, -19, 0, -10, -6, 14, 1, -11, -7, -1, 4, 17, 4, -3, -15, 6, 10, 2, 6, -16, -5, 5, 2, 0, 3, 0, 3, -8, 2, 5, -5, 0, 18, 5, -2, 7, -10, -16, 2, 4, -11, -8, 2, 6, 0, 4, 5, 2, -6, -1, 2, 1, -13, 26, -10, -17, -14, 1, -6, -5, 17, 26, 20, -19, 30, -17, 36, -1, 4, -4, -13, -22, 9, -21, 8, -19, 2, 19, -2, -9, -10, 11, 14, 21, -20, -5, 6, -13, -11, 0, 22, -14, 11, -8, 0, -13, -23, 4, 9, 27, -23, 21, 3, -29, -4, 0, 27, -14, -6, -5, 13, 9, 21, 7, 4, 20, 4, -29, -20, 27, -14, -19, -21, 28, -7, -18, 4, 16, 4, 1, -20, 4, 12, -13, 32, -8, 13, -14, -14, -40, 28, 9, -25, 18, -14, 13, 2, -22, 31, 17, 2, -20, -1, 5, 2, -12, 11, 8, -16, 22, 7, 0, 0, 3, -6, 1, 4, 4, 1, -1, 4, -3, -4, 2, -3, -4, 4, 0, 2, -2, 2, -10, -6, 18, -10, -10, 19, 17, -21, -4, -3, 8, 1, 0, -8, 15, 3, -1, 9, -19, 22, -19, -9, 10, -9, -6, 0, -11, 0, 14, 4, 24, 9, 1, -3, -12, 1, 5, 5, 1, -5, 0, 1, 0, -1, 0, 4, -1, 1, 0, 2, 3, 0, -9, 7, -3, 4, -8, -6, 0, 22, 0, 33, 6, -4, 2, -27, -17, 6, 7, 7, -10, -2, -1, 2, 6, 2, 5, 1, -3, -3, -4, 2, 8, 5, 5, 3, 7, -14, -7, 0, -9, -15, -13, 18, -3, 5, 15, 18, 8, -9, -19, -7, 1, -2, 5, -15, 13, 0, 1, -8, 13, 8, 15, -17, 5, 5, -12, 7, -16, 1, -5, -3, -13, 23, 30, 16, -18, 31, 5, -21, -33, 0, -3, 13, -12, 10, 10, -4, -9, 3, -14, 29, 20, 16, -9, -9, -25, -8, -17, -6, -4, 11, -4, 0, 1, 2, -1, -3, 0, -6, 7, 18, -11, 9, 8, -24, 0, -4, -3, -13, 15, -2, 9, -16, -21, 5, 1, -12, 0, 22, 8, 0, 18, -3, 7, -8, 5, 14, -16, 2, -22, -20, 9, 23, 7, -5, 23, -6, -36, 0, 2, 11, 9, -3, 16, 17, -24, 0, -7, -5, -23, 26, 5, -12, -17, -21, -21, -5, -3, 35, 7, 17, -31, 36, 32, 30, -16, -32, -25, -2, -10, 2, 4, 1, 3, 3, -6, 0, 2, 0, -5, 6, -28, 14, 4, -8, 20, -4, 10, 11, -22, -14, -34, 30, 2, 6, -12, 19, 9, -13, 10, -5, -3, 1, -3, 3, -4, 2, 0, -2, -3, -7, -7, 0, -20, 8, 25, 6, 1, 0, -6, 3, 2, -3, 2, 9, -8, 0, -2, -12, -1, -23, 25, 12, -16, -23, 16, 3, -16, -14, 34, 14, -2, -20, -4, 12, -4, -11, 0, 4, 16, -16, 17, -21, 4, -10, 2, -7, -15, 23, 13, 0, -15, 28, 22, 0, 3, 4, -3, 13, -36, 19, -13, -2, 22, -17, 24, 0, -13, -20, -2, 15, -17, -2, 34, -11, 37, -6, -6, -15, -33, 29, -31, 26, 21, -19, 42, -20, 31, -31, -50, -11, 3, -15, -2, 0, 19, 0, 25, -6, -14, -5, -8, 11, -1, 7, 21, 33, -7, -22, -17, -4, 0, -7, -5, 7, 8, 6, -5, -7, 10, -1, 17, -31, -12, -4, 0, 29, -16, 14, 14, 5, 5, 3, -7, 11, -5, 1, -3, -2, -6, -10, -2, 4, 0, 0, 0, 1, 1, 1, 18, 9, 1, 3, 0, -12, -5, -15, 19, 9, 12, 29, 14, -15, -16, -24, -4, -4, -12, 29, -1, 33, -7, -1, 0, -10, -6, 2, -6, 2, -13, 4, -2, 0, 0, 1, 1, 3, -6, -5, 6, 14, -11, 11, -2, -23, 10, 10, 9, -15, 8, 1, 7, 4, 6, 8, -1, -7, 2, -16, -7, -16, 0, -14, 12, -10, -11, 3, -6, 40, -1, 8, 12, -18, -34, 29, -21, 42, -21, -5, 4, 8, -12, -2, -7, -17, 5, 12, 0, -4, 5, 2, 1, 4, -2, 3, 15, -6, -7, 3, 0, 9, 5, -9, -8, -2, -5, -2, 5, 10, -4, 15, -14, 20, 6, 18, 0, -18, -10, 2, -21, -7, 23, 19, -2, -10, -1, -10, -5, -19, -2, 23, -2, -4, -23, 16, -26, -12, -31, 30, 21, -1, 2, -8, 5, 8, -6, -12, 8, -9, 20, -3, -3, 0, 3, 10, 0, -11, -7, -13, 17, 7, 5, -8, 5, 10, -4, -11, -1, 0, -1, 20, 0, -12, 1, 9, -11, -13, -18, 10, 14, 21, 22, -29, -1, 15, -11, 0, 1, -5, -1, -9, -16, -19, 9, 10, -15, 29, 30, -2, -10, -3, 4, 3, 10, -6, -6, -4, -6, 6, -1, -11, 4, -24, -1, -15, 2, 10, -7, 17, 13, -3, -9, 2, 0, -1, -5, 0, 8, 2, -10, -8, -17, -4, 28, -17, -21, 37, -1, -17, 11, 4, -10, -7, -1, 7, 3, 0, 0, -4, -1, -18, -1, 9, 9, 12, 3, -10, -13, -3, 14, 20, -6, 12, 0, -15, -25, 5, 17, -5, -6, -3, 26, -15, 17, -2, -22, -22, 6, -14, 27, 3, 5, -1, -5, 10, -8, -4, 6, -3, 0, 11, -9, 4, -23, -4, -26, -17, 59, 7, 4, 9, -2, 0, 1, -13, -1, 12, 9, -2, -1, 5, 0, -5, -5, -1, 4, -4, -3, 2, 0, -3, 15, 0, 1, 4, -1, -11, -2, 4, -11, -12, 8, 14, 2, -9, -9, 2, 18, 3, -1, -7, -1, 13, 14, 7, 0, 11, -32, 1, -4, -4, -2, 4, 2, -1, -1, 1, -4, -4, -1, -20, 9, 14, 11, -19, 14, 40, -21, -10, -7, 0, 1, 1, 1, -3, 12, 5, -7, -9, -4, 3, 0, -15, -3, -13, -18, -21, 1, 34, 23, -2, -24, -36, 16, 3, 28, 44, -21, -12, -6, -8, 30, 9, 1, -8, 1, -19, -1, 7, -12, 14, 2, 10, 22, 10, 17, 17, -38, -34, -22, -28, 7, -32, 0, 29, 12, -10, 37, 23, -18, -14, -15, 17, 1, -28, -11, 14, 2, 35, 1, -3, 6, -13, 9, 3, -10, -7, 12, -3, -12, 13, 23, 0, 9, -14, -1, -22, -16, 12, -12, 11, -5, -30, 24, 1, 7, 22, -10, -11, -13, 9, -1, -6, -16, -6, 3, 7, 2, 4, 1, 30, 5, -3, -12, 3, 1, 0, -14, -42, 33, -6, -17, 23, 7, 14, -10, 13, -12, -12, -6, 15, -28, 29, 4, 41, -14, -3, 5, -27, -21, 14, 5, 1, -17, -5, 0, -4, 9, -15, 1, -13, 8, 9, 3, 46, 3, -23, 0, -14, -25, 0, -6, 4, 0, 5, -4, 0, -3, -1, 5, -25, -12, -14, -16, 17, 6, -10, 1, 22, 22, 5, -13, 11, 4, 13, -4, -9, -4, -15, 5, 5, -22, 7, 23, -13, 10, 10, 17, -7, -24, 13, 8, 5, -10, -18, 9, 15, 8, 7, -13, 8, -1, -3, 9, -12, -10, 24, -12, 0, -16, 30, 4, -11, 7, -5, -18, 0, 27, -43, 6, 31, -2, -16, -1, -2, 12, -3, -6, -16, 1, 21, -15, 28, 11, -23, -12, -29, 31, -15, -11, 9, 13, 19, -20, -32, 32, 6, -27, 1, 6, 3, -6, 16, -13, 12, -3, 1, 9, 8, -18, 17, -8, -9, 11, -24, 0, 9, 16, -19, -1, -16, 2, 17, 10, 1, -20, -8, 8, 6, 0, -21, -4, 0, 11, 0, 7, 1, 3, 15, -5, 9, 5, 13, -10, -6, 8, 8, -7, -14, -2, -3, -8, 1, -9, -1, -6, 6, 1, 5, 8, -7, 2, -1, -6, -4, 1, -7, 3, 1, 0, -6, -39, 22, -1, 13, 0, 0, 18, -21, 7, -27, -3, 3, 10, 1, 1, 27, 7, -9, -5, -12, -24, 0, -5, 7, 13, 19, 15, -1, -11, 9, -6, 5, 24, -17, -17, 20, -26, -18, 14, -7, -21, 22, 8, -2, 13, 1, 26, -8, -21, 0, 15, -27, 7, 36, -21, -9, 3, -12, 12, -12, -2, -14, 7, 9, -1, -4, 10, 11, -2, 2, 31, -29, -30, -14, 29, 12, -4, 28, -30, -14, -3, -1, -2, 8, 10, -2, 8, -3, 2, -30, 22, 9, 12, -20, -4, 0, -8, 10, 7, -23, -1, 2, 11, 22, -26, -4, 3, 1, 10, -2, 12, -33, 18, 16, -13, 24, -5, 2, -9, 2, -6, 4, -21, 30, 5, 22, -21, 0, -15, 14, -5, 19, -2, 1, -3, -18, 20, -16, -1, 31, 0, -11, -3, -1, -6, -3, 13, -22, 10, 0, -5, -10, -14, 19, 14, -12, -2, 3, 6, -23, -13, 22, 6, 31, 7, -1, 23, -14, -28, 10, 6, 18, -34, 16, -29, 19, 0, -4, -14, 1, 0, -11, -1, -5, -23, -11, -7, 8, 31, 9, 23, -12, -9, -18, 0, -20, -21, 15, 27, -2, -6, -16, -10, 18, 11, -4, -9, -6, 12, 2, 0, -1, 5, 0, 2, 0, 2, -3, 1, 1, 0, -3, 27, -16, -10, -8, -10, 9, -1, -6, -6, 3, 0, 3, 0, -1, 4, 4, 7, 6, 1, -1, -4, -22, -4, 14, 20, -5, 12, -8, -21, 0, 30, 8, 11, -12, 6, -4, -18, -13, -14, 4, 15, -2, 7, -6, -8, 5, 4, 5, -4, 25, -10, 25, -5, 17, -1, -14, -29, -8, 0, -3, -11, 16, -3, -14, 4, 10, 20, 10, 1, 7, -5, 10, -7, -7, -6, -18, 0, 8, -22, 1, 16, 1, -17, 11, -11, 26, -14, -43, 27, 1, 10, -11, 31, 0, -18, 5, 15, -5, 15, 12, -26, 7, -4, 33, -19, -4, -14, 11, -9, -11, 5, 10, -19, 4, -9, 26, -3, 13, -9, 11, 8, 0, -14, 10, -13, 17, -7, -23, 15, 15, 15, 10, 6, -3, -8, -3, -27, -3, 0, 16, 19, -7, -14, -6, -5, -1, 3, -10, 3, 6, 1, -3, 7, -1, 2, 8, 2, -1, 11, -4, -3, -2, -18, -5, 9, 10, 19, 0, 0, 4, -3, -6, 7, 5, 0, 4, -2, -4, 5, -7, 22, -16, 13, -33, 14, -6, 5, -1, -3, -12, -8, 9, 5, 28, 11, -11, 6, -5, 1, 3, -5, -4, 6, 7, 6, 5, -5, -7, 1, 0, 0, -1, 6, 2, 0, 11, -8, 1, 20, -10, -10, 6, -13, -13, -2, 29, -2, -6, 3, -7, -9, -6, 18, -1, 13, 11, -16, -10, -20, -5, -14, 0, 1, 34, 35, -18, -1, -10, -9, -25, 18, -16, 12, -3, -18, 26, 26, -10, 0, 36, -9, 15, 7, -17, 7, -2, -14, -12, 20, -11, 17, 22, -3, -36, 20, 12, -19, -3, 28, 0, -11, 0, -4, -26, -12, 5, 34, -14, -15, 13, 7, 3, 4, -9, 13, -10, 15, 3, 7, 30, 9, 8, -1, -2, -37, -5, 14, -17, 11, 5, 0, -5, 1, 2, -5, -7, 0, 14, -6, 9, -8, -15, 14, 9, -7, 1, 1, 30, 0, 17, 1, -11, -18, -6, 10, 0, -7, -4, -2, -3, -9, 7, -4, 0, 5, 5, -5, 8, -2, -1, 6, 1, -6, 0, -2, 1, -5, -4, 2, 15, 16, 0, -28, 19, -3, -2, -7, -15, 20, 10, -16, -7, 1, -7, -7, 8, 19, -2, -6, -28, 15, 16, 15, -10, 1, 0, -5, 6, -1, 3, 8, -7, 6, -7, -5, -6, 2, -4, 4, -12, -4, -13, 23, -10, -18, 19, -8, 3, -7, 3, 0, 18, -6, 8, -6, -2, -3, -8, -35, 15, 18, 9, 0, -15, 25, 0, -4, -5, -1, 1, 0, 1, 22, -11, -18, 0, 7, 12, -5, -20, 2, -5, 4, 2, -12, 17, 0, 12, 15, 5, -20, 31, -2, -10, -13, -14, -8, -2, -15, 18, -9, -17, 7, 24, -19, 24, -9, 0, 3, -8, -1, 6, -1, -1, 8, 0, -2, 0, 24, 2, -3, -9, -14, -19, -12, -11, 30, 5, -7, 0, 0, -1, -20, 12, 4, 5, -2, 16, 23, -30, 0, 6, -16, 21, -13, 17, -12, 19, 17, 4, -9, -3, -13, -25, -13, -1, 15, -17, 18, -15, 19, -4, -21, 21, -12, 16, 3, 3, 1, 8, 17, -10, -2, -14, 18, -5, 0, 9, 19, 11, -12, 9, 0, 10, -25, -1, -12, -13, 1,
    -- filter=0 channel=8
    18, -9, -5, 16, -7, -11, -3, -4, 3, 0, 18, -10, -16, 0, -7, 13, -12, 10, -10, -14, -10, 30, -29, -6, 26, -5, 19, -5, -11, 20, 29, -13, -54, 17, 11, 17, -17, 9, 18, -10, 0, 1, 1, -13, 6, -3, 18, -2, -2, -3, 0, 35, -7, -21, 5, 5, -24, 16, -33, 0, -7, -10, -11, 2, -4, 37, 22, -12, 5, 0, 6, 10, -9, 4, 4, -4, 7, -9, -14, 20, 9, 6, 1, 5, -17, 1, 0, 0, 20, -23, 11, -41, 13, -7, 22, 29, -18, -3, 3, 0, -4, 1, -2, 4, 3, -1, 2, -1, 7, -9, 0, 8, 13, 20, -29, 5, -14, 4, -1, 7, 0, 17, 21, -31, 11, -12, -12, -1, -3, 3, -8, -6, 6, 22, -29, 5, 3, 10, -13, 10, -4, -4, 12, 2, 21, 1, -1, -18, 8, -2, -3, -4, -3, -3, 6, -7, 13, -7, 17, -20, -5, 19, 22, -15, 13, 7, -13, -22, 3, 1, 2, 7, 0, -7, -2, 0, 0, 5, -3, 26, 12, 9, -24, 9, -2, 0, -18, 6, -3, 13, 5, 4, 0, 4, -10, -8, -15, 5, 3, -14, 2, -31, 27, -4, 25, -15, 23, -29, -3, -45, 17, -1, 25, 6, -1, 22, -17, -9, 9, -19, 12, -9, 7, 18, -12, -4, -9, -2, -2, -24, 33, 5, -25, -12, 1, -14, 11, 24, 0, 20, 13, -3, -23, 14, -2, 4, -11, -16, -11, 34, 20, -16, -18, -29, 19, -3, 1, -4, 2, -4, -1, 12, 17, -9, -4, 15, -8, -13, 5, -7, 14, 7, -27, 9, 6, -13, 1, -5, 0, -2, 0, -6, -4, 8, 0, 0, -3, 5, 8, -12, -4, -2, 11, -11, 15, -5, 8, -11, 10, 23, -5, -5, -8, -21, -21, 25, 0, 1, 4, -13, -9, 8, -12, -7, 10, 14, 9, -15, 4, 13, -7, -5, -13, 7, 17, -4, 0, -8, 13, 19, -4, -7, -18, 21, -10, 0, -1, 2, 7, -2, 12, -11, 13, 20, -20, -17, 18, -6, 10, 2, -3, -31, 16, -16, 29, -10, -1, 3, -2, -21, -17, -2, -6, 25, 17, -20, 23, 6, 7, 7, -6, 16, 21, -25, -8, -5, -5, 3, 15, 7, -22, -9, 4, -4, -4, 0, -9, 17, 11, -2, 7, 0, 12, -17, -13, 35, -28, -18, 24, 7, 12, -12, -20, -29, 1, 10, 0, 1, 24, 15, -24, -22, 0, -9, 1, -27, 34, 22, -18, -1, 39, -1, -2, -11, 27, -26, -6, 11, 2, 10, 30, -13, 13, 0, -15, 7, -17, -10, -7, 8, 10, 0, -24, -4, 24, -1, -16, 18, -15, -41, 10, 8, 8, 24, 0, 24, -24, 15, 0, -8, -3, 0, 2, 5, -1, 2, -2, 0, -23, 16, 37, 11, 5, -7, -18, -15, -15, 11, 3, -8, 7, -20, -16, 14, -7, 12, 12, 1, -2, -4, -3, 1, -16, 1, 10, 8, 3, -8, -3, 5, -1, 17, 7, 34, -20, -27, -13, 1, 5, -6, -4, 4, 6, 0, -7, -2, -1, -3, -6, -16, -6, 10, 2, -11, 15, -7, 9, 13, -9, 7, -1, -12, -26, -9, 27, -11, 10, 13, -16, -23, -8, 20, -1, 22, 10, -25, 31, 0, -2, -24, -15, -3, -4, 23, 10, -14, 16, -2, -5, -7, -7, 12, 11, -17, 27, 10, -8, 11, -9, -9, 8, 0, -8, -11, -6, 6, 7, 8, 4, -6, 4, 7, -3, -6, -5, -2, 4, -5, 20, 32, 1, -5, -19, 5, -2, -15, -16, 4, -8, 5, 7, -6, 1, -1, 3, 11, -4, -5, -27, -39, 6, 32, 13, 37, -15, 31, 9, -48, 3, -15, 28, 5, -3, -12, -14, 21, -11, -8, -21, 12, 12, -1, -20, 36, -15, -15, -7, 27, 2, -5, 0, -8, -20, 22, 16, -3, -14, 19, -4, -17, 12, 12, 13, 26, -21, -39, 23, 0, 9, -11, -3, 12, -9, 0, 11, -4, -13, 0, 5, 31, 17, -6, 2, -2, -25, -7, 6, -24, 8, 31, -24, -8, 17, -37, -26, -11, 19, 27, -8, 0, 45, -27, -9, 7, 0, -16, -12, 7, -7, -30, 11, -6, 20, -14, 24, 7, 3, -7, 1, 6, 0, 0, 1, 2, -2, -1, -7, 1, 2, 3, 13, -19, -13, -5, 16, -2, 2, 1, -18, 33, -8, 29, -10, -13, 17, -14, -12, 1, -1, -8, -1, 9, 5, -3, -2, -2, 4, -1, 0, 15, 8, -12, -8, -9, 4, 2, -2, 1, 20, 2, -15, 2, 5, -17, -3, -9, 22, -18, -9, -17, -13, 10, -9, 1, 30, 0, 1, -4, -31, 14, -4, -6, -16, -4, 21, -7, 22, 5, 12, -4, -4, 9, -1, -6, -1, -6, 4, -1, -14, 14, -1, 2, -11, 6, 1, 4, -2, 3, -3, 3, 0, -12, -4, -7, -21, -1, 14, 41, 3, 0, -1, -1, 7, 1, 0, -5, -6, 0, 8, -2, -2, 0, 3, 7, -1, 0, 5, 0, -6, 3, -18, 6, -3, 21, -3, -2, 0, 12, 0, -9, -7, 19, 0, -3, 1, 13, -22, 14, 18, 7, -17, -24, 24, 2, 1, 38, -28, -16, 4, -4, 4, 5, 1, -9, 1, 1, -3, 3, 4, 5, 4, -2, -2, 14, -5, 0, -2, -10, 12, -19, 5, 8, -20, 10, 7, -8, 22, -13, -11, -1, 16, -3, 3, 3, -13, 28, -20, 1, 0, -3, 2, 10, -6, 0, -2, 4, -5, -7, -14, 5, -19, 9, -17, 19, 3, 14, 11, -5, -5, -3, 1, 20, 7, -21, 2, -13, -8, 16, 21, 0, -1, -13, 2, -4, 6, 3, 13, -12, -29, -2, 14, 16, -41, 19, 26, 6, -5, 9, 10, -12, 15, 1, -27, -15, 5, 10, -6, 7, 0, -1, 3, -1, -3, 9, -3, 2, -6, 6, -1, 2, -32, -1, 23, -26, -1, 1, 25, 17, 9, -9, -4, 5, 6, -6, -2, -7, -17, 7, 15, 19, 0, -23, -18, -8, -31, 21, 7, 17, -12, -2, -7, 16, -26, 30, -9, -8, -14, 25, 9, 5, 0, -5, -15, 8, 2, 16, -17, -7, -14, 1, 0, 27, -14, 17, 26, -3, -6, -10, 14, -37, 13, -18, 4, -12, 23, 20, -10, -8, -1, -7, 1, -6, -4, 7, -4, -3, 3, 2, 3, 8, -3, -7, -6, -19, 21, 10, -6, -9, 1, -4, -4, 2, -8, -1, 2, 12, -2, -8, 14, -8, -9, -10, 0, -15, 11, 28, -12, 11, 7, -14, 31, 5, 6, 0, -25, 22, -17, -9, 4, -18, -6, 14, -28, 14, 9, 3, 3, 7, 12, -6, 35, -22, 14, 9, -21, -10, -20, 5, -4, 5, 2, 7, -4, -10, 1, 0, 4, -4, 10, 28, -5, -2, 1, -19, -2, -12, 27, -8, -7, -15, -9, -8, 9, -12, 31, 6, -8, -1, -13, -19, 19, 9, 16, 23, -19, -26, 0, 18, 6, -4, -2, -4, 7, -15, 38, -16, -6, 2, -5, -2, 8, -2, -2, -13, -3, 3, -6, -10, 13, -17, 3, 0, 0, -20, 4, -15, 8, 5, 10, -26, 29, 5, 13, -27, -3, -22, 15, 16, -4, -5, -3, -1, 0, 6, 6, -8, -3, 7, 8, -18, 3, -26, 25, -14, 10, -4, -6, -3, 10, -6, 11, -8, 16, -23, 25, -13, -5, -8, -3, 0, -3, -1, 4, 0, -3, 0, 0, 0, 0, -31, 32, 0, 17, 21, -9, -31, 16, -15, -4, -6, -22, 0, -1, -7, 19, 5, 16, -10, 8, -14, 0, -6, 3, 4, -6, -3, 0, 10, 7, -7, 1, 1, -12, 3, 3, 1, 3, 6, -13, 1, -21, 6, -3, -9, 20, 0, -7, 24, -6, 3, 3, 1, -2, -6, 0, 2, 6, -1, -11, 15, -10, -5, 1, 27, -29, 0, -3, 3, 17, 17, -7, -12, -6, 40, -16, 0, -41, 7, 0, -8, -8, 2, 3, -1, 17, 13, -12, 0, -3, -1, -3, -9, 4, 12, 0, -2, 5, 0, 16, -3, 10, -18, 1, 31, 14, -14, -25, -9, -2, -6, 2, -5, 11, -2, 12, -4, 6, -7, 14, 6, 22, -4, -14, -12, -23, -22, 8, 25, -1, 22, -1, 7, 22, 4, -21, -11, -2, -17, -2, -3, -8, -21, 44, -21, -12, 3, -5, 19, 6, -2, 3, -6, -6, 7, -4, -1, 1, 0, 5, -22, -28, 36, -25, 24, 29, -23, 0, 9, 0, 2, 1, -3, 4, 0, 1, -2, 0, -1, 12, -3, 19, -35, -27, 11, 29, 16, -8, -11, -6, 21, 11, 13, -19, -2, 41, -20, -13, -26, 3, -7, -13, -8, -4, 24, 15, -4, 3, -12, 2, 0, -3, 14, -1, -16, -6, 3, 7, -6, 5, 0, -6, 13, -7, 0, -4, -1, -11, 3, 13, 31, -7, 2, -16, -28, -7, 5, -17, 18, -27, -9, 6, 31, -50, -9, 29, 17, 10, 3, 0, 1, 1, 0, 9, 2, -9, 0, 7, -11, 13, -6, 0, -15, -11, 41, -35, 30, -14, 0, -15, 17, 3, -7, -2, -3, -8, 2, 3, 19, -29, 15, -23, -14, -7, 10, 8, 0, -2, 41, -25, 0, -22, -15, 38, 55, -12, -2, -23, -9, 9, -5, 10, -16, 4, 5, -4, 16, -9, -6, -4, -37, 30, 14, -4, -23, -5, -7, 15, 15, 15, -7, 0, -5, -13, 3, 28, -21, 7, -20, -2, 3, 6, 20, -25, -19, 17, 4, 4, 10, 0, 41, -12, 14, 5, -40, -23, 25, 12, -24, 16, 29, 33, -28, -24, 17, 6, 4, -30, -17, -12, -19, -5, 4, 16, -10, 6, 11, 8, 3, -1, 14, -10, -7, 6, -12, -17, -4, 23, 26, -5, -8, 12, 4, 0, -8, 0, -5, 8, -1, -8, 1, 0, 5, -3, 2, -2, 1, 14, 4, 11, 12, 11, 5, -8, -22, -15, 8, 4, 3, -1, -4, 10, -18, 12, -31, -11, 34, 17, -7, -3, 2, 7, -10, -16, 7, 8, 0, -2, -7, -9, -10, -22, 18, -28, 21, 11, -14, 18, 4, -10, -9, 0, 11, -6, 8, 9, -14, -13, 26, -18, 9, 5, -4, -7, -10, -10, 11, 17, -2, -4, 19, -7, 10, -19, -11, 20, -6, -35, 27, 24, 4, -11, -8, -6, -17, -9, 6, 0, 7, 3, 5, 22, -6, -2, 18, -29, -3, -10, -14, 35, 7, -11, -9, -6, -1, -12, -8, 22, -4, -7, 0, -4, 7, 5, -10, 4, 0, 3, -5, -22, -35, 22, -1, 13, 30, 29, 25, -17, -46, -1, 22, 19, -14, -28, 2, 1, 8, -15, 10, 6, 0, -24, -3, -11, -14, 7, 17, 15, -2, -6, 8, -13, -9, 13, 1, -11, 6, 6, -3, 5, 2, -8, -1, 8, 0, 3, 3, -3, 5, 7, -6, -4, 22, -2, 17, -4, -21, 3, -10, -7, -6, 8, 28, 6, -8, 19, -19, 17, -30, -14, -1, -24, 11, -2, 14, -5, 7, 8, 13, 0, -2, 0, -4, 4, 0, -1, -1, 0, 8, 12, 11, 1, -7, 13, -19, -3, -11, 8, -6, -18, 4, -19, -1, 7, -7, 0, 19, 14, -3, -11, 10, -16, 0, 1, -4, 19, 16, -4, -23, 7, -1, 2, -3, -19, 9, 19, -11, -1, -4, -4, -11, 7, -13, -1, 11, -3, -5, -7, 6, 10, -15, 6, -14, 16, -11, -15, 23, 32, -36, 4, -2, -2, -4, -16, 14, -18, 18, 2, 10, 7, 0, -18, 10, -7, 7, -11, 10, -21, 20, -2, 6, -11, -5, -11, 0, 5, 4, 3, -6, -9, -15, 3, 2, -2, 17, -16, 5, -6, 16, 4, 3, 4, 0, 0, 0, -2, 3, -3, 0, 6, 28, 6, -4, -13, -17, 1, 11, -5, -13, -3, 11, 10, -18, 2, 15, -1, 3, -6, -11, 17, -10, 20, -12, -20, 3, 9, 23, -12, -12, -2, 17, -18, 5, 0, -17, -26, 3, 11, 31, -1, 5, 5, -7, 12, 4, -12, -10, -10, 4, -25, 3, -26, 17, -23, 31, 22, -20, 12, 25, 0, 4, 2, -2, 12, -2, 0, -3, -3, -16, 20, -10, -27, 4, 33, 7, -13, 13, -11, -11, -1, 1, 0, -3, -17, 1, 0, 20, 0, -4, -9, -9, -6, -12, -3, -5, 11, 16, 3, 4, 4, -2, -7, 2, 10, 0, -8, -10, -2, 3, 18, -6, -2, -1, -9, -2, -11, -9, 22, -4, 1, 6, 1, -13, -1, 6, 0, 3, -2, 1, -7, -3, -5, 10, -7, -5, 12, -6, 3, -1, 21, 27, -9, 28, -21, -5, -16, -18, 6, -2, 11, 1, -13, 18, 0, -15, -1, -3, 27, -20, -19, 5, -25, 12, 2, -1, -9, -3, 30, 3, 2, -5, 9, -7, -14, -1, 31, -7, 6, -6, -16, -2, -18, 4, 27, 12, -8, 9, 10, -4, 2, -15, 9, 14, 3, 13, 36, -20, -24, -17, 0, -2, 12, 3, -2, 0, 1, 3, 6, -2, -8, 7, -8, 21, -44, 15, 15, 9, 9, 1, -2, -18, -6, 24, 15, 7, -25, -9, 23, -18, 24, 5, 25, 6, -3, -21, 1, -21, -14, 13, 3, 13, -37, -12, 12, 0, 24, -14, 8, 0, 24, -16, -7, -18, -6, 10, 1, -5, 18, -2, 16, -22, 37, 17, 8, -8, -9, -35, 3, -4, -1, -27, 10, 7, -4, -17, 1, -1, 20, 18, -3, 4, 4, 4, -3, -9, 2, 11, -5, -5, 36, -8, 6, 38, 12, -16, -13, -9, -33, -13, -1, 11, -8, -12, 0, 7, 9, 1, -3, 8, 0, -9, 1, -4, 6, 1, -2, 5, 7, 1, 7, 4, -3, 0, 2, 3, 0, 5, -5, 0, 23, -32, 9, 6, 2, -5, 10, 13, -18, -2, -9, -14, 17, 10, -15, -4, -5, 8, -2, 6, 0, 2, 1, 3, -6, 19,
    -- filter=0 channel=9
    0, 15, -3, -11, 2, 3, 2, -12, -4, 10, 20, -7, 1, 0, -26, 6, 5, 8, 4, -4, -13, 14, 19, -6, 2, -9, 2, -4, -1, 12, 3, -8, 0, 1, 1, 8, 6, -1, 2, -6, -1, 0, 3, -4, -6, 5, -18, 17, 2, -1, -8, 8, 6, -12, 7, 7, 0, -2, -6, 4, 5, 4, 1, -8, 2, 31, -4, -15, -15, 18, -20, -20, -6, 19, -11, 4, -19, -3, -21, 37, -3, 7, 0, 5, -3, -13, 3, -2, -4, 12, 5, -9, 7, 5, -6, 19, 30, -7, -25, 17, -19, -3, -21, 21, 43, -8, -15, -15, -8, 11, 0, -18, 33, -5, -10, -25, -2, 15, 12, 21, -8, -22, 0, 14, 0, 15, 16, -18, 28, -5, -5, -14, -4, -3, -3, -13, 5, 5, 5, 4, 31, -26, 3, -13, 0, -10, -19, 6, -4, -5, 7, 10, 4, 1, 18, 12, 15, 5, -2, 2, -16, 3, -15, -15, 21, 28, 0, -20, 3, 5, 1, 0, -23, -21, 8, -8, 22, 2, -22, -11, -10, -7, 14, 13, 12, 34, -9, -5, -2, -14, -21, -22, 3, 18, -13, 20, -18, -24, 19, 7, 13, 0, -11, -2, -27, 18, -14, 0, -5, -3, 12, 21, -2, 2, -13, -25, -34, 0, 29, 28, -27, 9, 5, 26, 5, -11, -18, 7, -13, -17, 29, 31, -7, 1, 17, -12, 22, 16, -8, -21, -26, 30, -15, -9, 18, 20, 1, -25, 32, -24, 3, 10, -11, -37, -5, 2, -8, 4, -11, -12, -7, -5, 20, 16, 1, 21, -2, -7, -3, 1, 1, -35, 24, 19, 8, -4, -15, 6, 7, 14, 0, -11, -16, 7, -22, 5, -2, 1, -19, 2, 7, 3, 12, 2, 5, -15, 19, -4, 9, -4, 2, 4, -17, -8, 19, -1, 5, -31, 17, -16, -34, 36, 18, -28, -3, 36, 10, 19, 10, -33, 18, -20, -9, -18, -8, -12, -2, -21, 16, -4, 16, 15, 2, -1, -1, 3, -13, -34, 13, 9, 2, 27, -2, 4, -20, 9, -18, 26, 9, 13, 8, -13, -3, -14, -9, -11, 6, -13, -9, 2, 11, 11, 18, -7, -31, -6, 27, 5, 10, -1, 22, -2, -7, -17, 9, -3, -19, 5, -13, -2, -2, 1, 18, 13, -9, 25, 4, 2, -36, 11, 15, 3, -8, -12, -1, -17, 24, -7, 2, 5, 19, -4, -11, -4, -11, 11, -37, 15, 46, 10, -18, 10, 0, -4, 3, 3, 0, -8, -6, 9, 0, -1, 3, 4, -4, 5, -11, 18, -20, 7, 1, -18, -1, 16, -17, -15, 16, -2, 16, 7, 3, -16, 16, -24, 4, -17, 6, 27, -6, 10, -14, 0, -14, 5, 1, -8, -19, 13, 13, 1, -6, -4, 3, 12, -18, 17, 38, -33, 16, 12, -15, -5, -29, 0, -7, -13, 3, -13, -1, 25, -4, -18, 0, 10, 2, 1, -5, 6, 3, -11, 0, 0, 1, -5, 8, -9, -16, 13, -2, -20, 11, 22, -5, -9, -15, 0, -10, -1, 10, 0, -9, 12, 13, -1, -19, 24, 35, -21, -46, 17, 16, 11, -28, 8, 6, 11, 0, -17, 29, -18, -35, 28, 0, -1, -23, 10, 17, -20, -9, 30, -12, 2, -12, 18, -19, 2, -31, -10, 5, 13, 30, 39, -15, -21, 6, -11, 1, 10, 2, -9, -14, -5, 13, -1, -9, 26, -29, -14, 13, 1, -22, 8, -4, 26, 10, -5, 26, -13, -20, -1, 6, 14, -14, -6, -12, 24, -5, 1, 17, -10, -26, -4, 2, 19, -13, 7, 0, 16, -10, -13, -20, 37, -6, 0, -14, 4, -19, 5, 4, -19, 5, 22, 10, 14, 0, -7, 1, 20, -6, 1, -3, 2, -22, 21, -12, 3, -15, -9, -4, -11, -9, -9, 33, 30, -15, 3, -6, 2, -33, -10, 2, 8, -4, 37, 3, 18, -14, -8, 30, -6, 2, -14, 10, -14, 1, -5, -19, 8, -5, 3, 15, -6, 1, 0, 13, -8, -8, 1, 0, -12, -11, 40, -18, 8, -31, -9, -2, 28, 35, 2, 11, -11, -14, -17, -22, -8, -8, 6, -14, 5, -18, 4, 19, 23, 7, 13, -8, 5, -6, 5, -2, -7, -16, 17, 17, -10, 0, -4, 7, -28, 28, 0, -15, 7, 11, 2, -10, -7, -9, 0, -2, -11, 5, 0, 11, -8, 3, -15, 0, 5, -8, 4, 3, -6, 12, -15, -9, -11, 18, -3, 11, 15, 2, -13, 4, 8, 2, -1, -3, 4, -6, 4, -5, -3, 8, 30, -4, -4, -20, -17, -16, -18, 7, 36, 0, -6, -3, -6, -3, 9, 1, -5, 5, 0, -17, 0, 5, -6, 9, 3, -10, -5, 2, 8, -19, -3, 6, 11, -11, 10, -23, -5, -3, 15, 15, 5, 18, -38, 0, 5, -7, 27, -45, 4, 3, -16, 0, -19, 12, -5, 0, 1, 8, 5, 0, -1, 6, -2, 8, -2, 0, -2, 0, -5, 1, 5, -9, 7, 17, -6, 3, 4, 2, -12, 15, -22, -2, 16, -10, -2, -5, 22, -34, 8, -6, -3, 1, -2, 0, -4, -5, -1, 4, 5, 4, 3, -18, 10, 4, 2, 2, 11, 8, -5, -2, -16, -2, -13, 29, -7, 25, 7, -3, -7, 17, -13, 1, -8, -11, -7, -18, 25, 13, 2, -2, -4, -5, -17, 3, -3, 11, 21, -13, 12, 5, -9, 15, 0, -4, -2, 8, -13, -1, 0, 0, 1, 0, 2, 1, -8, 3, 8, 0, 0, 26, 7, 27, -21, 18, -7, -2, -5, -11, -25, 21, 9, 7, -24, -7, 23, 9, -30, 7, -8, 0, 0, 0, 1, 4, -2, -3, 1, 0, -5, 7, 3, 2, 0, 2, 2, 6, -5, 0, 3, -16, 22, -15, 18, 7, -10, 7, -2, 11, -17, 11, 2, 4, -9, -8, -13, 0, 4, 7, -5, 12, -7, -23, 7, 18, -5, -15, 25, -6, -5, 2, -5, 0, -4, 2, -2, 0, -4, -5, 5, -16, 11, -3, 3, 0, 0, -16, -3, 29, 16, -7, -2, 3, 0, 12, -3, -3, 7, 4, 2, 25, 0, 15, 0, -10, 22, -5, -9, -33, -4, 8, -7, 4, 13, -42, 9, -5, 6, 6, 13, 19, -9, -10, 31, -7, -17, -8, 4, -6, -10, 5, -48, 42, -15, -3, 5, -22, 8, -4, 34, -7, 1, -15, -1, 2, 6, -6, 19, -7, -4, 35, 0, 25, -13, 19, -23, -21, 10, -12, -13, 18, 16, 8, 27, 8, -27, -12, -18, 7, -17, 14, -5, -1, -12, -1, -1, 2, -6, 25, -11, -28, -16, -7, 11, 17, 11, 16, 3, -13, 6, 3, 8, -7, 20, -10, 21, -14, -19, 6, -10, -3, 1, 2, 6, 34, -9, -38, 30, -11, -26, 24, 10, -13, 17, 12, -21, 0, -6, -5, -13, -3, 0, -13, 7, -15, 0, 20, 7, 17, -21, -15, 7, 11, 7, 6, -5, 15, -11, -20, 14, 18, 5, 5, -5, -1, 5, 1, -2, -14, -7, 1, 6, 5, -28, 31, 10, -19, 19, -3, -20, 8, 4, 0, -4, -7, 0, 0, -1, 13, -10, 4, -6, -6, 0, 0, 3, 1, 0, -1, 1, -3, 9, 8, 0, -11, 4, 9, -15, -2, -3, 13, 22, 10, -9, -25, 12, -3, 5, -7, 3, 8, -5, -5, 2, 0, -3, 3, 2, -1, 4, 4, 3, -6, 0, 7, -3, 7, 0, -2, -6, -2, 2, -12, -4, -1, 9, -8, 1, -2, -5, 1, -7, 11, 5, -6, -17, 18, -9, 5, -3, -37, -19, 18, 21, 3, 15, -37, 19, -13, 31, 26, -7, -10, -9, -10, -8, 5, -7, 27, 7, 19, -13, 5, -14, 0, 0, 9, -14, 21, -29, 15, 11, -24, -3, 21, -20, -16, -27, 18, 26, 0, 0, 0, -3, 6, -7, 6, -7, -7, 7, 16, 8, -25, 0, 3, 14, -13, -19, 19, -5, -25, 4, 16, 6, 12, -2, 17, -15, -2, 0, -6, -6, -1, -4, 5, 9, 5, 1, 0, 0, 24, 1, 26, -44, 14, 15, 12, -5, -1, -29, 7, -13, 2, 13, 16, 2, -9, -5, -15, -5, -13, -8, -6, -19, -6, 14, -13, 24, 17, 0, -21, -4, 12, 15, 19, -3, -12, -9, 7, -3, 7, -20, 9, 19, 9, -27, 17, -8, 4, -9, -6, -5, -9, 23, -1, -5, -14, -6, -9, 14, 7, -5, 6, 12, -9, -3, 0, -6, 1, -5, 14, -11, 8, -9, 5, 10, 5, 7, -3, 0, -3, -14, -12, 10, 32, 1, -6, -10, 9, 2, -15, -2, 5, -33, 23, 25, 12, -2, -12, -4, -3, 3, -5, 2, 11, -11, -2, 5, 7, 3, 0, -9, 15, -5, 16, 2, 0, 5, -5, 0, 7, 8, 27, -22, 41, -17, 0, -25, -17, 5, 9, 26, -5, -7, -16, -9, 8, 8, -5, 5, -5, 5, 3, -1, 5, -1, 0, -4, 1, 2, 43, -6, 6, 16, 11, 1, -6, -14, -50, -16, 2, -8, -4, 12, -9, 11, -11, 14, -16, -3, 0, -2, -8, 5, 20, 6, -30, 24, -4, -8, 2, -5, 0, -6, 3, 5, 0, -5, 3, 3, 10, -20, 6, 0, -14, 19, -17, -2, 18, 5, -21, -1, -14, 4, -2, -7, 18, -1, 15, 18, 30, -21, 4, 18, -13, -15, -3, -14, 0, -6, -12, 11, -11, 1, -15, 38, 0, -21, 5, -2, 1, -5, -8, 21, 3, -11, -2, 0, 2, -4, 5, -4, 1, 0, -2, 10, -1, -6, 4, 5, 29, -9, 11, -24, -14, -6, -14, 27, 21, -8, -5, -4, 16, -1, 3, 0, 0, -9, -2, -1, -5, 1, -12, 7, -12, 2, 23, 24, -25, 10, 0, 5, 15, 9, 28, -1, -27, 11, 2, -19, -3, -13, -3, 14, 4, -13, 4, 8, -4, 2, -28, 13, -25, -4, -24, 17, -7, -21, 54, 10, -8, 22, 24, 0, -26, 14, -5, 2, 9, -28, 2, -5, -4, 2, 3, -1, 6, -2, 8, -9, 11, 29, 4, 6, -12, -10, -4, 6, -17, 3, 6, -7, -14, -2, -3, -14, -21, 0, 32, 26, 28, -5, 1, -33, 35, -4, -20, 41, -42, 3, -6, -2, 12, -25, 14, 21, 8, -9, -6, -11, -1, 3, -28, -4, -23, 1, 3, 31, -15, 28, 0, 17, -8, 4, -17, -24, -11, 25, -8, 29, 17, -21, 17, -4, 10, 0, -12, 2, -5, -16, 5, -3, -4, 9, 4, -14, -4, 7, -6, -2, 14, 0, 22, -17, -10, 19, 38, -46, -13, -9, 12, 0, 7, -13, -14, 19, -13, 14, -45, 32, -17, -3, -30, 11, -22, -11, 29, 22, 12, 8, -10, -1, 0, 17, -13, 5, 1, -2, -15, 13, -25, 28, -6, 18, 12, -10, -7, -9, 1, -13, -4, 4, 4, -2, 16, -26, 28, -9, -5, -15, 0, -32, 19, 13, 0, 12, -19, 4, 0, 3, 20, -8, -6, -23, -3, 5, -2, -21, 35, 16, 27, -20, -1, -10, -18, 0, 1, 7, 16, -2, 10, 22, 16, -10, -5, 3, 0, 2, -6, -23, 5, -4, -11, -31, 12, 15, 6, 25, -12, 10, -19, -22, -9, 3, -7, 22, -2, 32, 2, 2, 2, -7, 32, 4, -6, -6, -7, -1, -3, -12, 28, -12, -26, 4, 13, 13, -48, 39, -11, 0, 5, 1, 1, 9, 1, 0, -4, 0, -13, 10, 8, 5, 8, -10, -4, 8, 0, -12, -5, -1, 23, -14, 9, -1, -1, -4, -18, 8, 14, -8, 0, 2, 0, 6, 0, -2, 1, 2, 6, -5, -12, 21, 2, 9, 11, -4, 0, -12, -16, 10, 18, 11, 13, -6, 2, -29, -38, 4, 24, 3, -21, 38, -2, -2, -7, -16, 29, -27, 24, -18, 21, -23, 5, -26, 3, 1, 29, 16, -12, -19, -21, -14, -5, 10, -4, -1, -12, -3, 24, 19, -1, -4, -4, -30, 40, -12, 23, -4, 0, -9, -18, 39, -10, -3, -21, 10, -10, -21, -17, 36, 3, 4, -1, 0, -2, 1, -6, 0, -4, -2, -13, 3, -26, 23, 7, 6, 16, -8, -5, -9, 11, 22, 12, 0, -2, -11, -5, 2, -13, 4, 2, -11, 13, -26, -25, 15, 16, -15, 14, 16, -20, 1, 6, 9, -7, -21, 23, -7, 11, 6, 10, -28, -7, 5, -33, 22, -20, 34, -5, 8, 10, -23, -6, 25, -37, 8, 30, -7, -6, 9, -36, -3, -12, 8, 30, 11, 0, 15, -12, -2, 11, -6, 13, 33, -8, 26, -17, -34, 1, -4, -9, 7, -2, 20, -2, -15, -3, -15, -16, 25, 4, -14, -9, -10, 8, 5, 6, -9, 4, 3, -8, 7, 21, -13, -6, 2, -9, -2, 1, -11, -7, -6, 9, 9, -2, -22, 1, -5, 3, 16, -6, 30, -16, -20, 24, 10, -6, 6, -4, -9, 6, 5, -2, 2, 14, -4, -3, 6, -14, 4, 8, -7, -4, 17, 15, -27, 0, 10, -9, -12, -2, 3, 4, 7, -4, -7, 3, 2, -1, -3, -12, -14, 0, -3, 9, 7, -16, -7, 12, 26, -7, -5, 4, -9, 0, -4, -1, 5, -1, 7, -7, 1, 4, 2, 4, -6, -2, 3, -1, 2, -14, -22, -1, -7, 8, 18, 14, 29, -12, -20, -19, -2, -20, 19, 11, 8, 21, 0, -1, -9, 9, 4, 10, 5, 0, 11, -15, 6, -16, -1, -2, 3, 1, -14, 4, 11, -15, 9, 1, -7, -25, 25, -2, -18, -15, 4, 3, 8, 5, 18, 1, 39, -21, -32, 27, -9, -39, -28, 12, 48, -12, 20, -7, 1, -18, 0, 1, 34, 17, -31, 20, 26, -13, -5, 6, -16, -10, -18, 16, 4, -5, -5, 0, 0, 0, 5, 0, 2, 4, 1, 0, -6, 0, -5, 5, -2, 0, -2, -1, 16, 5, -17, 16, 16, 5, -10, -6, 22, -26, -1,

    -- ifmap
    -- channel=0
    0, 126, 276, 171, 3, 65, 0, 0, 0, 177, 193, 129, 0, 186, 0, 27, 60, 81, 0, 0, 38, 0, 0, 0, 136, 81, 129, 0, 265, 152, 203, 31, 81, 0, 0, 33, 65, 294, 124, 124, 181, 0, 0, 36, 72, 174, 0, 0, 142, 328, 0, 90, 0, 0, 78, 0, 368, 0, 0, 0, 0, 0, 213, 0, 0, 38, 101, 105, 0, 188, 0, 77, 0, 31, 41, 0, 77, 57, 0, 75, 0, 69, 0, 102, 0, 100, 0, 0, 0, 204, 73, 65, 48, 190, 208, 0, 156, 225, 0, 0, 0, 0, 0, 0, 0, 0, 15, 76, 0, 234, 0, 0, 0, 0, 0, 237, 0, 181, 37, 239, 199, 120, 0, 0, 153, 37, 41, 0, 11, 0, 196, 21, 56, 0, 196, 111, 28, 0, 60, 193, 0, 117, 0, 114, 484, 137, 136, 2, 0, 150, 211, 0, 76, 83, 0, 0, 0, 0, 0, 158, 171, 0, 0, 185, 182, 0, 0, 231, 0, 0, 419, 0, 0, 0, 0, 0, 97, 0, 0, 4, 0, 0, 38, 48, 0, 422, 3, 0, 407, 80, 0, 38, 17, 149, 121, 0, 0, 125, 163, 319, 161, 0, 24, 58, 0, 41, 71, 80, 0, 146, 0, 129, 0, 111, 43, 0, 32, 0, 44, 0, 0, 0, 0, 17, 70, 95, 0, 265, 155, 0, 0, 0, 69, 276, 64, 379, 279, 0, 0, 0, 0, 20, 29, 158, 328, 0, 0, 171, 0, 419, 0, 175, 0, 0, 100, 0, 0, 2, 79, 0, 0, 0, 0, 0, 51, 0, 0, 0, 123, 19, 0, 15, 85, 97, 0, 0, 80, 158, 300, 0, 146, 0, 18, 397, 0, 0, 245, 0, 445, 0, 41, 0, 0, 177, 0, 187, 9, 0, 0, 0, 0, 0, 276, 0, 137, 84, 234, 19, 2, 98, 121, 188, 147, 139, 159, 212, 0, 326, 0, 219, 17, 0, 0, 104, 51, 0, 0, 322, 0, 20, 0, 346, 243, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 66, 0, 23, 0, 94, 0, 131, 0, 0, 33, 267, 58, 137, 0, 26, 0, 92, 0, 0, 0, 0, 462, 38, 201, 0, 0, 256, 0, 0, 135, 312, 0, 0, 0, 0, 0, 238, 271, 0, 0, 141, 0, 102, 0, 50, 37, 184, 171, 15, 0, 0, 0, 10, 164, 0, 207, 85, 0, 41, 75, 56, 0, 0, 0, 0, 0, 68, 44, 26, 92, 22, 36, 297, 0, 88, 38, 0, 0, 40, 177, 59, 75, 0, 35, 341, 0, 79, 48, 142, 179, 157, 112, 0, 151, 274, 0, 106, 64, 17, 0, 146, 1, 0, 2, 22, 0, 124, 0, 41, 0, 0, 0, 214, 61, 129, 4, 83, 0, 0, 428, 0, 0, 0, 227, 0, 0, 0, 0, 0, 0, 60, 237, 318, 43, 120, 0, 141, 194, 129, 200, 28, 126, 0, 107, 16, 0, 0, 0, 0, 18, 0, 0, 372, 211, 71, 128, 0, 0, 0, 64, 32, 0, 0, 0, 67, 0, 0, 0, 0, 155, 169, 224, 0, 128, 0, 0, 108, 0, 239, 107, 0, 0, 0, 91, 93, 75, 0, 3, 43, 29, 20, 425, 0, 9, 0, 5, 0, 0, 113, 45, 0, 228, 0, 13, 39, 0, 0, 25, 0, 54, 79, 169, 95, 0, 36, 1, 81, 0, 34, 92, 97, 0, 171, 0, 297, 321, 90, 10, 0, 48, 0, 0, 34, 201, 253, 0, 406, 0, 253, 110, 0, 0, 280, 230, 0, 0, 0, 14, 23, 0, 0, 0, 0, 0, 227, 63, 321, 35, 0, 0, 0, 0, 0, 30, 66, 18, 0, 0, 87, 168, 103, 0, 0, 0, 46, 0, 0, 0, 49, 0, 15, 0, 269, 179, 132, 96, 83, 27, 0, 119, 39, 288, 285, 355, 0, 0, 0, 0, 0, 71, 0, 64, 0, 0, 58, 73, 36, 28, 0, 23, 26, 0, 65, 306, 0, 82, 45, 64, 106, 154, 69, 0, 0, 103, 0, 91, 134, 228, 0, 287, 0, 0, 11, 146, 31, 130, 0, 285, 0, 102, 141, 70, 0, 0, 230, 109, 0, 0, 27, 0, 0, 0, 80, 29, 0, 0, 124, 0, 0, 202, 84, 0, 23, 0, 0, 176, 61, 78, 0, 221, 0, 143, 367, 157, 0, 0, 14, 248, 0, 0, 94, 0, 0, 122, 208, 0, 314, 370, 5, 323, 115, 17, 115, 116, 176, 0, 0, 43, 0, 73, 0, 43, 0, 181, 0, 105, 280, 326, 50, 0, 257, 163, 83, 0, 36, 203, 177, 45, 0, 124, 152, 0, 0, 74, 77, 125, 0, 0, 55, 97, 0, 148, 39, 21, 4, 0, 32, 16, 21, 0, 57, 176, 0, 139, 3, 0, 284, 0, 0, 55, 301, 0, 0, 0, 94, 161, 0, 0, 63, 0, 58, 0, 0, 0, 0, 0, 0, 0, 100, 168, 0, 49, 0, 286, 0, 39, 96, 0, 0, 0, 178, 287, 0, 64, 84, 95, 0, 0, 0, 125, 134, 132, 0, 0, 0, 145, 0, 57, 118, 62, 0, 0, 0, 41, 0, 343, 0, 0, 0, 103, 0, 0, 0, 0, 273, 0, 141, 0, 0, 213, 0, 106, 43, 62, 180, 101, 0, 0, 11, 63, 98, 0, 0, 91, 210, 332, 0, 153, 25, 45, 215, 0, 0, 225, 20, 195, 106, 244, 9, 269, 75, 128, 17, 100, 162, 171, 0, 0, 50, 39, 0, 0, 17, 0, 23, 214, 0, 31, 218, 10, 0, 288, 0, 45, 60, 43, 82, 2, 43, 0, 0, 98, 364, 0, 0, 0, 0, 0, 12, 0, 0, 188, 0, 23, 10, 0, 0, 0, 0, 217, 0, 54, 9, 49, 40, 0, 36, 0, 296, 0, 0, 0, 112, 132, 0, 32, 0, 204, 206, 0, 0, 58, 222, 0, 13, 175, 30, 150, 332, 0, 180, 221, 0, 0, 0, 0, 0, 52, 207, 2, 0, 0, 47, 128, 0, 0, 0, 7, 0, 24, 0, 0, 0, 146, 0, 19, 190, 104, 252, 230, 76, 54, 0, 21, 25, 0, 0, 0, 321, 77, 241, 0, 250, 115, 0, 21, 212, 0, 17, 0, 283, 0, 114, 0, 0, 70, 343, 282, 162, 130, 0, 0, 89, 213, 94, 13, 91, 0, 123, 47, 455, 248, 112, 82, 0, 0, 55, 0, 83, 161, 0, 68, 0, 0, 57, 0, 5, 91, 75, 0, 108, 0, 0, 152, 0, 0, 0, 0, 132, 0, 35, 0, 265, 0, 0, 48, 394, 0, 0, 0, 176, 0, 71, 42, 0, 55, 0, 67, 77, 222, 44, 119, 39, 122, 0, 3, 0, 128, 18, 0, 0, 0, 94, 62, 214, 29, 0, 0, 176, 4, 0, 0, 35, 99, 119, 0, 11, 0, 80, 2, 146, 174, 0, 246, 6, 26, 118, 190, 0, 0, 64, 0, 0, 0, 342, 0, 61, 68, 0, 66, 0, 0, 141, 0, 0, 0, 221, 0, 40, 0, 142, 108, 85, 0, 339, 0, 157, 66, 122, 114, 115, 47, 89, 107, 0, 0, 243, 201, 0, 321, 5, 90, 34, 89, 104, 194, 0, 0, 19, 124, 22, 0, 0, 121, 68, 0, 0, 0, 5, 618, 127, 0, 0, 177, 56, 417, 0, 26, 0, 0, 184, 26, 230, 32, 4, 119, 0, 41, 0, 0, 0, 198, 305, 0, 56, 220, 22, 0, 113, 46, 0, 15, 0, 30, 49, 30, 262, 7, 0, 0, 186, 115, 0, 0, 0, 0, 0, 0, 76, 0, 0, 47, 38, 344, 0, 0, 23, 0, 130, 135, 0, 0, 0, 0, 22, 0, 64, 59, 0, 169, 397, 0, 0, 0, 32, 0, 62, 0, 95, 86, 0, 0, 0, 0, 117, 128, 97, 109, 91, 196, 60, 579, 0, 0, 0, 0, 176, 208, 65, 167, 0, 304, 273, 313, 0, 0, 0, 230, 118, 0, 0, 0, 0, 122, 0, 0, 0, 85, 0, 84, 82, 0, 0, 0, 0, 71, 0, 365, 10, 33, 108, 117, 0, 159, 8, 259, 45, 0, 0, 0, 22, 239, 78, 173, 234, 186, 0, 0, 0, 0, 181, 255, 0, 0, 10, 0, 0, 56, 0, 191, 0, 0, 182, 0, 14, 47, 85, 65, 95, 0, 147, 187, 0, 0, 0, 0, 86, 6, 0, 46, 0, 0, 0, 0, 0, 0, 186, 0, 0, 0, 410, 0, 110, 0, 26, 0, 0, 30, 0, 0, 0, 0, 79, 0, 0, 0, 0, 45, 0, 0, 85, 472, 0, 141, 0, 200, 0, 123, 30, 0, 0, 83, 30, 38, 111, 0, 0, 0, 73, 0, 9, 0, 62, 63, 0, 180, 80, 89, 232, 0, 0, 221, 43, 6, 0, 87, 121, 0, 98, 232, 79, 197, 80, 0, 35, 17, 160, 0, 165, 0, 95, 0, 81, 0, 0, 0, 0, 2, 0, 0, 0, 0, 121, 47, 0, 308, 146, 0, 0, 0, 130, 89, 0, 0, 92, 330, 95, 43, 149, 0, 0, 0, 0, 16, 0, 0, 0, 0, 65, 0, 397, 109, 0, 62, 0, 223, 148, 117, 0, 332, 89, 0, 131, 92, 0, 382, 96, 0, 0, 19, 82, 200, 141, 0, 0, 0, 121, 0, 228, 255, 21, 0, 52, 0, 167, 346, 143, 56, 0, 53, 0, 0, 0, 53, 0, 242, 115, 107, 288, 0, 41, 0, 107, 72, 30, 0, 0, 0, 162, 115, 53, 0, 0, 0, 190, 0, 382, 0, 235, 0, 0, 0, 161, 141, 284, 0, 136, 0, 52, 21, 33, 112, 0, 0, 52, 0, 88, 0, 0, 232, 100, 85, 0, 0, 26, 0, 4, 0, 0, 0, 75, 0, 10, 0, 424, 102, 0, 286, 0, 0, 0, 0, 316, 53, 81, 218, 150, 0, 235, 254, 0, 0, 187, 9, 26, 164, 19, 0, 0, 108, 0, 0, 0, 21, 229, 0, 0, 161, 0, 268, 91, 0, 160, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 169, 0, 0, 326, 0, 0, 0, 0, 0, 67, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167, 0, 0, 0, 0, 0, 0, 184, 33, 75, 201, 0, 201, 0, 0, 113, 0, 0, 26, 218, 273, 340, 416, 715, 65, 96, 0, 0, 0, 0, 146, 77, 0, 0, 185, 155, 103, 0, 0, 84, 13, 0, 6, 122, 68, 28, 0, 0, 0, 0, 0, 117, 0, 293, 0, 0, 50, 0, 0, 16, 0, 0, 0, 67, 321, 0, 298, 0, 115, 94, 0, 288, 119, 132, 0, 0, 57, 0, 0, 118, 0, 0, 0, 22, 269, 62, 276, 24, 0, 0, 0, 0, 61, 99, 0, 150, 112, 116, 174, 15, 0, 102, 200, 153, 274, 0, 49, 0, 114, 25, 0, 0, 0, 120, 0, 25, 100, 0, 162, 35, 84, 99, 122, 126, 70, 204, 257, 0, 187, 0, 256, 0, 0, 230, 0, 144, 159, 87, 28, 14, 253, 0, 38, 0, 0, 115, 28, 23, 57, 38, 39, 108, 19, 0, 132, 0, 75, 153, 0, 0, 92, 0, 0, 0, 441, 243, 71, 0, 379, 0, 0, 0, 0, 0, 0, 84, 0, 82, 0, 65, 0, 0, 199, 244, 0, 0, 77, 0, 142, 188, 91, 0, 9, 225, 0, 0, 0, 0, 325, 46, 83, 0, 0, 0, 168, 0, 0, 0, 63, 0, 0, 56, 0, 98, 38, 0, 0, 0, 0, 202, 0, 121, 467, 69, 93, 345, 56, 193, 138, 311, 0, 206, 92, 139, 87, 113, 0, 0, 464, 139, 0, 9, 476, 61, 0, 0, 0, 89, 0, 78, 75, 37, 0, 0, 0, 22, 84, 134, 0, 105, 0, 189, 159, 0, 0, 0, 150, 0, 95, 70, 136, 64, 235, 65, 87, 0, 63, 0, 261, 0, 187, 184, 0, 0, 0, 0, 239, 225, 0, 60, 0, 0, 39, 0, 0, 98, 385, 73, 0, 0, 31, 311, 0, 162, 0, 59, 105, 51, 0, 0, 108, 57, 0, 84, 0, 0, 22, 351, 0, 32, 108, 0, 121, 16, 0, 371, 0, 43, 0, 28, 0, 0, 250, 83, 279, 0, 0, 69, 38, 0, 208, 62, 0, 104, 248, 238, 0, 25, 89, 0, 0, 0, 0, 0, 175, 20, 0, 0, 274, 89, 7, 0, 0, 0, 294, 19, 69, 76, 0, 0, 124, 0, 0, 0, 88, 0, 0, 380, 14, 19, 153, 0, 0, 0, 0, 0, 24, 72, 137, 0, 111, 173, 0, 295, 319, 0, 0, 44, 406, 190, 0, 187, 0, 0, 0, 86, 0, 90, 63, 38, 62, 0, 51, 0, 0, 0, 139, 131, 0, 26, 0, 60, 98, 0, 0, 139, 0, 0, 0, 151, 119, 0, 0, 121, 130, 0, 19, 119, 0, 235, 0, 0, 154, 94, 100, 28, 0, 11, 0, 57, 218, 19, 313, 52, 0, 146, 33, 68, 0, 0, 0, 250, 0, 0, 0, 0, 63, 152, 89, 119, 0, 9, 0, 57, 18, 152, 149, 0, 124, 27, 81, 0, 0, 127, 0, 101, 397, 0, 8, 0, 0, 131, 0, 48, 0, 90, 0, 77, 5, 10, 0, 2, 0, 0, 0, 39, 0, 67, 0, 322, 248, 267, 100, 0, 0, 0, 0, 84, 159, 9, 0, 0, 0, 0, 0, 178, 0, 0, 0, 0, 0, 0, 0, 385, 93, 329, 111, 17, 205, 0, 0, 0, 70, 74, 0, 308, 86, 0, 0, 27, 0, 2, 0, 0, 0, 28, 243, 0, 25, 0, 41, 132, 0, 47, 121, 69, 0, 0, 0, 47, 136, 0, 293, 0, 0, 267, 0, 0, 30, 322, 0, 237, 141, 0, 0, 119, 0, 0, 320, 202, 0, 0, 40, 138, 0, 310, 0, 9, 91, 32, 0, 0, 0, 0, 116, 0, 0, 0, 63, 0, 205, 114, 191, 0, 148, 337, 103, 48, 0, 151, 0, 26, 0, 0, 77, 0, 0, 132, 0, 109, 0, 161, 0, 0, 0, 3, 0, 235, 
    
    
    others => 0);
end inmem_package;
