library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 
    0, 34, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 30, 
    0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 32, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 38, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 40, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 17, 0, 0, 0, 0, 0, 0, 0, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 25, 12, 0, 0, 0, 0, 0, 2, 11, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 12, 8, 1, 0, 0, 0, 0, 4, 7, 11, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 15, 13, 6, 2, 2, 7, 11, 10, 6, 4, 6, 10, 6, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 21, 14, 13, 14, 15, 17, 17, 14, 15, 13, 13, 15, 16, 17, 16, 13, 12, 16, 22, 18, 30, 
    5, 10, 0, 0, 0, 0, 0, 0, 0, 15, 33, 25, 16, 10, 10, 9, 10, 14, 16, 17, 18, 21, 21, 17, 12, 8, 8, 13, 19, 22, 15, 29, 
    2, 26, 6, 0, 0, 0, 0, 0, 3, 36, 26, 17, 10, 7, 9, 11, 12, 14, 16, 17, 16, 15, 16, 13, 9, 10, 15, 20, 18, 8, 5, 25, 
    3, 28, 27, 5, 0, 0, 0, 0, 27, 34, 15, 12, 13, 13, 12, 11, 11, 13, 13, 15, 15, 12, 11, 12, 15, 22, 27, 23, 10, 1, 12, 29, 
    2, 29, 28, 23, 0, 0, 0, 3, 21, 15, 4, 5, 8, 12, 13, 14, 15, 15, 15, 14, 14, 16, 16, 19, 24, 30, 29, 19, 14, 17, 24, 35, 
    0, 26, 24, 24, 19, 0, 0, 12, 35, 13, 9, 2, 0, 2, 5, 9, 13, 15, 15, 16, 16, 16, 18, 22, 28, 27, 15, 11, 14, 25, 26, 33, 
    0, 25, 22, 20, 22, 17, 0, 12, 36, 24, 18, 14, 10, 6, 3, 1, 0, 2, 5, 7, 8, 13, 17, 19, 14, 5, 1, 1, 8, 19, 23, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 50, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 52, 40, 9, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 66, 59, 56, 52, 20, 0, 0, 0, 0, 0, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 38, 42, 18, 29, 60, 60, 5, 0, 0, 0, 0, 33, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 34, 42, 10, 0, 0, 3, 31, 3, 0, 26, 61, 50, 0, 0, 0, 0, 44, 
    0, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 33, 28, 29, 14, 0, 0, 0, 22, 15, 0, 3, 51, 72, 22, 0, 0, 0, 51, 
    0, 148, 29, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 5, 23, 25, 36, 9, 0, 0, 0, 22, 39, 20, 13, 47, 80, 69, 0, 0, 0, 40, 
    0, 129, 14, 0, 0, 0, 0, 0, 0, 4, 32, 0, 0, 15, 24, 29, 52, 17, 0, 0, 0, 50, 55, 39, 15, 40, 72, 85, 38, 0, 0, 25, 
    0, 91, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 29, 15, 65, 33, 0, 0, 23, 63, 41, 29, 6, 20, 58, 86, 76, 4, 0, 20, 
    0, 74, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 50, 22, 67, 45, 0, 0, 25, 55, 35, 29, 2, 3, 32, 66, 76, 34, 34, 39, 
    0, 78, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 49, 32, 53, 32, 0, 0, 29, 63, 45, 38, 15, 1, 8, 41, 53, 17, 39, 51, 
    0, 81, 7, 109, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 38, 1, 0, 0, 20, 58, 62, 54, 32, 18, 13, 23, 20, 0, 17, 45, 
    0, 87, 17, 145, 97, 0, 0, 0, 0, 0, 0, 0, 43, 14, 0, 0, 0, 0, 0, 0, 0, 51, 61, 37, 18, 4, 0, 0, 0, 0, 0, 37, 
    0, 109, 36, 153, 171, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 62, 53, 10, 0, 0, 0, 0, 0, 0, 34, 
    0, 135, 65, 139, 199, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 46, 34, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 133, 79, 114, 193, 128, 0, 0, 45, 6, 0, 0, 0, 0, 0, 61, 17, 0, 0, 0, 0, 0, 8, 17, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 96, 70, 87, 168, 148, 20, 0, 65, 67, 12, 0, 0, 0, 2, 109, 84, 0, 0, 21, 40, 35, 35, 43, 16, 0, 0, 0, 0, 0, 0, 44, 
    0, 50, 65, 67, 136, 134, 29, 9, 117, 124, 63, 0, 0, 0, 32, 142, 162, 60, 0, 0, 26, 68, 92, 93, 69, 21, 0, 0, 0, 0, 9, 63, 
    0, 36, 88, 73, 117, 100, 0, 0, 169, 254, 200, 133, 87, 76, 90, 160, 205, 171, 112, 88, 103, 148, 186, 204, 192, 152, 101, 78, 83, 86, 131, 119, 
    0, 65, 118, 96, 121, 93, 0, 0, 171, 283, 278, 198, 111, 88, 96, 139, 187, 202, 203, 218, 239, 258, 273, 287, 292, 279, 253, 247, 257, 260, 271, 186, 
    0, 98, 120, 115, 129, 88, 0, 9, 143, 215, 220, 164, 128, 123, 130, 154, 199, 235, 258, 280, 295, 309, 313, 321, 334, 344, 343, 342, 349, 355, 351, 228, 
    67, 172, 121, 103, 101, 22, 0, 70, 169, 191, 222, 236, 236, 243, 244, 252, 275, 291, 297, 305, 319, 334, 342, 350, 361, 372, 376, 374, 379, 386, 378, 248, 
    165, 302, 203, 120, 67, 0, 0, 140, 202, 229, 266, 298, 314, 315, 306, 300, 303, 310, 317, 328, 343, 358, 369, 378, 385, 388, 383, 386, 401, 413, 399, 270, 
    193, 392, 313, 200, 86, 0, 50, 215, 254, 269, 282, 311, 329, 323, 310, 308, 313, 320, 330, 347, 361, 375, 388, 397, 396, 384, 378, 389, 417, 429, 398, 264, 
    192, 417, 392, 304, 159, 16, 80, 260, 313, 290, 292, 313, 332, 337, 321, 313, 317, 327, 341, 356, 372, 379, 379, 385, 391, 391, 397, 417, 443, 419, 363, 234, 
    189, 421, 421, 377, 264, 101, 104, 256, 315, 277, 290, 310, 332, 344, 337, 323, 317, 325, 340, 360, 374, 379, 373, 368, 374, 394, 425, 450, 448, 403, 344, 217, 
    184, 420, 420, 398, 345, 227, 171, 241, 293, 271, 274, 287, 309, 326, 329, 320, 318, 330, 348, 368, 378, 377, 363, 347, 350, 387, 435, 464, 455, 425, 356, 217, 
    154, 375, 368, 354, 343, 293, 241, 251, 277, 265, 256, 257, 261, 260, 261, 260, 264, 279, 304, 334, 347, 337, 318, 299, 292, 324, 379, 415, 409, 378, 318, 203, 
    71, 216, 212, 202, 202, 192, 174, 163, 169, 163, 153, 151, 152, 147, 134, 114, 109, 124, 151, 183, 199, 194, 180, 157, 136, 153, 199, 238, 238, 219, 196, 145, 
    
    -- channel=2
    131, 149, 142, 138, 138, 140, 143, 143, 144, 142, 140, 138, 140, 145, 147, 145, 143, 142, 142, 142, 140, 140, 139, 139, 138, 133, 132, 131, 131, 130, 103, 70, 
    111, 108, 98, 87, 89, 95, 99, 100, 102, 101, 92, 85, 90, 94, 96, 96, 95, 96, 96, 93, 96, 95, 97, 96, 97, 101, 102, 106, 106, 108, 75, 57, 
    86, 75, 74, 58, 56, 63, 69, 71, 73, 76, 68, 59, 63, 57, 59, 57, 55, 57, 64, 80, 82, 79, 73, 66, 66, 66, 78, 84, 88, 91, 55, 39, 
    85, 76, 77, 61, 59, 62, 67, 68, 72, 80, 77, 65, 61, 63, 57, 41, 34, 49, 76, 94, 106, 110, 109, 101, 90, 89, 90, 93, 92, 95, 54, 36, 
    71, 62, 78, 72, 74, 72, 66, 66, 71, 75, 57, 37, 36, 45, 39, 32, 42, 63, 81, 90, 110, 125, 128, 127, 122, 113, 101, 107, 96, 91, 53, 34, 
    52, 39, 60, 82, 82, 83, 70, 67, 72, 78, 62, 33, 30, 49, 64, 68, 84, 93, 102, 102, 107, 123, 124, 131, 131, 128, 117, 108, 103, 84, 48, 31, 
    45, 52, 77, 104, 96, 87, 71, 65, 65, 68, 71, 55, 60, 78, 96, 110, 128, 121, 105, 92, 91, 119, 121, 118, 118, 123, 124, 110, 106, 82, 41, 33, 
    44, 76, 112, 133, 117, 98, 76, 63, 52, 57, 69, 82, 80, 88, 101, 121, 142, 131, 94, 71, 69, 99, 109, 111, 114, 118, 129, 121, 105, 96, 40, 35, 
    47, 85, 134, 152, 123, 100, 86, 78, 72, 74, 89, 89, 79, 82, 93, 115, 131, 120, 92, 71, 53, 86, 106, 115, 114, 124, 139, 134, 107, 94, 44, 30, 
    37, 67, 139, 135, 118, 89, 79, 52, 32, 7, 64, 77, 70, 65, 80, 103, 119, 125, 96, 83, 57, 88, 99, 113, 124, 134, 138, 142, 122, 100, 59, 29, 
    33, 40, 118, 101, 107, 85, 79, 31, 0, 0, 10, 49, 48, 56, 72, 101, 113, 133, 98, 95, 60, 83, 89, 102, 122, 137, 136, 136, 132, 114, 72, 42, 
    40, 25, 99, 73, 90, 75, 74, 22, 0, 0, 0, 28, 49, 55, 79, 105, 113, 137, 89, 84, 45, 78, 82, 98, 117, 132, 131, 131, 141, 136, 98, 54, 
    47, 30, 88, 42, 69, 67, 69, 55, 2, 0, 18, 64, 61, 61, 84, 105, 109, 128, 72, 68, 33, 73, 76, 101, 120, 130, 136, 136, 142, 147, 119, 71, 
    50, 29, 84, 40, 65, 73, 60, 70, 37, 40, 57, 73, 65, 56, 67, 106, 101, 107, 60, 62, 28, 78, 97, 116, 135, 140, 139, 138, 143, 147, 112, 75, 
    48, 25, 76, 47, 78, 91, 78, 91, 84, 78, 61, 70, 62, 53, 66, 82, 97, 101, 63, 61, 43, 78, 91, 113, 129, 139, 136, 136, 139, 144, 106, 70, 
    37, 17, 74, 47, 90, 105, 101, 95, 111, 77, 48, 26, 36, 67, 78, 88, 99, 104, 85, 83, 60, 85, 108, 119, 112, 117, 113, 116, 129, 133, 90, 55, 
    25, 6, 76, 48, 86, 100, 112, 95, 126, 83, 40, 1, 23, 66, 85, 107, 113, 120, 98, 80, 59, 85, 85, 101, 104, 104, 105, 112, 122, 122, 71, 45, 
    17, 0, 84, 58, 82, 94, 103, 87, 114, 95, 59, 39, 49, 97, 113, 121, 124, 130, 114, 112, 89, 75, 72, 94, 101, 107, 114, 117, 119, 109, 56, 34, 
    19, 0, 97, 77, 77, 94, 96, 86, 89, 115, 100, 77, 91, 99, 117, 124, 124, 120, 116, 110, 107, 95, 89, 100, 111, 127, 129, 124, 114, 97, 44, 27, 
    24, 0, 105, 91, 77, 97, 100, 96, 63, 86, 103, 94, 113, 116, 109, 103, 111, 108, 90, 79, 88, 102, 103, 110, 125, 128, 133, 119, 104, 94, 48, 32, 
    22, 0, 95, 98, 75, 92, 93, 113, 95, 114, 125, 132, 120, 95, 80, 73, 107, 120, 108, 92, 99, 118, 141, 141, 131, 117, 110, 98, 97, 100, 66, 41, 
    4, 0, 71, 98, 81, 103, 92, 98, 59, 108, 123, 105, 96, 55, 38, 24, 44, 91, 125, 137, 141, 139, 147, 140, 130, 113, 106, 104, 106, 111, 94, 57, 
    0, 0, 31, 68, 80, 116, 87, 83, 30, 51, 64, 73, 61, 14, 3, 12, 38, 68, 101, 120, 135, 144, 140, 127, 119, 108, 104, 106, 113, 122, 119, 73, 
    0, 0, 1, 38, 53, 88, 78, 62, 21, 24, 48, 65, 59, 35, 32, 45, 68, 92, 113, 124, 128, 122, 116, 113, 111, 115, 116, 120, 121, 124, 133, 88, 
    15, 0, 2, 14, 36, 54, 52, 21, 25, 34, 67, 94, 105, 95, 92, 101, 110, 120, 124, 122, 120, 118, 117, 116, 117, 117, 119, 123, 123, 128, 146, 96, 
    56, 45, 45, 20, 18, 17, 14, 1, 43, 54, 94, 121, 122, 119, 119, 120, 125, 127, 128, 125, 122, 122, 119, 117, 114, 112, 112, 113, 117, 121, 128, 86, 
    71, 72, 95, 51, 2, 0, 0, 0, 79, 91, 127, 128, 124, 122, 121, 120, 121, 124, 123, 121, 118, 111, 109, 108, 109, 106, 103, 103, 104, 94, 106, 70, 
    68, 81, 119, 81, 16, 0, 0, 0, 80, 122, 132, 123, 126, 129, 131, 123, 118, 116, 116, 114, 111, 106, 101, 99, 105, 112, 112, 111, 107, 97, 106, 57, 
    68, 78, 126, 97, 50, 0, 0, 9, 83, 130, 119, 111, 115, 123, 127, 126, 123, 119, 117, 117, 118, 113, 106, 107, 116, 122, 125, 135, 141, 118, 109, 66, 
    67, 73, 125, 106, 79, 51, 41, 64, 101, 122, 109, 96, 95, 103, 110, 112, 112, 115, 122, 131, 133, 128, 119, 118, 116, 117, 128, 151, 163, 143, 137, 85, 
    55, 39, 90, 82, 76, 68, 72, 80, 94, 105, 93, 82, 76, 78, 77, 80, 82, 84, 90, 97, 102, 107, 100, 91, 82, 74, 86, 108, 120, 113, 121, 77, 
    32, 26, 55, 53, 52, 54, 58, 63, 65, 65, 61, 56, 52, 53, 50, 46, 40, 37, 42, 52, 60, 65, 60, 50, 35, 25, 36, 55, 69, 67, 74, 46, 
    
    -- channel=3
    0, 31, 27, 39, 42, 35, 36, 40, 39, 38, 34, 32, 33, 32, 35, 41, 46, 45, 40, 36, 35, 29, 24, 23, 29, 33, 33, 32, 35, 40, 50, 99, 
    0, 17, 14, 33, 39, 29, 31, 38, 39, 37, 30, 31, 28, 21, 28, 39, 46, 51, 44, 40, 37, 24, 8, 0, 7, 14, 22, 29, 36, 47, 87, 167, 
    0, 3, 0, 9, 16, 6, 10, 18, 19, 14, 5, 24, 27, 1, 2, 19, 30, 38, 30, 25, 23, 13, 0, 0, 0, 0, 0, 0, 13, 30, 89, 185, 
    0, 4, 0, 5, 15, 7, 11, 18, 16, 1, 0, 34, 71, 21, 1, 20, 32, 29, 17, 16, 26, 24, 9, 0, 0, 0, 0, 0, 0, 20, 86, 189, 
    0, 13, 0, 0, 3, 5, 10, 18, 12, 0, 0, 27, 104, 52, 19, 18, 25, 3, 0, 0, 17, 20, 17, 5, 0, 0, 0, 0, 0, 3, 81, 190, 
    0, 43, 0, 0, 0, 0, 9, 17, 15, 0, 0, 3, 84, 74, 52, 29, 21, 0, 0, 0, 10, 17, 9, 0, 11, 24, 0, 0, 0, 0, 75, 191, 
    0, 91, 0, 0, 0, 0, 8, 16, 20, 14, 0, 10, 53, 84, 84, 34, 3, 0, 0, 0, 14, 40, 13, 0, 20, 54, 23, 0, 0, 0, 64, 192, 
    0, 146, 0, 0, 0, 0, 0, 10, 31, 65, 48, 4, 18, 75, 90, 25, 0, 0, 0, 0, 10, 66, 33, 0, 19, 51, 42, 0, 0, 0, 45, 190, 
    0, 155, 0, 0, 0, 0, 0, 0, 16, 93, 89, 0, 0, 68, 79, 31, 0, 0, 0, 0, 0, 70, 58, 22, 10, 32, 43, 18, 0, 0, 15, 177, 
    0, 128, 0, 0, 6, 1, 0, 0, 0, 100, 112, 0, 0, 77, 76, 42, 16, 14, 0, 0, 0, 56, 76, 46, 0, 9, 40, 43, 0, 0, 0, 143, 
    0, 82, 0, 0, 32, 18, 0, 0, 0, 54, 96, 0, 0, 94, 82, 46, 41, 38, 0, 0, 0, 52, 80, 58, 0, 0, 29, 48, 32, 0, 0, 103, 
    0, 51, 0, 0, 38, 15, 9, 0, 0, 0, 76, 0, 0, 96, 102, 45, 51, 53, 0, 0, 2, 74, 80, 56, 0, 0, 14, 37, 38, 0, 3, 89, 
    0, 38, 0, 25, 39, 0, 12, 28, 0, 0, 27, 0, 0, 80, 113, 50, 51, 53, 0, 0, 29, 96, 89, 53, 0, 0, 0, 13, 25, 6, 22, 101, 
    0, 33, 0, 66, 58, 0, 0, 64, 0, 0, 0, 0, 0, 58, 89, 38, 47, 42, 0, 0, 47, 98, 77, 40, 0, 0, 0, 0, 15, 11, 38, 127, 
    0, 33, 0, 101, 101, 0, 0, 56, 0, 0, 0, 0, 17, 48, 51, 25, 43, 24, 0, 0, 44, 90, 75, 45, 0, 0, 0, 0, 8, 8, 45, 151, 
    0, 46, 0, 95, 135, 0, 0, 46, 24, 0, 0, 0, 66, 64, 10, 12, 31, 2, 0, 0, 14, 69, 78, 45, 0, 0, 0, 0, 0, 0, 49, 175, 
    0, 68, 0, 57, 146, 20, 0, 21, 42, 0, 0, 0, 53, 65, 10, 14, 11, 0, 0, 0, 0, 37, 85, 58, 0, 0, 0, 0, 0, 0, 56, 197, 
    0, 87, 0, 19, 132, 56, 0, 0, 51, 0, 0, 0, 6, 32, 8, 34, 14, 0, 0, 0, 0, 7, 75, 58, 0, 0, 0, 0, 0, 0, 70, 210, 
    0, 89, 0, 0, 107, 88, 0, 0, 43, 19, 6, 0, 0, 1, 0, 61, 44, 0, 0, 30, 13, 25, 57, 33, 0, 0, 0, 0, 0, 0, 80, 213, 
    0, 73, 0, 0, 82, 101, 0, 0, 55, 72, 58, 0, 0, 0, 0, 74, 91, 0, 0, 24, 34, 51, 41, 0, 0, 0, 0, 0, 0, 3, 77, 195, 
    0, 48, 9, 0, 69, 104, 0, 0, 53, 118, 76, 0, 0, 0, 0, 65, 108, 25, 0, 23, 43, 42, 14, 0, 0, 0, 0, 0, 6, 13, 69, 162, 
    0, 18, 22, 0, 62, 89, 0, 0, 35, 149, 110, 0, 0, 0, 0, 52, 102, 65, 26, 27, 21, 12, 0, 0, 0, 0, 0, 0, 19, 20, 58, 121, 
    0, 0, 7, 0, 50, 44, 0, 0, 28, 150, 131, 11, 0, 0, 0, 30, 69, 59, 37, 25, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 32, 81, 
    0, 0, 0, 0, 35, 0, 0, 0, 62, 157, 142, 30, 0, 0, 0, 10, 28, 27, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 78, 
    0, 0, 0, 0, 0, 0, 0, 0, 144, 174, 113, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 84, 
    0, 5, 0, 0, 0, 0, 0, 92, 200, 159, 49, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 95, 
    0, 38, 0, 0, 0, 0, 0, 168, 212, 103, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 101, 
    0, 49, 0, 0, 0, 0, 0, 182, 180, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 82, 
    0, 48, 0, 0, 0, 0, 0, 128, 132, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 25, 57, 
    0, 52, 0, 0, 0, 0, 0, 50, 75, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 12, 22, 37, 
    0, 47, 0, 0, 0, 0, 0, 5, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 31, 8, 19, 33, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 29, 24, 0, 11, 26, 
    
    -- channel=4
    71, 90, 93, 91, 90, 93, 94, 93, 93, 92, 89, 91, 93, 95, 97, 95, 92, 90, 88, 87, 84, 84, 85, 86, 85, 83, 79, 76, 74, 71, 60, 11, 
    48, 89, 89, 85, 86, 91, 95, 96, 97, 98, 96, 89, 82, 87, 95, 98, 97, 90, 85, 81, 74, 65, 62, 66, 73, 80, 87, 88, 87, 87, 77, 35, 
    55, 89, 90, 84, 85, 90, 95, 95, 98, 108, 121, 110, 85, 80, 90, 90, 83, 82, 83, 84, 81, 67, 53, 42, 43, 56, 71, 86, 94, 94, 78, 37, 
    57, 90, 95, 91, 88, 90, 93, 93, 94, 102, 121, 132, 108, 82, 76, 69, 57, 53, 74, 97, 103, 97, 83, 69, 55, 47, 58, 76, 93, 96, 77, 36, 
    47, 70, 83, 97, 101, 95, 91, 91, 92, 85, 81, 83, 75, 60, 44, 33, 29, 46, 73, 88, 87, 85, 86, 86, 80, 65, 44, 58, 79, 92, 77, 35, 
    34, 37, 40, 67, 98, 103, 97, 96, 98, 88, 62, 54, 63, 62, 51, 49, 58, 64, 69, 83, 78, 64, 55, 66, 75, 63, 43, 43, 59, 79, 74, 33, 
    44, 40, 39, 74, 93, 98, 98, 100, 102, 91, 75, 77, 94, 95, 81, 82, 90, 65, 44, 62, 79, 66, 45, 50, 54, 55, 47, 32, 46, 66, 69, 34, 
    66, 80, 83, 112, 103, 96, 102, 118, 125, 107, 78, 89, 105, 95, 75, 64, 66, 49, 27, 36, 59, 67, 56, 40, 43, 55, 58, 36, 29, 51, 63, 38, 
    67, 103, 119, 131, 101, 95, 103, 136, 170, 164, 127, 114, 95, 74, 61, 50, 49, 36, 21, 43, 65, 76, 67, 53, 55, 66, 71, 55, 26, 33, 44, 34, 
    54, 89, 112, 122, 98, 84, 79, 83, 112, 135, 121, 95, 83, 59, 53, 55, 52, 37, 36, 73, 89, 90, 73, 61, 64, 78, 74, 67, 39, 29, 33, 24, 
    51, 67, 86, 100, 95, 86, 72, 36, 24, 43, 57, 63, 87, 72, 59, 57, 62, 50, 44, 85, 98, 83, 62, 47, 54, 69, 72, 74, 62, 43, 36, 19, 
    59, 50, 71, 81, 80, 85, 84, 18, 2, 19, 30, 47, 90, 95, 74, 67, 76, 69, 48, 76, 83, 63, 46, 42, 48, 56, 65, 72, 75, 64, 49, 16, 
    67, 48, 77, 66, 49, 63, 94, 47, 19, 38, 59, 76, 90, 101, 96, 85, 74, 65, 41, 70, 76, 60, 46, 46, 46, 54, 65, 74, 75, 72, 61, 26, 
    75, 54, 85, 70, 37, 52, 85, 74, 39, 53, 95, 110, 79, 71, 70, 81, 72, 54, 23, 62, 78, 67, 63, 65, 66, 72, 77, 78, 74, 72, 70, 33, 
    81, 58, 84, 89, 58, 62, 86, 97, 64, 76, 93, 105, 93, 58, 47, 57, 55, 51, 30, 55, 67, 68, 59, 44, 50, 62, 65, 66, 69, 72, 75, 36, 
    83, 60, 83, 107, 86, 72, 88, 108, 84, 56, 38, 48, 49, 41, 45, 44, 52, 59, 35, 41, 63, 76, 68, 49, 37, 39, 45, 52, 64, 79, 79, 35, 
    84, 69, 85, 103, 94, 60, 73, 108, 97, 44, 16, 10, 26, 33, 47, 55, 59, 79, 65, 41, 27, 46, 51, 39, 25, 25, 41, 61, 79, 91, 81, 34, 
    76, 76, 90, 94, 100, 54, 56, 84, 103, 75, 23, 17, 46, 77, 101, 88, 58, 72, 90, 71, 52, 35, 19, 21, 28, 36, 59, 78, 89, 89, 74, 34, 
    65, 78, 91, 88, 102, 64, 53, 69, 83, 79, 55, 47, 66, 93, 116, 106, 65, 51, 64, 85, 79, 48, 27, 34, 47, 69, 86, 96, 92, 85, 73, 36, 
    58, 82, 92, 87, 90, 71, 64, 105, 97, 63, 50, 50, 81, 98, 113, 118, 82, 48, 26, 28, 29, 29, 38, 43, 47, 62, 73, 91, 93, 90, 76, 40, 
    53, 83, 96, 90, 80, 66, 65, 125, 167, 144, 106, 98, 109, 106, 100, 111, 111, 81, 56, 32, 25, 49, 70, 74, 67, 64, 67, 75, 83, 88, 73, 34, 
    34, 77, 103, 105, 92, 85, 84, 119, 155, 154, 138, 93, 64, 35, 28, 34, 49, 61, 70, 77, 85, 86, 84, 76, 71, 70, 72, 80, 88, 88, 73, 43, 
    0, 32, 66, 90, 100, 122, 110, 120, 104, 80, 46, 24, 0, 0, 0, 0, 7, 27, 45, 60, 73, 74, 65, 58, 56, 58, 65, 74, 79, 79, 77, 47, 
    0, 5, 9, 42, 74, 103, 95, 109, 74, 33, 19, 15, 15, 21, 22, 26, 37, 43, 50, 53, 54, 50, 47, 50, 53, 57, 60, 61, 63, 66, 75, 42, 
    15, 24, 1, 13, 47, 75, 88, 91, 45, 16, 40, 49, 51, 51, 47, 47, 49, 49, 48, 48, 51, 53, 54, 55, 57, 59, 55, 58, 67, 74, 91, 55, 
    32, 44, 18, 10, 23, 47, 89, 83, 40, 31, 46, 51, 50, 44, 40, 42, 47, 50, 51, 53, 53, 56, 58, 57, 51, 44, 42, 49, 62, 68, 82, 55, 
    36, 53, 36, 22, 2, 0, 63, 75, 63, 57, 59, 53, 51, 49, 42, 41, 45, 49, 51, 51, 49, 45, 43, 43, 43, 42, 43, 48, 54, 43, 48, 34, 
    37, 57, 51, 33, 0, 0, 11, 52, 62, 55, 49, 49, 58, 60, 55, 48, 43, 43, 45, 46, 44, 38, 33, 34, 43, 55, 60, 57, 48, 27, 30, 19, 
    40, 58, 54, 39, 11, 0, 0, 24, 33, 40, 26, 28, 41, 50, 52, 51, 51, 54, 56, 52, 49, 43, 35, 39, 55, 74, 79, 74, 69, 47, 34, 24, 
    39, 53, 48, 40, 28, 12, 25, 43, 36, 33, 24, 17, 19, 20, 25, 29, 38, 49, 60, 67, 65, 53, 42, 44, 58, 75, 85, 85, 80, 62, 48, 28, 
    1, 14, 2, 0, 0, 0, 2, 19, 16, 9, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 23, 16, 9, 1, 1, 11, 29, 37, 30, 14, 25, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    87, 64, 29, 25, 13, 14, 20, 16, 14, 15, 20, 23, 20, 22, 24, 23, 19, 16, 17, 17, 14, 16, 22, 27, 24, 16, 13, 14, 18, 15, 3, 0, 
    226, 262, 237, 235, 221, 219, 221, 217, 213, 209, 211, 213, 216, 224, 231, 228, 217, 207, 204, 208, 207, 205, 215, 226, 232, 224, 211, 199, 189, 174, 132, 20, 
    223, 246, 222, 225, 215, 216, 220, 216, 211, 208, 205, 189, 162, 174, 211, 219, 213, 203, 197, 189, 157, 123, 126, 160, 199, 225, 231, 216, 196, 176, 137, 25, 
    222, 244, 217, 225, 219, 221, 227, 223, 219, 227, 252, 235, 157, 145, 204, 228, 224, 213, 195, 153, 88, 33, 17, 40, 86, 137, 193, 224, 222, 197, 149, 28, 
    220, 248, 235, 254, 248, 233, 229, 224, 221, 240, 300, 333, 242, 167, 185, 204, 187, 160, 145, 129, 72, 30, 10, 10, 25, 50, 110, 197, 234, 219, 159, 29, 
    208, 218, 215, 273, 282, 245, 225, 218, 214, 232, 275, 312, 257, 155, 98, 75, 69, 68, 109, 127, 100, 61, 58, 67, 58, 41, 52, 133, 216, 235, 178, 32, 
    160, 113, 78, 194, 258, 246, 224, 221, 211, 198, 200, 208, 185, 103, 21, 0, 24, 47, 110, 175, 164, 91, 69, 99, 104, 55, 25, 68, 174, 235, 199, 42, 
    111, 0, 0, 78, 178, 215, 218, 219, 201, 142, 94, 115, 142, 103, 29, 14, 52, 81, 128, 209, 230, 136, 55, 72, 98, 62, 4, 14, 109, 214, 212, 59, 
    121, 0, 0, 53, 136, 174, 206, 235, 218, 105, 0, 22, 117, 112, 48, 23, 47, 77, 115, 181, 210, 132, 32, 15, 42, 43, 0, 0, 36, 159, 215, 86, 
    145, 38, 0, 95, 144, 151, 189, 270, 312, 237, 80, 59, 132, 104, 38, 7, 17, 30, 64, 128, 149, 85, 23, 0, 28, 52, 18, 0, 0, 71, 167, 94, 
    159, 74, 71, 156, 159, 134, 171, 264, 393, 396, 263, 162, 183, 104, 10, 0, 0, 0, 14, 116, 144, 90, 56, 33, 55, 90, 57, 2, 0, 0, 75, 56, 
    152, 68, 96, 174, 169, 148, 174, 199, 302, 376, 298, 218, 222, 135, 0, 0, 0, 0, 0, 137, 185, 124, 76, 50, 66, 104, 94, 41, 0, 0, 15, 0, 
    143, 52, 76, 143, 148, 180, 200, 166, 198, 300, 267, 221, 232, 185, 52, 6, 22, 0, 27, 169, 197, 122, 46, 24, 40, 81, 94, 63, 13, 0, 13, 0, 
    138, 47, 65, 103, 68, 151, 225, 174, 150, 242, 241, 201, 190, 191, 141, 98, 76, 48, 75, 198, 197, 108, 31, 11, 23, 53, 68, 68, 51, 49, 60, 0, 
    145, 60, 66, 74, 0, 52, 198, 176, 122, 198, 245, 244, 192, 168, 174, 170, 141, 93, 117, 220, 222, 125, 46, 22, 38, 75, 92, 110, 118, 114, 111, 16, 
    150, 65, 58, 62, 0, 0, 139, 165, 108, 181, 287, 319, 270, 185, 176, 185, 159, 118, 151, 236, 250, 186, 89, 35, 53, 111, 144, 161, 166, 156, 135, 22, 
    159, 66, 41, 65, 0, 0, 97, 166, 107, 136, 276, 326, 304, 204, 140, 131, 108, 115, 157, 209, 242, 232, 142, 66, 75, 129, 165, 176, 169, 164, 147, 24, 
    183, 94, 41, 72, 5, 0, 36, 163, 122, 73, 138, 201, 207, 152, 91, 53, 19, 95, 170, 145, 130, 170, 157, 99, 82, 102, 135, 171, 174, 178, 163, 32, 
    215, 151, 69, 82, 31, 0, 0, 121, 122, 70, 52, 95, 160, 143, 96, 29, 0, 47, 178, 160, 106, 102, 100, 66, 46, 72, 123, 185, 201, 197, 173, 38, 
    232, 202, 104, 98, 69, 0, 0, 58, 30, 0, 0, 8, 89, 100, 84, 23, 0, 0, 121, 186, 157, 105, 38, 1, 4, 59, 138, 209, 218, 199, 170, 42, 
    217, 208, 115, 99, 85, 3, 0, 38, 0, 0, 0, 0, 0, 42, 85, 71, 0, 0, 15, 61, 50, 2, 0, 0, 0, 0, 76, 142, 160, 134, 100, 0, 
    182, 186, 119, 95, 72, 0, 0, 57, 29, 0, 0, 0, 23, 127, 175, 177, 97, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    127, 150, 140, 118, 76, 0, 1, 119, 138, 85, 0, 7, 90, 134, 143, 129, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 33, 97, 142, 124, 86, 115, 185, 169, 101, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 77, 139, 141, 185, 195, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 67, 135, 189, 144, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 110, 200, 129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 176, 145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 42, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    51, 19, 0, 0, 0, 0, 6, 9, 4, 0, 0, 0, 0, 0, 0, 11, 31, 48, 58, 60, 45, 25, 18, 27, 59, 91, 101, 69, 16, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 136, 87, 94, 85, 75, 81, 78, 74, 66, 63, 76, 85, 82, 82, 77, 72, 73, 78, 90, 99, 101, 103, 104, 104, 90, 79, 63, 47, 36, 0, 0, 
    0, 95, 38, 48, 45, 41, 51, 49, 42, 28, 11, 31, 43, 27, 41, 54, 53, 53, 48, 34, 29, 25, 32, 45, 60, 67, 65, 52, 33, 15, 0, 0, 
    0, 96, 38, 50, 49, 46, 55, 56, 50, 52, 45, 82, 99, 47, 56, 81, 82, 64, 27, 18, 19, 9, 1, 0, 10, 37, 51, 60, 57, 39, 0, 0, 
    5, 123, 68, 77, 78, 57, 53, 53, 50, 80, 118, 182, 179, 85, 62, 59, 42, 9, 0, 50, 85, 84, 59, 29, 10, 20, 32, 42, 58, 60, 0, 0, 
    0, 126, 67, 78, 99, 72, 46, 43, 44, 70, 106, 155, 130, 46, 0, 0, 0, 0, 6, 82, 153, 154, 122, 95, 74, 53, 21, 14, 40, 66, 11, 0, 
    0, 74, 0, 19, 78, 81, 49, 42, 40, 43, 37, 48, 37, 5, 0, 0, 0, 22, 55, 116, 176, 167, 114, 100, 99, 60, 15, 0, 12, 55, 28, 6, 
    0, 52, 0, 0, 62, 71, 42, 28, 12, 10, 0, 0, 29, 68, 55, 30, 52, 80, 85, 121, 163, 163, 88, 66, 68, 43, 0, 0, 0, 29, 27, 30, 
    0, 122, 0, 39, 105, 72, 44, 27, 11, 30, 7, 0, 80, 127, 86, 49, 52, 72, 49, 57, 114, 135, 71, 32, 22, 25, 0, 0, 0, 1, 15, 48, 
    24, 218, 90, 162, 177, 83, 61, 69, 125, 216, 195, 107, 130, 152, 78, 33, 29, 34, 0, 0, 95, 135, 86, 54, 24, 40, 31, 0, 0, 0, 0, 31, 
    60, 264, 174, 252, 225, 79, 65, 104, 225, 346, 364, 209, 167, 169, 81, 29, 13, 15, 0, 7, 159, 207, 139, 94, 52, 72, 67, 17, 0, 0, 0, 0, 
    61, 260, 190, 286, 257, 96, 51, 57, 126, 258, 327, 214, 171, 197, 112, 36, 13, 27, 0, 75, 248, 262, 151, 91, 57, 82, 83, 51, 10, 0, 0, 0, 
    55, 242, 162, 298, 262, 112, 59, 49, 24, 147, 221, 180, 203, 245, 176, 81, 53, 68, 1, 130, 274, 243, 115, 58, 38, 68, 74, 63, 54, 18, 0, 0, 
    48, 248, 157, 286, 225, 82, 68, 69, 0, 81, 135, 169, 259, 288, 242, 150, 111, 107, 44, 157, 271, 224, 96, 52, 29, 42, 61, 74, 92, 59, 0, 0, 
    49, 277, 182, 262, 185, 48, 55, 81, 4, 44, 135, 223, 313, 295, 230, 184, 149, 115, 62, 165, 255, 210, 114, 81, 53, 63, 97, 115, 121, 85, 2, 0, 
    52, 309, 218, 263, 199, 56, 51, 98, 50, 58, 182, 309, 371, 294, 188, 161, 132, 106, 87, 161, 223, 208, 137, 79, 55, 82, 120, 134, 114, 69, 0, 8, 
    56, 346, 261, 293, 251, 105, 75, 116, 109, 73, 174, 280, 288, 209, 115, 103, 94, 79, 95, 154, 179, 169, 155, 97, 46, 65, 85, 89, 75, 41, 0, 13, 
    69, 385, 309, 325, 287, 158, 92, 138, 151, 65, 99, 118, 131, 105, 34, 74, 79, 64, 94, 102, 72, 117, 130, 70, 11, 22, 35, 48, 62, 53, 9, 19, 
    82, 401, 344, 341, 302, 197, 95, 153, 193, 107, 78, 43, 67, 96, 55, 102, 103, 75, 110, 123, 73, 76, 48, 0, 0, 0, 26, 56, 85, 74, 17, 20, 
    75, 380, 357, 335, 313, 236, 91, 108, 176, 123, 61, 14, 51, 100, 125, 163, 130, 65, 127, 156, 116, 69, 6, 0, 0, 36, 82, 105, 119, 91, 28, 26, 
    51, 336, 358, 314, 303, 249, 100, 108, 181, 133, 27, 0, 45, 143, 233, 274, 211, 92, 69, 58, 26, 0, 0, 0, 0, 52, 101, 125, 130, 97, 44, 46, 
    42, 311, 370, 312, 282, 224, 100, 196, 325, 316, 193, 140, 200, 311, 371, 380, 320, 190, 90, 21, 0, 0, 0, 34, 69, 95, 114, 121, 119, 98, 67, 72, 
    60, 312, 380, 348, 310, 231, 144, 324, 500, 520, 400, 300, 290, 311, 322, 307, 268, 197, 125, 81, 68, 89, 118, 143, 157, 164, 163, 165, 165, 150, 129, 122, 
    49, 278, 345, 363, 368, 303, 268, 425, 540, 484, 323, 189, 161, 147, 144, 137, 132, 129, 124, 124, 136, 157, 165, 168, 178, 191, 198, 201, 202, 194, 173, 163, 
    12, 210, 250, 300, 345, 309, 339, 468, 487, 332, 180, 119, 110, 117, 118, 119, 128, 133, 133, 137, 147, 161, 169, 178, 197, 216, 226, 221, 217, 214, 194, 192, 
    16, 199, 198, 223, 256, 266, 362, 466, 399, 196, 128, 145, 166, 173, 164, 156, 151, 148, 146, 150, 163, 179, 193, 211, 233, 247, 242, 234, 241, 260, 255, 241, 
    41, 229, 196, 187, 214, 260, 383, 475, 331, 126, 127, 162, 183, 175, 160, 156, 155, 156, 162, 174, 190, 208, 229, 247, 250, 235, 217, 224, 267, 316, 309, 259, 
    43, 240, 209, 186, 200, 262, 374, 459, 322, 138, 160, 179, 187, 183, 165, 156, 158, 167, 179, 192, 207, 219, 227, 234, 229, 209, 202, 236, 295, 316, 269, 210, 
    42, 248, 225, 208, 201, 227, 302, 355, 285, 153, 168, 189, 205, 207, 195, 175, 160, 164, 178, 196, 209, 212, 212, 205, 197, 201, 235, 283, 295, 256, 195, 150, 
    48, 259, 233, 219, 206, 191, 201, 216, 180, 129, 132, 159, 189, 208, 209, 196, 186, 191, 201, 216, 221, 213, 200, 186, 190, 232, 295, 331, 304, 237, 176, 131, 
    80, 272, 261, 246, 241, 216, 193, 181, 160, 134, 133, 145, 160, 172, 183, 192, 206, 228, 251, 275, 277, 251, 227, 221, 249, 313, 378, 394, 343, 263, 201, 138, 
    70, 205, 204, 191, 189, 179, 162, 140, 127, 109, 101, 101, 102, 101, 99, 100, 118, 156, 198, 228, 229, 205, 186, 188, 221, 280, 323, 314, 255, 189, 147, 84, 
    
    -- channel=7
    159, 128, 133, 126, 130, 135, 131, 130, 130, 129, 130, 132, 137, 141, 137, 130, 125, 121, 119, 113, 111, 113, 116, 117, 113, 111, 112, 112, 104, 94, 38, 0, 
    167, 116, 120, 109, 112, 120, 117, 115, 113, 116, 118, 119, 124, 127, 122, 114, 102, 94, 89, 81, 75, 80, 89, 94, 97, 97, 98, 99, 95, 84, 10, 0, 
    175, 115, 127, 117, 119, 125, 123, 119, 120, 135, 138, 130, 133, 139, 122, 105, 90, 77, 75, 69, 68, 75, 86, 93, 96, 103, 104, 103, 98, 90, 17, 0, 
    175, 116, 131, 122, 119, 123, 120, 117, 121, 152, 163, 128, 118, 130, 107, 75, 58, 58, 68, 75, 77, 78, 84, 91, 94, 107, 117, 116, 105, 92, 17, 0, 
    157, 102, 128, 127, 117, 119, 119, 116, 120, 143, 156, 90, 60, 70, 65, 43, 37, 74, 91, 85, 81, 81, 84, 89, 88, 85, 113, 127, 114, 100, 20, 0, 
    118, 56, 120, 133, 124, 118, 122, 119, 117, 115, 121, 84, 53, 38, 47, 60, 62, 99, 117, 88, 84, 85, 87, 81, 61, 55, 85, 128, 128, 108, 21, 0, 
    82, 19, 121, 161, 144, 129, 125, 121, 107, 101, 108, 107, 86, 54, 57, 77, 68, 93, 137, 108, 78, 81, 97, 85, 48, 30, 47, 104, 136, 115, 26, 0, 
    68, 24, 136, 184, 158, 149, 137, 136, 112, 93, 119, 138, 118, 72, 53, 65, 64, 78, 133, 122, 73, 65, 81, 84, 56, 27, 25, 66, 133, 127, 29, 0, 
    63, 34, 158, 190, 173, 159, 154, 174, 153, 118, 153, 175, 135, 79, 55, 62, 61, 66, 116, 131, 94, 68, 68, 84, 79, 48, 26, 39, 101, 136, 32, 0, 
    67, 50, 149, 177, 172, 148, 150, 203, 174, 119, 125, 163, 125, 91, 71, 61, 50, 63, 130, 140, 119, 92, 73, 79, 89, 61, 39, 26, 56, 123, 42, 0, 
    64, 76, 143, 161, 163, 141, 112, 178, 157, 78, 99, 160, 130, 91, 86, 66, 40, 65, 161, 154, 112, 105, 70, 66, 89, 68, 51, 31, 39, 88, 57, 0, 
    53, 89, 146, 139, 160, 146, 83, 118, 171, 89, 106, 173, 141, 86, 92, 96, 50, 70, 177, 159, 82, 92, 64, 62, 85, 78, 58, 42, 40, 73, 53, 0, 
    50, 103, 135, 108, 153, 155, 81, 79, 156, 112, 116, 190, 178, 109, 93, 107, 67, 72, 173, 148, 71, 79, 59, 56, 70, 84, 70, 58, 58, 84, 46, 0, 
    61, 118, 122, 61, 146, 174, 103, 62, 124, 150, 150, 170, 173, 118, 101, 92, 70, 81, 166, 137, 72, 82, 62, 64, 79, 95, 100, 87, 82, 101, 47, 0, 
    69, 121, 125, 34, 111, 185, 138, 75, 122, 177, 190, 160, 134, 133, 120, 90, 67, 90, 160, 135, 81, 77, 55, 56, 80, 89, 102, 98, 92, 112, 49, 0, 
    75, 112, 142, 43, 65, 173, 169, 101, 120, 170, 176, 108, 71, 94, 97, 88, 82, 101, 144, 138, 91, 71, 48, 57, 85, 90, 91, 100, 107, 124, 45, 0, 
    80, 94, 153, 71, 25, 135, 175, 111, 102, 154, 137, 79, 52, 67, 86, 86, 110, 122, 130, 114, 108, 58, 27, 38, 61, 80, 89, 111, 133, 139, 46, 0, 
    88, 74, 149, 98, 18, 91, 172, 124, 100, 112, 125, 102, 87, 98, 90, 71, 126, 149, 118, 98, 112, 70, 14, 17, 51, 93, 119, 133, 144, 138, 40, 0, 
    103, 65, 139, 122, 38, 57, 146, 117, 92, 84, 105, 140, 121, 127, 104, 48, 101, 167, 120, 94, 72, 47, 26, 31, 68, 119, 155, 155, 139, 128, 33, 0, 
    122, 69, 134, 135, 61, 53, 141, 107, 72, 74, 73, 120, 124, 143, 129, 48, 63, 128, 111, 50, 12, 5, 17, 24, 64, 113, 156, 148, 125, 115, 31, 0, 
    135, 71, 129, 136, 67, 60, 163, 142, 75, 73, 103, 147, 166, 175, 149, 77, 46, 75, 76, 34, 13, 3, 6, 20, 52, 86, 117, 103, 86, 75, 14, 0, 
    132, 63, 115, 128, 71, 84, 196, 195, 111, 78, 88, 122, 117, 111, 85, 38, 8, 11, 21, 21, 12, 8, 3, 2, 8, 24, 43, 36, 22, 17, 0, 0, 
    87, 46, 88, 109, 101, 133, 214, 200, 106, 34, 0, 33, 28, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 19, 71, 78, 99, 161, 202, 152, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 58, 55, 87, 176, 179, 90, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 49, 94, 174, 125, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 95, 157, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 45, 129, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 53, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 8, 13, 17, 15, 13, 14, 16, 16, 15, 13, 13, 13, 18, 20, 22, 22, 18, 18, 19, 17, 11, 9, 8, 10, 11, 11, 14, 17, 17, 41, 16, 
    0, 95, 117, 129, 126, 118, 120, 125, 122, 115, 111, 113, 121, 129, 130, 132, 132, 130, 126, 126, 118, 109, 103, 105, 108, 108, 106, 104, 107, 109, 155, 107, 
    0, 40, 52, 68, 67, 62, 67, 73, 71, 54, 41, 52, 64, 75, 74, 77, 87, 81, 59, 33, 22, 18, 16, 24, 30, 39, 45, 51, 55, 61, 123, 95, 
    0, 44, 55, 68, 66, 64, 71, 75, 69, 47, 48, 93, 101, 74, 73, 84, 82, 59, 22, 4, 10, 2, 0, 0, 0, 0, 20, 35, 45, 56, 128, 100, 
    0, 56, 58, 64, 56, 58, 72, 74, 65, 40, 59, 147, 157, 89, 63, 62, 41, 7, 0, 2, 32, 50, 37, 8, 0, 0, 0, 1, 23, 48, 124, 101, 
    0, 56, 42, 34, 45, 55, 69, 71, 60, 25, 32, 105, 131, 73, 32, 19, 0, 0, 0, 0, 51, 68, 70, 57, 48, 29, 0, 0, 0, 36, 122, 100, 
    0, 36, 0, 0, 18, 63, 71, 70, 67, 49, 31, 38, 51, 64, 46, 5, 0, 0, 0, 13, 65, 58, 49, 50, 68, 59, 13, 0, 0, 16, 119, 98, 
    0, 44, 0, 0, 1, 62, 66, 55, 56, 56, 39, 16, 38, 91, 86, 44, 28, 15, 0, 3, 74, 77, 35, 28, 49, 56, 26, 0, 0, 0, 107, 95, 
    0, 76, 0, 0, 28, 61, 49, 26, 32, 65, 40, 5, 51, 102, 91, 43, 28, 22, 0, 0, 29, 79, 55, 18, 22, 38, 35, 4, 0, 0, 90, 95, 
    0, 92, 2, 22, 77, 72, 41, 22, 77, 166, 102, 36, 68, 106, 90, 46, 24, 9, 0, 0, 0, 74, 95, 45, 15, 26, 52, 38, 0, 0, 56, 81, 
    0, 69, 16, 58, 96, 85, 33, 5, 54, 187, 173, 84, 80, 101, 86, 65, 47, 9, 0, 0, 29, 98, 118, 73, 24, 28, 53, 57, 15, 0, 14, 55, 
    0, 29, 0, 73, 103, 97, 48, 0, 0, 86, 106, 42, 63, 120, 92, 69, 74, 22, 0, 0, 80, 119, 114, 61, 14, 21, 49, 56, 36, 0, 16, 36, 
    0, 12, 0, 73, 94, 89, 81, 29, 0, 8, 37, 0, 44, 148, 121, 67, 95, 52, 0, 0, 91, 114, 91, 43, 1, 0, 17, 42, 48, 32, 58, 44, 
    0, 12, 0, 85, 60, 39, 87, 61, 0, 0, 0, 0, 35, 146, 148, 84, 98, 59, 0, 0, 92, 99, 76, 37, 0, 0, 0, 24, 52, 49, 89, 67, 
    0, 16, 15, 116, 47, 0, 52, 60, 4, 0, 0, 11, 67, 92, 103, 89, 95, 42, 0, 0, 95, 105, 88, 60, 20, 0, 0, 34, 58, 47, 98, 80, 
    0, 21, 20, 129, 72, 0, 15, 65, 14, 0, 4, 85, 142, 81, 39, 50, 68, 29, 0, 2, 87, 97, 75, 51, 25, 11, 19, 34, 42, 34, 98, 93, 
    0, 32, 7, 116, 111, 7, 0, 54, 24, 0, 0, 64, 111, 66, 17, 16, 22, 2, 0, 10, 62, 89, 109, 62, 13, 0, 0, 10, 14, 19, 116, 106, 
    0, 52, 0, 87, 126, 33, 0, 56, 48, 0, 0, 4, 25, 11, 2, 9, 7, 0, 6, 0, 0, 57, 103, 55, 0, 0, 0, 0, 11, 32, 139, 117, 
    0, 71, 0, 62, 124, 55, 0, 30, 65, 48, 8, 0, 0, 0, 6, 57, 23, 0, 49, 52, 6, 14, 41, 12, 0, 0, 0, 0, 37, 58, 150, 119, 
    0, 70, 10, 47, 119, 77, 0, 0, 35, 74, 48, 0, 0, 0, 28, 112, 62, 0, 46, 90, 81, 46, 4, 0, 0, 0, 0, 21, 58, 62, 136, 109, 
    0, 56, 16, 37, 111, 81, 0, 0, 25, 41, 14, 0, 0, 0, 30, 136, 104, 11, 0, 4, 21, 10, 0, 0, 0, 0, 0, 6, 35, 31, 104, 94, 
    0, 46, 19, 19, 84, 46, 0, 0, 122, 161, 85, 33, 13, 34, 71, 133, 141, 74, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 53, 
    0, 37, 25, 21, 71, 24, 0, 0, 159, 251, 184, 82, 33, 32, 31, 46, 55, 45, 35, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 29, 
    0, 0, 0, 26, 66, 17, 0, 17, 131, 167, 102, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 21, 
    0, 0, 0, 0, 20, 0, 0, 76, 143, 108, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 21, 
    0, 0, 0, 0, 0, 0, 0, 109, 135, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 37, 
    0, 5, 0, 0, 0, 0, 21, 151, 98, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 48, 
    0, 9, 0, 0, 0, 0, 30, 167, 85, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 33, 
    0, 6, 0, 0, 0, 0, 0, 96, 64, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 12, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 5, 4, 6, 0, 0, 0, 7, 0, 0, 0, 0, 1, 8, 13, 19, 23, 25, 29, 24, 16, 8, 0, 0, 18, 45, 45, 30, 17, 25, 9, 
    0, 67, 44, 40, 39, 40, 36, 33, 37, 35, 27, 26, 23, 18, 16, 15, 19, 32, 45, 60, 65, 55, 46, 36, 36, 52, 74, 82, 68, 47, 45, 33, 
    
    -- channel=9
    20, 72, 85, 84, 84, 85, 86, 87, 86, 86, 84, 82, 84, 88, 91, 90, 89, 87, 84, 80, 74, 69, 67, 68, 68, 69, 70, 68, 66, 64, 56, 29, 
    83, 101, 107, 99, 101, 108, 110, 109, 110, 111, 109, 109, 110, 109, 111, 110, 108, 108, 100, 90, 82, 77, 74, 73, 73, 76, 83, 89, 86, 81, 56, 11, 
    103, 124, 134, 125, 127, 133, 135, 135, 132, 133, 140, 148, 148, 134, 133, 131, 127, 115, 108, 100, 95, 92, 91, 89, 81, 82, 86, 97, 105, 105, 73, 16, 
    103, 123, 133, 127, 132, 136, 134, 135, 135, 140, 155, 152, 155, 153, 137, 121, 102, 82, 75, 82, 79, 74, 77, 80, 87, 89, 85, 88, 98, 106, 73, 13, 
    104, 116, 123, 116, 133, 140, 134, 132, 139, 161, 170, 128, 104, 127, 113, 82, 56, 57, 74, 80, 70, 53, 45, 56, 71, 87, 91, 93, 88, 98, 75, 14, 
    102, 99, 105, 95, 112, 138, 136, 133, 142, 173, 178, 106, 60, 83, 80, 54, 45, 68, 92, 85, 74, 56, 38, 42, 47, 53, 67, 91, 88, 85, 68, 15, 
    84, 72, 88, 104, 114, 131, 136, 135, 140, 149, 142, 99, 78, 66, 61, 59, 59, 75, 94, 81, 70, 69, 64, 53, 37, 21, 39, 70, 89, 79, 55, 13, 
    54, 25, 79, 133, 144, 140, 138, 133, 139, 135, 120, 111, 108, 83, 63, 65, 52, 57, 83, 89, 60, 58, 77, 68, 32, 11, 21, 46, 81, 81, 44, 9, 
    46, 0, 81, 140, 143, 154, 144, 143, 148, 149, 145, 158, 131, 82, 56, 63, 52, 39, 65, 92, 73, 56, 68, 65, 39, 22, 16, 30, 65, 84, 34, 0, 
    48, 4, 95, 120, 117, 152, 159, 176, 150, 122, 142, 162, 125, 66, 51, 51, 53, 28, 43, 94, 101, 70, 57, 58, 54, 37, 21, 18, 42, 78, 36, 0, 
    69, 22, 100, 91, 97, 140, 170, 193, 166, 90, 82, 115, 101, 72, 59, 49, 39, 27, 56, 110, 112, 80, 58, 50, 59, 46, 24, 10, 18, 57, 43, 0, 
    76, 31, 103, 76, 80, 121, 154, 173, 159, 85, 56, 110, 102, 77, 71, 60, 36, 31, 87, 133, 104, 70, 50, 47, 64, 50, 27, 14, 11, 35, 38, 3, 
    67, 31, 108, 76, 70, 105, 111, 132, 150, 101, 77, 141, 132, 77, 73, 87, 53, 37, 102, 142, 81, 52, 45, 48, 59, 49, 39, 25, 20, 28, 28, 9, 
    63, 36, 105, 58, 62, 108, 91, 103, 136, 106, 105, 171, 169, 84, 59, 92, 63, 47, 105, 124, 61, 48, 47, 46, 53, 56, 58, 50, 38, 39, 34, 12, 
    74, 49, 86, 18, 52, 124, 96, 94, 131, 135, 147, 178, 150, 103, 79, 80, 57, 50, 112, 118, 63, 50, 55, 44, 45, 56, 67, 65, 50, 61, 53, 15, 
    84, 53, 76, 0, 40, 114, 105, 93, 133, 159, 171, 141, 87, 80, 94, 75, 47, 57, 126, 129, 71, 62, 64, 51, 53, 59, 60, 60, 58, 77, 71, 16, 
    91, 49, 80, 6, 21, 84, 102, 85, 130, 155, 156, 100, 41, 47, 79, 74, 54, 72, 124, 127, 81, 56, 37, 44, 50, 48, 52, 58, 78, 106, 83, 17, 
    98, 42, 87, 21, 1, 59, 100, 66, 87, 137, 125, 77, 43, 55, 80, 87, 73, 86, 105, 119, 115, 75, 27, 16, 29, 36, 58, 81, 112, 133, 86, 13, 
    110, 44, 91, 39, 0, 38, 87, 65, 55, 90, 83, 90, 74, 80, 98, 80, 76, 98, 74, 81, 118, 78, 19, 8, 22, 47, 89, 123, 134, 132, 80, 11, 
    124, 58, 94, 63, 14, 23, 68, 70, 52, 50, 51, 72, 85, 92, 95, 47, 58, 101, 83, 57, 46, 19, 5, 11, 24, 55, 97, 126, 122, 116, 68, 5, 
    132, 67, 92, 85, 34, 15, 58, 70, 46, 33, 45, 80, 96, 120, 107, 31, 31, 78, 83, 56, 9, 0, 0, 0, 18, 40, 73, 94, 92, 95, 47, 0, 
    130, 57, 72, 89, 38, 21, 88, 106, 39, 21, 48, 90, 104, 102, 78, 12, 0, 5, 12, 2, 0, 0, 0, 0, 0, 0, 18, 30, 34, 35, 0, 0, 
    110, 31, 33, 62, 27, 40, 133, 178, 92, 25, 21, 42, 36, 21, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 0, 0, 26, 16, 64, 155, 183, 102, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 13, 77, 161, 140, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 73, 147, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 65, 84, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 24, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 1, 20, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 21, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 16, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 26, 26, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 23, 21, 17, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 13, 10, 11, 11, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 10, 11, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 17, 12, 11, 12, 12, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 6, 
    14, 6, 24, 23, 23, 25, 28, 30, 29, 36, 38, 34, 35, 33, 33, 31, 25, 18, 12, 10, 15, 22, 24, 25, 15, 0, 0, 5, 21, 31, 30, 31, 
    
    -- channel=11
    46, 165, 141, 155, 143, 135, 140, 140, 134, 127, 128, 139, 148, 149, 148, 146, 138, 126, 123, 124, 119, 114, 115, 120, 123, 119, 112, 106, 102, 93, 91, 5, 
    80, 259, 215, 242, 232, 221, 230, 230, 221, 210, 210, 230, 237, 230, 233, 236, 229, 212, 192, 183, 172, 154, 153, 167, 187, 197, 197, 189, 177, 163, 174, 53, 
    54, 239, 194, 226, 223, 216, 228, 228, 217, 205, 223, 271, 249, 199, 211, 229, 225, 198, 161, 139, 117, 92, 78, 92, 113, 138, 167, 179, 179, 169, 202, 72, 
    58, 247, 201, 232, 229, 219, 231, 231, 217, 202, 263, 380, 331, 206, 197, 213, 187, 144, 112, 127, 133, 101, 61, 34, 43, 70, 106, 144, 178, 184, 217, 80, 
    60, 245, 188, 222, 241, 225, 227, 226, 208, 186, 245, 392, 350, 187, 132, 118, 91, 48, 65, 135, 167, 147, 111, 73, 51, 36, 32, 67, 142, 194, 238, 89, 
    52, 203, 95, 143, 225, 235, 225, 225, 209, 163, 179, 278, 284, 174, 79, 31, 28, 7, 34, 144, 206, 172, 127, 109, 106, 57, 0, 0, 87, 186, 260, 100, 
    35, 155, 0, 49, 206, 236, 221, 225, 223, 182, 152, 187, 224, 200, 114, 30, 15, 8, 34, 160, 256, 201, 109, 104, 127, 77, 0, 0, 15, 144, 270, 114, 
    66, 175, 0, 28, 208, 227, 209, 222, 254, 234, 148, 126, 217, 260, 152, 37, 29, 35, 26, 121, 275, 246, 101, 65, 94, 74, 0, 0, 0, 75, 254, 131, 
    117, 246, 0, 126, 263, 220, 186, 222, 336, 387, 244, 153, 250, 285, 164, 46, 27, 27, 0, 46, 239, 278, 144, 55, 52, 69, 32, 0, 0, 0, 199, 131, 
    123, 301, 80, 246, 329, 223, 158, 198, 401, 566, 416, 225, 282, 307, 184, 74, 31, 1, 0, 19, 237, 303, 209, 93, 40, 73, 74, 9, 0, 0, 112, 100, 
    96, 285, 135, 347, 372, 236, 146, 133, 304, 550, 484, 301, 345, 356, 200, 101, 60, 0, 0, 49, 307, 345, 236, 105, 34, 86, 103, 55, 0, 0, 34, 43, 
    69, 253, 129, 392, 385, 258, 179, 103, 135, 414, 439, 286, 363, 418, 250, 118, 122, 29, 0, 98, 376, 356, 216, 90, 24, 74, 109, 88, 26, 0, 24, 2, 
    62, 244, 129, 387, 326, 228, 232, 141, 72, 264, 331, 245, 375, 485, 338, 165, 173, 81, 0, 135, 401, 343, 179, 59, 0, 32, 72, 93, 78, 41, 77, 8, 
    70, 265, 164, 385, 242, 144, 259, 187, 51, 161, 255, 263, 372, 440, 354, 225, 212, 105, 9, 173, 408, 328, 168, 68, 14, 24, 57, 111, 127, 98, 127, 37, 
    77, 297, 216, 413, 207, 60, 227, 218, 78, 113, 240, 361, 422, 367, 291, 240, 231, 114, 35, 195, 388, 306, 170, 76, 16, 36, 80, 134, 155, 124, 165, 69, 
    81, 337, 249, 439, 246, 37, 180, 264, 124, 89, 226, 390, 451, 303, 190, 182, 185, 114, 79, 191, 324, 305, 199, 75, 18, 45, 96, 140, 155, 132, 204, 94, 
    94, 382, 253, 437, 313, 60, 113, 275, 181, 73, 157, 292, 339, 234, 124, 128, 121, 98, 126, 159, 198, 247, 223, 82, 0, 11, 74, 132, 151, 155, 248, 118, 
    112, 430, 255, 407, 361, 106, 52, 263, 250, 106, 84, 142, 210, 175, 127, 141, 79, 75, 174, 149, 93, 158, 167, 32, 0, 0, 55, 140, 175, 183, 273, 128, 
    111, 461, 276, 372, 389, 164, 17, 190, 277, 187, 98, 69, 147, 168, 185, 224, 91, 41, 205, 215, 129, 89, 54, 0, 0, 0, 80, 171, 216, 206, 279, 129, 
    83, 459, 309, 343, 398, 220, 30, 128, 257, 201, 77, 0, 58, 143, 245, 335, 164, 9, 119, 160, 99, 46, 0, 0, 0, 9, 106, 197, 236, 208, 266, 124, 
    35, 429, 339, 319, 384, 233, 44, 161, 369, 274, 77, 12, 74, 186, 313, 419, 284, 90, 32, 22, 0, 0, 0, 0, 0, 0, 61, 141, 171, 132, 189, 89, 
    0, 377, 362, 319, 367, 215, 58, 245, 548, 518, 237, 96, 130, 212, 300, 369, 289, 133, 43, 0, 0, 0, 0, 0, 0, 0, 0, 36, 54, 23, 81, 28, 
    0, 278, 332, 327, 386, 252, 137, 331, 610, 564, 289, 83, 59, 112, 144, 165, 138, 61, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 
    0, 107, 204, 297, 370, 272, 239, 429, 568, 426, 154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 
    0, 0, 21, 163, 279, 245, 314, 511, 492, 243, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 7, 
    0, 0, 0, 8, 143, 213, 371, 548, 376, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 42, 
    0, 0, 0, 0, 14, 146, 392, 570, 274, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 94, 49, 
    0, 0, 0, 0, 0, 34, 314, 496, 193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 16, 
    0, 0, 0, 0, 0, 0, 110, 281, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 16, 0, 0, 0, 0, 
    0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 35, 51, 35, 0, 0, 0, 10, 79, 134, 111, 29, 0, 0, 0, 
    0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 30, 31, 8, 0, 0, 0, 40, 80, 80, 30, 0, 0, 0, 
    
    -- channel=12
    51, 70, 59, 60, 60, 59, 63, 63, 63, 63, 61, 60, 61, 65, 70, 71, 70, 66, 59, 51, 42, 38, 39, 42, 47, 47, 49, 54, 55, 53, 40, 17, 
    52, 112, 103, 106, 106, 103, 106, 108, 109, 110, 105, 98, 101, 110, 114, 118, 113, 103, 89, 73, 65, 59, 64, 67, 73, 80, 83, 88, 94, 97, 70, 66, 
    54, 133, 131, 134, 135, 131, 131, 132, 133, 142, 132, 117, 119, 123, 127, 125, 117, 108, 89, 81, 85, 78, 69, 68, 75, 83, 98, 107, 109, 113, 82, 84, 
    52, 131, 127, 129, 132, 131, 132, 133, 132, 140, 122, 104, 90, 79, 94, 96, 82, 86, 82, 67, 51, 42, 43, 51, 57, 60, 79, 96, 99, 106, 77, 84, 
    36, 105, 112, 117, 126, 132, 136, 137, 136, 136, 92, 79, 86, 60, 67, 81, 85, 92, 74, 32, 7, 0, 0, 2, 16, 30, 46, 79, 93, 98, 72, 82, 
    20, 80, 91, 112, 125, 137, 138, 141, 138, 139, 106, 89, 102, 85, 81, 78, 71, 70, 52, 16, 0, 0, 0, 0, 0, 13, 32, 56, 81, 88, 66, 79, 
    19, 99, 91, 90, 118, 139, 137, 141, 135, 133, 116, 85, 91, 79, 51, 22, 22, 40, 33, 7, 0, 0, 0, 0, 0, 9, 26, 45, 70, 82, 61, 79, 
    5, 83, 70, 59, 95, 124, 137, 144, 132, 123, 110, 87, 55, 31, 18, 0, 0, 21, 33, 17, 7, 9, 0, 0, 9, 19, 28, 38, 59, 79, 54, 77, 
    0, 54, 16, 20, 60, 88, 124, 139, 112, 96, 66, 31, 9, 8, 9, 0, 0, 18, 58, 46, 24, 30, 15, 6, 7, 13, 22, 33, 44, 67, 48, 76, 
    0, 29, 0, 0, 36, 65, 104, 119, 60, 7, 0, 0, 0, 0, 4, 4, 0, 26, 79, 51, 17, 16, 3, 0, 0, 1, 9, 26, 40, 49, 34, 76, 
    0, 30, 0, 0, 25, 63, 96, 104, 44, 0, 4, 0, 0, 0, 0, 9, 2, 28, 82, 36, 0, 0, 0, 0, 0, 0, 2, 12, 33, 34, 17, 66, 
    0, 34, 0, 0, 19, 58, 90, 118, 66, 23, 17, 5, 0, 11, 0, 0, 0, 35, 70, 12, 0, 0, 0, 4, 0, 0, 0, 0, 18, 26, 6, 44, 
    0, 45, 0, 0, 9, 54, 92, 121, 64, 39, 61, 28, 0, 0, 0, 0, 0, 39, 54, 0, 0, 0, 0, 11, 9, 7, 11, 5, 5, 17, 7, 30, 
    0, 39, 0, 0, 4, 38, 75, 123, 78, 51, 75, 28, 0, 0, 0, 0, 0, 32, 49, 0, 0, 0, 0, 0, 2, 7, 5, 0, 0, 11, 10, 40, 
    0, 32, 0, 0, 9, 18, 48, 107, 82, 64, 54, 0, 0, 0, 0, 0, 0, 33, 43, 0, 0, 0, 0, 0, 2, 5, 0, 0, 9, 27, 16, 57, 
    0, 22, 0, 0, 1, 0, 16, 62, 64, 61, 40, 0, 0, 0, 0, 0, 9, 38, 30, 8, 5, 0, 0, 0, 1, 8, 3, 0, 30, 54, 33, 68, 
    0, 9, 0, 0, 0, 0, 0, 31, 53, 37, 34, 0, 0, 24, 11, 12, 21, 43, 28, 11, 10, 9, 0, 0, 8, 20, 26, 34, 55, 74, 49, 73, 
    0, 0, 0, 0, 0, 0, 0, 3, 33, 11, 18, 33, 35, 57, 24, 15, 19, 21, 32, 42, 23, 11, 26, 31, 34, 40, 47, 58, 72, 80, 53, 80, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 8, 15, 29, 42, 8, 14, 6, 0, 13, 16, 0, 0, 29, 47, 42, 46, 48, 60, 84, 83, 53, 83, 
    0, 1, 0, 0, 0, 0, 0, 0, 12, 5, 34, 28, 37, 56, 1, 0, 4, 0, 0, 11, 19, 18, 23, 45, 45, 43, 42, 38, 62, 65, 38, 74, 
    0, 12, 0, 0, 0, 0, 3, 0, 0, 0, 5, 13, 2, 2, 0, 0, 0, 0, 0, 25, 38, 43, 34, 23, 24, 29, 34, 23, 41, 53, 28, 62, 
    13, 8, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 5, 0, 35, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 27, 49, 59, 48, 47, 56, 59, 53, 41, 38, 42, 45, 50, 59, 68, 65, 57, 53, 53, 42, 29, 26, 35, 50, 57, 57, 62, 73, 121, 191, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 21, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 25, 86, 221, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 84, 37, 0, 1, 13, 12, 0, 0, 12, 26, 10, 0, 0, 0, 0, 0, 0, 18, 85, 219, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 133, 101, 7, 0, 7, 0, 0, 0, 0, 47, 69, 43, 6, 0, 0, 0, 0, 0, 79, 223, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 147, 60, 16, 16, 0, 0, 0, 0, 13, 50, 57, 60, 56, 0, 0, 0, 0, 72, 228, 
    0, 6, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 26, 133, 131, 61, 22, 0, 0, 0, 0, 13, 10, 0, 40, 95, 70, 0, 0, 0, 51, 232, 
    0, 104, 35, 0, 0, 0, 0, 0, 5, 35, 2, 0, 0, 100, 158, 86, 6, 0, 0, 0, 0, 63, 45, 0, 3, 89, 112, 6, 0, 0, 10, 233, 
    0, 157, 93, 0, 0, 0, 0, 0, 0, 99, 101, 0, 0, 49, 137, 75, 0, 0, 0, 0, 0, 63, 113, 27, 0, 55, 106, 74, 0, 0, 0, 211, 
    0, 97, 61, 0, 0, 30, 0, 0, 0, 96, 191, 31, 0, 50, 141, 106, 13, 0, 0, 0, 0, 23, 152, 106, 14, 19, 80, 117, 34, 0, 0, 157, 
    0, 1, 0, 0, 48, 102, 0, 0, 0, 0, 169, 75, 0, 94, 155, 130, 80, 46, 0, 0, 0, 8, 149, 141, 21, 0, 45, 115, 113, 0, 0, 100, 
    0, 0, 0, 0, 83, 140, 49, 0, 0, 0, 54, 26, 0, 126, 188, 130, 117, 104, 0, 0, 0, 28, 144, 139, 11, 0, 3, 82, 126, 55, 0, 84, 
    0, 0, 0, 0, 76, 109, 87, 12, 0, 0, 0, 0, 0, 95, 233, 142, 111, 124, 0, 0, 0, 82, 163, 132, 11, 0, 0, 22, 81, 86, 59, 119, 
    0, 0, 0, 0, 92, 40, 41, 103, 0, 0, 0, 0, 0, 0, 203, 151, 97, 104, 0, 0, 0, 125, 181, 136, 24, 0, 0, 0, 30, 60, 91, 172, 
    0, 0, 0, 60, 180, 10, 0, 95, 0, 0, 0, 0, 0, 0, 103, 107, 83, 80, 0, 0, 0, 135, 174, 120, 25, 0, 0, 0, 0, 35, 77, 208, 
    0, 0, 0, 84, 275, 54, 0, 59, 46, 0, 0, 0, 0, 58, 39, 26, 47, 56, 0, 0, 0, 101, 154, 107, 9, 0, 0, 0, 0, 12, 59, 220, 
    0, 0, 0, 39, 301, 124, 0, 14, 81, 0, 0, 0, 0, 106, 42, 0, 0, 4, 0, 0, 0, 18, 142, 124, 9, 0, 0, 0, 0, 0, 53, 229, 
    0, 0, 0, 0, 250, 198, 0, 0, 100, 0, 0, 0, 0, 65, 33, 17, 0, 0, 0, 0, 0, 0, 87, 123, 25, 0, 0, 0, 0, 0, 50, 249, 
    0, 0, 0, 0, 181, 251, 0, 0, 47, 101, 0, 0, 0, 0, 0, 57, 42, 0, 0, 28, 5, 0, 38, 87, 12, 0, 0, 0, 0, 0, 58, 261, 
    0, 0, 0, 0, 110, 256, 0, 0, 0, 110, 98, 0, 0, 0, 0, 66, 147, 0, 0, 9, 74, 54, 64, 44, 0, 0, 0, 0, 0, 0, 71, 260, 
    0, 0, 0, 0, 56, 214, 28, 0, 0, 151, 153, 24, 0, 0, 0, 32, 241, 112, 0, 0, 30, 69, 63, 0, 0, 0, 0, 0, 0, 0, 68, 240, 
    0, 0, 0, 0, 35, 162, 0, 0, 0, 248, 260, 79, 0, 0, 0, 0, 203, 205, 82, 50, 25, 24, 14, 0, 0, 0, 0, 0, 0, 0, 48, 202, 
    0, 0, 0, 0, 32, 128, 0, 0, 0, 214, 300, 96, 0, 0, 0, 0, 68, 131, 106, 84, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 183, 
    0, 0, 0, 0, 0, 41, 0, 0, 0, 126, 246, 100, 0, 0, 0, 0, 0, 35, 26, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 187, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 192, 235, 127, 0, 0, 0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 217, 
    0, 0, 0, 0, 0, 0, 0, 0, 175, 268, 190, 78, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 249, 
    0, 0, 0, 0, 0, 0, 0, 15, 293, 276, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 251, 
    0, 0, 15, 0, 0, 0, 0, 102, 321, 219, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 224, 
    0, 0, 15, 0, 0, 0, 0, 47, 256, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 56, 188, 
    0, 0, 2, 0, 0, 0, 0, 0, 140, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 69, 80, 158, 
    0, 0, 2, 0, 0, 0, 0, 0, 64, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 6, 67, 74, 86, 150, 
    0, 0, 0, 0, 0, 4, 1, 0, 26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 12, 65, 48, 55, 122, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 57, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 19, 56, 59, 65, 65, 65, 69, 72, 72, 66, 57, 56, 60, 65, 71, 76, 78, 76, 75, 73, 65, 58, 55, 58, 63, 65, 67, 73, 81, 113, 138, 
    0, 0, 27, 30, 42, 42, 40, 49, 54, 55, 43, 32, 35, 40, 42, 49, 60, 66, 64, 58, 56, 49, 34, 22, 19, 28, 37, 47, 60, 78, 128, 202, 
    0, 0, 0, 0, 0, 0, 0, 5, 12, 11, 0, 0, 16, 22, 4, 3, 11, 22, 22, 20, 31, 34, 18, 0, 0, 0, 0, 0, 15, 39, 101, 189, 
    0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 0, 33, 44, 5, 0, 0, 8, 9, 16, 40, 67, 66, 45, 13, 0, 0, 0, 0, 19, 92, 190, 
    0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 38, 68, 27, 16, 18, 7, 0, 0, 26, 75, 96, 84, 66, 43, 0, 0, 0, 0, 74, 187, 
    0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 21, 76, 80, 68, 56, 25, 0, 0, 0, 57, 76, 76, 83, 92, 61, 0, 0, 0, 53, 181, 
    0, 18, 35, 0, 0, 0, 0, 4, 11, 16, 0, 0, 6, 86, 129, 115, 80, 43, 0, 0, 0, 44, 59, 42, 57, 107, 110, 25, 0, 0, 28, 173, 
    0, 83, 113, 0, 0, 0, 4, 0, 5, 46, 66, 35, 9, 58, 129, 122, 79, 45, 0, 0, 0, 37, 77, 46, 48, 97, 131, 85, 0, 0, 2, 156, 
    0, 99, 139, 0, 0, 9, 7, 0, 0, 40, 106, 51, 0, 38, 117, 111, 71, 49, 0, 0, 0, 19, 106, 86, 60, 82, 129, 128, 39, 0, 0, 134, 
    0, 53, 86, 0, 0, 41, 8, 0, 0, 0, 78, 48, 0, 35, 108, 118, 90, 73, 12, 0, 0, 10, 115, 118, 74, 66, 108, 149, 107, 0, 0, 110, 
    0, 0, 2, 0, 6, 64, 29, 0, 0, 0, 0, 7, 0, 32, 115, 126, 125, 111, 23, 0, 0, 12, 105, 121, 72, 40, 79, 134, 146, 66, 13, 101, 
    0, 0, 0, 0, 0, 53, 43, 0, 0, 0, 0, 0, 0, 25, 131, 133, 134, 132, 23, 0, 0, 31, 102, 110, 55, 13, 47, 98, 139, 115, 77, 116, 
    0, 0, 0, 0, 0, 21, 28, 35, 0, 0, 0, 0, 0, 0, 120, 122, 115, 129, 12, 0, 0, 47, 111, 115, 68, 16, 26, 67, 103, 115, 117, 149, 
    0, 0, 0, 0, 44, 2, 0, 57, 0, 0, 0, 0, 0, 0, 77, 91, 82, 96, 0, 0, 0, 57, 124, 117, 75, 30, 13, 30, 67, 85, 115, 176, 
    0, 0, 0, 11, 112, 32, 0, 46, 48, 0, 0, 0, 0, 0, 12, 26, 47, 66, 0, 0, 0, 50, 114, 115, 78, 30, 0, 0, 32, 54, 94, 177, 
    0, 0, 0, 19, 155, 85, 0, 16, 67, 0, 0, 0, 0, 7, 0, 0, 21, 44, 0, 0, 0, 17, 91, 110, 58, 0, 0, 0, 4, 27, 73, 177, 
    0, 0, 0, 0, 146, 135, 0, 0, 63, 0, 0, 0, 0, 6, 14, 13, 17, 18, 0, 0, 0, 0, 68, 98, 57, 0, 0, 0, 0, 4, 59, 185, 
    0, 0, 0, 0, 119, 159, 0, 0, 39, 48, 0, 0, 0, 0, 32, 45, 51, 4, 0, 0, 0, 0, 42, 92, 57, 0, 0, 0, 0, 0, 60, 194, 
    0, 0, 0, 0, 81, 164, 38, 0, 5, 82, 43, 0, 0, 0, 5, 68, 113, 9, 0, 19, 38, 24, 57, 75, 44, 0, 0, 0, 0, 0, 66, 195, 
    0, 0, 0, 0, 46, 146, 77, 0, 0, 97, 125, 56, 0, 0, 0, 59, 162, 83, 0, 5, 58, 76, 86, 79, 39, 0, 0, 0, 0, 6, 69, 185, 
    0, 0, 0, 0, 22, 116, 67, 0, 2, 145, 199, 118, 0, 0, 0, 14, 152, 135, 44, 37, 64, 100, 114, 97, 48, 0, 0, 0, 0, 22, 74, 170, 
    0, 0, 0, 0, 17, 101, 32, 0, 0, 157, 231, 129, 0, 0, 0, 0, 70, 130, 112, 106, 109, 110, 120, 113, 84, 47, 8, 0, 28, 55, 93, 162, 
    0, 0, 0, 0, 0, 68, 0, 0, 0, 96, 195, 116, 0, 0, 0, 0, 15, 79, 105, 127, 132, 122, 109, 107, 107, 95, 78, 72, 84, 103, 126, 177, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 157, 120, 30, 10, 10, 19, 53, 83, 97, 112, 120, 118, 114, 110, 111, 117, 117, 115, 121, 130, 146, 194, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 131, 162, 130, 101, 94, 91, 93, 102, 117, 123, 122, 122, 123, 126, 124, 119, 119, 122, 123, 127, 134, 155, 207, 
    23, 84, 20, 0, 0, 0, 0, 0, 124, 201, 168, 129, 119, 119, 117, 114, 119, 126, 129, 130, 129, 129, 127, 124, 120, 116, 113, 114, 119, 122, 139, 201, 
    20, 123, 127, 11, 0, 0, 0, 0, 191, 232, 150, 121, 122, 128, 124, 117, 117, 121, 124, 125, 127, 123, 119, 119, 121, 123, 117, 111, 108, 103, 117, 179, 
    17, 125, 164, 102, 0, 0, 0, 0, 190, 214, 133, 108, 118, 135, 134, 124, 117, 116, 119, 122, 127, 126, 118, 115, 124, 134, 134, 125, 123, 122, 123, 154, 
    14, 123, 167, 136, 70, 0, 0, 0, 155, 166, 108, 91, 95, 118, 129, 127, 121, 117, 120, 126, 137, 141, 130, 121, 123, 131, 138, 150, 169, 168, 149, 147, 
    7, 120, 166, 139, 120, 57, 0, 29, 131, 139, 109, 88, 83, 92, 102, 103, 98, 102, 114, 132, 147, 152, 143, 125, 102, 98, 120, 164, 196, 195, 175, 160, 
    0, 88, 124, 105, 99, 91, 65, 60, 101, 118, 99, 82, 75, 71, 68, 60, 50, 50, 60, 82, 107, 118, 106, 77, 39, 24, 58, 117, 156, 161, 150, 136, 
    0, 41, 59, 51, 47, 49, 49, 49, 56, 67, 60, 54, 53, 50, 44, 28, 12, 2, 3, 20, 42, 53, 46, 22, 0, 0, 0, 45, 77, 82, 79, 95, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 39, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 25, 
    0, 2, 26, 24, 20, 20, 20, 20, 19, 21, 35, 64, 60, 38, 24, 19, 12, 2, 1, 17, 41, 54, 45, 25, 0, 0, 0, 0, 4, 16, 48, 43, 
    0, 0, 18, 15, 14, 17, 17, 17, 13, 0, 0, 16, 15, 4, 0, 0, 0, 0, 0, 26, 54, 68, 72, 65, 53, 26, 0, 0, 0, 3, 43, 40, 
    0, 0, 0, 0, 0, 14, 22, 23, 21, 0, 0, 0, 0, 0, 5, 10, 13, 11, 18, 33, 28, 12, 5, 13, 37, 39, 10, 0, 0, 0, 38, 39, 
    2, 5, 0, 0, 0, 11, 24, 26, 28, 29, 27, 5, 1, 35, 64, 64, 57, 36, 23, 18, 6, 0, 0, 0, 0, 9, 10, 0, 0, 0, 26, 33, 
    48, 77, 44, 23, 18, 16, 19, 24, 31, 49, 53, 35, 29, 59, 58, 38, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 19, 29, 
    66, 96, 74, 67, 51, 23, 21, 29, 64, 102, 101, 64, 46, 36, 12, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 22, 31, 2, 0, 6, 20, 
    44, 41, 25, 49, 36, 6, 6, 2, 48, 104, 104, 63, 39, 16, 1, 3, 2, 0, 0, 0, 13, 21, 35, 33, 18, 16, 28, 42, 27, 0, 0, 4, 
    19, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 3, 11, 8, 17, 26, 19, 2, 30, 62, 40, 24, 2, 0, 0, 13, 29, 41, 22, 18, 2, 
    25, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 10, 20, 19, 36, 36, 5, 33, 48, 3, 0, 0, 0, 0, 0, 10, 34, 42, 46, 19, 
    34, 0, 0, 0, 0, 0, 18, 40, 0, 0, 0, 0, 0, 15, 26, 19, 34, 28, 3, 20, 20, 0, 0, 0, 0, 0, 0, 0, 12, 35, 54, 37, 
    36, 1, 12, 14, 0, 0, 0, 41, 21, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 11, 14, 0, 0, 4, 9, 2, 0, 2, 7, 5, 27, 24, 
    32, 0, 24, 40, 0, 0, 0, 21, 26, 5, 0, 15, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 6, 10, 7, 0, 0, 0, 13, 
    29, 0, 15, 38, 12, 0, 10, 19, 31, 1, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    35, 7, 4, 18, 21, 11, 2, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 32, 
    38, 14, 0, 0, 10, 0, 0, 0, 16, 12, 0, 0, 0, 0, 0, 16, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 33, 
    25, 0, 0, 0, 4, 0, 0, 0, 0, 34, 47, 7, 0, 0, 35, 64, 36, 0, 12, 33, 30, 17, 0, 0, 0, 2, 0, 0, 0, 0, 36, 31, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 21, 22, 0, 0, 0, 27, 76, 46, 0, 0, 0, 0, 3, 0, 0, 8, 14, 0, 0, 0, 0, 35, 30, 
    0, 0, 0, 0, 0, 0, 0, 36, 77, 88, 61, 40, 46, 37, 49, 69, 58, 36, 2, 0, 0, 0, 6, 36, 37, 7, 0, 0, 0, 0, 24, 21, 
    4, 0, 0, 0, 0, 0, 0, 37, 120, 151, 143, 113, 73, 35, 8, 0, 0, 12, 39, 49, 51, 61, 80, 95, 90, 59, 32, 21, 18, 19, 48, 34, 
    9, 11, 0, 0, 10, 9, 0, 27, 31, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 89, 94, 84, 75, 70, 65, 67, 72, 72, 78, 95, 55, 
    22, 6, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 29, 47, 57, 51, 46, 49, 56, 67, 71, 71, 74, 79, 37, 
    68, 55, 0, 0, 0, 0, 0, 5, 0, 0, 0, 5, 58, 86, 88, 85, 77, 66, 55, 49, 52, 50, 50, 55, 58, 62, 62, 60, 58, 59, 75, 41, 
    104, 116, 32, 0, 0, 0, 0, 30, 0, 0, 0, 50, 76, 70, 64, 63, 59, 56, 55, 59, 63, 64, 65, 65, 61, 49, 38, 37, 49, 63, 86, 48, 
    80, 108, 70, 35, 0, 0, 14, 45, 17, 5, 27, 53, 45, 36, 32, 35, 41, 47, 53, 58, 61, 59, 55, 54, 46, 31, 23, 30, 51, 54, 47, 3, 
    69, 85, 71, 63, 19, 0, 1, 5, 0, 10, 42, 48, 46, 45, 43, 41, 38, 40, 46, 51, 52, 46, 39, 36, 38, 41, 52, 65, 61, 25, 0, 0, 
    75, 86, 61, 69, 50, 9, 0, 0, 0, 0, 25, 26, 35, 43, 51, 50, 46, 46, 49, 50, 50, 49, 44, 36, 38, 56, 80, 87, 64, 30, 10, 0, 
    75, 83, 52, 59, 66, 52, 25, 0, 0, 1, 17, 11, 10, 11, 21, 33, 46, 55, 60, 61, 59, 53, 47, 43, 50, 69, 88, 86, 71, 55, 44, 12, 
    64, 73, 45, 48, 59, 75, 70, 58, 46, 50, 48, 38, 23, 7, 0, 0, 5, 21, 36, 48, 52, 48, 43, 40, 45, 55, 59, 50, 36, 35, 48, 20, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    43, 84, 90, 98, 98, 97, 99, 99, 96, 92, 94, 97, 98, 96, 95, 95, 93, 90, 85, 81, 75, 68, 66, 70, 79, 85, 85, 79, 74, 71, 88, 42, 
    33, 46, 67, 78, 84, 87, 88, 90, 90, 91, 101, 105, 98, 86, 86, 93, 95, 84, 63, 45, 36, 27, 17, 16, 25, 40, 57, 70, 74, 75, 112, 44, 
    27, 41, 62, 72, 77, 77, 76, 79, 80, 92, 128, 158, 137, 93, 77, 74, 58, 41, 30, 42, 62, 65, 43, 14, 0, 0, 10, 35, 58, 67, 118, 40, 
    33, 47, 68, 72, 76, 72, 70, 72, 71, 76, 103, 146, 132, 77, 38, 18, 0, 0, 22, 83, 123, 135, 114, 82, 47, 14, 0, 2, 31, 57, 117, 39, 
    25, 17, 19, 28, 56, 70, 71, 72, 67, 45, 21, 25, 35, 29, 4, 0, 0, 14, 68, 105, 126, 122, 113, 102, 83, 44, 0, 0, 0, 40, 117, 41, 
    24, 4, 0, 0, 22, 66, 76, 79, 75, 33, 0, 0, 24, 65, 66, 59, 66, 70, 78, 92, 98, 75, 48, 49, 65, 39, 3, 0, 0, 12, 105, 39, 
    76, 78, 30, 28, 39, 62, 76, 85, 92, 63, 38, 40, 79, 135, 127, 103, 74, 64, 48, 44, 55, 47, 13, 0, 15, 29, 19, 0, 0, 0, 87, 38, 
    163, 190, 148, 116, 98, 70, 80, 114, 165, 188, 155, 120, 132, 140, 103, 67, 32, 15, 0, 0, 22, 48, 35, 7, 8, 38, 51, 28, 0, 0, 60, 24, 
    196, 237, 206, 172, 127, 72, 74, 122, 231, 314, 279, 192, 138, 113, 79, 51, 22, 0, 0, 17, 73, 96, 93, 63, 46, 64, 84, 60, 19, 0, 31, 0, 
    172, 190, 167, 156, 123, 71, 57, 64, 141, 213, 212, 141, 117, 116, 93, 76, 48, 14, 38, 104, 158, 150, 118, 78, 50, 66, 91, 87, 56, 7, 30, 0, 
    140, 128, 105, 115, 100, 81, 46, 6, 0, 9, 40, 62, 102, 146, 126, 99, 93, 71, 100, 150, 178, 132, 76, 37, 26, 39, 70, 94, 92, 58, 57, 0, 
    125, 115, 72, 97, 57, 62, 50, 25, 0, 0, 0, 8, 92, 170, 163, 122, 132, 113, 144, 146, 135, 75, 37, 12, 8, 10, 37, 80, 102, 92, 94, 17, 
    128, 137, 98, 105, 17, 21, 52, 49, 0, 0, 0, 39, 97, 133, 141, 120, 127, 104, 129, 113, 112, 62, 51, 37, 26, 15, 33, 77, 100, 89, 108, 30, 
    144, 156, 127, 133, 31, 16, 61, 55, 27, 11, 52, 108, 106, 70, 42, 61, 86, 61, 92, 78, 95, 58, 67, 55, 46, 48, 63, 76, 70, 54, 87, 29, 
    155, 161, 143, 177, 98, 54, 72, 69, 57, 40, 76, 91, 82, 14, 0, 0, 22, 20, 59, 45, 51, 42, 59, 39, 24, 34, 36, 26, 12, 13, 77, 25, 
    168, 173, 146, 198, 153, 98, 81, 86, 71, 21, 0, 0, 0, 0, 0, 0, 0, 10, 22, 0, 0, 0, 42, 25, 4, 0, 0, 0, 0, 12, 96, 29, 
    180, 183, 136, 184, 165, 120, 75, 90, 84, 22, 0, 0, 0, 0, 0, 6, 18, 18, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 44, 116, 34, 
    168, 166, 108, 150, 157, 130, 73, 85, 84, 66, 0, 0, 0, 20, 87, 110, 75, 27, 36, 33, 4, 0, 0, 0, 0, 2, 14, 31, 43, 51, 114, 33, 
    132, 125, 74, 109, 142, 130, 87, 88, 87, 86, 36, 2, 24, 65, 145, 187, 126, 28, 9, 8, 4, 0, 0, 0, 29, 51, 51, 48, 46, 45, 110, 31, 
    99, 93, 58, 75, 115, 102, 112, 155, 211, 192, 120, 88, 102, 145, 205, 241, 185, 84, 0, 0, 0, 0, 7, 50, 84, 68, 42, 26, 31, 35, 99, 21, 
    95, 107, 71, 67, 101, 84, 133, 230, 354, 372, 296, 246, 201, 193, 170, 172, 152, 118, 41, 6, 17, 65, 124, 163, 168, 135, 87, 57, 51, 59, 117, 34, 
    97, 119, 79, 86, 131, 133, 196, 271, 345, 345, 252, 165, 91, 26, 0, 0, 4, 45, 75, 103, 144, 175, 193, 199, 190, 173, 143, 125, 115, 124, 160, 57, 
    89, 90, 38, 67, 135, 164, 227, 227, 194, 114, 39, 0, 0, 0, 0, 0, 0, 37, 96, 143, 171, 185, 180, 178, 183, 185, 183, 171, 159, 163, 189, 72, 
    111, 108, 24, 18, 70, 113, 171, 142, 78, 0, 0, 19, 60, 82, 78, 77, 88, 104, 122, 140, 162, 172, 179, 187, 199, 205, 204, 196, 192, 200, 226, 99, 
    161, 184, 85, 32, 34, 87, 140, 109, 31, 0, 23, 104, 142, 150, 144, 142, 139, 141, 153, 167, 181, 192, 204, 214, 213, 203, 192, 195, 213, 239, 273, 122, 
    181, 224, 149, 89, 70, 107, 125, 126, 46, 36, 97, 146, 156, 151, 145, 148, 156, 164, 175, 187, 198, 206, 212, 213, 198, 175, 169, 192, 227, 243, 256, 85, 
    177, 223, 183, 157, 127, 106, 89, 117, 63, 89, 137, 160, 163, 161, 157, 155, 158, 167, 180, 189, 195, 195, 190, 182, 173, 176, 196, 226, 227, 187, 165, 28, 
    182, 227, 193, 191, 164, 99, 34, 37, 24, 85, 128, 152, 167, 172, 173, 170, 169, 174, 182, 187, 186, 183, 175, 170, 179, 210, 249, 255, 205, 138, 121, 18, 
    188, 231, 194, 194, 181, 126, 42, 2, 0, 71, 101, 122, 131, 140, 152, 165, 180, 196, 204, 203, 193, 182, 174, 179, 209, 259, 286, 261, 202, 155, 147, 39, 
    177, 218, 186, 190, 183, 163, 115, 69, 61, 99, 117, 121, 113, 102, 103, 119, 145, 172, 193, 204, 196, 179, 175, 193, 233, 267, 265, 230, 183, 153, 155, 55, 
    78, 87, 52, 62, 58, 50, 45, 26, 12, 33, 45, 47, 38, 26, 16, 9, 13, 25, 37, 42, 37, 36, 48, 65, 75, 67, 47, 25, 12, 26, 56, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 147, 103, 123, 112, 98, 106, 107, 101, 95, 93, 104, 111, 113, 116, 118, 113, 98, 88, 85, 79, 71, 70, 75, 83, 81, 75, 70, 67, 59, 62, 19, 
    16, 207, 161, 194, 187, 171, 180, 181, 174, 163, 161, 180, 185, 178, 184, 189, 180, 161, 135, 121, 110, 92, 86, 97, 117, 130, 139, 135, 125, 113, 130, 52, 
    2, 177, 121, 154, 152, 144, 156, 155, 146, 138, 149, 196, 183, 124, 130, 147, 139, 117, 77, 49, 37, 14, 0, 0, 14, 37, 70, 91, 96, 91, 120, 38, 
    5, 181, 121, 151, 154, 147, 158, 159, 143, 128, 165, 292, 268, 123, 104, 123, 104, 57, 16, 32, 55, 44, 13, 0, 0, 0, 0, 40, 86, 101, 132, 45, 
    6, 173, 94, 126, 157, 150, 154, 155, 136, 107, 146, 301, 288, 121, 60, 39, 5, 0, 0, 57, 109, 100, 74, 34, 8, 0, 0, 0, 44, 109, 150, 51, 
    1, 140, 2, 36, 135, 155, 150, 153, 141, 102, 99, 184, 183, 100, 16, 0, 0, 0, 0, 85, 164, 131, 73, 54, 65, 31, 0, 0, 0, 92, 170, 62, 
    2, 125, 0, 0, 95, 150, 145, 154, 155, 124, 88, 86, 102, 110, 45, 0, 0, 0, 0, 102, 206, 156, 43, 28, 64, 35, 0, 0, 0, 46, 176, 77, 
    39, 186, 0, 0, 110, 134, 129, 150, 180, 181, 90, 29, 101, 167, 88, 0, 0, 0, 0, 56, 192, 191, 51, 0, 18, 10, 0, 0, 0, 0, 148, 95, 
    90, 270, 0, 94, 202, 133, 104, 130, 231, 318, 190, 68, 156, 216, 107, 0, 0, 0, 0, 0, 148, 201, 97, 9, 0, 0, 0, 0, 0, 0, 85, 89, 
    102, 306, 59, 239, 279, 144, 77, 99, 278, 492, 378, 176, 214, 245, 116, 26, 0, 0, 0, 0, 180, 228, 148, 50, 0, 10, 30, 0, 0, 0, 0, 33, 
    81, 277, 109, 327, 309, 156, 77, 59, 193, 444, 425, 228, 258, 290, 144, 48, 28, 0, 0, 5, 282, 293, 172, 53, 0, 23, 52, 21, 0, 0, 0, 0, 
    72, 255, 97, 346, 308, 166, 116, 55, 58, 277, 329, 174, 248, 353, 206, 63, 66, 21, 0, 74, 362, 307, 146, 22, 0, 8, 43, 38, 2, 0, 0, 0, 
    68, 249, 100, 358, 252, 120, 154, 99, 0, 145, 215, 131, 251, 385, 274, 103, 106, 64, 0, 126, 376, 271, 105, 0, 0, 0, 0, 29, 40, 14, 33, 0, 
    70, 268, 149, 382, 188, 30, 143, 124, 0, 70, 149, 176, 297, 337, 252, 144, 140, 69, 0, 154, 356, 241, 91, 11, 0, 0, 0, 44, 78, 49, 65, 14, 
    77, 305, 197, 399, 190, 0, 98, 137, 0, 23, 136, 287, 381, 273, 153, 134, 142, 57, 0, 148, 303, 215, 104, 26, 0, 0, 33, 74, 96, 60, 84, 44, 
    88, 357, 221, 395, 249, 16, 70, 161, 43, 3, 126, 325, 383, 219, 82, 74, 82, 35, 6, 117, 220, 199, 131, 19, 0, 0, 47, 80, 77, 52, 117, 71, 
    105, 412, 229, 381, 313, 69, 43, 181, 112, 0, 69, 194, 211, 128, 38, 41, 33, 10, 51, 94, 86, 122, 145, 25, 0, 0, 10, 52, 64, 69, 163, 94, 
    117, 453, 237, 356, 346, 119, 19, 174, 196, 46, 26, 32, 78, 78, 37, 91, 33, 0, 104, 88, 0, 46, 68, 0, 0, 0, 0, 47, 94, 109, 189, 99, 
    108, 457, 257, 322, 349, 172, 13, 125, 217, 133, 53, 0, 42, 88, 105, 207, 93, 0, 102, 131, 51, 22, 0, 0, 0, 0, 13, 83, 141, 136, 189, 94, 
    75, 426, 279, 286, 342, 209, 31, 102, 247, 205, 73, 0, 7, 76, 184, 322, 186, 2, 35, 58, 36, 0, 0, 0, 0, 0, 49, 111, 147, 115, 153, 68, 
    34, 389, 309, 261, 324, 213, 37, 156, 394, 326, 115, 1, 48, 156, 286, 381, 272, 92, 9, 0, 0, 0, 0, 0, 0, 2, 43, 89, 92, 45, 84, 35, 
    6, 355, 338, 271, 318, 199, 40, 229, 555, 540, 268, 114, 143, 236, 297, 322, 254, 130, 40, 0, 0, 0, 0, 0, 11, 27, 34, 45, 39, 11, 57, 39, 
    0, 293, 318, 303, 343, 222, 125, 341, 586, 547, 313, 114, 88, 134, 139, 124, 93, 42, 8, 0, 0, 0, 16, 35, 53, 57, 55, 55, 48, 31, 83, 75, 
    0, 184, 208, 273, 337, 248, 230, 451, 564, 387, 127, 0, 0, 5, 0, 0, 0, 0, 0, 0, 12, 34, 41, 43, 54, 69, 74, 70, 69, 62, 124, 122, 
    0, 118, 80, 170, 261, 222, 299, 526, 479, 199, 0, 0, 0, 14, 11, 6, 5, 4, 3, 8, 21, 36, 45, 55, 74, 92, 96, 90, 90, 90, 168, 166, 
    0, 140, 50, 77, 155, 202, 377, 567, 361, 33, 0, 10, 41, 44, 30, 26, 24, 21, 20, 26, 40, 55, 69, 87, 101, 103, 90, 86, 107, 132, 227, 203, 
    0, 154, 57, 56, 81, 167, 410, 567, 248, 0, 0, 33, 55, 42, 26, 26, 29, 32, 38, 48, 60, 72, 87, 101, 100, 81, 64, 79, 130, 169, 228, 173, 
    0, 158, 61, 65, 63, 111, 317, 448, 171, 0, 13, 48, 67, 59, 36, 29, 30, 38, 48, 59, 69, 71, 74, 82, 82, 68, 69, 104, 147, 138, 138, 100, 
    0, 169, 70, 72, 74, 72, 152, 226, 81, 0, 7, 42, 70, 76, 64, 47, 36, 45, 57, 68, 71, 66, 60, 56, 60, 82, 116, 148, 136, 84, 75, 61, 
    0, 179, 70, 74, 77, 64, 50, 53, 3, 0, 0, 9, 38, 51, 56, 52, 59, 76, 86, 95, 88, 67, 51, 45, 68, 129, 187, 194, 140, 69, 59, 54, 
    0, 166, 75, 76, 80, 68, 53, 29, 3, 0, 0, 0, 5, 7, 12, 17, 40, 74, 107, 135, 125, 86, 62, 60, 97, 175, 239, 222, 135, 58, 60, 34, 
    0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 0, 0, 0, 2, 43, 71, 60, 15, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 2, 3, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 4, 3, 2, 1, 2, 1, 0, 0, 4, 1, 8, 
    5, 5, 27, 25, 33, 33, 31, 32, 36, 39, 35, 21, 18, 28, 34, 36, 37, 37, 36, 34, 28, 23, 20, 21, 24, 26, 28, 30, 32, 33, 20, 33, 
    23, 25, 45, 41, 47, 48, 46, 49, 54, 63, 55, 25, 24, 45, 50, 49, 50, 57, 65, 48, 30, 21, 19, 20, 23, 29, 33, 40, 44, 46, 30, 39, 
    23, 25, 47, 43, 47, 47, 45, 50, 54, 61, 47, 19, 45, 66, 54, 47, 52, 61, 49, 30, 16, 14, 13, 14, 19, 18, 25, 38, 38, 39, 25, 38, 
    22, 22, 53, 51, 47, 47, 47, 50, 52, 52, 24, 7, 45, 65, 48, 41, 42, 38, 29, 2, 0, 0, 8, 20, 12, 14, 30, 35, 34, 32, 22, 39, 
    18, 15, 52, 48, 34, 41, 50, 52, 52, 48, 35, 24, 48, 51, 44, 35, 28, 22, 12, 0, 0, 0, 3, 5, 2, 15, 35, 40, 30, 22, 14, 38, 
    4, 8, 55, 39, 15, 32, 51, 52, 47, 41, 46, 54, 35, 20, 33, 38, 18, 5, 3, 0, 0, 0, 10, 2, 0, 13, 30, 34, 33, 22, 7, 35, 
    0, 3, 51, 21, 0, 30, 58, 62, 43, 22, 33, 29, 5, 0, 17, 19, 2, 0, 9, 3, 0, 0, 12, 3, 0, 9, 12, 22, 31, 27, 4, 31, 
    0, 0, 37, 0, 0, 40, 68, 74, 41, 13, 30, 26, 0, 0, 13, 15, 0, 3, 23, 22, 0, 0, 5, 13, 12, 4, 2, 11, 29, 29, 4, 24, 
    0, 0, 12, 0, 0, 50, 60, 50, 21, 0, 23, 22, 0, 0, 12, 13, 3, 8, 31, 27, 0, 0, 0, 26, 23, 0, 0, 3, 22, 33, 4, 18, 
    0, 0, 0, 0, 11, 52, 57, 35, 0, 0, 0, 29, 0, 0, 8, 10, 0, 16, 30, 3, 0, 0, 5, 28, 18, 0, 0, 4, 16, 25, 6, 11, 
    0, 0, 0, 0, 16, 56, 48, 51, 29, 0, 10, 30, 0, 0, 9, 16, 0, 20, 28, 0, 0, 0, 18, 33, 16, 0, 2, 5, 5, 9, 2, 13, 
    0, 0, 0, 0, 24, 53, 32, 47, 48, 1, 8, 17, 0, 0, 22, 29, 0, 15, 28, 0, 0, 0, 25, 22, 7, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 37, 51, 20, 37, 42, 16, 8, 0, 0, 0, 22, 25, 2, 24, 24, 0, 0, 13, 27, 26, 21, 12, 3, 0, 0, 8, 7, 20, 
    0, 0, 0, 0, 35, 51, 13, 25, 43, 28, 15, 0, 0, 20, 27, 16, 12, 31, 25, 0, 0, 5, 14, 12, 8, 2, 0, 0, 0, 26, 10, 23, 
    0, 0, 0, 0, 22, 44, 24, 15, 29, 20, 0, 0, 0, 34, 34, 11, 10, 23, 12, 0, 0, 24, 19, 23, 21, 7, 0, 0, 12, 26, 7, 27, 
    0, 0, 0, 0, 0, 34, 23, 0, 21, 17, 0, 0, 2, 29, 22, 4, 13, 14, 0, 0, 5, 0, 6, 35, 25, 14, 7, 10, 21, 24, 6, 33, 
    0, 0, 0, 0, 0, 27, 12, 0, 11, 20, 10, 7, 8, 27, 14, 0, 4, 12, 0, 18, 14, 0, 9, 32, 28, 15, 6, 4, 15, 22, 9, 38, 
    0, 0, 0, 0, 0, 17, 9, 0, 0, 0, 22, 30, 14, 16, 0, 0, 1, 7, 0, 26, 33, 21, 27, 35, 24, 11, 8, 0, 11, 30, 20, 43, 
    0, 0, 0, 0, 0, 11, 26, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 6, 0, 0, 8, 21, 25, 3, 0, 0, 0, 0, 15, 37, 21, 36, 
    0, 0, 0, 0, 0, 7, 19, 0, 0, 0, 6, 8, 0, 0, 0, 0, 10, 26, 14, 7, 7, 8, 1, 0, 0, 0, 0, 0, 12, 20, 4, 14, 
    3, 0, 0, 0, 0, 13, 9, 0, 0, 0, 17, 3, 0, 0, 0, 0, 2, 12, 14, 14, 3, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 
    0, 0, 0, 0, 0, 13, 10, 0, 0, 0, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    258, 307, 278, 272, 264, 269, 273, 271, 268, 268, 269, 272, 276, 280, 282, 279, 272, 268, 265, 258, 249, 245, 248, 253, 252, 247, 243, 241, 239, 230, 191, 93, 
    245, 251, 219, 213, 206, 214, 221, 216, 213, 212, 216, 217, 211, 211, 219, 219, 214, 203, 191, 183, 172, 167, 172, 184, 193, 199, 200, 200, 198, 193, 168, 56, 
    255, 285, 258, 253, 244, 253, 259, 254, 251, 256, 281, 276, 236, 225, 246, 249, 233, 211, 203, 206, 193, 172, 166, 175, 191, 210, 227, 236, 238, 232, 194, 71, 
    257, 286, 260, 258, 251, 256, 260, 253, 252, 269, 315, 301, 221, 196, 218, 211, 183, 175, 199, 219, 195, 165, 148, 149, 165, 181, 205, 231, 246, 239, 196, 69, 
    245, 262, 240, 259, 264, 260, 257, 250, 250, 260, 292, 267, 173, 142, 156, 155, 149, 162, 207, 225, 194, 145, 123, 130, 143, 147, 161, 205, 243, 248, 199, 66, 
    214, 198, 175, 242, 278, 273, 261, 256, 254, 248, 252, 223, 163, 136, 131, 137, 155, 168, 208, 228, 179, 119, 107, 123, 122, 97, 106, 157, 226, 251, 205, 64, 
    195, 145, 121, 232, 290, 274, 261, 260, 259, 240, 230, 237, 225, 191, 140, 144, 166, 163, 175, 211, 183, 121, 104, 128, 125, 90, 81, 118, 191, 243, 212, 67, 
    202, 129, 127, 248, 294, 262, 253, 268, 277, 238, 198, 225, 247, 192, 116, 114, 137, 127, 129, 186, 195, 134, 101, 120, 125, 107, 89, 93, 143, 222, 220, 77, 
    208, 131, 137, 245, 258, 229, 246, 303, 343, 279, 182, 198, 224, 159, 90, 91, 115, 105, 109, 182, 222, 161, 103, 102, 129, 135, 114, 88, 102, 176, 209, 84, 
    197, 130, 146, 220, 199, 185, 218, 278, 343, 279, 159, 153, 183, 126, 80, 91, 105, 94, 121, 223, 261, 187, 106, 89, 129, 155, 129, 90, 78, 126, 179, 86, 
    179, 118, 143, 195, 164, 165, 187, 204, 258, 214, 99, 117, 174, 132, 81, 94, 101, 83, 135, 258, 265, 162, 81, 71, 121, 157, 138, 103, 80, 103, 150, 83, 
    164, 110, 139, 178, 140, 168, 190, 164, 196, 202, 118, 152, 224, 159, 86, 95, 115, 83, 138, 257, 229, 108, 51, 65, 118, 153, 146, 125, 102, 106, 124, 71, 
    162, 113, 144, 144, 102, 166, 213, 168, 191, 226, 192, 214, 262, 182, 99, 106, 124, 82, 129, 236, 192, 78, 52, 75, 115, 145, 156, 151, 124, 114, 119, 54, 
    176, 133, 148, 106, 56, 160, 236, 176, 179, 238, 255, 274, 245, 150, 96, 115, 119, 75, 126, 213, 176, 84, 75, 90, 123, 151, 174, 176, 144, 130, 134, 52, 
    192, 146, 147, 91, 30, 142, 242, 201, 183, 235, 286, 279, 186, 98, 94, 124, 121, 90, 142, 214, 176, 100, 81, 84, 116, 153, 172, 172, 149, 150, 160, 60, 
    203, 150, 141, 106, 20, 97, 217, 212, 180, 211, 248, 222, 118, 61, 103, 138, 134, 129, 175, 212, 180, 133, 97, 76, 99, 133, 151, 159, 161, 184, 192, 65, 
    210, 148, 128, 119, 20, 39, 165, 209, 167, 159, 172, 153, 95, 82, 125, 146, 142, 170, 194, 181, 174, 161, 109, 70, 96, 128, 156, 182, 203, 228, 210, 63, 
    217, 147, 109, 117, 30, 8, 115, 189, 161, 146, 134, 155, 165, 167, 194, 165, 125, 171, 207, 180, 158, 145, 90, 65, 99, 142, 191, 232, 242, 242, 206, 54, 
    225, 163, 104, 114, 54, 3, 81, 165, 153, 122, 108, 147, 200, 217, 240, 170, 82, 132, 195, 177, 152, 126, 93, 97, 139, 188, 239, 271, 253, 232, 195, 53, 
    235, 194, 122, 119, 76, 9, 70, 167, 157, 95, 58, 115, 194, 229, 245, 157, 49, 73, 131, 118, 98, 82, 82, 111, 143, 173, 224, 256, 238, 219, 188, 57, 
    235, 216, 142, 128, 89, 17, 91, 214, 197, 94, 67, 119, 190, 225, 220, 144, 48, 54, 83, 88, 83, 88, 107, 119, 115, 124, 155, 188, 182, 171, 148, 33, 
    205, 202, 146, 136, 96, 40, 131, 261, 227, 95, 31, 82, 121, 115, 101, 61, 18, 29, 61, 83, 108, 116, 110, 95, 69, 64, 75, 101, 103, 100, 80, 0, 
    143, 126, 104, 129, 112, 87, 186, 267, 189, 2, 0, 0, 0, 0, 0, 0, 0, 0, 27, 48, 58, 55, 35, 15, 0, 0, 0, 10, 18, 19, 6, 0, 
    78, 24, 29, 88, 99, 113, 208, 222, 86, 0, 0, 0, 0, 0, 0, 5, 8, 9, 13, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 0, 0, 40, 72, 129, 217, 163, 0, 0, 0, 0, 17, 9, 7, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 0, 0, 0, 47, 142, 212, 103, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 0, 0, 0, 0, 97, 160, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 0, 0, 0, 0, 14, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 122, 107, 120, 104, 96, 102, 104, 100, 93, 91, 97, 103, 107, 111, 115, 111, 102, 100, 107, 107, 101, 99, 101, 101, 96, 87, 83, 86, 84, 124, 40, 
    4, 198, 168, 192, 170, 161, 174, 177, 167, 149, 146, 162, 164, 164, 175, 182, 182, 175, 169, 178, 170, 148, 135, 146, 160, 164, 163, 152, 145, 141, 236, 104, 
    0, 154, 108, 133, 120, 118, 137, 138, 126, 91, 99, 153, 126, 92, 120, 147, 158, 149, 123, 102, 84, 56, 36, 40, 53, 80, 103, 114, 119, 116, 227, 106, 
    0, 157, 109, 138, 129, 126, 145, 143, 125, 78, 139, 284, 241, 124, 130, 166, 165, 110, 66, 84, 99, 87, 47, 15, 7, 13, 42, 80, 120, 130, 241, 112, 
    0, 173, 106, 146, 154, 134, 141, 137, 116, 65, 169, 378, 328, 165, 115, 111, 67, 0, 3, 105, 181, 189, 149, 94, 66, 39, 0, 12, 84, 135, 255, 116, 
    8, 161, 36, 76, 146, 144, 134, 134, 120, 72, 119, 261, 258, 152, 55, 11, 0, 0, 0, 144, 256, 241, 184, 165, 175, 111, 3, 0, 26, 128, 277, 124, 
    37, 129, 0, 0, 104, 137, 130, 132, 138, 112, 83, 122, 157, 175, 91, 27, 38, 9, 14, 168, 311, 255, 151, 160, 203, 160, 29, 0, 0, 90, 289, 135, 
    86, 161, 0, 0, 99, 118, 102, 100, 140, 140, 42, 19, 149, 251, 175, 90, 104, 69, 14, 123, 306, 270, 139, 111, 150, 142, 60, 0, 0, 21, 285, 156, 
    152, 236, 0, 71, 174, 120, 66, 60, 184, 252, 102, 46, 212, 301, 202, 98, 102, 77, 0, 0, 226, 275, 164, 79, 90, 121, 105, 8, 0, 0, 240, 167, 
    186, 301, 83, 252, 271, 135, 44, 41, 270, 508, 354, 178, 282, 318, 201, 114, 108, 45, 0, 0, 197, 302, 242, 120, 77, 132, 154, 88, 0, 0, 151, 135, 
    164, 291, 165, 375, 321, 159, 51, 8, 231, 567, 458, 247, 326, 349, 214, 135, 142, 26, 0, 0, 303, 381, 302, 148, 84, 142, 174, 141, 18, 0, 74, 73, 
    149, 237, 167, 428, 331, 187, 124, 0, 44, 400, 368, 194, 317, 413, 253, 145, 191, 35, 0, 50, 431, 419, 282, 128, 68, 127, 170, 163, 90, 0, 74, 30, 
    149, 191, 175, 448, 282, 153, 204, 40, 0, 219, 233, 125, 309, 483, 337, 196, 245, 83, 0, 125, 477, 390, 232, 102, 43, 79, 115, 150, 137, 82, 136, 42, 
    142, 201, 233, 477, 204, 55, 212, 110, 0, 88, 131, 159, 341, 472, 364, 251, 283, 111, 0, 172, 476, 359, 214, 113, 54, 51, 81, 152, 177, 129, 198, 74, 
    135, 238, 289, 518, 197, 0, 163, 152, 0, 10, 118, 291, 441, 401, 302, 271, 282, 100, 0, 193, 427, 346, 242, 140, 73, 76, 115, 185, 202, 130, 227, 100, 
    134, 293, 304, 548, 279, 8, 121, 203, 53, 3, 148, 437, 533, 349, 218, 212, 213, 92, 15, 180, 357, 346, 260, 132, 66, 82, 131, 179, 156, 97, 242, 120, 
    142, 363, 307, 554, 404, 76, 86, 252, 127, 7, 108, 323, 394, 241, 139, 146, 113, 62, 87, 151, 216, 295, 298, 156, 51, 47, 84, 114, 93, 81, 271, 144, 
    153, 441, 322, 527, 491, 146, 60, 267, 218, 89, 57, 123, 194, 120, 122, 166, 72, 55, 157, 111, 81, 204, 233, 100, 0, 0, 16, 77, 95, 111, 304, 158, 
    138, 497, 349, 481, 533, 224, 46, 225, 299, 200, 92, 42, 104, 103, 179, 279, 111, 57, 198, 211, 154, 161, 125, 19, 0, 0, 8, 97, 141, 144, 314, 158, 
    82, 501, 367, 430, 536, 293, 33, 148, 313, 275, 92, 0, 19, 63, 233, 414, 208, 52, 152, 216, 196, 136, 35, 0, 0, 5, 56, 142, 178, 155, 297, 154, 
    7, 470, 378, 392, 514, 304, 23, 156, 402, 337, 115, 0, 25, 141, 338, 531, 381, 160, 112, 94, 65, 28, 0, 0, 0, 22, 72, 143, 161, 126, 258, 136, 
    0, 433, 406, 391, 475, 240, 0, 221, 628, 631, 366, 207, 236, 319, 439, 542, 457, 287, 172, 71, 23, 31, 57, 85, 96, 102, 105, 145, 154, 123, 240, 140, 
    0, 390, 411, 415, 472, 233, 42, 331, 758, 790, 529, 301, 243, 274, 311, 338, 305, 232, 180, 135, 114, 136, 162, 185, 196, 185, 180, 200, 209, 189, 293, 178, 
    0, 280, 322, 399, 463, 259, 183, 499, 766, 658, 376, 180, 117, 131, 134, 149, 172, 168, 165, 161, 178, 196, 197, 203, 218, 230, 236, 245, 252, 238, 338, 213, 
    0, 189, 177, 297, 345, 195, 286, 659, 714, 449, 240, 148, 145, 162, 158, 164, 177, 177, 173, 172, 188, 204, 208, 217, 242, 272, 278, 270, 264, 252, 379, 254, 
    66, 234, 134, 184, 197, 141, 408, 757, 586, 281, 171, 186, 218, 216, 201, 195, 195, 191, 187, 191, 207, 223, 239, 263, 289, 300, 285, 271, 283, 305, 463, 313, 
    109, 313, 180, 142, 98, 118, 517, 805, 479, 201, 171, 213, 233, 217, 197, 195, 199, 201, 207, 219, 238, 255, 274, 295, 298, 275, 241, 253, 320, 371, 491, 316, 
    112, 338, 241, 176, 83, 100, 500, 739, 426, 203, 198, 226, 248, 230, 204, 196, 198, 205, 218, 236, 252, 256, 268, 283, 274, 242, 229, 283, 364, 362, 398, 243, 
    112, 350, 273, 236, 139, 92, 344, 537, 326, 194, 200, 228, 261, 264, 241, 210, 196, 203, 222, 244, 258, 258, 248, 239, 229, 236, 282, 347, 373, 307, 301, 183, 
    123, 361, 277, 265, 217, 131, 200, 309, 226, 147, 157, 190, 232, 256, 252, 230, 227, 237, 252, 276, 281, 264, 236, 205, 211, 277, 376, 432, 400, 299, 280, 166, 
    147, 385, 305, 295, 291, 245, 222, 252, 220, 178, 165, 180, 196, 211, 218, 213, 231, 266, 310, 356, 351, 312, 270, 238, 264, 371, 491, 514, 424, 316, 293, 170, 
    104, 257, 203, 195, 197, 187, 161, 152, 143, 118, 104, 112, 112, 108, 96, 86, 107, 146, 197, 245, 243, 209, 175, 152, 179, 261, 342, 341, 265, 197, 178, 87, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 54, 58, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 103, 81, 50, 32, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 116, 83, 20, 5, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 1, 0, 19, 89, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 157, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 15, 63, 22, 0, 0, 0, 0, 0, 48, 74, 1, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    3, 234, 53, 77, 34, 0, 0, 0, 66, 197, 157, 48, 74, 89, 23, 0, 0, 0, 0, 0, 64, 100, 37, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    18, 250, 102, 147, 73, 0, 0, 0, 57, 226, 244, 102, 109, 116, 21, 0, 0, 0, 0, 0, 142, 151, 65, 13, 0, 6, 15, 0, 0, 0, 0, 0, 
    30, 228, 115, 179, 91, 0, 0, 0, 0, 137, 193, 84, 100, 148, 46, 0, 0, 0, 0, 37, 206, 171, 54, 4, 0, 4, 21, 7, 0, 0, 0, 0, 
    35, 225, 110, 199, 79, 0, 0, 0, 0, 39, 114, 63, 103, 187, 108, 15, 8, 24, 0, 70, 227, 155, 28, 0, 0, 0, 8, 12, 10, 0, 0, 0, 
    42, 239, 117, 221, 64, 0, 0, 0, 0, 0, 77, 91, 136, 181, 132, 55, 35, 38, 0, 88, 224, 137, 26, 0, 0, 0, 9, 24, 28, 0, 0, 0, 
    50, 265, 139, 249, 78, 0, 0, 0, 0, 0, 61, 160, 210, 167, 105, 62, 44, 26, 0, 66, 193, 124, 33, 4, 0, 3, 29, 37, 23, 0, 0, 0, 
    60, 303, 168, 269, 138, 0, 0, 4, 0, 0, 56, 184, 244, 145, 50, 30, 23, 1, 0, 31, 123, 100, 47, 2, 0, 0, 27, 18, 0, 0, 0, 0, 
    69, 356, 207, 281, 215, 18, 0, 50, 0, 0, 0, 108, 143, 70, 0, 0, 0, 0, 0, 0, 23, 53, 51, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    71, 396, 243, 284, 260, 83, 8, 82, 84, 0, 0, 0, 21, 19, 0, 18, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 398, 260, 277, 273, 145, 20, 99, 130, 41, 0, 0, 0, 33, 34, 90, 34, 0, 25, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 362, 259, 251, 257, 186, 43, 109, 168, 72, 3, 0, 0, 65, 103, 173, 101, 0, 0, 25, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    3, 323, 265, 225, 236, 188, 63, 143, 260, 164, 46, 0, 62, 151, 206, 269, 203, 49, 0, 0, 0, 0, 0, 0, 16, 39, 35, 22, 19, 0, 0, 37, 
    0, 313, 304, 234, 226, 174, 70, 203, 389, 367, 219, 135, 165, 240, 278, 298, 254, 144, 70, 37, 13, 34, 70, 106, 134, 134, 124, 115, 107, 85, 53, 92, 
    0, 302, 330, 274, 260, 211, 126, 274, 442, 429, 291, 185, 177, 204, 215, 212, 197, 155, 123, 112, 117, 143, 173, 199, 220, 225, 216, 210, 208, 198, 155, 156, 
    12, 265, 288, 290, 293, 240, 205, 349, 427, 347, 227, 136, 137, 150, 149, 149, 160, 157, 154, 164, 185, 211, 226, 238, 254, 267, 269, 269, 272, 268, 210, 198, 
    52, 258, 219, 240, 268, 229, 257, 375, 385, 246, 166, 148, 168, 186, 183, 176, 181, 185, 187, 198, 215, 236, 249, 261, 278, 294, 299, 299, 302, 305, 246, 234, 
    98, 306, 215, 202, 222, 222, 309, 386, 316, 159, 140, 189, 219, 221, 212, 205, 204, 205, 209, 221, 239, 261, 279, 294, 304, 309, 306, 308, 329, 350, 291, 274, 
    106, 344, 259, 211, 195, 209, 345, 419, 282, 123, 161, 217, 239, 230, 212, 209, 212, 219, 229, 245, 265, 282, 298, 313, 315, 304, 295, 313, 350, 370, 303, 270, 
    104, 355, 290, 256, 210, 190, 316, 406, 267, 133, 189, 233, 249, 243, 224, 215, 219, 230, 246, 263, 276, 286, 293, 302, 305, 300, 309, 334, 358, 350, 257, 219, 
    111, 361, 304, 293, 254, 194, 241, 310, 226, 138, 189, 222, 249, 255, 245, 232, 228, 241, 258, 271, 281, 281, 277, 276, 284, 312, 344, 370, 364, 316, 210, 173, 
    112, 365, 304, 301, 288, 227, 198, 226, 182, 137, 165, 191, 217, 230, 235, 234, 241, 258, 278, 292, 289, 275, 262, 258, 281, 337, 391, 407, 364, 301, 201, 160, 
    84, 322, 272, 265, 265, 240, 194, 182, 166, 136, 143, 155, 165, 169, 168, 165, 181, 214, 248, 276, 276, 252, 231, 223, 249, 314, 375, 382, 323, 264, 200, 159, 
    15, 173, 142, 136, 135, 126, 109, 91, 85, 74, 70, 77, 79, 73, 66, 55, 59, 80, 107, 135, 144, 129, 114, 106, 115, 152, 192, 199, 168, 132, 105, 82, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=24
    161, 103, 68, 58, 52, 56, 59, 55, 55, 60, 63, 62, 59, 62, 64, 63, 59, 58, 53, 47, 43, 46, 56, 60, 58, 52, 50, 54, 55, 50, 4, 0, 
    264, 259, 227, 213, 201, 203, 206, 199, 198, 205, 208, 196, 189, 203, 218, 216, 201, 187, 184, 182, 177, 178, 193, 209, 211, 203, 193, 186, 179, 168, 86, 24, 
    319, 323, 299, 291, 280, 281, 281, 275, 273, 287, 280, 228, 201, 235, 277, 277, 261, 257, 257, 235, 200, 174, 190, 226, 262, 283, 282, 271, 252, 232, 131, 56, 
    316, 317, 291, 289, 282, 285, 286, 280, 282, 310, 303, 216, 156, 190, 256, 274, 269, 271, 251, 184, 94, 38, 41, 95, 157, 212, 263, 291, 277, 248, 136, 56, 
    304, 300, 296, 319, 308, 295, 291, 286, 289, 330, 346, 277, 188, 183, 229, 252, 241, 243, 216, 131, 24, 0, 0, 0, 33, 96, 187, 285, 308, 269, 141, 54, 
    271, 259, 292, 358, 343, 308, 291, 287, 287, 325, 358, 329, 241, 156, 139, 144, 133, 150, 176, 121, 25, 0, 0, 3, 0, 20, 108, 237, 309, 288, 151, 54, 
    200, 143, 204, 322, 331, 307, 291, 291, 277, 279, 293, 282, 211, 89, 16, 15, 44, 92, 167, 165, 79, 21, 32, 64, 45, 12, 44, 156, 282, 309, 171, 57, 
    109, 0, 35, 190, 245, 274, 292, 304, 251, 176, 153, 176, 140, 40, 0, 0, 34, 83, 187, 244, 158, 56, 29, 69, 70, 23, 2, 73, 215, 310, 195, 71, 
    60, 0, 0, 71, 136, 219, 285, 325, 229, 59, 0, 51, 78, 21, 0, 0, 39, 83, 190, 272, 190, 55, 0, 11, 46, 18, 0, 0, 127, 273, 214, 101, 
    80, 0, 0, 32, 80, 167, 271, 361, 293, 76, 0, 3, 53, 3, 0, 0, 2, 48, 166, 228, 129, 6, 0, 0, 21, 26, 0, 0, 30, 187, 197, 124, 
    109, 14, 28, 43, 71, 140, 244, 371, 405, 231, 96, 86, 72, 0, 0, 0, 0, 0, 124, 187, 69, 0, 0, 0, 45, 55, 1, 0, 0, 72, 119, 105, 
    114, 46, 76, 57, 82, 149, 218, 317, 420, 326, 216, 190, 126, 0, 0, 0, 0, 0, 98, 178, 59, 0, 0, 18, 72, 94, 49, 0, 0, 0, 25, 48, 
    109, 40, 51, 35, 86, 189, 228, 243, 323, 329, 262, 230, 156, 14, 0, 0, 0, 0, 102, 187, 65, 0, 0, 2, 50, 92, 78, 15, 0, 0, 0, 3, 
    108, 30, 7, 0, 39, 192, 231, 216, 255, 309, 270, 199, 113, 37, 10, 0, 0, 15, 135, 190, 70, 0, 0, 0, 29, 73, 76, 35, 1, 22, 9, 1, 
    117, 29, 0, 0, 0, 115, 208, 196, 198, 289, 288, 183, 80, 60, 101, 96, 45, 76, 178, 208, 101, 19, 0, 0, 31, 75, 85, 75, 77, 106, 64, 23, 
    130, 16, 0, 0, 0, 6, 158, 155, 150, 258, 316, 231, 119, 103, 146, 151, 115, 126, 186, 230, 182, 92, 3, 2, 64, 126, 142, 143, 158, 176, 96, 32, 
    140, 0, 0, 0, 0, 0, 100, 120, 107, 191, 310, 288, 219, 165, 136, 116, 106, 146, 183, 227, 228, 167, 62, 38, 99, 174, 199, 198, 202, 207, 107, 34, 
    162, 0, 0, 0, 0, 0, 45, 104, 69, 92, 197, 243, 215, 165, 87, 26, 31, 128, 166, 167, 178, 164, 114, 99, 130, 175, 207, 211, 212, 216, 118, 40, 
    212, 27, 0, 0, 0, 0, 0, 76, 42, 8, 72, 164, 191, 158, 58, 0, 0, 76, 154, 131, 104, 117, 116, 109, 115, 155, 199, 225, 229, 226, 127, 46, 
    269, 91, 7, 0, 0, 0, 0, 40, 0, 0, 0, 43, 122, 111, 17, 0, 0, 0, 108, 150, 127, 84, 57, 48, 58, 112, 176, 222, 227, 218, 119, 48, 
    300, 131, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 14, 83, 65, 10, 0, 0, 0, 13, 105, 148, 151, 144, 54, 16, 
    288, 140, 37, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 62, 64, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    224, 120, 74, 23, 0, 0, 9, 27, 0, 0, 0, 0, 40, 91, 103, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    110, 53, 87, 69, 0, 29, 76, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 74, 85, 147, 134, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 98, 185, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 174, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 97, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 44, 46, 35, 13, 0, 0, 0, 12, 41, 49, 25, 0, 0, 0, 0, 0, 
    
    -- channel=25
    222, 253, 191, 181, 164, 168, 175, 171, 167, 169, 173, 176, 178, 183, 186, 181, 173, 167, 168, 169, 164, 166, 174, 179, 172, 159, 150, 148, 148, 140, 101, 0, 
    372, 403, 355, 339, 321, 330, 336, 327, 321, 320, 321, 316, 313, 329, 344, 340, 327, 313, 308, 306, 294, 287, 301, 325, 334, 328, 317, 303, 286, 266, 189, 0, 
    391, 408, 367, 353, 338, 351, 361, 351, 343, 343, 351, 320, 263, 279, 339, 351, 335, 320, 311, 291, 249, 209, 213, 252, 298, 335, 352, 346, 324, 295, 209, 0, 
    389, 405, 368, 361, 348, 359, 368, 358, 354, 377, 427, 394, 270, 246, 323, 346, 321, 296, 289, 272, 202, 136, 112, 132, 181, 243, 309, 358, 362, 325, 219, 0, 
    385, 395, 379, 407, 397, 376, 367, 356, 357, 403, 494, 472, 313, 236, 261, 262, 239, 230, 264, 263, 192, 127, 102, 113, 130, 156, 220, 319, 376, 355, 234, 0, 
    349, 318, 316, 418, 441, 399, 365, 354, 352, 381, 455, 432, 303, 200, 145, 127, 145, 174, 243, 275, 223, 144, 125, 149, 146, 114, 142, 250, 356, 374, 256, 0, 
    276, 159, 153, 348, 427, 399, 365, 356, 346, 332, 346, 339, 274, 174, 78, 78, 129, 168, 248, 316, 283, 176, 135, 181, 176, 106, 86, 174, 305, 375, 282, 0, 
    228, 44, 22, 264, 354, 351, 353, 359, 326, 238, 171, 217, 266, 181, 64, 77, 148, 186, 252, 342, 328, 203, 119, 146, 159, 106, 58, 100, 228, 351, 306, 25, 
    229, 38, 27, 257, 302, 293, 339, 398, 380, 219, 67, 137, 247, 172, 64, 72, 131, 157, 211, 322, 331, 196, 83, 83, 118, 112, 62, 49, 137, 285, 304, 61, 
    263, 95, 123, 295, 269, 243, 319, 442, 513, 361, 144, 145, 234, 149, 43, 53, 88, 98, 154, 297, 318, 180, 65, 53, 113, 148, 91, 29, 55, 188, 251, 68, 
    282, 147, 218, 335, 248, 209, 284, 423, 553, 478, 276, 231, 277, 153, 19, 25, 52, 36, 113, 309, 334, 193, 76, 60, 135, 193, 141, 54, 19, 99, 163, 31, 
    271, 164, 248, 332, 245, 228, 270, 323, 451, 477, 340, 295, 333, 187, 19, 13, 47, 15, 111, 347, 345, 191, 77, 72, 153, 214, 186, 112, 40, 62, 95, 0, 
    256, 156, 241, 283, 198, 255, 306, 262, 344, 419, 349, 356, 394, 256, 89, 62, 73, 29, 145, 378, 330, 158, 50, 50, 122, 190, 193, 154, 90, 76, 80, 0, 
    259, 163, 224, 204, 106, 228, 339, 245, 274, 382, 371, 391, 374, 252, 160, 155, 139, 71, 187, 390, 318, 145, 55, 63, 119, 180, 202, 190, 149, 135, 117, 0, 
    276, 187, 218, 145, 19, 151, 315, 249, 237, 355, 423, 441, 365, 240, 210, 234, 198, 132, 236, 393, 322, 172, 72, 63, 117, 191, 231, 237, 213, 211, 179, 0, 
    295, 201, 210, 132, 0, 75, 278, 259, 214, 318, 461, 477, 357, 243, 235, 259, 219, 185, 280, 395, 361, 257, 136, 75, 132, 220, 265, 277, 259, 262, 220, 0, 
    317, 208, 198, 156, 0, 8, 229, 271, 202, 255, 403, 437, 336, 238, 222, 222, 194, 218, 306, 345, 338, 305, 192, 103, 144, 228, 273, 294, 285, 292, 240, 0, 
    348, 232, 199, 190, 22, 0, 164, 286, 215, 198, 247, 279, 286, 235, 211, 167, 119, 218, 308, 260, 236, 251, 175, 111, 142, 209, 265, 307, 315, 316, 246, 0, 
    387, 284, 221, 219, 71, 0, 91, 261, 211, 149, 148, 200, 282, 270, 235, 131, 39, 169, 308, 274, 226, 193, 127, 108, 145, 211, 289, 347, 348, 331, 248, 0, 
    417, 343, 254, 239, 132, 0, 58, 218, 163, 23, 0, 89, 208, 245, 255, 112, 0, 61, 216, 234, 200, 144, 80, 63, 113, 199, 305, 372, 357, 323, 237, 0, 
    415, 372, 269, 241, 162, 14, 62, 224, 135, 0, 0, 0, 158, 252, 290, 177, 22, 27, 104, 111, 89, 47, 20, 18, 57, 137, 239, 297, 276, 243, 167, 0, 
    381, 371, 285, 248, 156, 17, 89, 295, 216, 2, 0, 1, 184, 287, 319, 245, 114, 53, 57, 33, 1, 0, 0, 0, 0, 36, 101, 141, 129, 106, 52, 0, 
    303, 314, 286, 280, 184, 78, 187, 385, 316, 102, 0, 35, 161, 204, 204, 164, 90, 33, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    181, 181, 214, 285, 245, 185, 320, 433, 303, 73, 0, 0, 27, 22, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 18, 78, 202, 253, 286, 411, 393, 160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 80, 182, 318, 433, 285, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 89, 279, 408, 214, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 191, 322, 178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50, 171, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 24, 34, 31, 11, 0, 0, 0, 0, 18, 48, 38, 0, 0, 0, 0, 0, 
    47, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 2, 21, 38, 51, 56, 44, 22, 7, 7, 29, 68, 92, 73, 21, 0, 0, 0, 0, 
    
    -- channel=26
    127, 124, 139, 137, 146, 151, 149, 152, 153, 152, 147, 143, 148, 153, 154, 154, 155, 152, 144, 132, 126, 124, 123, 126, 129, 136, 144, 149, 149, 146, 127, 105, 
    206, 193, 207, 198, 207, 214, 213, 215, 219, 221, 215, 216, 227, 231, 227, 224, 218, 211, 197, 178, 170, 172, 172, 165, 159, 165, 178, 196, 205, 203, 153, 99, 
    243, 234, 255, 244, 247, 248, 246, 248, 249, 249, 242, 250, 285, 290, 260, 237, 222, 206, 200, 201, 204, 221, 231, 229, 217, 202, 203, 213, 223, 228, 174, 107, 
    238, 226, 249, 242, 247, 248, 244, 246, 249, 244, 206, 170, 217, 260, 228, 195, 183, 181, 175, 150, 155, 176, 210, 230, 234, 236, 223, 209, 207, 218, 170, 107, 
    217, 199, 225, 217, 231, 251, 251, 253, 258, 254, 202, 124, 152, 207, 215, 199, 195, 196, 163, 114, 97, 98, 116, 146, 179, 208, 239, 225, 201, 201, 164, 107, 
    200, 194, 244, 226, 219, 246, 256, 255, 260, 274, 256, 189, 164, 198, 228, 221, 194, 197, 162, 93, 70, 91, 96, 88, 97, 149, 209, 234, 209, 189, 147, 102, 
    178, 202, 295, 271, 250, 255, 258, 251, 249, 259, 257, 222, 187, 163, 180, 180, 155, 160, 154, 84, 48, 99, 131, 106, 81, 102, 161, 229, 229, 191, 133, 97, 
    117, 156, 280, 287, 276, 280, 268, 250, 245, 265, 290, 257, 178, 131, 137, 132, 111, 128, 163, 118, 58, 91, 154, 154, 120, 105, 138, 202, 244, 209, 121, 80, 
    49, 75, 190, 222, 264, 280, 265, 227, 182, 185, 257, 243, 162, 121, 131, 141, 128, 134, 186, 175, 107, 108, 156, 179, 150, 114, 120, 174, 241, 236, 127, 64, 
    14, 21, 112, 139, 222, 276, 267, 217, 74, 0, 93, 164, 122, 116, 136, 141, 138, 160, 195, 173, 120, 117, 125, 146, 140, 105, 97, 132, 208, 255, 159, 71, 
    27, 36, 68, 97, 193, 262, 261, 243, 111, 0, 16, 100, 83, 102, 149, 144, 131, 162, 208, 135, 66, 94, 105, 125, 123, 97, 90, 101, 156, 231, 189, 100, 
    28, 67, 79, 78, 176, 230, 240, 274, 205, 56, 73, 124, 80, 73, 154, 159, 116, 154, 203, 108, 35, 86, 112, 132, 132, 107, 82, 83, 112, 179, 182, 121, 
    25, 77, 90, 80, 191, 222, 199, 229, 238, 123, 121, 155, 97, 50, 103, 137, 100, 127, 181, 94, 41, 96, 131, 147, 151, 139, 115, 91, 100, 148, 146, 117, 
    22, 65, 67, 71, 219, 251, 198, 212, 238, 173, 140, 134, 123, 83, 79, 96, 87, 123, 162, 83, 36, 95, 123, 130, 138, 141, 126, 101, 106, 145, 129, 105, 
    20, 53, 45, 38, 199, 274, 219, 205, 240, 204, 132, 70, 76, 113, 105, 81, 81, 134, 161, 97, 50, 80, 100, 118, 120, 107, 104, 98, 113, 157, 138, 102, 
    15, 34, 45, 5, 124, 248, 211, 180, 224, 215, 120, 1, 0, 91, 123, 120, 109, 141, 176, 134, 61, 55, 96, 128, 129, 109, 101, 119, 152, 190, 152, 106, 
    2, 2, 41, 0, 50, 190, 188, 151, 199, 247, 179, 97, 66, 114, 152, 150, 162, 170, 183, 181, 140, 69, 50, 99, 126, 127, 134, 155, 191, 214, 157, 104, 
    0, 0, 29, 0, 12, 142, 175, 110, 137, 213, 227, 186, 139, 142, 144, 142, 189, 183, 167, 211, 210, 139, 106, 117, 138, 168, 183, 188, 206, 222, 159, 100, 
    8, 0, 15, 0, 0, 94, 163, 100, 92, 142, 189, 191, 139, 130, 103, 90, 178, 198, 129, 103, 136, 146, 131, 128, 147, 173, 201, 201, 212, 227, 160, 99, 
    53, 0, 18, 14, 0, 61, 134, 101, 99, 147, 199, 215, 175, 155, 86, 49, 148, 220, 171, 114, 80, 100, 128, 135, 139, 160, 191, 190, 195, 209, 150, 97, 
    93, 0, 32, 43, 3, 58, 107, 39, 31, 145, 219, 212, 167, 102, 27, 0, 23, 135, 187, 174, 146, 120, 119, 122, 126, 157, 178, 177, 175, 184, 131, 99, 
    96, 0, 10, 39, 26, 96, 136, 4, 0, 0, 38, 57, 25, 0, 0, 0, 0, 0, 64, 108, 109, 84, 45, 20, 26, 61, 97, 109, 110, 114, 85, 95, 
    64, 0, 0, 0, 0, 70, 104, 3, 0, 0, 0, 0, 3, 10, 13, 0, 0, 4, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 
    27, 3, 1, 0, 0, 35, 42, 0, 0, 0, 0, 17, 46, 57, 61, 42, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 
    0, 7, 56, 9, 7, 62, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 
    0, 0, 32, 44, 52, 58, 0, 0, 4, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 19, 76, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 45, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 63, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 57, 55, 34, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 64, 45, 48, 55, 42, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 45, 5, 5, 42, 55, 16, 0, 0, 0, 0, 0, 
    0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 29, 26, 0, 0, 0, 20, 0, 0, 7, 38, 48, 0, 0, 0, 0, 0, 
    8, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 26, 21, 0, 0, 0, 0, 10, 0, 0, 30, 60, 42, 0, 0, 0, 0, 
    0, 93, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 40, 14, 0, 0, 0, 8, 25, 13, 2, 35, 68, 73, 16, 0, 0, 0, 
    0, 84, 17, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 8, 59, 22, 0, 0, 0, 55, 33, 12, 0, 25, 60, 78, 54, 0, 0, 0, 
    11, 81, 18, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 14, 0, 51, 35, 0, 0, 19, 70, 21, 1, 0, 9, 36, 71, 71, 28, 16, 0, 
    15, 86, 41, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 2, 42, 31, 0, 0, 23, 60, 19, 9, 4, 6, 13, 50, 65, 31, 39, 4, 
    8, 88, 73, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 15, 0, 0, 20, 50, 21, 24, 21, 16, 13, 32, 41, 0, 20, 0, 
    0, 89, 84, 142, 33, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 3, 0, 0, 0, 0, 42, 35, 31, 24, 20, 16, 12, 0, 0, 0, 0, 
    0, 98, 85, 164, 101, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 6, 32, 23, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 124, 102, 178, 170, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 140, 130, 179, 206, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 116, 138, 169, 209, 137, 38, 9, 16, 16, 0, 0, 0, 0, 0, 90, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 59, 111, 135, 183, 147, 58, 67, 98, 84, 23, 0, 0, 0, 24, 134, 116, 7, 0, 0, 0, 32, 33, 41, 24, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 90, 106, 159, 124, 45, 81, 191, 195, 98, 26, 29, 28, 73, 151, 159, 92, 54, 22, 28, 61, 103, 141, 129, 73, 0, 0, 0, 0, 0, 0, 
    0, 16, 98, 110, 150, 94, 21, 57, 212, 298, 225, 156, 131, 125, 122, 147, 173, 156, 142, 141, 143, 182, 232, 274, 286, 248, 188, 142, 130, 135, 152, 85, 
    3, 60, 107, 123, 143, 89, 26, 69, 188, 281, 258, 218, 183, 158, 145, 153, 183, 204, 224, 254, 292, 326, 351, 373, 391, 390, 369, 344, 339, 350, 336, 194, 
    131, 156, 124, 122, 121, 72, 28, 112, 202, 237, 224, 219, 239, 221, 215, 227, 259, 293, 319, 346, 376, 400, 416, 425, 438, 454, 458, 454, 453, 461, 441, 255, 
    237, 299, 210, 123, 83, 33, 26, 152, 234, 229, 244, 298, 339, 344, 344, 345, 356, 371, 385, 401, 418, 436, 451, 463, 474, 483, 488, 492, 496, 505, 486, 289, 
    302, 433, 356, 210, 82, 20, 71, 200, 256, 238, 294, 373, 403, 404, 395, 390, 393, 401, 414, 432, 452, 469, 484, 498, 501, 501, 495, 502, 519, 535, 511, 313, 
    320, 490, 468, 338, 169, 43, 107, 249, 279, 271, 354, 404, 422, 419, 405, 398, 403, 415, 430, 453, 475, 492, 503, 512, 513, 504, 501, 515, 537, 544, 498, 291, 
    321, 506, 523, 449, 308, 140, 110, 244, 303, 303, 379, 408, 421, 431, 423, 413, 414, 426, 444, 466, 485, 499, 499, 501, 506, 514, 535, 557, 568, 538, 449, 249, 
    319, 514, 548, 506, 428, 279, 181, 214, 311, 326, 374, 393, 410, 425, 431, 425, 422, 434, 454, 475, 492, 499, 495, 485, 488, 523, 570, 599, 588, 528, 427, 233, 
    312, 512, 548, 522, 484, 397, 297, 270, 314, 349, 363, 373, 387, 397, 404, 405, 412, 429, 456, 482, 495, 495, 482, 466, 468, 510, 575, 615, 597, 542, 442, 240, 
    253, 431, 471, 454, 437, 401, 346, 308, 315, 331, 334, 331, 331, 326, 317, 309, 313, 333, 365, 404, 427, 423, 404, 382, 372, 401, 465, 520, 514, 477, 401, 238, 
    142, 233, 272, 264, 254, 239, 220, 202, 198, 201, 204, 201, 199, 192, 179, 163, 156, 163, 185, 210, 229, 235, 227, 217, 204, 210, 236, 270, 285, 276, 234, 147, 
    
    -- channel=28
    74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    278, 111, 148, 124, 139, 147, 126, 121, 127, 139, 137, 121, 140, 163, 155, 146, 132, 131, 141, 124, 114, 136, 159, 158, 141, 126, 111, 113, 114, 105, 0, 0, 
    331, 181, 240, 224, 240, 240, 213, 210, 218, 236, 185, 102, 171, 273, 255, 231, 225, 222, 207, 167, 138, 165, 214, 247, 262, 249, 217, 191, 173, 163, 46, 1, 
    329, 176, 240, 222, 235, 244, 220, 218, 235, 275, 195, 0, 38, 222, 254, 234, 239, 248, 207, 93, 18, 4, 56, 131, 181, 232, 253, 223, 174, 146, 38, 0, 
    322, 186, 279, 237, 204, 228, 229, 228, 246, 311, 287, 69, 26, 170, 246, 246, 245, 271, 208, 50, 0, 0, 0, 0, 9, 93, 228, 275, 215, 141, 20, 0, 
    281, 181, 361, 319, 211, 197, 229, 227, 233, 280, 318, 207, 91, 89, 159, 201, 163, 208, 206, 32, 0, 0, 0, 0, 0, 0, 142, 283, 269, 168, 1, 0, 
    190, 89, 376, 344, 215, 189, 233, 231, 205, 213, 266, 226, 94, 0, 16, 82, 44, 110, 211, 94, 0, 0, 0, 0, 0, 0, 47, 242, 313, 225, 1, 0, 
    88, 0, 244, 218, 149, 186, 250, 237, 137, 92, 203, 230, 60, 0, 0, 35, 4, 52, 232, 212, 0, 0, 0, 56, 6, 0, 0, 144, 315, 293, 36, 0, 
    58, 0, 76, 13, 24, 162, 273, 256, 29, 0, 14, 139, 3, 0, 0, 22, 25, 51, 240, 278, 55, 0, 0, 38, 46, 0, 0, 22, 251, 347, 115, 0, 
    118, 0, 3, 0, 0, 121, 291, 376, 128, 0, 0, 34, 0, 0, 0, 0, 0, 60, 259, 235, 14, 0, 0, 0, 42, 0, 0, 0, 125, 322, 179, 4, 
    166, 0, 23, 0, 0, 84, 238, 466, 370, 0, 0, 29, 0, 0, 0, 0, 0, 34, 306, 201, 0, 0, 0, 0, 58, 0, 0, 0, 0, 191, 151, 43, 
    151, 68, 78, 0, 0, 87, 126, 399, 501, 177, 8, 103, 0, 0, 0, 0, 0, 0, 330, 195, 0, 0, 0, 9, 82, 25, 0, 0, 0, 34, 40, 31, 
    130, 70, 62, 0, 13, 171, 75, 220, 438, 232, 78, 106, 0, 0, 0, 0, 0, 0, 328, 174, 0, 0, 0, 13, 81, 68, 13, 0, 0, 0, 0, 0, 
    126, 43, 3, 0, 40, 253, 104, 110, 346, 253, 107, 8, 0, 0, 0, 0, 0, 4, 318, 156, 0, 0, 0, 0, 27, 37, 15, 0, 0, 0, 0, 0, 
    136, 18, 0, 0, 0, 249, 128, 33, 238, 272, 154, 0, 0, 0, 0, 0, 0, 32, 283, 142, 0, 0, 0, 0, 46, 37, 17, 0, 0, 0, 0, 0, 
    154, 0, 0, 0, 0, 175, 123, 0, 123, 295, 261, 48, 0, 0, 29, 12, 0, 44, 197, 158, 0, 0, 0, 0, 89, 93, 63, 22, 11, 53, 0, 0, 
    178, 0, 0, 0, 0, 80, 144, 0, 0, 255, 302, 193, 11, 0, 30, 6, 51, 68, 88, 135, 140, 0, 0, 0, 120, 155, 122, 63, 56, 86, 0, 0, 
    219, 0, 0, 0, 0, 0, 169, 0, 0, 56, 201, 227, 86, 24, 0, 0, 62, 110, 0, 18, 146, 83, 6, 61, 143, 169, 148, 76, 60, 107, 0, 0, 
    289, 0, 0, 0, 0, 0, 158, 30, 0, 0, 50, 179, 104, 45, 0, 0, 0, 161, 26, 0, 0, 42, 72, 109, 142, 137, 128, 72, 66, 126, 2, 0, 
    363, 0, 0, 0, 0, 0, 117, 0, 0, 0, 25, 186, 135, 79, 0, 0, 0, 120, 126, 63, 22, 23, 80, 129, 152, 153, 146, 98, 80, 131, 18, 0, 
    422, 0, 0, 0, 0, 0, 140, 0, 0, 0, 0, 66, 62, 21, 0, 0, 0, 0, 43, 92, 98, 47, 22, 38, 80, 132, 154, 119, 92, 123, 18, 0, 
    470, 44, 0, 0, 0, 0, 183, 3, 0, 0, 0, 0, 32, 62, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 66, 53, 19, 25, 0, 0, 
    482, 206, 5, 0, 0, 0, 119, 0, 0, 0, 0, 19, 130, 186, 176, 106, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    390, 319, 225, 29, 0, 0, 76, 0, 0, 0, 0, 32, 87, 117, 121, 93, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    202, 212, 309, 212, 80, 126, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 9, 176, 259, 267, 272, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    72, 0, 6, 155, 346, 431, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 19, 261, 485, 201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 0, 0, 0, 93, 342, 281, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    77, 0, 0, 0, 0, 100, 157, 26, 0, 0, 32, 41, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    140, 0, 0, 0, 0, 0, 17, 0, 0, 0, 32, 47, 52, 50, 52, 63, 52, 17, 0, 0, 0, 0, 0, 10, 37, 0, 0, 0, 0, 0, 0, 0, 
    200, 108, 74, 87, 84, 78, 79, 79, 68, 76, 96, 102, 103, 105, 120, 150, 170, 174, 151, 100, 62, 61, 91, 149, 200, 192, 114, 34, 20, 47, 26, 6, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    82, 36, 36, 30, 22, 24, 23, 19, 18, 20, 27, 28, 28, 32, 34, 33, 29, 24, 22, 20, 19, 22, 27, 30, 25, 18, 14, 14, 14, 7, 0, 0, 
    188, 180, 174, 174, 164, 162, 159, 154, 148, 146, 149, 152, 154, 165, 174, 172, 159, 149, 143, 142, 137, 134, 145, 159, 167, 164, 151, 138, 124, 107, 73, 0, 
    211, 218, 215, 221, 214, 215, 213, 208, 202, 197, 190, 169, 152, 181, 217, 225, 221, 203, 178, 144, 102, 86, 100, 138, 170, 191, 199, 188, 173, 152, 115, 0, 
    212, 218, 216, 228, 223, 224, 222, 216, 212, 220, 240, 210, 155, 175, 220, 235, 226, 195, 148, 87, 32, 0, 0, 12, 57, 111, 157, 187, 187, 163, 123, 0, 
    214, 229, 233, 253, 241, 227, 223, 217, 212, 234, 300, 296, 215, 169, 179, 176, 149, 123, 104, 67, 15, 0, 0, 0, 0, 10, 86, 157, 189, 173, 130, 0, 
    192, 189, 202, 250, 246, 224, 221, 217, 208, 211, 260, 269, 200, 115, 60, 47, 36, 54, 86, 74, 28, 1, 0, 1, 0, 0, 11, 106, 182, 191, 144, 5, 
    128, 70, 80, 167, 214, 211, 219, 222, 205, 184, 191, 190, 149, 55, 0, 0, 0, 17, 105, 134, 81, 19, 14, 36, 25, 0, 0, 48, 148, 199, 158, 8, 
    83, 0, 0, 64, 142, 178, 209, 212, 177, 110, 76, 93, 97, 46, 0, 0, 0, 23, 120, 186, 156, 50, 1, 21, 24, 0, 0, 0, 98, 192, 176, 18, 
    100, 0, 0, 21, 90, 145, 197, 221, 176, 57, 0, 25, 81, 51, 0, 0, 0, 13, 93, 160, 154, 54, 0, 0, 0, 0, 0, 0, 23, 152, 188, 38, 
    143, 26, 0, 45, 76, 123, 185, 285, 308, 195, 60, 56, 86, 49, 0, 0, 0, 0, 51, 116, 108, 38, 0, 0, 0, 0, 0, 0, 0, 69, 149, 47, 
    147, 93, 66, 106, 90, 110, 153, 294, 405, 346, 198, 148, 135, 52, 0, 0, 0, 0, 39, 118, 104, 50, 12, 0, 11, 15, 0, 0, 0, 0, 59, 22, 
    127, 110, 99, 140, 123, 143, 146, 221, 335, 354, 250, 199, 180, 64, 0, 0, 0, 0, 51, 155, 137, 65, 23, 1, 22, 39, 17, 0, 0, 0, 0, 0, 
    108, 99, 90, 123, 124, 177, 172, 155, 251, 286, 216, 180, 195, 117, 17, 0, 0, 0, 91, 174, 145, 58, 4, 0, 0, 20, 19, 0, 0, 0, 0, 0, 
    109, 99, 84, 72, 65, 150, 194, 129, 171, 212, 183, 149, 159, 142, 90, 44, 23, 2, 129, 191, 142, 48, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 
    125, 106, 86, 42, 0, 66, 162, 100, 109, 171, 208, 178, 122, 115, 124, 105, 71, 38, 134, 193, 155, 61, 3, 0, 0, 19, 35, 47, 38, 41, 40, 0, 
    148, 107, 83, 44, 0, 0, 111, 90, 71, 169, 288, 288, 210, 143, 117, 108, 82, 59, 136, 197, 185, 104, 18, 0, 17, 67, 85, 90, 79, 78, 71, 0, 
    175, 104, 69, 64, 0, 0, 74, 87, 28, 118, 246, 282, 220, 123, 70, 50, 47, 52, 107, 151, 187, 152, 68, 18, 47, 87, 103, 94, 89, 102, 100, 0, 
    212, 117, 57, 72, 0, 0, 48, 105, 34, 39, 112, 162, 152, 80, 26, 0, 0, 50, 80, 53, 79, 112, 86, 30, 28, 59, 81, 98, 108, 132, 128, 0, 
    250, 149, 62, 75, 0, 0, 16, 101, 56, 15, 12, 84, 118, 86, 47, 0, 0, 38, 116, 77, 59, 50, 39, 17, 18, 35, 73, 117, 140, 157, 147, 6, 
    272, 180, 74, 78, 32, 0, 0, 45, 0, 0, 0, 2, 41, 60, 57, 0, 0, 0, 81, 118, 81, 29, 0, 0, 5, 51, 107, 153, 163, 165, 147, 12, 
    273, 199, 82, 77, 52, 0, 19, 43, 0, 0, 0, 0, 0, 55, 91, 50, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 62, 107, 110, 102, 85, 0, 
    270, 219, 102, 74, 37, 0, 29, 98, 55, 0, 0, 0, 81, 171, 198, 171, 84, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    251, 251, 169, 107, 47, 0, 72, 144, 157, 70, 3, 42, 109, 168, 175, 142, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    151, 187, 203, 180, 119, 97, 162, 180, 147, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 27, 111, 173, 165, 175, 203, 178, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 84, 169, 243, 226, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 123, 282, 266, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 233, 279, 131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 86, 167, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 2, 14, 0, 0, 0, 0, 0, 0, 
    67, 55, 30, 30, 30, 28, 25, 16, 7, 2, 6, 10, 10, 9, 18, 38, 62, 82, 88, 74, 52, 37, 42, 67, 109, 137, 115, 62, 22, 6, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 2, 4, 5, 4, 3, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 7, 20, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 3, 2, 0, 0, 0, 0, 0, 0, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 9, 0, 
    0, 3, 2, 0, 0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 6, 0, 
    1, 10, 8, 7, 6, 0, 0, 0, 4, 15, 9, 7, 6, 4, 5, 5, 3, 2, 0, 0, 3, 5, 7, 2, 0, 0, 0, 0, 5, 10, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
