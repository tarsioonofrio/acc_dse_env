library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=2
    -7789, -6336, 3831, 3759, 9293, -10212, 14756, -10861, 8263, -7640,

    -- weights
    -- layer=2 filter=0 channel=0
    7, 27, -17, 13, 37, 7, 8, 24, -5, -93, 4, -9, 6, -34, 12, -59, -19, 37, -2, 4, -32, -23, -31, -52, -24, 3, -43, 15, -2, -22, 77, 11, -13, -61, -24, 5, -3, 10, 13, -1, -30, -19, -9, -23, 33, -8, 24, 9, 0, 50, 10, 45, -7, -67, 9, -64, -7, -23, -26, 0, -7, -18, 0, 22, 47, 17, -10, 32, 11, 0, -19, 8, 0, -53, -3, 0, -55, -10, 22, -18, -15, 37, -5, -44, 6, -12, -1, -46, -42, -14, -35, 5, -8, 14, 30, 13, 16, 6, -28, 15, -19, 23, 2, 34, -1, -21, 17, 40, -57, 6, 13, 2, 31, 32, 15, -14, -1, -49, 14, -6, -34, 18, -60, 11, 6, -6, 1, -6, 54, 45, -49, 19, -11, -8, -12, 6, 1, -50, 19, 11, -12, -63, 11, 7, 67, 50, -22, 14, -6, -21, 0, -65, -64, 22, -14, 0, 2, -34, -19, 9, 37, 11, -13, 8, -97, 20, 2, -69, 30, -23, 5, -54, -16, -92, 11, -55, 63, 27, -42, -25, -22, 11, 25, -45, -68, -22, -37, -2, -2, 5, -22, -2, 36, 43, -44, 24, -98, -1, -1, -20, 6, 5, -4, -4, -56, -90, 27, -26, 10, -7, -9, -32, -21, -3, -12, -14, -48, -8, -5, 4, 10, 17, 33, 20, -35, -6, -33, -2, 78, -5, 17, 13, -22, 20, 12, -3, 0, -17, 16, -51, -21, 28, -16, -22, -22, 18, -16, -25, 0, -38, -26, -18, 11, 27, 20, -7, -48, -7, -2, 17, 57, -8, 11, 30, -28, -51, 6, 36, -2, 47, 26, -7, -98, 12, 7, 4, -12, -40, 3, -19, -3, 16, -12, 0, 7, 33, 35, -17, -34, -1, -17, 18, 30, -7, 0, 84, -7, 11, -8, 11, -22, 67, 13, -44, -48, 43, 5, -14, -7, -36, -15, -15, 10, -28, -24, -17, 25, -19, 15, 4, -10, 11, 3, 15, 6, 10, 20, 15, 8, -4, 14, 6, -28, 52, -7, 0, -1, 54, 5, -33, -8, -43, -17, -21, 8, 10, -22, 10, 12, -6, 17, 6, 0, 27, 0, 3, -14, 0, -15, -24, 5, 7, -11, -4, -7, -42, -18, 20, 4, 43, -10, 11, -6, -22, -1, 4, -12, 44, -13, 8, 13, -25, -12, 22, 51, 43, -17, 0, -79, -15, -17, -39, -5, -22, 0, 4, 0, -123, -3, -51, 55, 47, -13, 0, 25, 28, -8, 16, 10, 21, -1, -1, 3, 26, -14, -6, 0, 26, -51, 5, -71, -8, -8, -36, 26, 7, -12, 9, -34, -126, -5, 32, 46, -17, -2, -16, -22, 2, -13, 11, 18, 6, -3, -29, -12, -43, 2, -4, -43, 0, -19, 3, 108, -13, 4, 16, -40, 14, -16, 16, 33, 3, -19, 10, -133, 24, -18, 4, -7, 30, 15, -14, 14, 0, -2, -26, -12, 12, -5, 21, -37, -24, -1, 2, 66, 18, 15, 48, -38, -28, -12, 37, 69, 64, -30, 0, -80, 28, 25, 23, -19, -34, -7, 8, 23, 32, 22, -2, -23, -20, 18, 11, -29, 12, -6, 0, 25, -1, 7, 28, -6, -29, 39, 23, 11, 20, 21, -101, -25, 47, 7, 2, 3, -59, -30, -22, 14, -6, -10, 2, 0, -51, -6, 18, -14, -3, 42, -12, -27, -1, 7, 38, 14, -23, 31, 5, 11, 37, 17, -37, 26, 67, -3, 7, -32, -32, 13, 9, -41, 2, -22, 38, 21, -45, -27, 14, -18, 13, 17, -22, -21, -6, -6, 11, 8, -48, 0, 3, 9, 22, -1, -9, 14, 76, 10, 21, -33, -30, -1, -13, -43, 38, -12, 16, -7, -20, -16, 13, -11, 37, 11, -6, -76, 11, -14, -49, 36, -28, -12, 7, 30, -24, 18, 12, 58, 10, -10, 6, -20, 54, 13, 35, -8, 33, 0, 16, 14, 0, 27, 1, 53, 60, -37, -7, -54, 18, 7, -57, 9, 18, -13, -13, 10, -16, -17, -18, 13, -19, -22, 0, -24, 68, -14, 12, 3, 72, -5, -23, -22, 11, 14, 16, -36, -27, -37, -30, 68, -8, 11, -34, -17, 0, -17, -4, -31, -52, -14, 15, -91, 27, 43, 37, -23, -4, -18, -1, -26, -23, 27, 10, 16, 4, 7, -16, -9, 4, -25, 7, 58, -8, 3, 7, -26, -49, -29, 2, 67, -57, -2, 15, 2, -5, -7, 66, -9, 30, -6, 31, -13, 12, 43, -28, -41, 17, 16, -19, -21, 30, -18, -6, 18, 1, -4, 8, -14, -40, 0, 11, 84, -22, 6, -36, 3, -22, 2, 50, -52, 20, -49, -5, -6, 26, 18, 47, -28, -75, -23, -11, 25, 25, 16, -54, 30, -12, 21, 9, -10, -15, 20, 15, 17, 6, -6, 14, 3, 6, 13, -1, -42, 9, -43, 24, -18, 33, 0, 62, -9, -34, 3, 16, -30, 28, -2, -49, 1, 24, 10, 16, -10, -46, -8, 8, 20, 10, 13, 51, 17, 15, 23, 26, -46, 1, -28, -7, -50, 38, 29, 39, -5, -58, 13, -6, 5, 0, -8, 0, -19, -21, -19, -30, -13, -44, -21, 20, 83, -4, 12, 35, 35, -27, 13, 21, -35, 34, -37, 9, -34, 48, 27, 12, -7, -35, 27, -4, 8, -6, -43, 13, -54, 19, -22, -30, 23, -8, -24, 14, 41, -63, -17, -13, 13, -49, -28, 26, -10, 30, -7, -4, -41, 62, 33, -19, -16, 14, 8, -16, -18, 5, -22, 12, -7, 22, 25, -74, 21, -48, 20, 0, 6, -50, 8, 60, -55, 6, 34, 45, 4, 2, 16, -21, -24, 15, -2, -2, 21, 3, 15, 1, -24, 2, -6, -8, 10, -8, -5, -1, 3, -3, 0, -27, 62, -141, 4, -17, -27, -23, -30, 43, -25, 12, -6, -7, -51, 23, 35, 4, -24, 8, 37, -26, -43, 11, 18, -22, 2, 0, -8, -49, 0, -41, -37, -30, 48, -47, 0, 27, -36, -13, -4, 4, -40, 25, -44, 12, -43, 27, 25, 11, -26, -31, 6, -22, -20, 13, 35, -33, 30, 25, -10, 6, -3, -8, 8, -21, 37, -15, 26, 7, 6, 25, 28, 23, -47, -28, -13, 1, -37, 22, 27, 4, -8, -48, 1, -23, -23, 0, 40, -24, 15, 15, -2, 42, -2, -42, -8, -32, 7, -1, 0, 35, -21, -11, 41, -14, -36, -13, 2, 10, -21, 29, 28, 13, -13, -41, -2, -6, -24, -4, 8, -2, -33, 20, -12, -14, 9, -44, 9, -9, 30, -48, 28, -34, -12, 12, 31, 11, -56, -33, -14, -33, -5, 39, 17, 25, 4, -52, 5, -17, -66, -25, -27, 17, -42, -8, 10, 0, -21, -59, 0, -13, 16, -41, 21, 9, 27, 34, -15, 67, -17, 31, -11, -48, -37, -8, 14, -2, -9, 1, 35, 4, -28, -24, -32, -20, -24, 22, 21, -35, 76, 5, 24, 11, -4, -87, 28, 105, -16, -22, 2, 1, 12, 12, -27, 35, -51, 4, 32, -36, 22, 27, 39, 21, -16, 19, -34, -9, -43, 15, -12, -31, 23, -16, -3, 24, -1, -96, -26, 13, -4, -9, -10, 14, 10, 31, 0, -13, -57, -3, 27, -7, 22, -5, 5, 15, -4, 27, 36, 8, 11, 15, -11, -52, 44, -3, 7, 11, -23, -82, 18, -11, -22, 7, -17, 12, 27, 46, 7, 20, -5, 20, 10, -18, 24, -17, 5, -9, -39, 11, 42, 14, 0, 35, -12, 41, 34, -8, 15, 12, 10, -16, 20, -46, 2, 34, 18, 23, -1, -13, 13, 16, -14, 24, 28, 5, 19, -4, 2, 12, -13, -25, 18, 11, 21, 1, -21, -13, 6, -41, 16, 31, -2, -41, 19, -94, -18, -4, 42, -7, -2, -1, -1, 11, 9, 27, 7, 0, -5, -19, 10, -1, -40, -45, -8, 6, 82, -32, -3, -2, 1, -52, 24, 0, 10, -42, 15, -67, 1, 10, 24, -12, 5, -13, -36, -31, -42, -8, 19, -14, -7, -15, -4, -15, -30, -92, -28, 23, 30, 12, -2, -22, -32, -87, 26, 41, -2, 1, 11, 0, -31, 27, 18, -4, -33, -8, -6, -29, 3, -20, 6, -19, -2, -25, 3, 18, -20, -5, -17, 26, -101, 16, -9, -45, 33, 3, 23, -6, -25, -43, -13, 43, 13, -7, -17, 4, 18, 13, -19, -16, -109, 14, 4, -40, 6, 1, 36, 4, -31, 61, 4, 20, -97, 10, -5, -28, 41, -2, 28, 12, -12, -128, 38, 39, -8, 7, -9, 6, 5, 15, -14, -30, -69, 13, -8, -8, 3, 5, 20, 33, 4, 8, 29, -6, -14, -10, -5, -27, 30, 23, 30, 31, -4, 13, 36, -11, 4, 31, 0, 16, 14, 21, 2, -35, -42, -6, -13, -4, 34, 21, 6, 48, 2, 21, 4, 24, -28, 7, 40, -13, 8, 13, 71, 53, -24, -4, 16, -54, -17, 36, 2, 5, 1, -25, 8, -10, -72, -22, -17, 19, 22, -10, 17, 56, -4, 10, 12, 17, 28, -3, 18, 15, -4, 29, 34, 24, 12, -15, 44, -98, 8, 24, -7, 24, 12, -31, -1, 8, -29, 0, -11, 0, 15, 14, 18, 30, -45, -38, 2, 7, 47, -10, -3, 11, -7, 2, 43, 13, -22, 23, 44, 4, -58, -2, 21, -13, -4, -28, -3, -17, -34, -15, 3, -19, -13, -4, 5, 27, -122, -43, -4, 45, 78, 12, 5, 15, 21, -49, 10, -6, -1, -17, 33, -9, -59, 11, -6, -13, 19, -22, -4, -22, -13, -59, 26, -34, 0, -5, 7, 9,
    -- layer=2 filter=0 channel=1
    -21, -48, -21, 1, -2, 5, 3, 6, -2, 102, 15, 9, 50, 10, -13, -8, -33, -32, -1, 28, 5, 3, -1, 27, -35, 25, 29, -24, 21, 16, 59, -9, 17, 2, -14, -1, 7, 8, 5, -10, -14, 48, 6, -9, -58, 1, -7, 57, -33, 15, -21, -52, 37, -4, 2, 47, -23, 20, -1, -28, -15, 20, 21, -1, -30, 14, 4, -3, -11, 7, 3, 3, 29, 57, 3, -9, -1, -30, 10, -26, 33, -30, -22, -14, 21, -1, 0, 25, -19, -52, 8, -13, 1, 24, 11, 18, -10, 42, 1, -15, 7, 5, -2, -3, 10, 2, -15, -20, -5, -46, 18, -39, 14, -17, -3, 14, -34, -2, -1, 45, -17, 25, 3, -9, 6, -2, 18, -22, -5, -21, -8, 13, 37, 0, -14, 15, -13, 8, -12, 38, 0, 20, 1, -37, -25, -18, 7, 1, 0, -33, -16, 35, 18, 11, -6, -9, 13, -15, -19, -22, -20, -31, -15, 18, 18, 30, -11, -18, -6, 32, -5, 5, 32, 33, -10, 24, -28, -14, 15, -37, 15, 7, -7, -4, 17, 31, -4, -21, 3, 15, -33, -11, -5, 9, -46, 0, 11, -14, -1, -30, -8, 41, 18, -10, 9, 17, -9, 21, 15, -28, -15, -19, 28, 42, -2, 28, 23, 13, 23, -38, 0, 26, -13, -32, -28, -8, 0, 10, -15, 11, 6, -13, 13, -3, -5, -25, 24, -29, -1, 8, -19, -25, -53, 3, 21, -3, 9, -25, -38, 38, 3, -26, 13, 28, 21, -20, -15, 15, 8, 2, -20, -13, 0, 5, 10, 33, -10, 10, -11, -38, -13, 24, -36, -3, -35, -14, 6, 8, -2, -17, -15, 10, -2, -20, -23, -1, -48, -8, -28, 45, 3, -14, -13, -27, 8, -41, -20, -41, -21, -21, 31, -16, -3, -75, 36, -6, -10, 42, -14, -36, -8, 12, -8, 7, -18, 6, -12, 9, -32, 1, -36, 51, 1, -22, 7, -21, -16, -25, -4, -40, -8, -2, 10, -62, 20, -33, 6, -64, 25, 28, -27, -12, -40, 14, -25, -2, -11, 34, -39, -50, -39, 26, -50, 17, 11, -6, 41, -1, -7, -9, -21, -10, -42, 28, 0, -6, 15, -27, -13, 0, 50, 43, -31, -32, -2, 28, -2, -8, -20, 10, -35, -5, -53, 17, -25, -28, 12, 20, 22, -15, -13, -26, 0, -11, -26, 18, 14, -6, -4, -1, 5, 19, 31, -13, -21, -31, -16, -9, -5, 26, 1, 11, -2, 10, -29, 22, -15, -8, -17, 19, 20, 0, -14, 5, -26, 6, 21, -14, -7, 5, -17, -37, 0, -10, -42, -4, 0, 50, 9, 15, -21, 18, -1, -31, -18, 35, -17, -9, -8, -28, 34, 12, -33, 11, 9, 33, 10, -2, -31, -27, 25, -34, -12, -92, 8, -7, -25, -10, -9, 20, 2, -36, -14, 35, -6, -43, 1, 29, 15, 12, -18, -5, 40, 23, -24, -6, 8, 25, 10, -28, -17, -18, 30, 29, 25, -38, -9, 1, 12, 51, 0, 10, 6, -27, -33, 22, 5, 11, -15, 36, -18, 9, 3, -7, 39, -14, -82, -27, 14, -8, 16, -43, -18, 21, 47, 37, 58, 52, 7, 9, 17, 39, -20, -2, -10, -41, -54, 30, 3, 37, -21, 14, -31, 25, -29, 49, 46, -45, -30, -25, 31, -12, -7, -90, -9, -15, 88, 7, 54, -28, 35, -2, 32, 67, -57, 8, -29, -16, -19, -4, -6, 68, -64, -15, -42, 42, -50, 2, -4, -3, 35, -6, 0, 2, -10, -65, -12, 5, 33, -63, 33, -60, -5, -22, 33, 43, -21, -6, -32, -43, -65, 10, 12, 37, -29, -34, -27, 27, -1, 1, 10, 27, 23, -5, -4, 2, -19, -47, -25, -27, 39, -27, 13, -94, 17, 0, 30, 45, 17, 13, -8, -40, -29, 3, 16, 22, -16, -15, -7, 28, -1, -71, -9, 17, 37, 23, -39, 62, 25, -18, -11, -4, 28, -15, -40, -89, 1, -11, -6, -10, -13, 20, -13, -26, -1, 18, 32, -51, -19, 2, -15, -11, 41, 19, 23, -2, 37, 4, 10, 14, -16, -22, 0, -25, 33, -33, -17, -62, 35, -35, -64, -35, -11, -8, -22, -23, 14, 44, -15, -70, -16, 13, -42, -1, -2, -55, 0, -6, -44, -10, 28, 15, -7, -79, -20, -5, 12, 63, 11, -54, -15, -49, 16, -10, -48, 28, -48, -66, -57, 11, 38, 23, -23, 0, 43, 40, 0, -11, 32, -2, -11, 2, 34, 35, 35, -74, -11, 18, 46, 14, 6, -64, 21, -4, 20, 19, -82, 15, -26, -87, -93, 17, 23, 43, -24, -33, -1, 54, 21, 5, 28, -29, -16, 1, 26, 32, 30, -72, -21, -23, 83, -51, 36, -29, 81, -7, 17, 31, -88, 49, -18, -38, 3, 7, 53, 71, -65, -39, 14, 39, -2, -12, 44, 17, -40, 2, -9, 22, 45, -67, -56, 2, 76, -90, 32, -157, 87, 31, -35, 23, -60, 18, 1, -92, -64, -25, 9, 45, -80, -40, 23, 38, 3, -10, 40, -1, -24, 27, 3, 5, 17, -42, -37, -4, 13, -85, 19, -11, 34, -7, -19, 0, -39, -10, -36, -71, -61, 2, 5, 43, -49, -48, 23, 42, -16, -15, -11, -5, 2, 15, 6, 66, 29, 1, -18, -11, -1, -75, 7, -118, 37, -25, -41, -70, -8, -12, -28, -4, 9, 50, 37, -23, -10, -7, -6, 3, -7, -4, -21, -13, 40, -28, -56, 58, -23, 44, 7, -13, -12, -45, -29, -121, -30, -16, -92, -12, 2, 2, -26, -27, -18, 5, 18, -42, 0, -20, -22, -18, 20, -56, -9, -27, 35, -59, -8, 99, -34, -57, 13, 58, 71, -28, 23, -36, -21, -13, 21, -29, -35, 32, -59, -17, -18, 48, 63, 42, -63, -36, 36, 62, 42, -31, 29, 27, 17, 10, -10, 33, 21, -35, -14, 34, 10, 15, 4, 7, 51, -16, 0, -51, -29, -4, -35, -9, -67, 12, -4, 41, -33, -42, 18, 56, 36, 8, 18, 14, 29, 2, -11, 9, 8, -14, -22, 34, 68, -32, 18, -13, 24, 0, -13, -50, -27, 27, -25, -1, -5, 12, 22, 54, -47, -55, 49, 35, 7, 16, 23, -11, 19, 6, 3, 40, 8, -33, -2, 68, 34, -17, -14, -16, -4, 55, 1, -76, -62, 9, -57, 5, -1, 14, 32, 58, -51, -55, 33, 22, 25, 14, 29, 3, -37, -29, 13, -9, 5, -53, -28, -21, 4, -21, 21, 34, 56, -21, -23, -37, -40, 28, -37, -51, -81, -4, 9, 37, -54, -44, 57, 15, 26, 28, -9, -38, 12, -48, -16, -29, 6, -9, -36, -27, 16, -43, -11, -45, 47, -95, -24, -6, -2, 5, -40, -2, -45, 68, 24, -38, -37, -11, -23, 40, -10, 34, -26, 23, 89, -12, -7, -17, -76, -21, -9, 0, -11, 14, -36, -174, -99, 19, -42, -45, 2, -46, 3, -34, -2, -40, -5, -35, 3, -32, -63, 21, -1, 14, -9, -5, 17, 15, 28, 69, -40, 37, -1, 9, 47, -1, 37, -64, -7, 30, 52, 51, -40, -4, -18, -41, -7, 25, 37, 7, -46, -13, 36, 5, 24, -9, 17, -14, 19, -2, -20, 53, -25, 2, -26, -8, 55, 21, -9, -15, 41, 15, 30, 12, -5, -21, -63, 21, 12, 15, 8, 30, -57, -14, 62, 9, 13, 62, 13, -16, 13, -8, 26, -1, -42, 29, -22, 35, -19, -41, -24, -10, 9, 27, 11, -14, 7, -5, -43, 41, -87, -13, 2, -4, -23, -37, 39, -22, 5, 36, 21, -16, -14, 3, 14, 0, 5, 17, -4, 24, -3, 0, 11, -35, 15, -2, 6, 20, -16, 4, -27, 12, -74, 18, 9, -2, -36, -47, 53, -6, 26, 77, 40, -20, -26, 10, 34, 6, 24, -65, -12, 27, 27, -48, 19, -21, 58, -22, -24, 25, -23, 7, -31, -13, -92, 37, 34, -3, -20, -24, 58, -27, 6, 82, 12, -34, 13, -23, 12, -35, 16, 40, -18, -44, 0, -64, -13, -12, 20, -5, -46, -19, -19, 4, 9, 3, -112, 76, 6, -52, 21, -20, -1, -8, -26, 20, -27, 24, 128, 4, -13, -33, -35, -28, 23, 28, -63, -10, -34, -108, -120, 51, -18, 3, -26, -90, -10, -83, 38, -69, -41, -24, 29, -35, -65, -17, -35, -5, -39, 5, 56, 23, 8, 42, -11, -28, -2, -41, 34, 34, -13, -55, 8, 40, 12, 57, -11, -27, -11, -32, -3, 2, 2, -3, 4, -25, 41, -42, -29, 38, -28, -5, 75, 10, 1, 4, -44, -40, -18, 6, 19, 2, -1, -29, -20, 62, 50, 36, -23, -13, -26, -42, -31, -8, 24, -17, -11, -34, 65, -46, -28, 68, -3, -20, 14, 44, 18, 0, 15, -31, 1, -14, 30, 15, -13, -53, 16, 53, 39, 16, 6, -5, -29, -18, -51, 2, 11, -19, -1, -11, 21, -25, 8, 85, -18, 1, 30, 16, -22, 0, 7, -7, -15, -6, 12, 18, -1, 9, 31, 27, 7, 51, -16, 13, -31, -15, -111, 5, 8, -23, -9, -3, 9, -27, 0, 73, -14, 13, -96, 10, -7, -6, 40, -42, 16, -74, 0, -15, -3, 2, 53, 81, -84, 40, -40, 4, -20, -39, -116, 14, 17, -27, 29, -11, 18, -52, 46, 45, -24, 16, 14, 25, 24, -55, 13, 17, 25, -19, -5, -56, -8, -36, 12, 77, -83, 36, -18, -14, 1, 12, -87, 66, -46, -30, 59, -2, -22, -18,
    -- layer=2 filter=0 channel=2
    -37, 22, 22, 4, -18, -18, -9, -37, -12, 35, -14, -24, -77, 28, -11, -33, -52, -31, 0, -42, 20, 6, -2, -28, 14, -56, -15, 0, -15, 34, 4, -16, 26, 15, 13, -10, -5, -4, -53, 14, 3, -30, -38, 0, -21, -46, 6, -31, -25, -6, 0, -23, 29, 25, 12, -19, 13, 23, 13, -17, -29, 54, 5, -15, -22, 6, -15, -25, -66, 0, -16, -8, 22, -47, 2, -10, -15, -45, 4, 23, 34, 7, 2, 17, 2, 0, -2, 2, 0, -6, -3, -5, 2, 45, -6, -3, -14, 13, -30, -24, -23, -9, -16, -6, -21, -12, 17, -15, -47, -58, 4, -13, 21, 9, 20, 1, 5, 0, -6, -32, 3, -18, -23, -5, 16, 22, 13, -5, -56, -63, -4, -21, 17, -17, -5, 1, -5, -51, -4, -18, -21, -18, -17, 4, 7, 4, 1, 8, 7, -18, 6, -29, 23, 10, -13, -9, 15, 1, -39, -4, -64, -39, -6, -23, 42, -1, 16, -22, -54, -38, -16, 16, -9, -22, 8, -41, -39, 18, 46, 15, 8, -6, 0, -30, 33, 8, -19, -4, 7, 22, -7, -3, -21, -34, 19, 2, 39, -26, -4, -7, -10, -37, -4, 9, -25, -14, -20, -1, -1, -3, 0, -27, 9, -1, 15, 3, 21, -20, -27, -4, -8, 42, 17, -1, -60, 34, -6, -6, -18, -17, 5, -7, -20, -1, -23, 22, -37, 33, 26, 24, -53, 24, 25, -20, 20, -37, 0, 22, 41, -25, -39, -1, 14, 25, 0, 9, 14, 14, -14, -4, -7, -1, -22, -65, -31, -1, -10, 4, 0, -43, 26, 7, -11, 37, 23, 2, -6, 10, -15, -17, 0, 18, -13, 24, -7, 30, -25, 14, 33, -12, 11, 17, -14, 13, -6, -31, 31, -15, -7, 26, 15, -35, 15, 17, 28, 40, 15, 1, -11, 30, 8, -9, 36, 27, -12, -7, 27, -6, 18, -18, 12, -27, -7, 3, 4, -15, -20, -16, -5, -13, -37, -7, -8, -29, 40, 22, 21, 9, -3, -2, -11, -13, -11, 2, 64, 46, -19, -39, 8, 5, -36, -18, -30, 5, -16, 9, 24, 27, 16, -12, 3, -13, 13, 2, -19, 42, 42, 17, -15, 6, 22, -11, -28, 0, -22, -7, 52, 13, -23, -11, 2, 3, -26, -30, -3, 28, -9, -17, 15, 9, 12, -23, 1, 13, -8, 3, -29, 2, -9, -44, -6, 8, -6, -3, -2, 38, 13, 38, 22, -21, -38, 3, -4, 4, -15, 13, -25, 11, 7, 19, -16, -2, 5, -43, 14, -8, 9, 7, -31, 40, 11, -100, 2, 6, -37, -51, 11, -12, 24, 10, -2, -19, -21, 14, 13, 29, 21, 13, -45, -20, 8, 30, -41, 21, -1, -9, 12, -2, 15, 31, -30, 36, 17, -33, -31, 26, 42, -68, 7, -12, 9, 11, 27, -17, -60, 1, 10, 21, 7, 21, 10, 14, -10, -12, -34, 4, 24, -42, 10, 27, 15, 19, -6, -12, 21, -1, -19, 53, 11, -43, -7, 16, 0, -9, 27, -7, -34, 23, 27, -8, 27, 9, 40, 30, 26, 6, -32, 3, -21, -62, 33, -8, -9, 12, 21, -22, 45, -49, 18, 53, 17, -51, -40, -16, 11, 29, 58, 10, 12, 4, 23, -3, -3, -16, 8, 22, -34, 38, 13, -3, -50, 9, 21, -4, -43, 7, 29, -28, -1, -89, 13, 16, 17, -1, -31, -6, 19, 38, 91, 45, 3, -70, 3, 17, -17, 3, -30, -24, -16, 5, 20, 5, -9, -4, -13, -20, -20, -3, -13, 11, 26, -73, -11, 37, 39, -36, -23, -11, 1, 28, 79, 42, -13, -28, -4, 0, -18, 6, -50, 31, 12, -17, -15, 24, 16, -28, 19, -13, 17, 10, -9, 17, 28, -53, -11, 25, 21, -40, -25, -35, -3, 7, 13, -4, -19, 14, -1, -13, -26, 19, -25, 43, 10, 29, -42, 3, 9, -92, 23, 0, 0, 12, -42, 28, -21, -19, 7, 14, -21, -16, 25, 33, 18, 5, 6, -43, -70, 0, 9, 13, -12, -4, -22, -10, 1, 18, -19, 14, -7, 8, -17, 5, 27, 33, -32, 60, 12, -53, -44, 44, -7, -14, 35, -17, 5, -45, -20, 0, -42, -22, 12, 17, -12, -2, -17, 16, 0, -3, -41, 9, 10, -19, -2, 3, 22, 9, -1, 55, 15, -17, -61, 35, 24, -30, 1, -21, 15, -7, 5, -6, -65, 21, 43, 1, -42, 9, -1, 15, 15, -3, -29, 0, -23, -11, -7, -14, -32, -18, 41, -21, 16, -14, 35, 35, 24, 6, 6, 0, -7, 8, 84, -19, -12, -28, -7, -23, 10, -40, 0, 17, 36, 13, -9, 8, -48, 40, -2, -43, -38, -2, 29, -27, 27, -13, 49, 6, 30, 20, -22, 0, 20, 25, 96, 26, -6, -34, -18, -8, 0, 28, -25, -17, -11, 26, 42, -11, -27, 0, 13, -19, -21, -7, 3, -7, 37, -2, 54, 0, 18, -24, -26, -69, 15, 35, 65, 7, -10, -29, 8, -13, -10, 31, -45, 22, 1, -2, 6, 1, 29, -15, 13, -16, 16, 19, -60, 22, 53, -132, 40, 18, 18, -17, -20, -35, 17, 29, 54, 31, -33, 28, 22, -29, -9, 14, -23, -3, 10, 38, 10, 40, 2, -70, 48, -27, 11, -9, -57, 38, 34, 32, 24, 22, -22, -20, 1, 4, 29, -1, -9, -23, -78, 24, 15, 24, -15, 5, -28, 5, 22, 10, -23, 7, -5, -14, 6, -26, 32, 55, -48, 49, -2, -61, -22, 19, 23, 4, 19, -4, 17, -32, -45, -16, -60, 1, 2, 16, 15, 30, -22, 1, 20, -5, -7, -4, 12, -31, 4, -13, 9, 36, 15, 41, -14, -32, -21, 57, 23, 44, 0, -19, 18, -52, -14, 43, -61, 3, -10, -10, -39, 22, -3, -36, 12, 0, -9, -14, -4, 23, -20, -65, -7, -21, 72, 13, 0, -25, 26, 45, 30, 49, 14, -13, 0, -44, 19, 47, -24, -19, -32, -23, 8, -12, 19, -17, 9, 15, -29, 12, -25, -11, -11, -38, -14, -15, 30, 6, 49, 5, 44, 13, 11, -8, -2, -5, -3, -7, 48, 11, -5, -44, -2, 18, 1, 18, -44, 5, -15, -3, -6, 0, 14, -53, -15, -43, -32, -21, 8, -5, 26, -90, 71, 16, -26, 45, -22, 5, 7, 4, 26, 27, -30, -10, -8, -17, -25, 2, -47, 28, 11, -2, 12, 5, -16, -30, 12, -18, -3, -13, -1, -2, 29, 29, 38, 20, -8, 17, -18, -9, -6, 1, -10, 11, -53, 1, 12, 6, -50, 4, -17, 23, 24, 11, -33, 17, 29, -64, 19, -64, 7, -36, -60, 36, 23, -45, 19, 25, -33, -21, 9, -6, 6, 2, -22, -24, -48, 6, 10, 13, -14, -7, -61, -14, 7, 0, -81, 22, 30, -29, 34, 17, 25, 20, 2, 0, 4, -53, 18, 22, 21, 36, 24, -2, -9, -3, -28, -10, -3, 6, 18, 3, -13, 24, -41, -6, 8, 8, -44, 8, 29, -39, -1, -66, 5, 13, 9, 14, -2, 45, 1, 24, -10, 10, 17, -3, 0, -43, -61, -2, -64, 8, 9, -4, -33, 27, -14, -3, 21, -7, -10, 20, 13, -18, -13, -51, -15, 6, 32, 5, 14, -30, -25, 36, -7, 1, 1, 12, -14, -30, 8, 7, -43, 24, 10, 16, -27, 35, -4, -59, 23, 2, -45, -11, 0, 3, -23, -30, 1, 10, 11, -2, -3, 31, 18, -18, 1, 24, -22, 11, -1, -42, 37, -38, 5, -17, 26, 15, -9, 14, -31, -81, 9, 13, -15, 3, -2, 0, 2, -19, -20, 25, 17, 0, 42, -62, 23, -27, -4, 7, -6, -18, 1, -26, 27, -2, -21, -7, 29, -2, -31, 27, -22, -56, 16, 3, -7, 13, 9, -62, 14, -26, 1, -24, -24, 1, 4, -5, 16, 30, -4, -9, 3, -17, 3, -28, -15, 0, -16, 29, 30, -3, -20, 34, -63, 9, 14, 0, -12, 33, 25, -77, -20, -50, 26, 39, 1, 32, -6, -46, -25, 30, 7, -20, 8, -21, 7, -45, -42, -40, -6, 9, 12, -7, -17, 13, -9, 2, 15, -2, -66, 13, 5, 8, 26, 19, -18, 1, 49, 33, -3, 3, 39, -55, -33, -3, 31, 73, 7, 65, -33, 57, 22, -20, -44, 32, -15, -13, -4, 4, 5, -39, -55, -9, 11, -19, 21, -26, -4, 17, -9, 4, 16, 2, 31, -44, -3, -52, -7, 39, 0, 18, 38, 33, -39, -24, 14, 1, -8, -7, 23, -13, -20, -5, -36, -37, -20, 0, -9, 75, 0, 46, -44, 23, -18, -12, -16, -48, -43, -70, -14, 36, 17, 26, 33, -27, -37, -11, -20, -4, -65, 27, 43, -35, -41, -11, -19, -35, -16, -6, -20, 16, 13, 4, -55, 39, -6, 18, -28, -83, -62, -55, 11, 23, 10, 37, 64, 18, -15, -35, 9, -6, -44, 8, 16, -40, -11, -7, 15, -13, -12, -10, -39, 62, 32, 47, -30, 31, 13, -31, -49, -64, 8, -64, 20, 0, -2, 32, 74, 18, 5, -31, -11, 11, -28, 17, -43, -31, 6, -5, 45, 4, 1, 18, -41, 33, -2, 12, 10, 8, 6, 2, -36, -53, 11, -25, 7, 10, 0, 10, 73, -17, -9, -6, -15, -20, -21, 24, -95, -38, 2, 19, 18, -13, 3, 24, -36, -16, 9, 22, 29, 45, 1, 8, -38, -20, -16, 16, 23, -21, -13, -18, 14, -25, 0, 9, -32, -7, 8, 3,
    -- layer=2 filter=0 channel=3
    1, -15, -39, -5, 10, 4, -34, 25, -17, 17, -31, -39, 0, 28, -46, -36, -40, 30, 10, -13, 4, 16, -5, 20, 8, -3, 17, 7, -3, 1, -17, -54, 29, -44, -25, 9, 11, -8, -24, 3, 1, 30, 13, 9, -33, 38, -34, -50, -28, 16, 34, -13, 10, 0, -5, 28, 73, -16, -1, -28, -3, -19, -4, -41, 5, -5, 21, -6, 21, 17, -17, -16, -5, 3, 13, 0, 3, 38, -21, -69, -29, 37, 43, 13, 5, 7, 15, 1, 5, -8, 28, -25, 17, -9, -16, -29, 45, 16, 0, 3, -3, 3, -27, 7, 5, 12, 0, -2, 0, 19, 6, -59, -33, 13, 17, 0, 18, 19, 20, 11, 0, -10, 30, -19, 19, -5, -1, -18, 43, -3, -7, -32, -40, -11, 14, -10, 0, 20, -13, -54, -23, 41, 6, -33, -18, 19, 49, -1, 12, 10, 12, 24, 26, -36, -2, -4, 13, -7, 13, -14, 34, -18, -1, -5, -19, -20, -12, -2, 3, 17, -39, -42, -27, 12, -16, -69, 8, -15, -8, -5, 1, 48, 20, 30, -24, 23, -9, -39, 17, 25, -3, -11, 42, 60, -21, 2, -41, 9, -6, -3, -19, 15, -24, -29, -44, -5, -41, -36, 12, 0, -8, -23, -23, 15, -9, 44, 20, -10, 5, -9, -17, -3, -6, -31, 17, -11, -51, 2, 6, -13, 0, 44, -21, -3, -3, 5, -10, 26, 7, -39, -5, 4, 31, 29, -5, 16, -10, 2, 36, -4, 1, 21, -6, 1, 22, -3, 7, -8, -9, 3, 36, 23, 6, 9, 7, 28, 2, -14, -38, 18, 17, -17, 15, 11, 2, 23, 25, -13, -9, 25, 26, -4, -24, -13, 9, -19, 7, -52, 18, 25, -8, 0, 7, 5, -25, 5, -6, 2, -9, -7, -26, -21, 17, -65, -21, 7, 15, -26, 0, -23, 0, 22, 56, -3, 0, -22, 20, 16, 0, 6, 4, 13, -39, -4, -14, -8, 14, 16, 7, 24, 11, -22, -24, -34, 20, -7, -19, -32, 34, 2, -2, -9, 16, -3, -1, -18, 0, -3, 0, 24, -10, -33, 34, 8, -14, 6, 22, 33, 15, -11, 15, -1, -11, -61, -22, -7, 43, 17, -5, -28, 36, -34, 19, -17, 25, 4, -13, -3, -17, 7, 8, 8, -8, -34, 20, 10, -15, 7, -22, 32, 3, -32, -11, 30, 29, -8, -44, -29, -12, -71, -34, 9, 13, -7, -15, 2, 11, 18, 22, -9, -27, -3, 39, -1, 15, 1, 23, 19, -30, -6, -8, 18, 13, 31, 14, 12, 0, -26, -41, -10, 2, 10, -25, -2, 24, 7, -2, 9, -7, 12, 29, -1, 13, 10, -1, -2, -5, -6, 23, -11, -30, 6, 0, 6, 13, 0, -4, 3, 4, -28, -13, -5, 12, -71, -13, -7, 28, -34, 23, 5, 4, -8, 35, 12, 11, 29, 11, -14, 8, -7, -23, 24, -14, 0, -15, 0, 6, -11, 17, 5, 3, 8, -57, 13, -25, -45, -6, -33, -23, -43, -11, -15, -10, 21, 9, -4, -3, -26, -12, 10, 34, -39, -4, 18, 18, 8, 9, 15, -33, -17, 0, -9, -14, 7, -78, -21, -10, 6, -8, 38, -52, -22, -10, -29, 24, 17, 41, 0, -5, -61, 3, -2, 3, -53, -17, -1, -14, -24, 6, -8, 2, 22, -5, 24, 24, 2, -80, 14, 76, 16, 13, -41, -14, -30, 28, -21, 47, 12, 28, 19, -19, -59, 34, 16, 0, -42, -5, -3, 22, -5, 19, 27, 34, 12, 0, -3, 34, -6, -43, 35, 7, 11, -30, -14, 15, -39, 20, -42, 19, -4, 22, 53, -51, -48, 16, 15, -2, -4, 8, -19, 12, 1, -2, 6, -14, 19, 0, 0, -17, 3, -24, 17, -13, 16, -30, -11, 24, -8, 24, -4, 35, -20, 11, -13, -35, -24, 15, 3, -14, -15, -18, -4, -25, -2, -5, 19, -11, 18, 5, 10, 21, 12, -54, 53, 34, -3, -81, 8, 39, -41, -6, -10, 3, 23, 20, 9, -25, 25, -15, 0, -26, 18, 18, -1, 5, -23, -18, -24, -21, 20, 28, 0, -9, 22, 1, -24, 58, -19, 32, 4, 38, -51, 5, -3, 4, 28, 18, 0, 4, 4, 4, 7, 14, 25, -15, 22, 10, -26, -34, -7, -1, 0, 2, 14, -3, 18, -91, 15, 17, -9, -37, -7, -5, -42, 0, 9, 19, 16, 27, 0, -31, -15, 30, 8, -4, -11, -40, 6, -7, -5, 0, 0, -14, -12, 14, 0, 3, 28, -76, 4, 7, 14, 9, -34, -59, 2, -1, -30, 3, 21, 39, -18, -46, -48, 16, 1, -29, -7, -34, -29, 2, -2, 18, -14, 5, -19, 20, 6, 15, 37, -31, 12, 27, 44, -39, -40, -20, -32, 15, -39, 12, 17, 11, 15, -57, -67, 14, 15, -37, -28, -47, -18, 16, -6, 12, -7, 36, 7, -32, 12, 29, 26, -37, 36, 9, 23, -60, -38, 12, -76, 25, 5, 5, 22, 34, 0, -37, -37, 26, 14, -46, -13, -11, 25, -5, 0, 6, 21, -8, 14, 0, 8, -4, 9, -66, 29, 30, 63, -57, 19, -2, -15, -6, 4, 42, 2, 22, -33, -33, -23, 27, 16, -15, -17, -17, -1, 0, -4, 34, -27, -5, -4, -14, 1, 46, -1, -42, 18, 4, -57, -40, -23, 21, -43, 15, -21, 12, 31, 22, -35, 5, -3, 13, 15, 12, 20, 4, -20, -9, -11, -38, -9, 12, -47, 0, -35, -4, -8, -24, 25, 0, -18, 16, -31, -14, -19, -14, 0, -22, 14, 38, 14, -2, 16, 25, 13, 1, -9, -35, -36, -15, 0, -14, -7, 13, -16, -4, -30, -22, 34, -37, 17, -2, 8, -25, -4, -21, -32, -8, -44, 2, 5, 29, 0, -58, -13, -2, 20, -12, 9, -28, -34, -18, -3, -14, -15, 15, -12, 32, 6, 3, 28, -82, 23, -52, 38, 17, -34, -28, -31, 1, -14, 12, 10, 58, -25, -20, -28, 11, 8, -42, -11, -23, -49, -38, 5, -6, -18, 13, 12, -12, 11, 13, 74, -40, 47, -41, -81, 17, -51, -46, -29, -20, -14, 0, -11, 43, -26, -23, -21, 5, 4, -4, 2, -17, -12, -20, -4, -21, -9, 2, 4, -13, -11, 12, 27, -8, 15, -16, -17, -34, 5, -30, 8, 5, 13, 2, 9, 46, -9, -56, -1, 16, 20, -22, -3, -23, -9, -6, -4, -8, 14, 0, 7, 1, -9, -15, 19, -56, -8, -28, 14, -21, -15, -3, -17, 19, -29, 8, 11, 30, -40, -41, -26, -10, 17, -32, -28, -18, 0, -18, 30, -37, 25, 3, 14, 17, -3, 37, 11, -21, -2, -14, -53, -26, -5, -8, -22, 0, 17, 19, -14, 40, -16, -1, -9, 23, 11, -10, 16, -1, -10, 15, 0, -17, 3, 15, 18, 31, -11, 1, 9, -3, 36, 38, 22, 48, -4, 32, -28, -28, -7, 0, 0, 27, 10, -6, 38, -5, 13, 43, 36, -13, -55, -1, 10, -10, 0, -9, 15, 13, 2, -18, 17, -40, 25, -27, 59, 2, 9, -30, 0, 5, -10, -7, 16, 62, -4, -45, -1, 2, -1, -14, -13, -2, -72, -8, 19, -3, -9, 19, 17, -17, 5, 12, 44, -7, -7, 14, -39, -9, 1, 16, 4, 9, -12, 3, -4, 44, -5, -15, -30, -11, 17, 3, 12, -10, -24, -44, 0, -17, -8, 11, -12, 28, -22, 17, 3, -5, -3, 26, 26, 11, -17, 17, -10, 10, 11, 1, 8, 52, -8, -8, 20, -13, 16, -17, 4, -4, -5, -10, -12, -17, -4, 15, 6, 10, -16, 15, 1, 4, 18, 6, -8, 19, 30, -49, -23, -7, 9, 4, -16, 33, -14, -27, -11, 2, 2, -22, 10, -26, -28, -8, 16, -68, 3, 12, -47, -6, 6, -7, 40, -4, 1, -43, 34, -34, 18, -17, -12, 1, -15, 25, 10, 52, -1, -54, -26, 23, 4, -14, -7, 9, 6, -10, 12, -22, 5, 3, 12, 1, -8, 31, 0, -31, -7, -6, 46, 0, 8, 8, 0, -22, -6, 7, 14, 23, -4, -41, -1, -14, 15, 16, 26, 0, -11, 0, -10, -35, -24, -8, 36, 21, -6, 23, -3, 23, 44, 27, 37, 15, -5, 32, -17, -22, 46, -4, 55, 18, 42, 27, 35, -18, 8, 44, 25, 20, -39, -21, -16, 23, -3, -1, 19, -4, -13, -3, -6, -17, 27, -24, 2, 1, 11, -2, -16, -9, 8, 2, 18, 41, 28, -7, -1, -18, -4, -5, 10, 5, -67, -23, 39, 4, 21, 33, 7, 6, -26, 11, -39, -33, -7, -8, -18, 14, -13, 13, 0, 10, -22, 21, 10, 47, -9, -19, -5, -6, -10, -67, -48, -11, -29, -14, 1, -22, 14, 13, 22, -7, -12, -16, 3, -5, -26, 30, -5, 6, 0, 34, -16, -18, -4, 18, -30, -14, 12, -19, 5, -16, 14, -11, -5, 1, 17, -12, -18, -38, 14, -3, 24, 46, 4, -6, 25, -4, -18, 27, 61, 8, -7, 3, 8, 0, 19, 29, -42, 17, -3, -15, 8, -24, -11, -25, -16, 6, 33, -7, -8, -40, 18, 25, -35, 23, -14, 0, 22, 3, 6, -8, -14, 14, -3, -13, -28, -21, 24, -5, 11, 23, -24, 4, -3, -3, 4, 15, -7, 7, -3, -33, -14, -25, 1, 12, 35, 15, -12, 4, 0, 3, 17, -24, -5, 14, 19, 48, -21, -16, 23, -7, 48, 70, -28, 34, 37, -15, -24, 9, 23,
    -- layer=2 filter=0 channel=4
    -54, 10, 9, -6, 24, 12, -6, 30, -10, 11, -34, -22, 38, 30, -11, 31, -16, -58, -25, 23, -24, 11, 0, 29, -58, -48, 30, -28, -28, 3, -17, -7, -16, 10, 0, -18, 12, -2, 3, -9, -9, 4, -25, -15, 15, 25, 18, -19, -48, -20, 5, 40, 7, -5, 10, 21, -34, -41, -4, -4, 5, -8, -38, 6, -17, -12, 0, -35, -3, -28, 1, -17, -49, 59, -9, -18, -15, 26, -17, -20, -44, -14, -47, -12, 20, -15, -1, 1, -36, -38, -40, 13, 2, 10, -52, 13, 6, -29, 23, -9, 21, -13, -13, -36, 0, 39, -24, 22, -31, -2, 3, 26, -47, -22, -16, -27, 2, -6, 3, 29, -58, -44, -13, 19, 7, -4, -47, 24, 3, 61, 23, -25, -47, 11, -10, -17, -21, 34, -25, 25, 1, 23, 12, -6, -17, -18, -10, 9, 0, 13, 14, 16, -72, -78, -8, 17, 3, 11, -46, 0, 17, 64, 22, -30, -44, -19, -10, -50, -14, 31, -21, 1, 9, -23, -35, 37, 20, -21, -44, 4, 13, 14, -1, -44, -27, -49, -16, 15, -10, 1, -58, -5, 4, 40, 6, -45, 5, -22, -36, 18, -42, 70, 11, -13, 52, -20, -32, -66, 0, -12, -42, 47, 21, 33, 10, -34, 10, -27, 6, -21, -30, 2, -9, -5, 8, -1, -4, -31, 42, 20, -6, 20, 21, -10, 1, 1, 14, 69, -28, -63, -5, -43, 47, 29, 3, -23, -1, 16, -21, -49, 15, -10, -2, -14, -12, -9, -26, -17, -15, -6, 29, 18, 16, 13, -10, -3, 0, 34, -2, 21, -17, -53, -34, -33, -9, -23, -1, -11, 5, 5, -36, -65, -6, -3, 18, -4, -5, 9, -2, -34, 2, 9, 29, -33, -5, -35, -15, 12, 48, 43, -17, -4, 10, -46, -35, -34, -43, 4, 23, 6, 13, -16, -69, -60, 0, 20, 30, 0, -16, 18, -10, 7, 25, 3, -10, -14, -18, -68, 5, 35, 48, 3, -39, -33, -2, -50, -18, 9, -15, -39, 9, -4, 18, 13, -86, -39, -9, 10, 37, -5, 8, 22, 17, -5, 29, -20, -23, -30, -26, -104, -16, 40, 43, 41, -19, -51, -61, -22, -23, 19, -54, -30, 10, 1, 17, -11, -58, -73, -35, 13, 20, -9, 12, 17, 16, 36, 9, -14, -86, 1, -31, -22, 10, 16, 23, 27, -17, -27, 19, 21, 24, -7, -1, -21, 18, 51, 15, -23, -70, -33, -17, 10, 4, -16, -6, 26, 57, 34, -14, -5, -82, -12, -10, -15, -13, 31, 4, 9, 10, -12, 10, 28, 29, -24, 9, 41, -6, 24, -14, -3, -2, -45, -19, -12, -29, 2, -35, -6, -30, 13, 17, 10, 20, 30, 26, 0, 16, -9, -8, 0, -15, 29, 7, 68, -45, -5, 56, 32, -13, -19, 8, -13, -3, -58, -13, 25, 9, -6, -33, -12, -20, -17, 2, 49, 56, 1, 13, 15, -2, -24, -14, 12, -14, -34, 2, 22, -9, -14, 17, 27, 10, -3, 6, -23, -29, -24, -2, 21, -14, 13, -12, 8, -32, -11, 27, 17, 43, 5, 6, -14, 2, 9, 19, 26, -32, -28, -10, -75, -44, 21, 14, -22, -9, -16, 0, -40, -34, -14, 12, 1, -7, -2, 18, -8, -42, -14, 46, 8, -14, -18, 9, -54, 0, -26, 21, -8, -2, -13, -23, 19, -20, 41, 16, 5, 21, -2, 6, -27, -10, -3, -3, -23, 0, 28, 28, 16, -1, 12, 35, 2, -54, -31, 0, -65, 35, -8, 39, -22, 26, -11, -14, -13, 5, 10, -28, 25, -2, 7, 20, -27, -81, -29, 11, 15, 2, 34, 9, 0, 26, 32, 26, 5, -31, -14, 18, 7, 21, -20, 19, -20, -13, -14, -7, 20, 3, 0, -45, 56, -6, 43, 3, -28, -35, -12, -22, 1, 7, 8, -6, -8, 5, 11, 30, -20, -74, -1, 3, -21, -14, -17, 4, -16, 12, 26, 3, -15, 47, 8, 3, 21, -9, 0, 2, -18, -50, -22, -50, 24, 4, -23, -11, -28, -41, -25, 15, -30, -1, -11, 43, -38, 20, -25, 31, 4, -15, 21, 25, -12, 30, -27, 58, 3, -7, -16, -2, -8, -3, -65, -31, 58, 17, -15, -1, 5, 22, -5, -12, 21, 34, 39, 26, 39, 35, 12, -10, -11, -23, 3, 17, -24, 8, 16, 31, -23, -2, -24, 21, -52, 17, -25, 10, 7, -25, 8, 0, -10, -5, -24, -7, 27, 30, -7, 9, 53, 33, 25, 31, -44, -14, -2, 4, -51, -8, 39, 10, -1, 29, 15, 9, -25, 14, -6, 28, -43, -15, 25, -12, -10, 23, 21, -27, 16, 2, -16, -8, 60, -7, -5, -40, -45, -16, -5, -16, -99, 2, 6, -83, -21, 13, -29, -1, -35, 15, 27, 17, -147, -17, 34, -23, -25, 24, 4, -6, 16, -2, -7, -19, 5, 0, -1, -6, -53, 15, -11, 5, -58, -17, 11, -21, -12, 0, -4, 5, -29, -5, -7, 25, -50, 10, 33, -1, 16, -4, -4, -12, 2, -21, 0, 47, 37, 42, -6, -1, -22, 13, 33, 23, 17, 37, 22, 14, 17, 21, 0, -5, -9, -7, -9, -1, 0, -9, 38, -21, -8, 3, -15, 26, -11, -89, 7, 23, -35, 38, -17, -4, -16, 20, 76, 25, -19, 49, 29, 43, 12, -4, -28, 23, -4, -5, -82, -20, 43, 1, -11, -23, 12, -43, 37, -4, -6, -25, 13, 12, 28, -8, 1, 15, -12, 21, -9, 2, -13, 27, -2, 36, -12, -6, -17, 16, -18, -10, -56, -34, 22, 8, -6, -5, 12, 18, 17, 2, 18, -15, 14, 19, -19, 18, 0, 47, -48, -22, 8, 0, -40, 32, 1, 11, -33, 4, -6, 34, -26, -4, -62, -3, 12, 20, 34, -13, -5, 22, -10, -28, 12, -7, -14, -7, 50, 9, 18, 34, -35, -14, 3, 32, -46, -11, 22, -25, -6, 25, -23, -2, -1, 27, -56, 26, -14, 30, 28, 3, -50, 30, -8, -33, -9, 21, -12, -36, 29, 12, 47, 19, -36, -48, 10, -12, -2, -21, 38, -90, -59, 28, -25, 7, 18, 80, -10, 19, -72, 14, 22, -60, -87, 19, 1, -40, 7, -7, -26, -27, 21, 20, 51, 20, -37, -20, 3, 26, -21, 3, 22, -46, -73, 26, -11, 6, 16, 42, -21, 20, -63, 19, 6, -51, -16, -4, -14, -24, 8, -41, 3, -8, 27, 24, 12, 25, -10, -10, -37, 37, -49, 7, 16, -25, -28, 14, -4, 4, -25, -47, -17, -2, -20, 30, 4, 9, 6, 1, -47, 6, 2, -19, 6, -3, -13, -26, 38, 16, 49, -8, 3, -10, 8, -46, 41, 26, -31, 6, -16, 1, -6, -9, -15, -24, 34, -10, 7, -22, 16, 32, -10, 13, -16, -57, 6, 13, 37, -4, 0, 33, -12, 44, -27, -30, -16, 35, -33, 16, 6, 24, -2, 3, -27, -21, -43, -16, 30, -8, 18, 17, -9, 64, 27, 8, 7, -59, -1, 0, 17, 10, 33, 20, -26, -14, 5, -27, 17, 37, -7, 2, -31, 40, 11, 23, -7, -43, -66, -20, 29, -5, 23, 20, -7, 25, 5, -18, 4, -42, 34, 28, 28, 7, 58, 61, -2, -8, 6, -8, 24, 16, -2, -14, -46, -1, 1, 0, -3, 6, -72, -22, 65, 24, 8, -13, 0, 70, -15, -19, -12, -9, 20, 1, 14, -14, 69, 43, -37, -28, 17, 4, -30, -41, -2, -30, -104, 14, -20, 28, 9, 5, -49, -12, 6, 35, -5, -31, -7, 26, -15, -23, -23, -18, 9, -12, -14, 21, 71, 44, -5, -50, 32, 13, -78, 6, 18, -18, -60, 4, -5, 0, 31, 8, -24, -26, 34, 13, 0, -38, 11, 23, -60, -19, 13, -5, 4, 10, 60, -21, 40, 33, 39, 0, 27, -7, -36, -11, -10, -40, -25, 19, 35, 0, -9, -16, -51, -11, 17, 2, -8, -15, 8, -24, -65, 11, 12, 49, 4, -11, 8, 0, 54, -8, 20, -1, 0, -11, -75, -50, -4, -7, -25, 13, -7, 1, -29, 8, -108, 5, 13, -6, 0, 22, -16, 11, 51, 38, 9, -39, -7, -1, 10, -19, -1, -4, -56, 31, -23, 9, -67, 79, -48, 4, 29, 29, 5, 10, -13, -6, -68, 28, -1, -4, 34, 13, -1, 3, 20, 45, 35, -67, -5, -30, 22, -16, 30, -1, -15, -9, -33, -21, -7, -22, -31, 12, -5, 16, 11, 37, -12, -2, -61, -49, 25, -20, 30, -2, -46, 20, -29, 31, 2, -84, -8, -25, -11, -43, 55, 10, -30, 2, 15, 0, -9, -3, -22, 11, -23, 36, -5, 26, 14, 8, -53, -32, 22, 10, 42, -16, 10, 26, -1, 13, 4, -22, 24, -42, -27, -53, 80, -2, -2, -13, 17, -20, -5, -31, -1, -30, -35, 41, -13, 12, -9, -30, -54, -21, 7, 36, 4, 20, -24, 16, -48, 21, 21, -11, -19, -23, -32, -30, 40, 17, -6, -25, -8, -11, 20, -17, 4, -31, -21, 17, -6, 27, 59, -30, -72, -47, 31, -4, 1, -10, -15, 7, -48, 31, 13, -5, -1, -3, 14, -41, 27, 5, -4, -19, -27, 14, -116, -24, -7, -2, -31, 34, -18, 12, -6, -62, -22, 15, 0, 0, 18, -5, -39, 23, -33, 26, 32, 8, -12, -75, -16, -39, 32, 0, 51, -10, 47, 31, -30, 4, -17, 14, -7, 31, 13, 15, -59, -54, -42, 43, -17, -29, 8, 36, -23,
    -- layer=2 filter=0 channel=5
    74, 30, 16, -50, -61, -71, -66, 4, -50, 15, 0, 11, -37, -46, -28, -16, 19, 57, 35, -52, 10, 23, 31, 10, 39, -33, -21, -19, 24, 7, -27, -12, 30, 26, 8, -18, -71, -22, -33, 28, -5, -50, -14, 19, 0, -43, -42, -12, 46, 1, 4, 0, -18, 34, 6, 0, 9, 30, 40, -35, -1, -10, 11, -11, 39, 22, -2, 14, -40, 6, -2, -15, 32, 0, -18, -29, -9, 1, -58, -96, 39, -3, -23, 6, 5, 37, 2, 5, 26, 49, 2, -4, -15, -6, 10, -6, -14, 9, 11, 46, -14, 42, 30, 33, 6, -57, -2, -38, 57, -39, -27, -84, 23, 34, 14, 8, 8, 15, 18, -1, 40, 41, 4, -1, 7, -13, -21, 15, -32, -9, -4, 60, -11, 51, 7, 40, -21, -23, 9, -8, -22, -18, 1, -5, -36, 7, 4, -34, 13, -1, -9, -7, 57, -6, 6, -19, -8, 0, 14, -18, 10, 12, -6, 6, 52, 33, 16, 59, -19, -16, 4, 0, 10, -19, 10, -8, -14, 29, 56, -11, 3, -24, -10, 3, 63, 11, 41, -12, -31, -37, 13, -49, 40, -48, 30, -6, 12, -2, -7, 50, -37, -25, 0, -45, 13, 38, 19, -46, -1, 55, 47, -18, 17, -16, 4, -8, 50, -11, 5, 3, -4, -18, 17, -37, 53, 31, 0, 2, -53, -24, -26, -50, -30, -13, -21, 0, -52, -35, -2, -12, 1, 22, 23, -43, -37, 4, -14, 18, 18, 7, 25, -11, 0, -38, -33, -5, 15, 34, -21, -19, -38, -35, -24, -24, -11, 1, -5, -29, 13, 20, -36, -88, 32, -37, -19, -34, -20, 20, -3, 28, 35, 20, 0, -24, -19, 18, -19, 5, -6, 23, -12, 14, -31, 30, -2, 31, 13, 7, 5, -13, 19, 27, -85, -107, 44, 2, -3, -26, -7, 2, 5, 30, 8, 41, 3, -28, -42, 52, -4, -3, -6, 25, 4, -3, -16, 30, 20, 18, 32, -7, 16, -16, 18, 53, -91, 8, 37, -9, -33, -13, 3, 18, -12, 18, 21, 13, 19, -18, -42, 16, -5, 12, -29, -16, 21, 26, 31, 25, 27, 7, 19, 0, 27, 22, 24, 4, -44, 19, 26, -14, 7, -5, 9, 16, -16, 3, 45, -3, 23, 13, -11, 27, 36, -21, -10, -18, 1, 4, 35, 31, 33, 49, 18, -6, 0, -3, 13, 55, -16, -37, -39, 3, 0, -36, -16, 6, -2, 13, 25, 9, 11, -21, -18, -17, -2, -60, 6, -22, 1, -8, 14, -11, -6, 11, 4, 0, 4, 28, -4, -6, -10, -45, -56, 9, 48, -52, -9, -17, 0, 18, 44, -1, 7, 8, 26, -10, -34, -11, 24, 0, 29, -16, -52, -44, -6, -45, -15, 1, 1, 4, -62, 3, 44, -48, -10, 52, -8, -73, -28, -22, 9, -9, 35, 18, 1, -7, 8, 4, 35, 24, 9, 19, 10, -35, -45, -24, 0, -21, -5, 15, 8, -42, -29, -4, -40, -41, -26, 13, -49, -62, 13, -3, 7, 37, 16, -25, -27, -16, -6, 1, -11, -3, 19, 21, -49, -50, 17, -1, -6, -18, -6, 30, 2, -62, 7, 16, -61, 14, 6, -40, -21, 5, 9, 17, -8, 38, 2, 17, -22, -19, -19, 28, -30, 20, -3, 42, -62, -37, 41, 0, -6, -26, -42, 40, -19, -36, 23, 14, -95, 29, -22, -45, -49, 16, 14, 14, -17, 39, 8, -37, 5, -47, -6, -3, -11, -44, 20, -2, -27, -23, 12, 25, -6, 11, 14, 19, -14, -7, -8, 61, -67, 8, -9, -74, -45, -14, -11, -4, 3, 30, -12, 30, -14, -15, -48, 0, 17, -48, 26, -23, -24, 6, 45, 1, 11, -42, -3, 29, 0, 10, -24, 17, -19, -37, -82, -2, -17, -11, 18, -34, 0, 31, 32, -1, -12, -40, -3, 31, -20, -24, 57, -44, -3, 14, 24, 0, -5, -30, 5, -3, -22, -12, -16, -14, 28, -76, 27, 40, 7, -15, 8, -24, 5, 20, 33, 15, -3, 2, 26, 28, -17, 1, 37, -24, 11, 5, -18, -36, 8, 2, -5, 6, -5, -4, -83, -8, -7, -7, -26, 53, 0, -41, -19, -9, -15, -12, 35, 28, -36, -8, 22, -15, 37, -6, 29, -6, -18, 10, -23, 6, -31, 2, 13, 16, -6, -4, -11, 37, 0, -72, -22, 0, -50, -35, -32, 1, -3, 4, 47, 12, -32, -26, 6, -14, -40, -16, 4, 14, -33, -16, 5, 35, -20, -29, 8, 42, 9, -44, -27, 34, -57, -36, -40, 17, -70, -11, 4, -7, 6, 23, 9, 13, -47, -60, 12, 30, -36, -20, 0, 13, -41, -41, 39, 10, 1, -39, 28, 37, -3, 5, 32, 32, -81, 27, -33, -1, -35, 10, 11, -7, -19, 57, 23, 12, -8, -54, 20, -12, -49, -25, 17, 6, -34, -25, 70, 24, 13, 9, 3, 18, 1, -26, 17, 16, -41, 1, -37, -7, 0, 34, 0, 9, -3, 9, 31, -10, -11, -17, 14, 13, -48, -4, 38, -36, -13, 6, 29, 18, 14, 14, 8, 39, 44, -16, -66, 37, -44, -31, -41, -48, -22, -71, 2, -24, 4, 20, 14, -15, -50, -20, 1, 19, -49, -16, 12, 0, 7, -12, 7, -4, 16, 41, -8, 30, 4, 11, -82, -10, 38, -3, -22, 31, 67, -42, 11, -29, 8, 10, 33, -22, -15, 12, 26, 24, -31, 18, -13, -21, 17, 24, -38, -27, -6, 19, 6, -20, 0, 13, -33, -24, -3, 6, 10, 37, 31, -72, -14, -45, -9, 15, 24, 3, -42, 12, 6, 14, 8, 15, -7, 6, -6, 5, -11, 6, 11, 18, 12, 14, 10, -2, -75, 28, -34, -5, -3, 0, -10, -54, -2, -17, -5, 40, 39, -21, -31, -26, 17, -13, -43, -9, -25, 18, -47, -3, -43, 33, -19, 19, 10, 41, 16, -10, -32, 2, -42, -7, -53, 2, -21, -8, 13, -28, 15, 12, 21, -43, -30, -10, 29, 8, -48, -7, -14, -12, -46, -5, 13, 22, 17, -30, 36, 4, 23, -4, 10, 31, 3, 1, -5, -21, -42, 24, -6, -31, 5, -41, -5, -19, -36, -16, 30, 1, -62, -31, 9, -2, -37, -13, 9, 27, 15, 3, 50, 18, 16, 3, -6, 31, -18, -2, 14, -43, -25, -36, -3, -18, 21, 19, 13, -14, -43, -36, 7, 19, -50, -13, 6, -22, -12, 19, 13, 41, 33, 27, 5, 24, -1, -4, -15, 44, -38, -65, -34, 9, 2, -38, 29, -40, -2, 5, 70, -20, -55, -34, 25, 16, -16, 8, 20, 1, 5, 1, 24, 1, 0, 14, 3, 7, 0, -6, -33, -9, 26, -127, -19, 40, 67, -27, -17, -35, -9, 22, 46, -17, -29, 48, 13, -28, -16, 19, 26, 21, 18, -3, -12, -20, -11, -9, -23, -5, -23, 7, -42, -15, 14, -55, 74, 27, 9, -92, -29, 2, 0, 16, 31, 30, -40, 8, -3, -15, 13, -5, 5, -27, -13, -7, -25, 3, -17, 41, -4, 1, 4, 22, -52, 0, -16, -66, -14, -43, 0, -29, -29, -14, 24, 30, 32, 38, -36, -30, 4, -13, -36, 8, 1, -25, -35, -8, 3, 8, -6, 8, -3, 15, -29, 37, -42, 38, -47, 66, -35, -44, -46, -36, 20, -31, -17, 39, 23, 3, -45, -16, -13, 0, -16, 26, 6, -14, -21, 4, 26, 22, -1, 12, 12, 2, -31, 12, 23, -9, -22, 30, -4, -55, -25, -5, -2, -24, -18, 8, 14, 3, -41, -9, 10, -16, -12, -12, 5, -14, -31, -14, -23, -3, -7, 10, 0, -6, -1, -9, -4, -31, -73, 15, -15, -13, -32, 1, -2, -16, -13, 0, 41, -11, -9, -23, 10, -20, -26, -28, 24, -66, -19, 4, -6, 4, -9, 39, 17, 13, -38, 10, -52, 9, -14, -24, 0, -13, 3, -71, 7, -13, 6, 15, 52, 16, -31, -45, -20, 40, -32, -31, -14, -48, 18, 0, 14, 9, 34, 28, -12, -30, 4, 0, -50, -7, 34, -50, -24, -7, 39, -30, -5, -2, 4, -1, 57, -8, -13, 18, -8, -32, 13, -18, 48, -39, 21, 5, -55, -55, -3, -13, -28, -16, 4, 26, -10, -33, 71, -58, 21, 41, 20, -25, -45, 3, -8, 0, 23, -7, -7, 15, 31, 10, 54, 27, 42, -56, 19, 17, -31, 11, -8, 26, 12, -9, 0, 6, -36, 43, -7, -8, 0, 6, 4, -59, 6, 12, -29, 15, 11, 6, -24, 32, -1, 17, -15, -7, 30, -59, -12, 20, -14, 7, 8, 29, 30, 36, 0, 6, -9, -30, 34, -34, -27, 34, -7, -50, 0, 15, 9, 0, 4, -24, -11, -9, 4, 1, 10, 0, 18, -31, 22, 28, 5, -14, -7, 30, 36, -4, -3, 13, -27, -6, 23, -37, 21, -20, 27, -21, 2, -7, -9, 24, 51, 0, 6, -17, -11, -6, -26, -5, 9, -33, 5, 30, -17, -2, -23, 30, 20, 17, -23, -2, -5, -3, -1, -17, 9, -21, 52, -37, 2, 6, -11, 5, 26, -16, -26, 18, -2, -15, -39, -1, 40, -79, 17, -1, 38, -20, -26, 35, -9, 48, -10, 10, -67, -1, 24, -23, 17, 3, 34, -58, 3, -23, 17, 30, 56, -3, -37, 26, -13, -5, -56, 3, 5, -58, 10, 23, -7, -9, 22, 43, 0, -27, 0, -14, -36, -19, 40, -26, -25, -17, 62, -38, -15, -24, -2, 3, 55, 5, -19, 24, 15, 8, 12, 46,
    -- layer=2 filter=0 channel=6
    14, -16, 25, 6, -62, -4, -60, -62, 16, -27, -40, -45, -33, -5, -53, -33, -14, -19, -16, -26, 35, 23, 29, -18, -27, -17, -18, -28, 19, -5, 8, -78, 7, 54, 20, -11, 24, -17, -28, -23, -2, 41, -9, -40, -10, -14, -10, -21, -38, -2, -2, 12, 28, 58, 28, 11, -79, -25, 3, -13, 12, -1, 18, -74, 4, 6, 2, -4, 6, -2, -27, 0, 18, -3, -14, -21, -25, -1, 17, 66, -21, 9, 21, 4, -12, -2, 13, -1, -39, -7, 8, 11, 20, -7, -3, -58, 17, -53, 14, 5, -50, -10, -17, 2, -9, -7, -32, -22, 8, 69, -6, 54, -46, -1, 30, 10, 3, -6, 12, 15, -21, -20, 25, 12, 28, 16, 7, -35, 32, -28, 6, 4, -15, -5, 0, -5, 30, -16, 1, -47, 18, 30, 23, 4, 5, -37, -4, -2, 30, 65, 4, 29, -35, 17, 8, -4, 6, 27, 24, -40, 3, -68, 18, 1, 21, -37, -9, 7, 0, 9, 14, -26, 8, 33, -42, 8, -73, -21, 10, 19, 17, -10, -5, -26, -26, 7, 5, 19, 17, 30, 20, -24, -32, -97, 18, -9, 58, -1, -45, -41, -6, 21, -23, -62, -8, -18, -44, 83, -58, 21, 9, -24, 21, -10, 12, -23, 6, 3, 27, 9, 27, -6, 19, -48, 31, 10, 5, 22, -26, 15, -17, -50, 33, 9, 14, -12, -7, -13, 19, 8, -15, 9, -9, -12, 12, 26, 18, -1, 3, 18, 4, 9, 20, -3, -17, -24, 18, 14, 7, -36, -21, -22, 9, -13, -7, -2, 8, 12, -10, -12, 18, -17, -20, -24, -15, 5, 13, 11, 0, 7, -18, 20, 21, 10, -7, 8, -25, 11, 8, 0, 6, 4, -32, -9, -7, -30, -18, -32, -71, 5, 12, -8, -5, -20, -19, -75, -28, -27, 27, 30, 15, -42, -104, -10, 22, 23, 1, 2, -23, -23, -1, -59, 15, 64, -34, -16, 1, -9, -22, -93, -74, -29, -16, 0, 37, -93, -16, -11, 23, 2, -3, 43, 26, -51, -30, 14, 13, -15, 10, 31, 40, -15, 7, -93, 25, 28, 0, -52, -35, 72, -59, -58, -50, -50, 13, -30, 34, -24, -66, -44, -16, 20, 31, -2, 14, -98, -51, -8, 19, -33, -4, 41, -8, -5, -34, -89, 14, 20, 38, -28, -2, -33, -51, -9, -7, -57, 15, -5, -21, -4, -35, -35, -8, 0, 26, -12, 5, -38, 14, 26, 15, -3, 27, 10, 2, 10, -30, -34, 3, -10, 62, -19, -7, 16, -4, -22, 24, 3, 30, 16, -74, -8, -89, 10, 3, -31, 2, 2, 0, -20, -13, 26, -9, 49, 18, -25, -10, 7, 9, -32, -15, -14, -6, 32, 13, -58, 33, -52, 18, -27, -45, -18, -14, -48, -34, 3, -15, -40, 10, 21, -8, -1, -8, 8, 36, 14, 46, -9, -54, -44, -23, -33, 18, -13, 3, -3, -11, -31, 24, -12, -21, -16, 11, -25, 48, 2, -26, -58, -15, -17, -22, 3, -6, 4, 18, 15, 9, 1, 17, 6, -45, 58, 8, -26, 19, 14, -7, -13, 17, 30, -55, -20, -80, 6, -20, -83, 33, -30, -49, -70, 0, 0, 28, 13, 30, -18, -55, 28, 2, -23, -12, 27, 5, 63, -1, -43, 72, 19, -61, -17, -2, 34, -45, -90, -88, 2, -38, -116, -4, -176, -79, 12, 43, -15, 16, -1, 31, -50, -44, -8, 2, 3, 8, 32, 20, -48, -19, -40, 30, 37, -36, 23, -19, 59, -55, -13, -66, -9, -19, -64, 8, -3, -92, 14, -14, 3, 27, -8, 26, -47, 11, 5, 14, -18, 7, 43, 17, -1, -37, 14, -3, -18, 7, -30, -30, 24, -42, 10, -5, -8, 6, -14, -73, -10, -76, -14, 0, -15, 23, 3, -4, 18, 27, 52, 35, -21, -5, 19, -38, 28, 1, 17, -30, -21, 34, -13, 46, -36, 17, -11, 30, -8, 4, -12, -49, -49, -13, -44, 39, -6, -15, -6, -8, 28, -26, 28, 11, 42, 23, 0, -29, 7, 26, 10, -29, -5, 0, 15, 41, -77, 33, -21, 18, -31, -32, -1, 28, -49, -48, -19, 7, -38, -20, 20, -14, -16, 12, 27, 13, 24, 7, -40, -22, -8, -46, -61, 8, -15, 81, 5, 3, -53, -15, 0, -8, -24, -52, -32, -39, -100, -59, -34, -8, 47, 13, -6, 9, 25, 25, 37, 8, 15, 5, 8, -58, 48, -62, -39, 70, -20, 31, -43, -21, -18, -55, -47, -56, 6, -56, -46, -27, -64, -76, -12, 18, -37, 7, -5, 32, 0, 3, 18, -29, 1, 20, 17, -34, 24, -108, -67, 98, 34, -64, -16, -24, -32, -23, -46, -42, -14, -95, -92, 44, -218, -77, 55, 18, -62, 18, -17, 64, -77, -41, -32, -30, -6, 42, 30, -20, -9, -39, 25, 83, 23, -39, 5, -27, -11, -22, -32, -29, 14, -35, -89, -58, -42, -99, 52, -54, -21, 40, -10, 35, 13, -6, -2, 12, -30, 5, 23, -15, -23, -7, 24, 17, -34, -9, -30, 11, -88, -26, 0, -41, -12, 38, -49, -39, -20, -66, -11, -45, -6, 30, 6, -5, 35, 43, 0, 7, -14, 2, -1, -37, 30, 9, 7, -34, -10, 7, -4, 40, -6, 11, -42, -2, -25, 3, -29, -64, -50, -38, -39, -9, 7, -20, 12, -17, 9, 10, 59, 13, 18, -11, -10, -35, -5, 16, -34, -18, 17, 16, 35, 19, -62, 34, 0, -27, -21, -33, 9, -36, -22, -122, -12, 8, -61, -7, 14, 18, 30, -1, -21, -9, 32, 16, -7, -22, 9, -2, -16, -4, 7, 69, 6, 7, -50, 4, 1, -47, -35, -31, 59, -7, 4, -47, -62, -70, 39, 10, 20, 17, 6, 0, 9, 10, 2, 7, 24, -43, 19, -16, -28, 15, -11, 46, -18, 8, -35, -6, 14, -38, -3, -18, -28, 30, -49, -72, -26, -8, 14, 26, 16, 7, 10, 29, 35, 32, -32, 0, 30, -24, 53, -71, -11, 49, -3, 32, -23, -44, -73, -43, -12, -16, -4, -60, -1, -78, 17, -119, 8, -64, -21, 21, 12, 17, -13, -26, -2, -7, 23, 4, 19, -28, 67, -16, -2, 31, 8, 5, 42, 23, -70, 11, 14, -53, -30, 8, -84, -39, -127, -43, 10, -38, 54, 36, 29, 25, 25, 3, 45, -3, -3, -23, 30, -26, -3, 28, -17, 21, -11, 11, -14, -3, -74, -14, -7, -38, -22, 41, -4, -34, -110, -27, -19, -16, 39, 18, 36, 4, 5, -12, 42, -24, -16, -17, 28, -38, 22, 5, -40, 5, -3, -9, -30, 56, -13, 34, 1, -6, -13, 2, 37, -45, 29, -72, -72, -17, -60, 25, 14, 11, 14, 26, 22, -36, 19, -4, 7, -23, 15, -23, -38, 6, -20, 76, 37, 18, -45, 6, 12, 0, -24, -26, 55, -12, -40, -164, -29, 8, -67, 0, 13, -1, 26, 21, 11, -51, 16, -9, 1, -51, 1, -30, -78, -9, 0, 82, 0, 19, -23, -35, -18, 0, -39, -49, 12, -18, -55, -87, -23, 25, -9, 28, -5, 2, -8, 9, -37, 0, 27, -10, 16, -70, 43, -18, -55, 12, 8, 50, 3, -18, -29, -8, 0, -9, -72, 22, 16, -75, -74, -46, -64, -53, 30, 14, 6, -6, 12, 2, 21, 14, -17, -2, 3, -20, -11, -12, 4, -23, 2, 57, -1, -13, -29, 42, 29, -42, 1, -23, 42, -61, -29, -17, -53, -43, -11, 9, 44, -21, 36, 38, 49, 15, -31, -31, 9, -31, -3, -2, 1, 12, -6, 30, 0, 50, 6, -24, 14, -12, -19, 32, 32, -36, 37, -23, -51, -48, 11, 26, 50, -15, 18, 25, 59, 0, -13, -8, 34, -9, 41, 12, -26, 8, -10, -4, -19, 26, -17, 37, 5, 1, -55, -10, -13, -59, 15, 9, -27, -16, -4, 20, 7, 12, -11, -6, 24, 11, -2, -5, 14, -37, 21, 18, 26, 3, -31, -71, -24, 29, -39, 23, 2, 24, -54, -22, 15, -46, -36, 19, -50, -12, -27, 18, 18, 15, -10, 6, 8, -24, 18, -4, 36, -24, 17, 23, -84, 33, -8, 23, 5, 30, -1, 27, 41, 73, -24, -6, 19, -44, -72, -71, -39, 53, -33, 4, 33, 14, 41, -11, 12, -13, 19, 12, -13, -14, -19, -15, -58, -7, 0, 42, 11, 39, -31, -4, -7, 63, -35, -2, 19, -36, -5, -88, -32, 27, -53, -8, -21, -6, 9, 4, -19, 6, 25, -3, -15, -27, -1, -14, 2, -20, -27, 23, 11, -1, -10, 53, -11, 30, -36, 23, -33, -58, -12, -10, -5, -9, -27, 0, 22, -12, -15, 11, 33, 0, 29, -21, -15, -23, 31, 33, -62, -3, -18, 14, 0, 34, -34, 16, -37, -2, -79, 6, -7, -35, -71, -10, -46, 3, 8, -13, 31, -6, -8, -8, 22, -6, 19, -15, 4, -16, 6, 0, -27, -9, -26, -7, 4, 31, 7, 12, -58, 21, -92, -11, -31, -10, -40, -22, -47, -35, -33, 11, 30, 6, -10, -16, 24, 2, 15, -4, 8, -10, -4, 28, 6, 14, -15, -19, 0, 28, -69, 27, -40, 38, -55, -13, -26, -65, -16, 2, -52, 4, -6, 1, 11, 17, 25, 7, 40, -37, 25, 10, 2, -35, 6, 27, 9, 39, -32, -39, -2, 40, -48, 35, 26, 20, -101, 10, -29, -39, -58, -10, -33, 0, -33, 25, 22, 22, 18, -25, 12, -37, 43, 11, 12, -37, 9,
    -- layer=2 filter=0 channel=7
    -12, -17, -2, -6, -12, 10, 6, 2, 21, 11, 29, 20, 22, -36, -2, -11, 54, 15, 1, 16, -35, -34, -45, -4, -6, -6, -14, 21, -21, -28, -76, 29, -51, -18, 13, 9, 34, 4, 34, 39, -7, -36, 7, -6, 19, -30, 26, 4, 46, -4, 30, -2, -38, -22, -46, -42, 0, 25, 8, -6, -22, -33, -35, 7, -23, -47, 32, -13, 63, 0, 15, 55, -13, 13, 23, -13, 20, 0, -3, 58, -11, -4, 29, -12, -17, -33, -25, -1, 62, 18, -20, 4, 0, -57, -15, 8, 0, 2, 35, -45, 27, -50, 3, 14, -24, 73, 36, 25, 10, -80, 4, 10, 7, -27, -21, -35, 7, -21, -29, 36, 3, 18, -7, 12, -12, -16, -32, 21, 14, 30, 41, -43, -41, -20, -22, 38, 0, 11, 25, 33, 3, -71, -30, -43, 34, -13, -24, -7, -4, -3, -38, 30, 0, 9, -15, 25, -17, -31, -12, 27, -23, 38, 24, -8, 0, -8, 2, 5, 33, -66, 2, 16, 25, -44, 11, 17, 27, -15, -22, 25, -35, 8, -49, 6, -44, 22, -11, 22, 8, -25, 23, 19, -23, 8, 16, 33, 32, -17, 12, -22, 2, -47, -25, 37, 50, -58, 54, 41, -43, -10, -12, 31, -29, -27, -27, -32, -65, 42, -65, 19, -20, -13, -55, 11, 32, 8, 19, -37, -33, -10, -16, -46, 0, -10, 7, 13, 40, -113, -39, -55, 45, 8, -8, 0, 1, 16, 8, -18, 0, -20, -3, 13, -8, -6, -17, 11, 19, -42, 19, 1, 16, -14, -3, 19, 0, -2, 7, 3, 17, 0, -17, 18, 38, 23, 21, 36, -11, 24, -9, -2, -1, -18, 33, -29, -45, 0, 32, -15, -9, -52, 8, 25, 57, -20, 36, 73, -21, -27, -12, -22, -1, -29, 4, 78, -45, 29, 26, 9, 4, -44, -19, -23, 64, 9, -32, -14, -45, -7, -19, 0, 43, -18, -2, -1, 1, -24, 6, 38, 4, 22, 4, -4, -18, 34, -26, -45, -50, 10, 2, -25, -6, -16, -16, 31, 75, -34, 23, -2, -4, -6, -26, 7, 63, 31, 4, -14, -51, 4, -29, 13, 40, -2, 8, -20, -8, 28, -3, -76, 49, -39, -64, -26, -31, 13, 0, 18, 50, 18, 13, -43, -21, -13, -51, -22, 16, -15, 13, 27, 8, 0, 43, 65, 33, -25, 20, -17, -5, -32, -10, 25, 45, 22, 5, 9, -21, -9, -8, -22, 10, 0, -37, -2, -33, 16, 2, 8, -25, -17, 0, -26, 44, -42, 15, 12, -31, 6, -18, -5, 24, -22, 18, 21, -11, -9, 39, 19, 13, -53, -6, 0, 0, 18, 42, -25, -33, 10, 13, -1, 56, 26, 14, -32, -34, -10, -50, -11, -5, 9, -15, 17, 68, -70, -47, 10, 89, -46, 9, 83, 30, 26, 12, -4, -22, -16, 20, -16, -15, -28, -52, 15, 44, 28, 7, -14, -4, 7, -32, 64, -7, 27, -5, 10, 9, 0, -20, 30, 40, -28, -8, 32, -7, 34, 16, 20, 13, -21, 11, -35, -19, 11, -17, -1, -7, -27, -123, 19, 25, 11, 42, 77, 6, 12, 15, -32, -56, 54, -61, -31, -5, -81, -57, -31, -2, 0, -26, -6, 30, -35, 6, -5, -43, 19, -24, -3, 45, -16, -134, 30, 17, 18, 40, 53, 30, 20, 79, 22, -56, 6, -42, -85, -43, -32, -56, -55, -14, -22, -69, 22, 51, -10, 23, 8, -6, 4, -12, 33, 43, 0, -113, -4, -38, 35, 24, 19, 69, -5, 63, -8, -77, -65, -68, -74, 71, -53, -69, -59, -16, -12, -26, -7, 58, -24, -1, -26, 12, 5, -32, -4, 25, -13, -47, -2, -8, 10, 47, 38, 16, 26, 11, -17, -71, 3, 4, -56, 52, -28, -13, -76, 5, -31, -22, 12, 27, -31, -1, -13, -14, 8, -1, 26, -56, -4, 6, -3, 61, -32, 28, 46, -52, 39, 2, -34, 41, -42, 14, 50, -26, -36, 44, 53, 1, -24, -10, 1, 24, -10, 20, 7, -37, 15, -24, 13, 18, 71, 23, 13, -57, -3, -48, 30, -21, 11, -23, 12, 57, -57, -27, -17, 13, 45, 12, 38, 21, -3, 13, -30, -1, -43, -3, -7, 23, 0, -33, 7, 55, 40, -13, -15, -40, 2, -13, 4, 0, 58, -14, -30, -4, -57, -70, 69, 74, 5, -55, -46, 27, -13, 11, 35, 29, 33, -31, -26, 0, 1, -53, -27, 37, -16, -95, -4, 32, 23, 12, 63, 3, 29, 22, 25, -59, 75, -68, -23, 23, -41, -20, -29, 14, -25, -11, 26, 33, -41, 3, -34, -60, -10, -1, 17, 33, -21, -124, 22, -9, 36, 63, 27, 22, 35, 33, 26, -20, 71, -59, -62, -4, -61, -54, -20, -1, -25, -61, -25, -30, -25, -3, -49, -45, -29, 30, 12, 48, 11, -90, 11, -57, 34, 56, 35, 45, 27, 0, -1, -74, 48, -7, -68, 63, -117, -53, -75, 5, -18, -38, -21, -28, -32, -33, -40, -43, 23, 7, 23, 2, 9, -50, -1, 20, -4, 16, 89, -42, 13, -20, 12, -44, -2, -20, -53, -16, 7, 2, -61, -3, -15, -23, 5, 24, -2, 8, 0, -28, 7, -29, -13, 1, -27, 20, 2, 53, -28, 16, -3, -59, 4, -5, 4, 17, 25, -16, -12, -82, 17, 35, 0, 19, -19, 12, 1, 14, -39, -23, -13, 4, 20, -13, -27, 31, 41, 21, 14, -48, 26, -45, 2, 29, 22, -24, -2, 27, -20, 16, 27, 61, 38, 0, 31, 28, -20, 30, -19, -15, -19, -4, 18, 1, -21, -13, -3, 54, 59, 34, -2, -74, -12, -8, -32, 43, 41, 19, -12, -60, 1, -22, 10, 55, 9, -47, -88, 13, -4, 28, 49, 8, -45, -71, -1, 45, 9, -59, -28, 38, 47, 29, 9, -11, -28, 7, 9, -34, 39, 19, -17, -58, -26, -22, -79, 57, 9, 6, -72, 2, -17, 20, 26, -63, -37, -44, -10, -15, 8, -39, -10, 12, 58, 24, -2, 19, -22, -3, 72, -46, 42, 10, -23, 5, -6, 28, -35, 46, -8, 38, 29, 33, -11, -1, 20, -40, -13, -15, -38, -60, 24, -3, 0, 37, 20, 4, 4, -3, -13, -16, 43, -46, 62, 24, 21, -10, 31, -42, -23, 15, 15, -41, 5, 3, 7, 0, -9, -64, -21, -8, -28, -2, 19, 26, -7, 2, -7, 22, -14, 49, -37, 28, 52, -45, 34, 14, 27, -62, 41, -54, -6, -83, 22, -6, -60, -8, -9, -5, 40, 4, -18, -36, 8, -6, -2, 6, -1, -21, -35, -2, 14, 49, 9, 18, -7, -31, 7, 18, 47, -32, 53, -15, -15, -92, 12, 6, -33, 16, -2, 22, -4, -32, -70, -35, 12, -1, 11, -8, 36, 51, 42, -2, 26, -71, 33, -28, 33, 19, 21, 11, -8, 27, -42, 34, -44, 34, 26, -17, 63, 31, 37, 8, -3, -31, -4, 14, -18, 3, 0, 12, -24, 36, 46, 7, -25, -76, -1, -3, -30, 35, 58, 32, -33, -31, -71, 16, -76, 29, -14, -39, -19, -4, -7, 14, 3, -47, -19, -16, 28, 30, 1, -35, -23, 25, 53, 44, -21, -24, -22, -11, -33, 5, 49, 28, -20, -43, -65, 15, -91, 23, 10, -17, -30, -1, 6, 34, 11, -68, -35, -49, 30, 28, 7, -62, 16, -18, 35, 78, 4, 0, -13, -31, 2, -49, 17, 17, 17, -24, -33, 53, -95, -16, 18, 24, -23, 12, -16, 41, 33, -60, -58, -31, 13, 0, 39, -33, -6, 0, 1, 32, 14, 44, -32, -5, 1, -69, 41, 40, 11, -11, -17, -1, -23, -102, 26, 62, -3, 21, -7, 16, 0, -61, -43, -49, 19, 42, 6, -12, -33, -25, 25, 5, -13, 36, 7, -29, 16, -38, 59, 20, 10, -28, 67, -12, -65, -66, -5, -3, -43, -8, -3, 19, 33, -55, -100, -48, 22, 5, -23, -42, -19, 14, -7, -22, 37, 40, 31, 18, 20, -7, 44, 25, 15, -7, 49, 11, -111, -34, -18, -6, 2, 19, 33, 16, 6, -79, -22, 1, -28, 16, 9, 25, -18, 43, -22, -13, 35, 0, 52, -13, 29, 43, 14, -38, 9, 8, -15, -10, 41, 8, 17, -34, 28, 50, -8, -2, -45, -55, -5, 28, -63, -12, 13, 16, -11, 47, 17, -6, 28, -55, 12, 14, -40, 18, 37, -17, 51, -16, -67, 17, 51, 7, -40, -66, -13, 15, 25, 20, -27, -70, -28, -13, -45, 22, 13, -29, -2, -6, 20, 7, 16, -5, -7, -16, -35, -20, 11, 2, 5, -19, -67, -21, -71, -6, -7, -47, -6, 31, 16, 2, 2, -26, -27, -67, -35, 13, -3, 24, -30, 5, 0, 12, -4, 9, -18, 10, -23, -32, 49, -18, 51, -13, -49, -19, 40, -35, -33, -16, -12, 12, 35, 8, 22, -4, -39, -39, -8, 4, 0, -1, -4, 24, -37, 16, 32, 40, -39, 13, -7, -64, 57, -34, 18, -10, -41, -14, -22, -85, -11, -14, 19, 29, 10, 15, 18, -42, -61, -39, -11, 11, 26, 33, -21, -17, -28, 10, 35, 51, -23, -10, -1, -66, 23, 7, 80, 1, 7, -34, 20, -115, 14, 20, -6, 12, -13, 9, 0, -66, -62, -13, 2, 7, -17, -13, -37, 31, -6, -11, 50, 22, 24, 13, 17, -7, 45, -25, 6, 9, -3, 1, -77, -64, -22, -3, 4, 24, 41, 29, -6, -64, -24, 15, -79, -18, 11, 42, -45,
    -- layer=2 filter=0 channel=8
    -37, 31, -25, 5, 24, 21, 20, 53, 10, -120, 9, 7, 12, 15, 19, -81, 67, -14, 7, 55, -18, -28, -32, -56, -106, 27, 27, 21, -16, -1, -26, 23, -54, 31, -39, 18, -20, 19, 37, 38, 31, -20, 23, 2, -10, 25, 8, -84, 6, 4, -25, 7, 9, -28, -15, -14, -26, 22, 0, 15, 12, -11, -7, 31, -21, 0, 7, 2, -15, 23, 21, -77, 23, -28, 16, 28, -28, -9, 6, -66, -11, 10, -11, -2, -13, -68, -15, -52, -54, -10, -22, 26, 10, -10, -34, 15, -55, -2, 1, -6, -5, 11, 9, -70, 13, 38, 1, 26, -48, -12, -21, -23, -19, -6, -25, -15, -5, -20, 1, -32, -38, -29, -30, -1, 16, -14, 14, 18, -38, 37, -22, 2, 37, 27, -15, -57, 29, 10, 21, 4, -55, -1, -10, -12, 32, -5, -35, -16, -24, -16, -5, -41, -57, -47, -10, 4, 17, -17, 25, 1, 5, 41, -19, 11, 5, 39, 14, -12, 18, 6, 18, 24, -72, -20, -9, -88, 70, -1, -29, 8, -8, -28, 7, -57, -55, 0, 3, -13, 28, 23, 13, 8, -8, 32, -27, 9, -2, 44, 10, 30, 31, -48, 18, -9, -58, -1, 23, -104, 40, -6, -12, 0, 1, -38, -5, -45, -66, 0, 30, 11, 6, 4, 32, 25, -87, -12, -10, 5, -39, 42, 10, 37, 10, -29, 4, -16, -8, -5, 21, -47, 23, 25, 15, -5, -30, -52, 10, -4, -37, 27, 19, -1, 2, -13, -6, 7, -15, 17, 18, 3, -21, 12, -2, 2, 1, -10, 16, 16, -3, -4, 2, -58, 23, 14, 1, 0, 26, -18, 15, -10, -48, -6, -11, -6, 19, 13, 35, 35, -27, 12, 24, -32, -25, -3, 9, -25, -6, 8, 18, 5, -9, -28, -21, -8, 9, 28, 6, 4, 24, -6, 0, 1, -13, -45, -8, 12, 12, -42, -11, 6, -11, -26, -3, -14, 46, -22, -6, -27, -18, 14, 13, 5, 29, -9, -21, 26, 14, 5, 16, 48, 8, 6, 0, -14, -37, -37, -13, -3, 13, -39, -31, -12, -32, -40, -9, -20, -26, -11, -12, -26, -16, 10, 35, 24, -3, 8, -37, 0, -4, 32, -4, 34, 23, -14, 12, -36, -30, -22, -5, 9, 19, -25, 11, -8, 13, 15, 14, -16, -11, 11, 8, -32, 0, 11, 7, -12, 23, -3, 2, 5, 18, -18, -33, 3, 2, 38, -6, -42, -105, -56, 20, -9, 2, -37, 20, 11, -56, 48, -5, -8, -12, 20, 0, 8, 3, -54, 32, -27, -7, 21, 6, -1, 70, 30, -22, 24, -24, -20, 12, -43, -75, -26, 4, 21, 21, -18, 29, 16, -51, -25, -24, -5, -33, 3, -15, 69, -3, -33, 44, -1, -3, 33, -8, -31, 82, 0, 6, 15, -23, -33, -4, -42, -67, 2, -10, 7, 15, -31, 14, 24, -8, -21, 0, -10, 0, -1, -21, -21, -27, -23, 19, -30, -41, -84, 0, -29, 11, 5, -15, 11, 27, -3, 17, -39, -107, -1, 16, -4, 14, -25, 19, -3, -2, -23, -29, 6, -6, -7, -10, -56, -7, -18, 22, 23, 6, -26, -9, -47, 30, -26, 18, 7, 18, 37, 13, -2, -8, -30, 2, -5, 7, -43, -3, -26, -3, -4, -55, -11, 13, -13, -27, -19, -29, 35, 14, 46, -21, -55, -8, 90, 0, -24, 9, 37, 28, 30, -17, -3, -54, -19, 5, 3, -6, -47, 14, -19, -2, 8, -19, 0, 21, -37, -24, -16, -15, 59, 27, 24, 22, -62, 9, 4, 2, 17, -1, 36, 8, 23, 10, 24, -22, -58, 17, -5, 23, -34, 13, -5, -24, -13, 13, 0, -29, -5, 4, 36, -16, 11, 11, -5, 4, -66, 0, -16, -19, 51, 0, 8, 24, 19, 16, -23, -50, -24, 1, 6, 20, -35, 9, -16, -61, 43, 8, 13, -58, 7, 16, 24, 37, -50, 37, 17, -12, -84, 17, -13, 49, 30, -22, 25, 29, -6, 34, -49, -77, -16, 20, 14, 33, -18, 6, 7, -24, -18, -29, -20, -4, 12, 24, 15, 16, -19, -3, 22, -2, -3, 36, -79, 61, -6, -5, 27, -4, -15, -13, -11, -1, -5, 5, -3, -8, -56, -8, 17, -22, -13, -3, 4, 13, 25, 0, 22, -2, -9, 8, 18, 2, 36, 19, 11, 30, -19, -8, -6, 27, -1, 7, -17, -31, -22, 8, -26, 18, -8, -3, -11, -39, -32, -17, -9, -5, -6, -12, -13, -17, 3, 7, -3, -6, -24, 13, 24, 10, -25, 29, 0, 4, 11, 0, -21, -47, 0, 25, -9, 3, -28, 19, -16, -15, -5, -31, -21, 5, -25, -51, -21, -32, 18, -16, 0, 9, -59, 40, -2, -36, -29, 26, 38, 3, 0, -10, -14, -55, -25, 26, 2, -4, -36, 26, -5, -24, -9, -40, 2, -2, -35, 2, -4, -59, 15, 6, 5, 34, -83, 2, 32, -37, 13, 7, 62, 19, 13, -1, -7, -43, -6, 7, -14, -6, -28, 31, -26, -16, -8, -8, 4, -43, -6, 6, 5, -32, 14, 11, -19, 44, -65, -2, -64, -26, 4, -25, 65, 29, 10, 26, -32, -41, -14, 13, -18, -19, -28, 37, -41, -35, 24, -12, -37, -71, 9, 8, 44, 6, 15, 32, 19, 32, -58, 6, 16, 15, 13, -10, 84, -33, 6, 21, -19, 7, -24, 8, 8, 15, -28, -6, -16, -1, 13, -55, -20, 33, -18, -6, 13, -39, -51, -14, -10, 27, 0, 39, -44, 92, -35, 34, 25, -51, 11, -8, 21, 46, 36, 0, 14, 5, -56, -17, -15, -40, -41, -23, 42, 11, 17, -22, -3, -16, -22, -42, 28, -4, 32, 21, -99, 23, 36, 32, 59, -14, -11, 21, -5, 27, -8, 31, -29, 0, -3, 18, -16, -64, -18, -24, 16, -21, -9, 18, -48, -24, -47, -9, 11, 26, 3, 27, -32, 4, -40, 39, 68, 11, 0, 13, -35, 16, -8, 25, 9, -11, -4, 45, -25, -28, -24, -11, 29, -43, 8, 37, -33, -9, -96, -7, 4, 38, -35, 30, 28, -39, -10, 35, 31, -16, 32, -19, -32, -82, 9, 29, 32, 23, -14, 41, -20, -34, -11, -22, 14, -64, -25, 35, -11, 4, -46, -3, 2, 24, -72, 30, 78, -12, 22, 9, 61, -3, 34, 17, -53, -51, -42, 33, 12, 13, -6, 41, -20, -19, -2, -8, 6, -30, -11, 5, 41, -23, -32, -26, -8, 52, -7, 6, 67, -3, -1, 6, 61, 36, 25, 29, 3, 23, -4, 36, -13, -24, 9, 20, -24, 5, 12, -60, -18, -34, 16, 7, 89, 6, -10, 5, 17, 65, 9, -11, 99, 9, -22, -10, 39, -33, -20, -3, 32, 21, -25, 30, 0, 23, -42, -12, -30, -11, -9, -60, -49, 29, -34, -8, -33, -34, -34, -9, -33, 20, 15, 3, 14, 30, 7, 33, 5, -110, 26, -38, 46, 56, 23, 2, 36, -27, -59, -14, -7, -58, -12, -6, 18, 33, -12, -25, 4, 19, -72, -46, 28, 60, 48, 6, -3, -8, 36, 8, -1, -24, -20, 6, 2, 87, 25, 16, 0, -21, -21, 32, -37, -48, -28, -4, 27, -22, 17, -10, 8, 28, -131, -30, -4, 21, 54, 21, 41, 38, 72, 15, 28, -29, -3, -6, -70, 52, 24, 53, -7, -44, -8, 69, -25, -54, -48, 32, 58, -77, 8, 25, -10, 33, -180, -34, -17, 39, 49, 49, 17, 24, 37, 40, 39, -33, -13, -23, -115, -19, -12, 32, 21, -40, -6, 57, -10, -21, -34, -15, 52, -42, -11, 15, -40, 30, -133, -40, -40, 46, -29, 58, 73, 34, 4, 9, 28, -24, 17, 0, -50, 28, -17, 43, 28, 0, -1, -3, -39, -34, 3, -27, 71, -87, 30, 8, 16, 27, -62, -35, -27, 48, 8, 2, -1, 10, 1, 2, 52, -20, 18, -1, -22, 63, 18, 51, 0, -17, -8, 30, -13, -24, 9, -71, -45, -57, -9, -27, 38, 51, 8, -34, -17, 21, 4, -4, 40, 13, -22, 14, 29, -32, -7, -28, 43, 91, -24, 26, 27, 10, -22, -22, 0, 9, -30, -71, -98, 36, -37, -15, -57, -22, 22, -41, 37, -48, -35, 6, -39, 61, 40, 52, -41, -81, -16, -45, 57, 69, 37, -13, 95, -2, -59, -120, 29, -6, -14, -18, 0, -1, -22, -25, 1, -15, -55, -47, 40, -16, 60, 4, -46, 27, 54, 13, -28, -31, -26, -13, 25, 54, 20, 45, 12, -35, 24, 3, 21, -52, -20, 8, 13, -36, -26, 0, 9, 8, -123, -58, 46, 3, 43, -8, -13, 17, 62, 47, -14, -6, -52, -11, -15, 79, 43, 67, 26, -31, 22, 4, 0, -53, -13, 38, 21, -52, -20, -7, 22, 41, -158, -49, -40, 20, -4, 17, -22, 71, 42, 17, 2, -53, -14, -16, -36, 66, 45, 50, 12, -17, 12, 36, -11, -37, -45, 21, 5, -34, 9, -3, 20, 46, -168, -56, 4, 17, 5, 28, -14, 29, 16, 17, -5, -19, -41, -3, -26, 73, -6, 38, 21, 6, 4, 40, 7, -7, 0, -12, -13, -46, 1, -22, 31, 49, -68, -49, -8, 0, -30, 33, -11, 58, 61, -4, -21, -20, -29, 6, -17, 98, 0, 56, 21, 9, -22, 33, 10, -14, 39, -110, -115, -90, -21, 2, 41, 0, -25, -11, 28, -42, -15, 6, -22, 42, -21, 30, -42, -64, -94, -56, 29, 90, -23, -1, 82, 8, -70, -79, 30,
    -- layer=2 filter=0 channel=9
    1, -23, 3, 43, 3, 7, 52, -68, 33, -24, 25, 7, -22, -49, 52, 23, -24, 4, -7, 0, -50, -14, -15, -3, 46, 42, -13, 13, 13, -39, -70, 18, -22, 5, 20, 35, -35, 9, 18, -67, 11, -6, 29, 25, 16, -40, 18, -36, 10, 18, -30, -59, -23, -6, -4, 32, 80, -26, -2, 6, 0, -1, -39, 4, -20, -17, 3, -8, -4, 1, 35, 9, -3, -30, -20, 16, 64, -55, 1, -37, -9, -20, 2, -12, -16, 3, -20, 4, 21, 38, 23, -7, -21, -23, -38, -2, -30, -17, 4, 37, 7, 11, 11, 3, 10, -37, -17, -9, 68, 6, 3, -6, 33, -48, 4, 1, -10, 43, 4, -8, 17, -1, 45, -3, -43, 11, 13, 4, -47, -12, 31, 41, 22, -5, 37, -44, 2, 9, -19, 6, 38, -33, 16, -47, -28, 18, 10, 8, -8, -13, -10, 11, 39, 53, 27, -18, -33, 9, -18, -9, -67, -15, 20, 19, 19, 3, 21, 26, 0, -5, -4, 13, 48, -15, 32, -64, -36, -2, 3, -30, -6, -51, 9, 54, 70, 6, -13, 11, -10, -9, -48, 25, -57, -30, 14, 8, 17, 5, 44, -13, 38, 16, 12, 71, 0, -6, 22, -117, -24, -35, 3, -13, -26, -27, -22, 37, 24, -1, -12, 11, 18, -2, -49, 27, -44, -6, 26, -5, 1, -5, -7, 53, -2, 4, 34, 1, 7, 0, -15, 72, -42, -24, -5, -20, -5, -6, 3, 10, 1, 30, 12, -5, -8, 6, -6, -2, -21, 7, 43, -10, -1, 1, 23, 12, 0, 18, -1, 5, 5, -42, 4, 11, -15, 31, -5, 7, -28, -9, -21, 30, -2, -25, 6, 2, 2, -4, -9, 10, 0, 14, 1, 2, -42, 0, 17, 8, 0, 30, -8, 7, -7, -17, 9, 6, 16, -27, 14, 4, -28, 18, -3, 10, -18, -24, 31, -15, -15, -33, 17, -8, -1, -13, 16, -32, -19, 5, 18, 0, 8, 19, -4, 30, 5, -41, 12, 39, 7, 18, -5, -14, 1, -9, 6, 0, -25, -27, 40, 10, -18, -26, -16, 12, -12, 25, -20, -22, -17, -13, -1, 37, -12, -12, -5, 14, 32, -50, 28, -126, 2, 5, 3, 10, -13, -16, -23, 1, 0, -15, 29, -9, -19, -37, 0, 12, -43, -9, 14, -12, 1, 14, -13, 19, 1, -2, -5, 17, 29, 1, 1, 28, -39, 9, 14, -4, -13, -15, -17, 6, 39, -1, 0, -3, -4, -38, -24, 25, -12, -4, 67, 30, -3, -6, 0, -11, 27, -2, -3, 21, 24, -12, 25, -58, 9, 8, 30, -30, 12, -27, -8, -2, 6, -31, 28, -3, 12, 15, 19, 34, -35, 17, 6, -19, 8, 14, 0, -10, -9, 20, -14, -18, 1, 11, -10, 26, -29, -67, -32, 23, -8, 7, 5, 72, 6, 17, 23, -21, -48, 5, -2, -18, -15, -2, -21, -23, 11, 25, 11, -51, -2, 5, 4, 5, -2, -48, 14, -31, 16, -18, 6, -7, -18, -1, -3, 7, -5, 0, 10, 2, 10, -13, -28, -8, 0, 13, 10, -24, -5, 9, -7, 11, -15, 20, -17, -3, 23, -33, -23, -70, 16, 13, 34, -43, -13, -11, -17, 14, -27, 0, 16, 32, 0, -20, 18, -13, 24, -22, -4, -4, 8, 36, -29, -40, -2, 68, -5, 16, -12, 1, 7, -63, -16, -3, -3, -66, 17, 9, -10, 4, -21, 0, -8, 37, 18, -30, -15, -12, 63, 11, 23, -11, -2, 8, -14, -69, 12, 45, 30, -5, -1, 13, 13, -123, -30, 37, 13, -51, 0, 10, -7, 19, -23, -26, 0, 27, 29, -42, 2, 5, -13, 8, -15, 1, -4, 0, -16, -12, -9, 15, 12, 30, -10, -32, 14, -3, -57, -18, 28, -28, -48, -8, -24, -4, 6, -37, 12, 26, 3, -49, 22, 10, 2, -55, -36, 13, -11, -25, -34, 20, -12, 22, -6, 38, -9, -22, 8, 39, 7, -30, 17, -16, 0, -38, -23, -16, 2, -38, 19, -10, -33, -22, 22, -4, -29, -29, -34, -16, -14, -20, -72, 19, -9, 25, -30, -28, 28, 19, -29, 52, -8, -102, -30, 53, -10, 10, -21, 46, -15, -12, 27, -8, -67, 20, -15, 9, 21, 26, -1, -8, -25, 0, 3, -73, -28, 19, 45, 11, 6, -71, -8, -74, -21, 18, 20, 20, -13, 18, -31, 7, -60, -62, 14, 39, 33, -18, 11, 31, 45, 37, 29, 41, -52, 9, 8, -29, -6, 33, 16, -21, -51, -56, -16, -82, -28, 41, 34, -34, 20, 2, -14, 33, -81, -8, -16, 29, 20, 15, 57, 2, 47, 13, 38, 20, -22, -6, 2, -66, -36, 56, 35, 29, -35, -28, 0, -117, -48, 60, 60, -24, 50, 34, -21, 20, -59, -18, 0, 46, 31, -3, 44, -12, 40, 34, 19, 31, 6, -28, -19, -46, -9, 49, 76, -8, -52, 41, 11, -85, -39, 28, 37, -42, -5, 10, -19, -8, -1, -25, 9, 25, 61, -22, 46, -7, 31, 0, 29, 17, 3, -6, 19, -61, -17, 12, 43, 5, 12, -25, 13, -69, -27, 33, 56, 7, 5, 12, -36, -33, -30, -53, 4, 18, 20, -41, 30, 7, 25, -15, -18, 27, 10, -31, -31, -5, -25, 26, 0, -17, 15, -35, -4, 31, 6, -44, 4, 10, 22, 22, -5, -31, 9, 0, 19, -26, -21, -24, 15, -60, -1, -20, -50, -19, 19, -12, -60, 46, -16, 18, -46, 3, 20, 35, -17, -93, -8, -49, -33, 60, 12, 10, -38, 23, 22, 26, 42, -71, -88, 4, -10, -26, 16, 36, -12, -7, 16, -18, 18, -13, -22, 18, -4, 14, 15, -46, -14, -64, 9, -42, 14, 14, -34, 14, -42, 14, -33, 9, 10, 2, 3, -20, 32, -19, 28, 65, 16, -17, -3, -5, 19, -50, 5, 0, 31, 23, -36, -43, -7, -63, 2, 35, 6, 16, -1, 22, -31, -12, -78, 32, 8, -3, 22, 37, 19, 0, 25, 23, 19, 18, 13, 9, -22, -38, 0, 17, -15, 27, -77, -71, -2, -174, -50, 37, 49, -36, -6, 37, -40, -1, -50, -17, 12, 39, 14, 7, 19, 7, 29, 3, 11, 6, 11, -12, -6, -47, -20, 10, 24, -2, -60, -21, -3, -105, -66, -4, 31, 10, 21, -12, -41, -27, -47, 0, 14, 13, -9, -27, 18, 16, 13, 0, 5, -18, 24, -35, -18, -29, -15, 21, 40, -27, -34, -46, -7, -149, 1, -29, 30, 44, -9, -17, -30, -26, -33, 12, 27, -8, 14, -29, 4, 27, 39, 28, -13, 11, 46, -15, -65, 6, 6, 26, -65, -38, -24, -85, -8, 10, 58, -116, 33, -8, 13, 15, -12, 1, -34, 20, 34, -65, 10, 13, 15, -79, -8, 8, -17, 3, 46, -19, -45, 51, -29, 15, -47, 1, 25, -50, -62, -59, -43, -14, -49, 52, 19, -55, -7, -23, 5, -3, 32, -85, -5, 2, -43, -39, 2, 43, -26, -35, 33, -39, -18, 13, -30, 25, 23, -38, 21, -2, 8, -73, -15, -27, -8, 22, -48, -40, -40, -15, -28, 13, 34, -25, 0, -17, -26, 6, 16, 93, -42, -59, 19, -15, -10, 30, 8, 1, 20, -75, -14, -25, -19, -112, -11, -1, -3, 17, -24, -4, -9, 0, -54, 24, 44, -19, 4, 5, -39, -16, 24, 29, -15, -28, 42, -15, 15, -4, -20, -23, 12, -15, -38, -60, -12, -124, -47, 71, -2, 11, -26, 15, -24, -7, -15, 52, 2, -33, -16, 20, -45, -25, -13, 49, -16, 16, 38, 5, -36, 8, -12, -38, 8, -16, 1, 22, -20, -85, -18, 73, -11, 13, -20, 2, -31, -13, -76, 30, 18, -2, -1, -20, -20, 0, 6, 69, -24, -34, 38, 5, -21, 5, -30, 1, 16, -30, 6, -31, 16, -54, 2, 25, -9, 27, -16, -23, -26, -34, -79, 16, 31, 2, -8, -22, -16, 36, 41, 33, -8, 11, 22, 3, -21, 18, -11, 13, -27, -35, 0, -36, -27, -9, 41, -10, -16, 52, 30, 15, 4, -14, -22, 22, 22, -86, 13, 22, -20, -20, -61, 63, -9, 5, 60, 17, -3, 10, -29, -68, -26, 26, 0, -6, -32, -21, -53, 66, -120, 39, 38, -107, 4, -115, 16, -3, -7, -65, 2, -7, -40, -45, 0, 68, -25, -53, 71, 11, -19, 4, -47, 27, -7, -56, 26, -36, 0, -191, 0, 51, -9, 41, -21, -52, -19, -54, -28, -6, 49, -45, 10, -13, -17, 13, -2, 58, -45, -46, 52, 16, -10, 23, 23, -7, 3, -61, 16, -31, 15, -6, -8, 36, -28, 37, -28, 0, -18, -39, -67, 51, 13, -7, 8, 5, -8, -1, -50, 87, -27, -37, 19, 34, 20, 9, -1, -46, 1, -20, 35, -5, -27, -29, 23, 62, -23, 26, -51, -3, -18, 0, -6, 19, 0, -1, 10, -7, -42, -29, -7, 62, -41, -27, 19, 34, -6, -32, 12, -14, 29, -24, 9, 22, -52, -87, 0, 74, -31, 28, -33, 3, -26, -27, -5, 21, 13, -38, 33, -26, -5, -19, -22, 95, -42, -33, 10, 46, 15, 8, 20, -14, 10, -2, 15, -39, -41, -71, 11, 51, 3, 22, -16, -15, -24, -34, -73, 48, 17, -26, -1, 0, 4, -20, 2, 56, -4, 8, -21, 0, -42, -6, -1, -52, -40, 0, 22, -51, -82, 2, 33, 61, -77, 42, -7, 15, -8, 6, -95, 62, -8, -83, 5, 25, -36, -60,

    others => 0);
end iwght_package;
