LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias

					-- weights

			324, 249, 301, 
			153, 153, 66, 
			79, 244, 268, 
			

			0, 0, 0, 
			20, 0, 0, 
			100, 179, 158, 
			

			120, 27, 81, 
			352, 153, 283, 
			323, 324, 138, 
			

			372, 449, 297, 
			278, 294, 269, 
			126, 0, 0, 
			

			405, 324, 240, 
			235, 159, 72, 
			73, 0, 6, 
			

			250, 399, 531, 
			402, 533, 410, 
			378, 62, 85, 
			

			84, 13, 0, 
			0, 0, 0, 
			0, 0, 12, 
			

			348, 180, 151, 
			250, 220, 86, 
			541, 338, 265, 
			

			302, 547, 351, 
			585, 525, 346, 
			521, 435, 391, 
			

			0, 0, 0, 
			0, 76, 0, 
			23, 119, 105, 
			

			272, 394, 518, 
			364, 281, 388, 
			253, 58, 20, 
			

			57, 0, 0, 
			0, 0, 0, 
			0, 196, 121, 
			

			102, 0, 0, 
			50, 101, 86, 
			268, 382, 347, 
			

			215, 335, 292, 
			257, 278, 249, 
			313, 240, 221, 
			

			0, 113, 190, 
			232, 243, 55, 
			447, 111, 50, 
			

			0, 0, 4, 
			0, 0, 102, 
			0, 0, 0, 
			
