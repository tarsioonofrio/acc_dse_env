library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    47, 47, 52, 47, 47, 45, 54, 54, 41, 24, 23, 39, 43, 41, 35, 
    52, 52, 53, 46, 53, 64, 27, 29, 5, 24, 2, 6, 26, 43, 38, 
    2, 65, 53, 50, 51, 22, 2, 0, 12, 41, 0, 5, 0, 21, 54, 
    0, 80, 48, 53, 26, 38, 4, 0, 1, 41, 0, 0, 0, 0, 66, 
    0, 44, 26, 67, 28, 14, 0, 0, 0, 71, 2, 0, 8, 0, 26, 
    0, 26, 25, 11, 41, 12, 0, 0, 0, 107, 0, 0, 11, 0, 2, 
    0, 0, 33, 4, 46, 50, 0, 0, 0, 80, 0, 0, 9, 13, 0, 
    0, 0, 0, 12, 32, 34, 0, 0, 0, 59, 0, 0, 14, 10, 32, 
    0, 1, 0, 37, 0, 7, 0, 0, 34, 0, 0, 0, 17, 48, 48, 
    0, 0, 0, 37, 0, 13, 42, 0, 0, 0, 0, 0, 38, 59, 29, 
    34, 0, 0, 96, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    26, 31, 30, 31, 31, 31, 32, 33, 35, 27, 15, 14, 20, 29, 30, 
    28, 39, 33, 34, 28, 40, 39, 35, 15, 1, 12, 16, 7, 8, 26, 
    30, 0, 32, 33, 34, 19, 8, 4, 5, 0, 3, 0, 11, 1, 10, 
    32, 4, 31, 32, 41, 4, 27, 6, 0, 0, 0, 3, 0, 6, 0, 
    0, 15, 27, 0, 31, 28, 13, 8, 3, 0, 9, 17, 1, 6, 7, 
    0, 0, 16, 44, 0, 0, 13, 9, 22, 0, 2, 0, 0, 0, 7, 
    0, 10, 0, 41, 1, 0, 1, 0, 10, 0, 0, 4, 0, 0, 5, 
    0, 0, 0, 17, 6, 1, 0, 0, 0, 1, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 16, 0, 21, 5, 0, 0, 0, 30, 
    0, 0, 0, 0, 5, 0, 0, 19, 10, 0, 0, 0, 0, 20, 20, 
    0, 0, 0, 0, 9, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    9, 6, 8, 5, 7, 10, 5, 6, 8, 7, 7, 13, 10, 5, 8, 
    12, 9, 8, 3, 12, 17, 0, 1, 2, 34, 14, 16, 26, 25, 9, 
    0, 36, 10, 6, 12, 23, 0, 22, 27, 47, 0, 2, 0, 31, 27, 
    0, 67, 9, 15, 0, 31, 3, 0, 10, 53, 0, 8, 3, 8, 59, 
    0, 30, 0, 48, 0, 0, 0, 0, 3, 76, 3, 0, 17, 0, 32, 
    0, 13, 0, 0, 55, 0, 0, 0, 0, 106, 0, 0, 25, 3, 5, 
    0, 0, 12, 0, 56, 32, 0, 0, 0, 89, 0, 0, 25, 29, 0, 
    0, 0, 0, 1, 39, 27, 0, 2, 0, 54, 0, 0, 32, 8, 4, 
    0, 4, 0, 37, 0, 24, 10, 13, 34, 6, 31, 0, 35, 33, 13, 
    0, 1, 0, 59, 0, 0, 36, 0, 0, 0, 0, 28, 41, 29, 3, 
    55, 0, 0, 90, 0, 0, 9, 0, 0, 3, 35, 28, 28, 40, 26, 
    59, 28, 0, 49, 0, 0, 36, 35, 22, 27, 27, 29, 29, 26, 19, 
    12, 55, 54, 0, 0, 20, 17, 23, 26, 29, 33, 27, 17, 24, 31, 
    11, 29, 72, 0, 2, 26, 15, 22, 25, 24, 24, 27, 25, 38, 2, 
    0, 26, 30, 37, 21, 36, 25, 19, 24, 23, 14, 31, 47, 2, 0, 
    
    -- channel=3
    5, 6, 0, 0, 0, 2, 1, 2, 2, 16, 27, 20, 5, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 17, 35, 0, 0, 0, 18, 16, 1, 
    36, 36, 1, 0, 0, 34, 23, 15, 0, 0, 0, 0, 0, 20, 6, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 14, 0, 9, 5, 6, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 13, 
    12, 0, 0, 15, 52, 22, 0, 0, 0, 0, 5, 14, 1, 0, 0, 
    0, 0, 28, 0, 10, 0, 9, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 30, 25, 6, 0, 6, 0, 4, 8, 0, 
    0, 0, 0, 0, 0, 34, 2, 0, 0, 0, 28, 36, 12, 0, 0, 
    7, 0, 0, 0, 6, 13, 0, 0, 0, 45, 33, 9, 0, 0, 7, 
    2, 0, 0, 0, 0, 0, 4, 36, 23, 0, 0, 0, 0, 18, 20, 
    49, 27, 0, 0, 52, 57, 27, 25, 16, 4, 0, 0, 0, 0, 0, 
    0, 36, 10, 7, 52, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 40, 46, 13, 0, 0, 0, 0, 0, 0, 7, 0, 0, 24, 
    0, 0, 3, 31, 11, 16, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    14, 17, 20, 18, 16, 19, 19, 18, 16, 12, 6, 10, 14, 8, 5, 
    16, 21, 23, 18, 25, 51, 14, 16, 0, 11, 3, 0, 0, 10, 10, 
    0, 24, 20, 18, 19, 8, 0, 0, 0, 31, 0, 0, 0, 0, 15, 
    0, 29, 16, 25, 14, 25, 17, 0, 0, 23, 0, 0, 0, 0, 16, 
    0, 45, 7, 63, 82, 42, 0, 0, 0, 30, 14, 0, 0, 0, 0, 
    0, 28, 4, 0, 25, 16, 16, 0, 0, 78, 0, 0, 0, 0, 0, 
    0, 1, 1, 0, 29, 47, 28, 8, 0, 67, 0, 0, 0, 4, 0, 
    8, 18, 0, 14, 30, 66, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    15, 33, 0, 27, 0, 0, 0, 0, 18, 0, 0, 0, 0, 3, 18, 
    22, 24, 0, 31, 0, 0, 28, 25, 0, 0, 0, 0, 12, 29, 12, 
    49, 26, 0, 91, 43, 25, 53, 19, 0, 0, 0, 5, 1, 9, 0, 
    4, 33, 23, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 50, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 10, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 9, 14, 0, 0, 
    19, 19, 0, 0, 0, 0, 26, 13, 4, 0, 0, 0, 0, 0, 0, 
    33, 53, 9, 18, 89, 53, 0, 0, 0, 0, 16, 15, 6, 15, 0, 
    0, 0, 3, 0, 0, 0, 14, 11, 11, 27, 0, 0, 0, 9, 21, 
    0, 0, 0, 0, 0, 6, 4, 7, 6, 10, 0, 0, 0, 8, 11, 
    1, 9, 20, 17, 14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 2, 0, 9, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 2, 7, 0, 0, 40, 0, 0, 0, 0, 27, 18, 0, 
    0, 0, 0, 31, 94, 73, 33, 0, 8, 4, 17, 42, 20, 0, 0, 
    0, 0, 21, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 10, 2, 0, 13, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 23, 16, 3, 
    
    -- channel=6
    22, 21, 25, 26, 26, 21, 28, 26, 24, 17, 5, 4, 11, 20, 18, 
    24, 26, 30, 28, 26, 32, 34, 17, 4, 0, 5, 0, 0, 0, 17, 
    9, 0, 26, 25, 32, 12, 0, 0, 0, 12, 15, 0, 15, 0, 1, 
    10, 12, 26, 23, 23, 0, 24, 13, 5, 7, 4, 7, 0, 0, 0, 
    4, 46, 33, 14, 46, 64, 14, 1, 0, 0, 15, 18, 0, 0, 5, 
    9, 6, 22, 48, 0, 0, 17, 9, 8, 22, 25, 0, 0, 0, 3, 
    2, 30, 0, 15, 14, 15, 21, 12, 0, 31, 0, 0, 0, 1, 12, 
    16, 1, 19, 6, 32, 35, 6, 0, 0, 32, 1, 0, 0, 9, 0, 
    17, 12, 12, 0, 30, 0, 0, 9, 0, 29, 0, 0, 0, 0, 35, 
    1, 17, 1, 8, 3, 8, 0, 30, 25, 0, 0, 0, 3, 33, 19, 
    0, 16, 0, 16, 54, 49, 44, 0, 0, 0, 0, 5, 3, 0, 0, 
    0, 0, 4, 73, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    
    -- channel=7
    38, 41, 37, 39, 38, 35, 44, 41, 37, 45, 45, 41, 34, 33, 32, 
    35, 38, 40, 43, 35, 34, 40, 51, 49, 10, 11, 14, 22, 34, 37, 
    61, 46, 40, 39, 39, 60, 29, 4, 0, 10, 24, 11, 24, 18, 36, 
    29, 3, 42, 37, 46, 9, 29, 14, 16, 20, 30, 21, 11, 11, 22, 
    11, 33, 42, 5, 52, 21, 32, 14, 22, 0, 15, 18, 12, 15, 8, 
    1, 41, 38, 23, 41, 15, 34, 14, 23, 0, 43, 16, 16, 12, 0, 
    0, 61, 29, 46, 33, 9, 68, 22, 32, 22, 28, 8, 1, 3, 16, 
    0, 33, 4, 37, 13, 67, 53, 32, 20, 27, 25, 11, 8, 29, 13, 
    15, 30, 11, 26, 14, 15, 8, 19, 8, 24, 29, 26, 3, 9, 31, 
    29, 24, 31, 0, 34, 8, 0, 34, 13, 48, 37, 2, 16, 39, 43, 
    38, 23, 30, 0, 27, 18, 52, 66, 42, 7, 0, 0, 9, 27, 22, 
    39, 30, 19, 44, 82, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 
    1, 17, 0, 85, 9, 0, 1, 0, 0, 0, 0, 0, 9, 1, 0, 
    0, 0, 7, 92, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 30, 
    1, 0, 0, 22, 1, 0, 9, 0, 0, 0, 0, 0, 0, 7, 0, 
    
    -- channel=8
    0, 2, 0, 2, 1, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 4, 0, 22, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 4, 0, 0, 7, 0, 0, 0, 7, 6, 3, 0, 0, 
    29, 0, 5, 0, 8, 0, 8, 0, 0, 0, 30, 0, 0, 0, 0, 
    36, 8, 24, 0, 45, 23, 34, 12, 0, 0, 18, 16, 0, 3, 0, 
    14, 22, 38, 0, 0, 10, 48, 15, 23, 0, 37, 18, 0, 0, 0, 
    22, 38, 5, 17, 0, 0, 24, 29, 23, 0, 38, 11, 0, 0, 6, 
    26, 45, 11, 18, 0, 0, 46, 0, 12, 0, 22, 13, 0, 0, 10, 
    39, 18, 38, 0, 1, 0, 8, 1, 0, 10, 0, 7, 0, 0, 0, 
    25, 16, 55, 0, 16, 0, 0, 30, 1, 0, 3, 0, 0, 0, 2, 
    0, 19, 50, 0, 88, 14, 0, 17, 26, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 46, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 34, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 48, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 5, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 0, 4, 0, 8, 0, 0, 0, 0, 0, 
    0, 8, 0, 13, 0, 0, 0, 0, 0, 0, 11, 0, 1, 0, 0, 
    15, 6, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    38, 1, 0, 23, 0, 0, 27, 27, 3, 0, 0, 1, 4, 6, 0, 
    53, 44, 0, 16, 7, 27, 20, 20, 21, 17, 22, 21, 23, 20, 22, 
    21, 44, 33, 21, 1, 19, 17, 17, 15, 18, 18, 21, 27, 28, 24, 
    26, 25, 54, 42, 18, 16, 11, 16, 21, 23, 25, 34, 26, 37, 42, 
    23, 31, 29, 21, 16, 33, 35, 23, 18, 15, 16, 20, 23, 16, 15, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 3, 7, 6, 3, 6, 2, 0, 2, 0, 0, 0, 2, 0, 0, 
    5, 8, 6, 3, 11, 72, 5, 0, 0, 12, 21, 0, 0, 0, 0, 
    0, 0, 3, 4, 0, 0, 0, 0, 3, 41, 25, 31, 0, 0, 0, 
    0, 30, 0, 8, 5, 19, 35, 14, 6, 5, 27, 0, 0, 0, 0, 
    52, 63, 8, 42, 116, 72, 30, 20, 0, 39, 48, 18, 17, 6, 0, 
    30, 52, 21, 0, 8, 37, 66, 28, 8, 78, 32, 3, 7, 16, 16, 
    62, 24, 0, 0, 0, 74, 31, 47, 6, 49, 24, 17, 10, 29, 17, 
    71, 64, 25, 15, 16, 47, 16, 0, 11, 29, 28, 3, 7, 2, 16, 
    76, 62, 30, 40, 22, 0, 9, 23, 31, 0, 0, 0, 0, 20, 18, 
    63, 60, 38, 45, 15, 16, 52, 63, 11, 0, 0, 0, 13, 20, 0, 
    52, 59, 23, 129, 146, 72, 50, 22, 16, 3, 18, 36, 18, 0, 0, 
    0, 45, 67, 105, 0, 0, 0, 0, 0, 4, 11, 13, 27, 24, 23, 
    17, 0, 79, 39, 0, 23, 13, 12, 13, 20, 29, 36, 20, 21, 57, 
    21, 16, 9, 2, 15, 24, 25, 13, 17, 24, 17, 10, 18, 44, 0, 
    24, 23, 5, 0, 0, 0, 1, 23, 35, 40, 19, 24, 69, 49, 15, 
    
    -- channel=12
    1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 4, 0, 4, 4, 0, 0, 0, 1, 0, 0, 7, 4, 0, 
    0, 11, 1, 0, 6, 0, 0, 0, 10, 35, 0, 0, 0, 16, 7, 
    0, 64, 0, 1, 0, 3, 0, 0, 0, 55, 0, 0, 0, 0, 43, 
    0, 35, 0, 44, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 31, 
    0, 0, 0, 14, 32, 0, 0, 0, 0, 134, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 46, 34, 0, 0, 0, 101, 0, 0, 2, 9, 0, 
    0, 0, 0, 0, 37, 51, 0, 0, 0, 66, 0, 0, 16, 3, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 15, 0, 18, 0, 17, 14, 16, 
    0, 0, 0, 38, 0, 1, 14, 0, 3, 0, 0, 0, 29, 25, 0, 
    28, 0, 0, 113, 0, 0, 32, 0, 0, 0, 3, 9, 9, 0, 0, 
    42, 2, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 45, 47, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 4, 0, 0, 6, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
    
    -- channel=13
    36, 42, 41, 39, 38, 41, 44, 46, 40, 28, 23, 30, 36, 34, 33, 
    41, 49, 44, 41, 43, 50, 25, 32, 24, 21, 4, 2, 13, 31, 31, 
    11, 41, 43, 44, 43, 33, 17, 7, 7, 20, 0, 0, 0, 5, 37, 
    0, 26, 38, 45, 30, 30, 13, 0, 0, 17, 0, 0, 0, 0, 35, 
    0, 14, 18, 43, 27, 3, 0, 0, 0, 29, 6, 0, 1, 0, 1, 
    0, 5, 16, 23, 39, 13, 12, 0, 0, 43, 0, 0, 2, 0, 0, 
    0, 0, 19, 29, 34, 29, 5, 0, 0, 35, 0, 0, 0, 6, 0, 
    0, 0, 0, 21, 22, 20, 0, 0, 0, 26, 0, 0, 3, 1, 13, 
    0, 0, 0, 21, 0, 10, 7, 4, 8, 9, 10, 0, 6, 24, 30, 
    0, 0, 0, 17, 0, 0, 16, 9, 0, 0, 0, 0, 13, 33, 25, 
    21, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    70, 70, 71, 70, 71, 67, 74, 80, 75, 66, 59, 60, 60, 60, 61, 
    72, 72, 73, 72, 72, 57, 59, 68, 59, 37, 13, 20, 40, 58, 59, 
    55, 77, 74, 76, 76, 70, 53, 36, 19, 10, 0, 0, 0, 30, 55, 
    0, 31, 68, 77, 64, 53, 18, 2, 4, 20, 8, 11, 6, 5, 47, 
    0, 0, 49, 66, 14, 2, 6, 3, 4, 23, 5, 0, 4, 0, 20, 
    0, 8, 45, 54, 48, 26, 9, 2, 0, 21, 3, 6, 7, 0, 0, 
    0, 0, 50, 55, 36, 29, 16, 8, 0, 18, 3, 0, 4, 4, 0, 
    0, 0, 3, 36, 28, 21, 5, 18, 9, 22, 13, 1, 7, 9, 26, 
    0, 0, 0, 17, 17, 27, 19, 9, 14, 24, 28, 13, 12, 25, 45, 
    7, 0, 0, 1, 0, 10, 18, 0, 0, 26, 12, 6, 8, 42, 58, 
    14, 0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 4, 6, 
    0, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 6, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 
    22, 10, 0, 0, 10, 0, 0, 0, 1, 0, 5, 7, 4, 8, 0, 
    16, 17, 0, 0, 0, 0, 14, 1, 11, 1, 15, 2, 0, 4, 0, 
    14, 32, 0, 0, 0, 7, 16, 5, 1, 0, 6, 3, 6, 0, 0, 
    27, 32, 13, 6, 0, 4, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    26, 25, 28, 17, 12, 0, 1, 12, 0, 3, 17, 13, 0, 0, 0, 
    37, 20, 29, 7, 25, 13, 29, 50, 39, 24, 30, 38, 42, 44, 43, 
    74, 53, 32, 8, 55, 65, 58, 58, 62, 64, 70, 73, 76, 73, 77, 
    83, 59, 32, 30, 72, 65, 66, 62, 65, 68, 76, 77, 80, 86, 86, 
    96, 79, 46, 77, 65, 66, 65, 64, 70, 74, 81, 87, 88, 89, 95, 
    92, 87, 67, 78, 65, 68, 74, 70, 67, 71, 76, 77, 78, 90, 92, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 4, 14, 16, 0, 0, 
    5, 0, 0, 0, 0, 16, 30, 35, 0, 0, 0, 0, 0, 6, 0, 
    7, 0, 0, 0, 6, 6, 0, 0, 0, 0, 2, 0, 10, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 
    2, 0, 0, 11, 15, 0, 0, 0, 4, 0, 0, 13, 0, 0, 0, 
    0, 2, 12, 2, 0, 0, 0, 0, 0, 0, 12, 8, 5, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 9, 0, 0, 8, 18, 0, 0, 0, 
    0, 0, 10, 0, 0, 25, 22, 4, 0, 30, 7, 21, 7, 0, 0, 
    0, 0, 8, 1, 0, 0, 0, 0, 0, 0, 11, 5, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 17, 23, 
    0, 0, 0, 0, 30, 57, 41, 39, 16, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 2, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 8, 33, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=17
    39, 39, 38, 36, 37, 34, 44, 49, 35, 25, 27, 34, 33, 35, 32, 
    39, 42, 41, 39, 35, 3, 23, 28, 30, 0, 0, 0, 19, 30, 29, 
    18, 50, 42, 42, 42, 51, 15, 9, 0, 0, 0, 0, 0, 15, 31, 
    0, 9, 36, 38, 20, 10, 0, 0, 0, 7, 0, 0, 0, 0, 35, 
    0, 0, 21, 11, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 19, 
    0, 0, 19, 33, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 18, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 1, 0, 11, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 25, 0, 0, 0, 14, 0, 7, 10, 10, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 22, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 32, 10, 0, 0, 0, 25, 13, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 4, 29, 24, 31, 0, 3, 
    57, 0, 8, 0, 7, 0, 32, 10, 14, 0, 41, 4, 17, 12, 0, 
    60, 45, 22, 0, 72, 24, 42, 24, 15, 0, 38, 34, 15, 30, 0, 
    16, 47, 31, 0, 0, 4, 65, 32, 49, 0, 43, 26, 5, 21, 20, 
    17, 71, 10, 19, 0, 5, 48, 38, 48, 0, 50, 28, 8, 12, 27, 
    26, 68, 21, 37, 0, 6, 38, 12, 28, 0, 37, 30, 0, 10, 14, 
    47, 41, 44, 27, 3, 0, 23, 25, 11, 23, 0, 12, 0, 12, 8, 
    36, 34, 75, 11, 39, 0, 0, 66, 8, 0, 17, 0, 11, 5, 3, 
    27, 32, 68, 0, 119, 47, 9, 35, 45, 21, 13, 18, 14, 15, 16, 
    0, 20, 47, 25, 64, 18, 7, 6, 20, 13, 21, 19, 28, 28, 27, 
    40, 0, 0, 60, 36, 24, 25, 22, 21, 21, 25, 28, 29, 22, 35, 
    41, 30, 0, 84, 23, 21, 33, 23, 18, 22, 22, 24, 29, 22, 36, 
    44, 30, 21, 27, 15, 7, 14, 24, 25, 34, 32, 22, 25, 56, 55, 
    
    -- channel=20
    40, 33, 39, 36, 37, 36, 39, 40, 36, 28, 23, 28, 28, 32, 29, 
    38, 38, 41, 36, 42, 21, 31, 26, 13, 14, 2, 13, 25, 29, 28, 
    13, 35, 41, 37, 45, 29, 0, 10, 22, 26, 1, 0, 0, 33, 25, 
    0, 55, 36, 41, 20, 30, 3, 10, 5, 48, 0, 13, 0, 5, 43, 
    0, 25, 24, 68, 0, 32, 0, 0, 0, 59, 2, 0, 4, 0, 45, 
    10, 2, 17, 56, 16, 17, 0, 0, 0, 85, 0, 0, 13, 0, 5, 
    15, 0, 23, 0, 36, 34, 0, 0, 0, 62, 0, 0, 13, 13, 5, 
    14, 0, 24, 0, 50, 33, 0, 2, 0, 53, 0, 0, 19, 16, 16, 
    0, 0, 0, 4, 31, 18, 0, 0, 23, 9, 19, 0, 22, 22, 38, 
    0, 7, 0, 26, 0, 33, 26, 0, 31, 2, 0, 2, 21, 38, 24, 
    4, 9, 0, 69, 0, 6, 26, 0, 0, 0, 1, 2, 6, 0, 0, 
    19, 2, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=21
    9, 14, 12, 10, 10, 13, 12, 11, 9, 9, 11, 13, 14, 13, 12, 
    9, 15, 14, 11, 12, 12, 8, 13, 17, 7, 6, 8, 9, 8, 10, 
    10, 10, 9, 10, 10, 20, 0, 5, 8, 21, 5, 8, 11, 8, 13, 
    3, 12, 5, 12, 8, 9, 10, 8, 9, 20, 2, 11, 3, 5, 20, 
    0, 14, 2, 18, 16, 25, 8, 4, 10, 17, 5, 5, 11, 9, 18, 
    0, 0, 0, 19, 8, 4, 1, 7, 8, 27, 0, 0, 11, 10, 10, 
    0, 4, 0, 12, 32, 4, 4, 0, 4, 32, 0, 0, 8, 7, 4, 
    0, 0, 0, 2, 23, 18, 1, 6, 0, 27, 0, 0, 11, 11, 3, 
    0, 1, 0, 3, 1, 11, 0, 4, 4, 17, 0, 4, 13, 8, 13, 
    0, 0, 0, 19, 0, 14, 9, 8, 5, 4, 10, 13, 17, 19, 8, 
    2, 0, 0, 13, 0, 3, 21, 4, 0, 11, 3, 11, 7, 0, 0, 
    5, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 2, 0, 2, 4, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 1, 3, 0, 0, 2, 4, 0, 0, 0, 0, 1, 3, 
    6, 4, 0, 0, 1, 31, 0, 0, 0, 9, 13, 11, 0, 0, 0, 
    0, 0, 3, 4, 3, 0, 1, 12, 8, 9, 0, 0, 0, 0, 0, 
    5, 27, 1, 5, 2, 9, 9, 0, 0, 0, 0, 0, 1, 1, 0, 
    0, 10, 0, 0, 0, 0, 0, 3, 0, 20, 15, 0, 5, 1, 0, 
    0, 0, 0, 3, 0, 0, 15, 7, 12, 15, 0, 0, 0, 0, 9, 
    2, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 11, 12, 12, 0, 
    1, 4, 0, 0, 0, 0, 0, 0, 0, 3, 0, 11, 0, 0, 4, 
    0, 0, 2, 0, 4, 0, 17, 17, 0, 16, 0, 0, 1, 14, 5, 
    0, 0, 0, 20, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 18, 0, 0, 0, 0, 1, 17, 1, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 8, 7, 0, 0, 0, 0, 3, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 10, 0, 4, 14, 2, 0, 
    
    -- channel=23
    52, 50, 52, 52, 53, 43, 59, 67, 53, 32, 22, 27, 31, 43, 43, 
    52, 55, 56, 55, 51, 5, 43, 33, 16, 0, 0, 0, 3, 25, 37, 
    17, 32, 58, 59, 61, 44, 8, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 53, 52, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 38, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 33, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    7, 5, 2, 6, 7, 4, 7, 7, 10, 22, 18, 3, 0, 12, 12, 
    0, 5, 5, 10, 0, 0, 38, 22, 35, 0, 7, 19, 5, 0, 8, 
    45, 0, 3, 5, 7, 26, 19, 19, 0, 0, 23, 0, 37, 7, 0, 
    76, 0, 12, 0, 22, 0, 14, 22, 5, 0, 21, 22, 12, 22, 0, 
    32, 0, 35, 0, 0, 27, 40, 24, 25, 0, 8, 45, 0, 21, 11, 
    42, 0, 27, 38, 0, 0, 10, 25, 45, 0, 51, 33, 0, 9, 10, 
    15, 41, 0, 40, 0, 0, 28, 9, 50, 0, 41, 26, 0, 0, 20, 
    13, 2, 30, 14, 0, 0, 52, 12, 9, 0, 11, 35, 0, 8, 0, 
    16, 0, 58, 0, 27, 4, 6, 8, 0, 42, 11, 36, 0, 0, 0, 
    0, 0, 51, 0, 47, 6, 0, 12, 37, 16, 37, 2, 0, 0, 18, 
    0, 0, 55, 0, 14, 39, 0, 18, 38, 20, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 121, 15, 3, 2, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 49, 53, 0, 4, 0, 0, 0, 0, 0, 1, 0, 0, 
    4, 0, 0, 40, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 32, 
    15, 0, 0, 10, 11, 0, 0, 0, 0, 0, 9, 0, 0, 14, 23, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 3, 3, 0, 0, 5, 3, 1, 0, 0, 0, 0, 1, 0, 0, 
    3, 10, 7, 0, 8, 29, 0, 0, 0, 4, 0, 0, 0, 8, 0, 
    0, 17, 3, 0, 3, 15, 0, 0, 0, 46, 0, 0, 0, 4, 20, 
    0, 63, 3, 8, 0, 7, 0, 0, 0, 53, 0, 0, 0, 0, 51, 
    0, 59, 0, 46, 27, 0, 0, 0, 0, 56, 0, 0, 3, 0, 8, 
    0, 19, 0, 0, 45, 0, 0, 0, 0, 125, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 61, 24, 0, 0, 0, 107, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 36, 62, 0, 0, 0, 67, 0, 0, 16, 0, 0, 
    0, 2, 0, 33, 0, 0, 0, 0, 27, 0, 9, 0, 5, 27, 16, 
    0, 0, 0, 49, 0, 0, 19, 6, 0, 0, 0, 0, 45, 38, 0, 
    50, 0, 0, 118, 0, 0, 22, 0, 0, 0, 5, 9, 3, 0, 0, 
    37, 8, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 27, 32, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 6, 
    0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 30, 0, 0, 
    
    -- channel=28
    9, 21, 14, 16, 12, 13, 14, 19, 11, 5, 8, 12, 18, 10, 14, 
    15, 17, 13, 16, 15, 43, 0, 5, 10, 12, 0, 0, 0, 17, 15, 
    0, 36, 14, 19, 8, 7, 18, 0, 0, 7, 0, 16, 0, 0, 30, 
    7, 0, 8, 14, 6, 10, 9, 0, 1, 0, 26, 0, 17, 0, 8, 
    31, 0, 0, 0, 53, 0, 4, 0, 0, 0, 5, 0, 6, 14, 0, 
    0, 28, 13, 0, 40, 7, 46, 6, 12, 0, 0, 9, 1, 9, 0, 
    0, 17, 9, 31, 6, 6, 29, 17, 21, 0, 17, 0, 0, 3, 0, 
    0, 46, 0, 30, 0, 4, 16, 7, 30, 0, 29, 0, 0, 0, 24, 
    0, 9, 0, 36, 0, 0, 12, 1, 10, 0, 0, 15, 0, 26, 2, 
    30, 1, 29, 0, 0, 0, 9, 31, 0, 13, 25, 2, 11, 7, 11, 
    36, 0, 23, 0, 61, 0, 0, 29, 27, 0, 0, 0, 0, 0, 0, 
    0, 30, 27, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 83, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    13, 16, 12, 17, 16, 15, 17, 18, 16, 15, 13, 6, 13, 20, 19, 
    13, 19, 11, 20, 9, 11, 40, 20, 21, 0, 23, 19, 0, 1, 18, 
    22, 0, 16, 19, 10, 0, 31, 16, 0, 0, 22, 13, 36, 0, 0, 
    83, 0, 24, 10, 27, 0, 28, 20, 10, 0, 42, 7, 23, 19, 0, 
    68, 0, 48, 0, 39, 31, 48, 32, 19, 0, 25, 50, 5, 35, 0, 
    35, 0, 55, 4, 0, 6, 49, 37, 57, 0, 50, 44, 0, 21, 24, 
    32, 39, 13, 56, 0, 0, 25, 36, 58, 0, 58, 35, 0, 0, 27, 
    27, 37, 27, 45, 0, 0, 54, 6, 30, 0, 30, 40, 0, 1, 14, 
    34, 1, 66, 0, 23, 0, 21, 15, 0, 38, 0, 35, 0, 0, 7, 
    2, 0, 79, 0, 43, 0, 0, 41, 13, 1, 36, 2, 0, 0, 20, 
    0, 5, 73, 0, 91, 39, 0, 13, 48, 30, 0, 0, 0, 0, 7, 
    0, 0, 27, 0, 80, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 23, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 53, 9, 0, 5, 0, 0, 0, 0, 0, 0, 0, 2, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 29, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 13, 6, 3, 28, 25, 25, 0, 0, 
    45, 0, 0, 0, 0, 0, 12, 17, 15, 0, 32, 12, 27, 13, 0, 
    60, 3, 0, 0, 19, 14, 36, 27, 21, 0, 28, 32, 16, 27, 0, 
    46, 19, 0, 0, 0, 21, 38, 32, 37, 0, 38, 39, 12, 26, 21, 
    48, 39, 0, 0, 0, 0, 29, 30, 43, 0, 51, 33, 16, 15, 20, 
    42, 56, 22, 14, 0, 0, 44, 20, 28, 0, 32, 36, 10, 8, 0, 
    52, 42, 53, 11, 5, 16, 26, 18, 7, 17, 2, 31, 4, 0, 0, 
    35, 34, 67, 17, 39, 6, 11, 39, 14, 7, 31, 21, 0, 0, 0, 
    21, 34, 67, 0, 72, 39, 8, 44, 53, 43, 36, 33, 32, 31, 37, 
    31, 33, 49, 0, 77, 68, 51, 53, 55, 49, 51, 54, 59, 57, 62, 
    67, 26, 14, 39, 92, 54, 55, 53, 53, 53, 57, 59, 59, 62, 65, 
    78, 59, 1, 78, 57, 53, 60, 54, 53, 56, 60, 62, 68, 58, 68, 
    78, 64, 52, 64, 52, 45, 50, 53, 52, 61, 64, 59, 53, 77, 84, 
    
    -- channel=32
    4, 2, 5, 0, 0, 4, 2, 0, 0, 0, 0, 6, 2, 0, 0, 
    3, 4, 7, 0, 10, 3, 0, 0, 0, 12, 0, 0, 6, 17, 0, 
    0, 46, 3, 0, 6, 16, 0, 0, 7, 50, 0, 0, 0, 19, 23, 
    0, 68, 0, 9, 0, 19, 0, 0, 0, 82, 0, 0, 0, 0, 71, 
    0, 27, 0, 80, 0, 0, 0, 0, 0, 104, 0, 0, 0, 0, 27, 
    0, 13, 0, 0, 80, 4, 0, 0, 0, 166, 0, 0, 14, 0, 0, 
    0, 0, 4, 0, 73, 47, 0, 0, 0, 133, 0, 0, 4, 14, 0, 
    0, 0, 0, 0, 54, 65, 0, 0, 0, 84, 0, 0, 27, 4, 0, 
    0, 1, 0, 36, 0, 23, 0, 0, 35, 0, 15, 0, 25, 33, 13, 
    0, 4, 0, 63, 0, 0, 42, 0, 0, 0, 0, 2, 40, 31, 0, 
    59, 0, 0, 143, 0, 0, 39, 0, 0, 0, 0, 5, 9, 8, 0, 
    69, 46, 0, 91, 0, 0, 3, 1, 0, 0, 0, 3, 1, 0, 0, 
    0, 66, 95, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 3, 7, 
    0, 2, 125, 0, 0, 4, 0, 0, 3, 1, 0, 1, 0, 17, 0, 
    0, 1, 8, 0, 0, 15, 8, 0, 5, 0, 0, 6, 36, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 10, 12, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 4, 8, 0, 23, 5, 16, 6, 0, 
    29, 0, 0, 0, 0, 0, 18, 15, 16, 0, 5, 16, 3, 13, 0, 
    31, 11, 0, 0, 0, 0, 19, 10, 27, 0, 29, 24, 0, 10, 3, 
    25, 36, 0, 0, 0, 0, 12, 16, 26, 0, 34, 19, 4, 0, 13, 
    21, 30, 0, 0, 0, 0, 42, 13, 18, 0, 23, 25, 0, 9, 1, 
    32, 18, 45, 0, 0, 5, 10, 7, 0, 6, 0, 26, 0, 0, 0, 
    27, 23, 52, 0, 17, 0, 0, 16, 12, 1, 22, 0, 0, 0, 0, 
    2, 16, 52, 0, 41, 8, 0, 25, 31, 15, 6, 5, 7, 0, 2, 
    20, 14, 22, 0, 76, 55, 35, 34, 36, 30, 35, 39, 44, 47, 50, 
    61, 20, 0, 39, 72, 38, 40, 38, 41, 40, 42, 43, 48, 45, 45, 
    67, 44, 0, 73, 45, 38, 45, 39, 38, 42, 51, 53, 55, 45, 72, 
    71, 52, 45, 47, 46, 39, 42, 41, 37, 46, 54, 48, 35, 68, 72, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 28, 13, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 24, 16, 6, 0, 5, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 28, 0, 0, 0, 0, 0, 36, 11, 0, 0, 
    5, 0, 0, 0, 0, 2, 0, 0, 0, 22, 32, 9, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 22, 17, 0, 0, 0, 0, 5, 10, 
    32, 30, 0, 0, 34, 76, 39, 39, 29, 17, 15, 16, 14, 10, 16, 
    14, 28, 15, 0, 71, 13, 13, 14, 12, 9, 7, 2, 13, 22, 4, 
    24, 16, 18, 49, 31, 10, 8, 9, 15, 12, 19, 26, 26, 6, 38, 
    22, 20, 22, 40, 28, 29, 32, 20, 3, 0, 10, 17, 0, 0, 23, 
    
    -- channel=37
    10, 16, 13, 13, 10, 16, 14, 13, 14, 16, 16, 15, 13, 7, 5, 
    9, 16, 15, 14, 14, 23, 12, 23, 20, 9, 0, 0, 4, 8, 6, 
    21, 16, 13, 13, 13, 30, 14, 0, 0, 11, 7, 0, 0, 0, 7, 
    0, 0, 8, 16, 19, 12, 11, 0, 0, 15, 11, 6, 0, 0, 1, 
    5, 6, 5, 24, 38, 22, 20, 3, 0, 3, 12, 0, 0, 0, 0, 
    16, 24, 9, 26, 57, 41, 27, 3, 0, 22, 26, 4, 1, 0, 0, 
    13, 22, 12, 15, 24, 34, 42, 15, 0, 27, 17, 0, 0, 0, 0, 
    28, 24, 0, 9, 9, 52, 28, 18, 3, 20, 19, 0, 1, 6, 0, 
    35, 37, 7, 17, 12, 17, 6, 6, 0, 1, 20, 1, 0, 0, 3, 
    41, 32, 12, 12, 14, 9, 13, 15, 1, 23, 1, 0, 0, 10, 15, 
    42, 35, 13, 33, 18, 8, 39, 44, 15, 0, 0, 0, 0, 4, 3, 
    21, 40, 20, 52, 52, 11, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 31, 60, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    18, 5, 0, 0, 5, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 
    2, 18, 0, 0, 0, 0, 16, 0, 7, 0, 9, 0, 0, 0, 0, 
    5, 11, 0, 0, 0, 17, 28, 6, 0, 0, 0, 0, 0, 4, 0, 
    17, 19, 14, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    14, 14, 21, 0, 16, 0, 0, 0, 0, 15, 18, 1, 0, 0, 0, 
    16, 8, 20, 0, 0, 10, 35, 49, 37, 7, 7, 19, 27, 32, 32, 
    67, 34, 14, 0, 67, 46, 37, 37, 42, 47, 50, 51, 51, 49, 53, 
    63, 50, 3, 41, 56, 44, 47, 43, 42, 44, 48, 51, 61, 61, 52, 
    69, 55, 43, 73, 46, 43, 42, 44, 48, 52, 59, 65, 60, 62, 88, 
    70, 61, 50, 55, 49, 52, 58, 48, 44, 44, 54, 49, 41, 66, 67, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    23, 21, 23, 26, 26, 20, 22, 26, 27, 22, 17, 15, 20, 23, 27, 
    25, 23, 24, 26, 27, 13, 27, 15, 17, 11, 13, 7, 3, 15, 24, 
    8, 15, 23, 26, 23, 8, 16, 16, 13, 2, 12, 21, 18, 7, 13, 
    31, 0, 22, 24, 16, 22, 15, 19, 14, 0, 17, 6, 17, 11, 5, 
    41, 0, 30, 30, 23, 18, 12, 13, 9, 0, 14, 22, 13, 24, 1, 
    17, 0, 29, 0, 0, 7, 10, 24, 20, 0, 13, 22, 10, 23, 20, 
    24, 0, 10, 31, 0, 0, 5, 18, 26, 0, 19, 15, 8, 10, 18, 
    7, 12, 18, 26, 16, 0, 21, 3, 20, 0, 12, 14, 5, 5, 24, 
    7, 0, 13, 0, 7, 2, 11, 5, 13, 11, 0, 19, 2, 12, 17, 
    0, 0, 21, 0, 13, 11, 11, 14, 2, 9, 22, 17, 6, 10, 24, 
    0, 0, 18, 0, 34, 20, 0, 2, 21, 21, 12, 10, 0, 0, 4, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 5, 3, 1, 0, 0, 2, 
    2, 0, 0, 0, 26, 3, 4, 3, 6, 5, 4, 2, 0, 3, 3, 
    6, 0, 0, 0, 13, 4, 6, 2, 3, 1, 0, 0, 3, 0, 0, 
    6, 0, 0, 0, 5, 0, 2, 8, 5, 3, 4, 5, 2, 3, 15, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 0, 1, 41, 10, 0, 0, 0, 16, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 7, 9, 0, 0, 
    24, 19, 3, 0, 3, 0, 31, 9, 1, 0, 0, 0, 0, 0, 0, 
    26, 55, 9, 3, 94, 45, 3, 1, 0, 0, 19, 16, 8, 16, 0, 
    0, 1, 6, 0, 0, 0, 22, 14, 20, 22, 0, 0, 0, 8, 19, 
    0, 0, 0, 4, 0, 5, 4, 7, 10, 5, 0, 0, 0, 8, 14, 
    0, 15, 5, 24, 2, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 1, 0, 0, 6, 6, 0, 0, 0, 0, 0, 15, 
    0, 0, 5, 0, 8, 0, 0, 48, 0, 0, 0, 0, 20, 19, 0, 
    0, 0, 0, 32, 92, 71, 22, 0, 0, 0, 16, 35, 8, 0, 0, 
    0, 0, 14, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 20, 17, 0, 
    
    -- channel=42
    95, 97, 100, 100, 99, 93, 103, 107, 99, 82, 67, 70, 77, 87, 83, 
    98, 102, 105, 103, 100, 105, 95, 87, 57, 35, 31, 33, 43, 64, 81, 
    68, 68, 102, 103, 107, 86, 47, 23, 26, 43, 34, 24, 31, 36, 67, 
    25, 63, 95, 102, 89, 55, 53, 33, 26, 45, 34, 34, 12, 20, 55, 
    14, 72, 86, 85, 81, 77, 41, 27, 19, 36, 43, 33, 27, 18, 40, 
    17, 47, 78, 90, 42, 46, 51, 35, 23, 68, 45, 13, 28, 20, 22, 
    16, 47, 50, 70, 66, 64, 54, 37, 20, 67, 23, 21, 24, 27, 35, 
    31, 25, 41, 48, 66, 76, 33, 33, 20, 74, 33, 17, 24, 37, 49, 
    32, 35, 17, 38, 51, 26, 26, 36, 34, 52, 34, 6, 19, 49, 92, 
    34, 40, 12, 32, 25, 38, 33, 44, 43, 32, 8, 0, 36, 86, 81, 
    30, 40, 10, 60, 49, 43, 53, 21, 5, 0, 0, 0, 4, 0, 0, 
    0, 10, 23, 95, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 4, 4, 0, 0, 1, 5, 4, 0, 0, 0, 8, 10, 
    0, 0, 0, 5, 0, 0, 34, 6, 4, 0, 24, 23, 0, 0, 6, 
    18, 0, 0, 3, 0, 0, 25, 15, 0, 0, 28, 14, 43, 0, 0, 
    94, 0, 8, 0, 20, 0, 26, 28, 12, 0, 42, 9, 24, 27, 0, 
    70, 0, 43, 0, 19, 37, 49, 40, 25, 0, 25, 60, 7, 40, 0, 
    54, 0, 47, 14, 0, 0, 43, 40, 69, 0, 59, 50, 0, 24, 31, 
    49, 40, 0, 46, 0, 0, 12, 37, 61, 0, 61, 46, 3, 0, 34, 
    40, 29, 40, 31, 0, 0, 61, 1, 27, 0, 28, 50, 0, 0, 7, 
    44, 0, 91, 0, 39, 0, 17, 20, 0, 43, 0, 38, 0, 0, 0, 
    0, 0, 89, 0, 45, 6, 0, 36, 34, 0, 33, 0, 0, 0, 9, 
    0, 4, 81, 0, 98, 56, 0, 0, 47, 38, 10, 4, 0, 0, 14, 
    0, 0, 20, 0, 91, 27, 0, 0, 9, 5, 3, 2, 3, 6, 13, 
    32, 0, 0, 27, 80, 7, 13, 8, 10, 6, 2, 6, 7, 0, 0, 
    29, 7, 0, 44, 23, 3, 23, 12, 0, 3, 7, 1, 10, 0, 23, 
    41, 5, 4, 0, 18, 0, 0, 3, 2, 13, 24, 2, 0, 38, 51, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 32, 12, 7, 2, 16, 0, 
    0, 36, 0, 0, 0, 0, 0, 7, 19, 45, 0, 14, 4, 13, 21, 
    0, 29, 0, 0, 0, 0, 0, 0, 13, 45, 0, 0, 14, 0, 27, 
    6, 29, 0, 0, 35, 0, 0, 0, 0, 82, 0, 0, 21, 5, 6, 
    0, 14, 0, 0, 26, 22, 0, 0, 0, 74, 0, 0, 21, 22, 8, 
    8, 0, 0, 0, 13, 42, 0, 13, 0, 50, 0, 0, 28, 26, 0, 
    5, 25, 0, 25, 9, 13, 0, 8, 19, 0, 22, 0, 31, 12, 0, 
    18, 28, 0, 41, 0, 18, 14, 0, 22, 12, 0, 14, 31, 4, 0, 
    53, 20, 0, 72, 0, 7, 57, 22, 1, 5, 30, 43, 50, 42, 30, 
    95, 54, 3, 65, 0, 29, 51, 50, 48, 56, 64, 66, 68, 69, 63, 
    75, 92, 62, 31, 0, 56, 56, 58, 58, 65, 68, 71, 71, 70, 73, 
    69, 73, 115, 14, 41, 61, 53, 58, 63, 67, 74, 77, 71, 89, 84, 
    67, 76, 80, 46, 59, 74, 69, 60, 63, 62, 64, 70, 79, 67, 53, 
    
    -- channel=45
    0, 0, 0, 2, 3, 0, 0, 1, 5, 5, 4, 0, 0, 5, 7, 
    0, 0, 0, 3, 0, 0, 30, 7, 11, 0, 8, 12, 0, 0, 2, 
    20, 0, 0, 1, 0, 0, 35, 13, 1, 0, 18, 8, 29, 0, 0, 
    63, 0, 3, 0, 15, 0, 3, 28, 8, 0, 37, 9, 24, 27, 0, 
    61, 0, 41, 0, 0, 25, 37, 39, 19, 0, 5, 52, 0, 27, 0, 
    77, 0, 54, 34, 0, 22, 24, 26, 42, 0, 59, 58, 0, 16, 24, 
    78, 11, 10, 35, 0, 0, 0, 35, 42, 0, 61, 42, 0, 0, 26, 
    65, 2, 47, 10, 0, 0, 68, 9, 25, 0, 33, 44, 0, 0, 12, 
    51, 0, 104, 0, 47, 0, 17, 5, 0, 21, 0, 49, 0, 0, 0, 
    2, 0, 79, 0, 41, 27, 0, 0, 36, 10, 37, 0, 0, 0, 11, 
    0, 4, 68, 0, 68, 37, 0, 5, 55, 29, 0, 0, 0, 0, 9, 
    0, 0, 19, 0, 92, 57, 0, 2, 13, 0, 0, 0, 0, 0, 9, 
    23, 0, 0, 3, 104, 3, 6, 3, 3, 0, 0, 0, 0, 0, 0, 
    23, 1, 0, 27, 31, 0, 14, 5, 0, 0, 1, 0, 6, 0, 18, 
    33, 0, 4, 0, 16, 0, 0, 1, 0, 0, 14, 0, 0, 14, 41, 
    
    -- channel=46
    12, 9, 10, 12, 14, 10, 9, 15, 16, 13, 10, 7, 8, 9, 13, 
    14, 10, 10, 13, 12, 1, 9, 8, 15, 9, 4, 1, 1, 10, 13, 
    4, 14, 14, 14, 13, 4, 13, 13, 1, 0, 0, 0, 0, 2, 6, 
    10, 0, 12, 14, 10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    28, 29, 26, 30, 30, 23, 31, 33, 30, 35, 40, 32, 30, 30, 29, 
    29, 23, 23, 33, 21, 10, 45, 37, 48, 11, 23, 22, 20, 28, 31, 
    49, 34, 28, 32, 21, 18, 62, 32, 1, 0, 23, 28, 40, 12, 21, 
    74, 0, 34, 23, 38, 12, 18, 22, 21, 0, 61, 14, 39, 30, 0, 
    78, 0, 60, 0, 26, 8, 51, 38, 31, 0, 19, 46, 10, 40, 0, 
    51, 25, 74, 0, 0, 36, 54, 34, 51, 0, 67, 69, 4, 30, 23, 
    45, 50, 53, 59, 0, 0, 46, 52, 63, 0, 80, 39, 5, 0, 31, 
    36, 50, 39, 54, 0, 0, 98, 36, 51, 0, 55, 46, 0, 14, 37, 
    48, 15, 77, 8, 17, 21, 36, 12, 6, 31, 0, 73, 0, 4, 7, 
    34, 13, 94, 0, 51, 17, 0, 24, 12, 41, 76, 16, 0, 0, 44, 
    0, 17, 90, 0, 85, 13, 0, 61, 92, 43, 0, 0, 0, 23, 39, 
    0, 18, 49, 0, 113, 76, 10, 11, 25, 6, 5, 0, 0, 0, 7, 
    20, 0, 0, 32, 121, 7, 9, 6, 4, 0, 0, 0, 7, 6, 0, 
    26, 4, 0, 121, 40, 0, 13, 1, 0, 0, 0, 4, 11, 0, 28, 
    29, 0, 0, 30, 17, 0, 10, 12, 0, 0, 7, 0, 0, 8, 49, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 44, 2, 0, 0, 1, 21, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 
    9, 36, 0, 0, 1, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 37, 0, 0, 50, 21, 0, 0, 0, 8, 13, 6, 3, 8, 0, 
    0, 0, 0, 0, 0, 0, 14, 4, 13, 29, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 3, 0, 10, 4, 
    2, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 11, 1, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 4, 0, 0, 2, 26, 0, 0, 0, 0, 7, 8, 0, 
    0, 0, 0, 42, 74, 45, 0, 0, 0, 0, 26, 31, 7, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 0, 22, 5, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 3, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 0, 2, 0, 0, 0, 
    0, 33, 0, 0, 0, 0, 8, 0, 0, 15, 0, 0, 0, 0, 0, 
    1, 40, 0, 28, 37, 19, 0, 0, 0, 48, 13, 0, 6, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 90, 0, 0, 3, 0, 10, 
    6, 0, 0, 0, 11, 33, 0, 0, 0, 55, 0, 0, 7, 22, 0, 
    9, 0, 0, 0, 26, 18, 0, 0, 0, 22, 0, 0, 10, 0, 0, 
    2, 9, 0, 15, 0, 0, 0, 4, 18, 0, 0, 0, 0, 8, 0, 
    0, 7, 0, 40, 0, 0, 22, 18, 0, 0, 0, 0, 25, 0, 0, 
    20, 4, 0, 103, 32, 39, 20, 0, 0, 0, 31, 42, 23, 0, 0, 
    0, 0, 7, 59, 0, 0, 0, 0, 4, 12, 17, 18, 27, 24, 19, 
    14, 2, 37, 0, 0, 19, 14, 15, 18, 26, 33, 34, 16, 19, 42, 
    13, 22, 29, 0, 0, 22, 19, 19, 21, 24, 19, 14, 17, 45, 0, 
    8, 26, 15, 0, 0, 10, 4, 15, 32, 32, 19, 27, 63, 28, 4, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 2, 6, 4, 10, 5, 1, 0, 0, 
    7, 0, 0, 0, 0, 9, 10, 8, 0, 3, 19, 15, 10, 0, 0, 
    24, 0, 0, 0, 0, 1, 12, 7, 4, 3, 24, 9, 9, 0, 0, 
    40, 11, 0, 0, 38, 21, 33, 14, 7, 0, 23, 16, 5, 7, 0, 
    35, 32, 7, 0, 34, 34, 34, 20, 12, 0, 37, 24, 7, 10, 2, 
    34, 37, 11, 1, 7, 12, 44, 24, 26, 0, 39, 15, 3, 5, 6, 
    38, 46, 20, 11, 0, 26, 43, 21, 16, 0, 27, 18, 6, 7, 0, 
    49, 43, 31, 19, 2, 19, 17, 9, 10, 6, 10, 19, 0, 0, 0, 
    41, 37, 44, 15, 34, 8, 14, 27, 11, 17, 20, 3, 0, 0, 0, 
    31, 37, 45, 8, 51, 27, 25, 51, 43, 15, 7, 8, 16, 21, 21, 
    31, 39, 42, 24, 69, 40, 25, 24, 24, 16, 17, 19, 20, 20, 23, 
    23, 20, 25, 50, 58, 21, 21, 17, 15, 14, 18, 21, 26, 27, 27, 
    29, 22, 15, 65, 25, 20, 20, 18, 18, 20, 21, 24, 24, 21, 32, 
    29, 23, 16, 33, 15, 14, 20, 20, 18, 21, 22, 18, 17, 33, 32, 
    
    -- channel=51
    7, 7, 9, 11, 11, 7, 6, 4, 11, 11, 2, 0, 3, 5, 7, 
    8, 5, 9, 11, 11, 44, 17, 12, 0, 7, 27, 13, 0, 0, 8, 
    16, 0, 7, 7, 10, 1, 1, 0, 5, 31, 35, 25, 29, 0, 0, 
    30, 20, 6, 9, 22, 6, 38, 28, 24, 10, 29, 14, 8, 9, 0, 
    36, 56, 18, 13, 76, 61, 31, 24, 15, 4, 32, 31, 22, 21, 2, 
    31, 38, 13, 25, 0, 8, 44, 25, 32, 39, 46, 11, 15, 24, 19, 
    29, 53, 0, 12, 14, 37, 42, 35, 23, 43, 25, 22, 16, 23, 25, 
    43, 39, 30, 14, 24, 52, 37, 13, 7, 36, 27, 15, 12, 18, 2, 
    56, 45, 41, 20, 38, 0, 0, 33, 14, 22, 0, 0, 0, 6, 25, 
    41, 45, 41, 28, 23, 24, 14, 53, 34, 10, 6, 0, 12, 22, 10, 
    33, 41, 30, 53, 101, 73, 70, 37, 30, 21, 21, 43, 44, 30, 27, 
    20, 26, 34, 90, 46, 0, 1, 0, 15, 29, 35, 35, 37, 41, 37, 
    52, 20, 20, 79, 3, 33, 33, 29, 31, 36, 41, 48, 46, 39, 50, 
    44, 38, 26, 40, 29, 36, 38, 32, 33, 39, 42, 36, 37, 54, 46, 
    49, 40, 35, 0, 25, 23, 27, 34, 44, 47, 42, 34, 53, 71, 40, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 4, 0, 0, 
    0, 4, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 10, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    2, 1, 0, 0, 0, 0, 0, 0, 0, 4, 13, 14, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 15, 0, 0, 20, 18, 0, 
    6, 51, 0, 0, 1, 52, 16, 23, 1, 5, 0, 0, 0, 18, 14, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 42, 0, 5, 2, 0, 39, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 9, 
    0, 3, 0, 13, 109, 21, 0, 0, 0, 35, 0, 0, 8, 0, 0, 
    0, 0, 21, 0, 46, 7, 0, 0, 0, 39, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 18, 0, 27, 0, 32, 0, 0, 16, 4, 0, 
    0, 0, 0, 15, 0, 58, 11, 0, 4, 0, 44, 19, 29, 10, 0, 
    17, 3, 0, 17, 0, 0, 14, 0, 0, 31, 12, 13, 0, 0, 0, 
    45, 0, 0, 20, 0, 0, 0, 17, 0, 0, 0, 0, 0, 19, 13, 
    78, 50, 0, 0, 9, 64, 54, 52, 23, 9, 4, 7, 1, 0, 0, 
    0, 62, 51, 0, 27, 0, 0, 2, 1, 0, 0, 0, 0, 10, 0, 
    0, 0, 76, 31, 8, 1, 0, 0, 4, 0, 5, 17, 8, 1, 12, 
    0, 3, 11, 59, 15, 31, 25, 2, 0, 0, 0, 5, 0, 0, 0, 
    
    -- channel=54
    20, 20, 20, 23, 21, 19, 24, 21, 18, 19, 15, 12, 15, 17, 13, 
    19, 20, 21, 25, 20, 30, 35, 22, 12, 0, 14, 9, 1, 6, 17, 
    22, 3, 22, 21, 21, 21, 9, 0, 0, 11, 33, 18, 21, 0, 8, 
    32, 2, 27, 18, 25, 5, 32, 20, 14, 9, 34, 15, 4, 0, 0, 
    41, 47, 42, 7, 71, 64, 44, 20, 9, 0, 34, 32, 10, 11, 0, 
    43, 43, 46, 20, 3, 27, 46, 27, 24, 0, 61, 20, 9, 14, 7, 
    37, 57, 16, 24, 7, 22, 59, 40, 29, 16, 44, 19, 5, 9, 24, 
    48, 47, 33, 32, 14, 51, 60, 20, 17, 20, 31, 18, 3, 25, 12, 
    57, 50, 46, 14, 37, 6, 10, 18, 10, 31, 4, 9, 0, 1, 23, 
    45, 49, 50, 11, 41, 18, 6, 49, 34, 17, 13, 0, 4, 24, 23, 
    28, 49, 48, 15, 86, 60, 54, 52, 39, 10, 0, 8, 10, 13, 10, 
    19, 29, 48, 69, 82, 0, 0, 0, 0, 5, 9, 9, 11, 16, 15, 
    25, 13, 13, 88, 21, 10, 13, 8, 7, 8, 10, 17, 23, 15, 18, 
    19, 12, 13, 59, 13, 12, 14, 10, 8, 12, 14, 13, 10, 14, 36, 
    28, 10, 11, 4, 7, 1, 8, 11, 15, 18, 19, 8, 15, 43, 22, 
    
    -- channel=55
    26, 25, 25, 25, 25, 23, 31, 34, 27, 22, 21, 23, 21, 24, 23, 
    25, 31, 26, 27, 21, 0, 25, 28, 22, 0, 0, 2, 17, 20, 22, 
    26, 25, 31, 29, 30, 24, 13, 12, 0, 0, 0, 0, 0, 10, 15, 
    0, 0, 30, 26, 24, 1, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 13, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    54, 55, 55, 60, 61, 52, 59, 65, 65, 57, 47, 40, 46, 55, 57, 
    57, 58, 56, 63, 53, 44, 76, 61, 57, 17, 31, 29, 20, 31, 53, 
    58, 18, 60, 63, 60, 29, 63, 31, 14, 0, 22, 11, 40, 11, 24, 
    77, 0, 59, 56, 70, 26, 38, 32, 18, 0, 45, 19, 28, 28, 0, 
    57, 0, 76, 2, 35, 44, 46, 39, 24, 0, 24, 53, 9, 34, 6, 
    43, 0, 77, 68, 0, 24, 48, 35, 50, 0, 56, 47, 0, 22, 26, 
    38, 34, 30, 82, 0, 0, 26, 43, 47, 0, 56, 38, 6, 0, 29, 
    38, 16, 38, 50, 4, 0, 56, 15, 30, 0, 40, 40, 0, 8, 27, 
    36, 0, 72, 0, 52, 1, 27, 25, 0, 51, 2, 39, 0, 0, 38, 
    9, 0, 66, 0, 35, 19, 0, 30, 25, 19, 38, 4, 0, 19, 57, 
    0, 8, 59, 0, 77, 35, 0, 6, 40, 27, 0, 0, 0, 0, 14, 
    0, 0, 15, 0, 78, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 5, 1, 0, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 1, 40, 44, 30, 15, 5, 0, 
    4, 12, 0, 0, 0, 0, 18, 17, 23, 50, 30, 28, 19, 6, 7, 
    27, 51, 0, 0, 34, 28, 36, 20, 22, 26, 37, 16, 24, 9, 4, 
    46, 71, 0, 0, 78, 37, 40, 24, 16, 56, 47, 20, 32, 20, 5, 
    40, 70, 8, 0, 41, 41, 65, 32, 25, 74, 41, 23, 26, 31, 22, 
    50, 68, 17, 3, 20, 81, 50, 42, 25, 61, 39, 27, 33, 40, 12, 
    66, 82, 34, 46, 17, 41, 28, 30, 29, 17, 40, 17, 24, 18, 0, 
    78, 83, 45, 60, 39, 18, 31, 50, 36, 30, 15, 8, 20, 9, 0, 
    89, 73, 50, 86, 50, 41, 73, 76, 37, 16, 26, 33, 46, 44, 32, 
    109, 88, 60, 109, 93, 61, 68, 66, 58, 58, 66, 72, 78, 82, 79, 
    83, 95, 76, 110, 56, 66, 66, 65, 65, 69, 76, 81, 85, 83, 90, 
    88, 76, 103, 99, 58, 72, 66, 66, 69, 76, 84, 90, 82, 96, 103, 
    89, 85, 77, 86, 64, 74, 76, 69, 72, 78, 80, 79, 91, 103, 77, 
    
    -- channel=58
    8, 12, 4, 6, 7, 6, 9, 11, 9, 16, 22, 18, 9, 6, 6, 
    3, 7, 4, 9, 1, 0, 6, 19, 38, 1, 0, 4, 16, 10, 5, 
    34, 25, 7, 9, 6, 61, 37, 26, 0, 0, 0, 0, 4, 4, 8, 
    12, 0, 8, 6, 17, 0, 0, 0, 0, 0, 23, 11, 15, 0, 1, 
    0, 0, 10, 0, 0, 0, 22, 4, 18, 0, 0, 0, 0, 0, 0, 
    5, 12, 12, 18, 56, 19, 12, 0, 9, 0, 27, 25, 0, 0, 0, 
    0, 41, 21, 28, 15, 0, 33, 8, 18, 0, 32, 3, 0, 0, 0, 
    0, 24, 0, 11, 0, 0, 58, 36, 13, 0, 24, 18, 0, 9, 4, 
    7, 12, 11, 0, 0, 46, 20, 2, 0, 34, 19, 48, 6, 0, 0, 
    27, 12, 28, 0, 6, 0, 0, 0, 0, 31, 46, 1, 0, 0, 17, 
    17, 12, 41, 0, 0, 0, 0, 47, 23, 11, 0, 0, 0, 14, 13, 
    36, 26, 0, 0, 105, 62, 39, 34, 8, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 56, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 105, 6, 0, 0, 0, 0, 0, 0, 2, 0, 0, 27, 
    0, 0, 0, 55, 10, 3, 6, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 10, 6, 0, 0, 0, 12, 20, 7, 0, 0, 0, 14, 7, 6, 
    49, 23, 3, 0, 49, 43, 35, 36, 31, 28, 30, 35, 37, 40, 40, 
    49, 45, 16, 26, 43, 30, 31, 29, 29, 31, 35, 39, 44, 45, 41, 
    54, 42, 51, 31, 28, 32, 30, 31, 33, 37, 46, 50, 47, 51, 64, 
    54, 48, 45, 34, 33, 38, 39, 31, 30, 34, 42, 40, 36, 51, 47, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 
    9, 0, 0, 0, 0, 18, 6, 10, 0, 5, 21, 12, 3, 3, 0, 
    1, 0, 0, 0, 0, 0, 0, 9, 8, 18, 17, 19, 14, 6, 0, 
    6, 0, 0, 0, 0, 4, 23, 17, 19, 1, 8, 8, 7, 0, 7, 
    43, 24, 0, 19, 55, 34, 12, 9, 5, 0, 34, 24, 13, 7, 0, 
    35, 29, 1, 0, 17, 10, 27, 13, 13, 13, 28, 16, 11, 5, 6, 
    37, 24, 7, 0, 0, 28, 50, 33, 15, 21, 25, 22, 15, 20, 0, 
    42, 37, 35, 5, 13, 35, 16, 11, 0, 6, 29, 32, 20, 0, 0, 
    44, 41, 28, 16, 23, 23, 9, 0, 28, 29, 22, 7, 0, 0, 0, 
    28, 35, 34, 13, 0, 3, 28, 47, 27, 10, 5, 3, 18, 19, 17, 
    64, 43, 19, 23, 79, 65, 54, 53, 40, 33, 33, 38, 38, 39, 41, 
    41, 58, 32, 58, 72, 35, 36, 34, 32, 31, 33, 36, 42, 43, 37, 
    46, 38, 63, 63, 38, 36, 32, 35, 36, 39, 46, 49, 43, 45, 63, 
    48, 44, 43, 53, 40, 45, 44, 34, 31, 35, 41, 39, 29, 47, 39, 
    
    -- channel=61
    99, 105, 103, 105, 103, 99, 108, 116, 105, 85, 72, 76, 85, 92, 92, 
    101, 111, 109, 109, 106, 94, 95, 88, 72, 40, 26, 27, 41, 72, 88, 
    63, 79, 107, 111, 109, 96, 59, 38, 25, 27, 25, 23, 25, 32, 74, 
    39, 35, 102, 107, 89, 65, 50, 25, 18, 31, 34, 28, 20, 14, 54, 
    29, 39, 89, 85, 74, 50, 42, 23, 16, 18, 41, 30, 23, 21, 21, 
    4, 28, 85, 64, 43, 45, 48, 40, 24, 19, 32, 22, 24, 20, 16, 
    6, 26, 59, 92, 53, 38, 53, 33, 34, 24, 31, 19, 15, 20, 28, 
    7, 32, 20, 65, 55, 48, 29, 28, 33, 42, 34, 22, 17, 29, 57, 
    11, 17, 1, 31, 27, 34, 38, 27, 29, 48, 35, 20, 16, 50, 81, 
    24, 20, 17, 13, 27, 14, 27, 43, 13, 33, 19, 10, 24, 70, 83, 
    14, 22, 20, 15, 31, 14, 5, 13, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 34, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    1, 0, 0, 0, 2, 0, 5, 0, 0, 5, 0, 0, 1, 3, 0, 
    0, 4, 0, 0, 0, 0, 4, 2, 26, 0, 0, 3, 0, 10, 0, 
    0, 11, 0, 0, 0, 19, 0, 15, 0, 0, 0, 0, 0, 4, 0, 
    12, 0, 11, 53, 0, 22, 0, 3, 0, 52, 0, 0, 0, 0, 20, 
    65, 0, 26, 19, 0, 45, 0, 0, 0, 21, 0, 16, 0, 0, 15, 
    98, 0, 25, 0, 0, 21, 0, 10, 0, 0, 0, 4, 2, 0, 0, 
    73, 0, 49, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    24, 0, 41, 0, 37, 0, 0, 0, 15, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 56, 36, 0, 20, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 24, 0, 10, 0, 0, 6, 0, 9, 10, 2, 0, 5, 
    0, 3, 17, 0, 0, 28, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 76, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 36, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 4, 7, 0, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 13, 15, 15, 2, 0, 
    0, 7, 0, 0, 0, 6, 22, 41, 7, 1, 0, 0, 0, 2, 0, 
    2, 13, 0, 2, 0, 29, 0, 0, 0, 0, 0, 0, 8, 0, 5, 
    6, 0, 0, 13, 0, 0, 0, 0, 0, 25, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 2, 0, 0, 0, 8, 0, 0, 0, 
    10, 0, 10, 0, 0, 0, 0, 1, 0, 0, 7, 5, 11, 0, 0, 
    0, 9, 5, 12, 0, 0, 0, 0, 0, 0, 3, 10, 0, 0, 3, 
    0, 0, 0, 0, 0, 25, 22, 0, 4, 33, 0, 10, 6, 1, 0, 
    0, 0, 0, 24, 0, 0, 30, 0, 0, 0, 5, 10, 0, 0, 0, 
    4, 0, 11, 0, 0, 0, 0, 0, 0, 28, 15, 0, 0, 26, 28, 
    0, 5, 0, 0, 0, 43, 35, 34, 13, 4, 0, 4, 3, 1, 0, 
    0, 0, 21, 0, 38, 1, 0, 2, 4, 0, 4, 0, 0, 0, 7, 
    1, 3, 0, 0, 3, 3, 4, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 2, 30, 7, 0, 0, 0, 0, 3, 0, 7, 0, 0, 0, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 18, 0, 0, 0, 
    0, 0, 27, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 23, 2, 
    4, 17, 1, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 34, 1, 
    0, 0, 0, 20, 0, 0, 0, 28, 29, 0, 0, 0, 0, 0, 8, 
    34, 25, 0, 28, 2, 0, 21, 0, 0, 0, 0, 0, 4, 6, 0, 
    113, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 12, 
    0, 23, 0, 0, 0, 5, 61, 0, 0, 3, 20, 12, 4, 12, 24, 
    0, 7, 7, 0, 0, 4, 82, 37, 37, 21, 8, 20, 19, 18, 22, 
    0, 3, 7, 2, 4, 5, 70, 80, 36, 40, 37, 24, 8, 14, 15, 
    0, 3, 3, 4, 7, 6, 28, 42, 37, 43, 11, 4, 11, 13, 14, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 8, 1, 0, 32, 12, 9, 9, 19, 2, 0, 0, 
    25, 3, 0, 1, 2, 7, 0, 11, 30, 28, 7, 0, 1, 0, 0, 
    18, 8, 9, 7, 7, 7, 12, 79, 63, 17, 19, 16, 0, 0, 0, 
    0, 13, 11, 8, 10, 10, 14, 28, 24, 20, 6, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 18, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 13, 0, 0, 0, 6, 28, 0, 0, 0, 
    30, 40, 33, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 43, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 36, 0, 
    18, 47, 22, 9, 0, 0, 55, 71, 47, 0, 0, 0, 0, 0, 24, 
    64, 28, 5, 52, 16, 0, 0, 0, 7, 18, 19, 30, 33, 24, 9, 
    117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 
    23, 2, 12, 11, 13, 14, 8, 15, 18, 0, 14, 8, 17, 14, 21, 
    31, 55, 29, 32, 34, 35, 23, 19, 14, 12, 20, 28, 37, 17, 20, 
    9, 52, 0, 0, 18, 35, 80, 12, 34, 35, 35, 7, 0, 9, 31, 
    0, 39, 38, 18, 26, 32, 96, 0, 0, 0, 0, 22, 26, 24, 31, 
    0, 31, 33, 28, 31, 32, 56, 0, 0, 22, 33, 23, 16, 28, 29, 
    0, 26, 32, 33, 34, 36, 47, 44, 30, 30, 10, 17, 23, 22, 24, 
    
    -- channel=67
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 17, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 9, 33, 24, 24, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 64, 17, 1, 0, 0, 0, 0, 0, 0, 34, 55, 65, 42, 0, 
    0, 0, 0, 29, 29, 82, 94, 80, 45, 0, 0, 0, 0, 0, 0, 
    82, 74, 47, 0, 0, 0, 0, 0, 0, 13, 49, 68, 64, 56, 48, 
    7, 0, 1, 5, 0, 0, 0, 0, 37, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 36, 34, 3, 26, 26, 38, 55, 56, 36, 
    30, 74, 67, 65, 54, 41, 24, 8, 13, 11, 20, 19, 6, 8, 2, 
    32, 29, 39, 60, 74, 81, 82, 78, 64, 54, 38, 20, 0, 0, 0, 
    12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 26, 17, 5, 0, 34, 26, 4, 15, 41, 22, 0, 0, 0, 
    0, 0, 2, 3, 0, 0, 12, 21, 41, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=68
    49, 50, 50, 50, 50, 50, 50, 50, 50, 48, 50, 50, 50, 50, 51, 
    48, 50, 50, 49, 49, 49, 49, 49, 46, 16, 38, 50, 49, 49, 50, 
    48, 49, 50, 49, 50, 47, 50, 30, 14, 7, 34, 58, 49, 50, 50, 
    51, 50, 51, 51, 51, 29, 49, 29, 41, 34, 39, 58, 49, 51, 51, 
    0, 0, 52, 48, 49, 43, 58, 49, 54, 39, 20, 1, 0, 39, 51, 
    63, 73, 51, 23, 33, 0, 15, 25, 45, 36, 38, 49, 32, 67, 52, 
    0, 0, 10, 52, 29, 0, 0, 15, 52, 37, 21, 6, 18, 10, 29, 
    2, 34, 0, 26, 28, 47, 77, 21, 0, 0, 0, 2, 18, 34, 39, 
    81, 55, 66, 74, 60, 35, 32, 25, 43, 30, 36, 16, 8, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 1, 12, 8, 1, 27, 
    0, 0, 0, 0, 0, 0, 18, 0, 6, 0, 0, 0, 7, 26, 40, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 3, 22, 28, 12, 22, 38, 
    0, 0, 0, 0, 0, 0, 0, 3, 17, 31, 14, 7, 19, 29, 41, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 28, 33, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 7, 0, 0, 0, 0, 0, 0, 
    81, 80, 14, 0, 0, 0, 0, 0, 0, 0, 22, 52, 52, 32, 0, 
    0, 0, 0, 5, 12, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 
    0, 43, 0, 0, 0, 64, 90, 8, 0, 0, 0, 0, 9, 27, 21, 
    49, 42, 71, 57, 15, 0, 0, 0, 27, 14, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 
    0, 0, 25, 21, 2, 0, 48, 56, 27, 31, 43, 52, 21, 0, 10, 
    10, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 14, 12, 
    11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 26, 33, 0, 0, 0, 
    0, 15, 11, 8, 9, 10, 0, 0, 34, 42, 12, 0, 4, 6, 4, 
    
    -- channel=70
    28, 28, 28, 28, 28, 28, 28, 28, 28, 29, 25, 28, 28, 28, 28, 
    27, 28, 28, 28, 27, 27, 27, 27, 27, 21, 0, 17, 28, 27, 28, 
    25, 26, 27, 27, 28, 28, 24, 28, 0, 0, 16, 9, 28, 28, 27, 
    22, 26, 27, 28, 28, 28, 14, 17, 25, 31, 34, 42, 26, 27, 28, 
    0, 0, 0, 25, 26, 17, 41, 24, 37, 29, 23, 0, 0, 0, 24, 
    51, 64, 56, 15, 6, 5, 0, 0, 0, 13, 18, 40, 43, 55, 27, 
    0, 0, 0, 2, 38, 0, 0, 0, 34, 32, 15, 0, 0, 5, 0, 
    0, 42, 4, 9, 0, 30, 74, 63, 0, 0, 0, 0, 10, 15, 44, 
    12, 36, 41, 55, 41, 22, 10, 0, 24, 27, 10, 17, 1, 0, 0, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 
    0, 0, 0, 1, 0, 0, 0, 29, 2, 0, 10, 29, 34, 0, 13, 
    3, 0, 0, 0, 0, 0, 0, 0, 18, 20, 1, 0, 0, 21, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 14, 15, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 29, 7, 13, 21, 26, 
    
    -- channel=71
    38, 38, 38, 38, 38, 39, 38, 39, 37, 39, 39, 40, 39, 38, 38, 
    38, 38, 38, 38, 37, 37, 37, 37, 40, 55, 31, 31, 37, 37, 37, 
    40, 39, 37, 37, 36, 41, 37, 50, 43, 38, 45, 38, 39, 38, 38, 
    32, 36, 39, 38, 38, 52, 29, 34, 13, 10, 0, 14, 40, 39, 39, 
    18, 17, 36, 38, 38, 41, 34, 38, 33, 44, 65, 55, 45, 22, 39, 
    27, 25, 52, 45, 53, 79, 81, 75, 53, 36, 8, 10, 13, 11, 39, 
    31, 13, 32, 20, 56, 0, 0, 0, 0, 58, 70, 68, 65, 66, 34, 
    0, 6, 4, 11, 12, 1, 17, 56, 28, 0, 0, 0, 0, 0, 19, 
    0, 59, 30, 49, 55, 59, 61, 60, 48, 63, 61, 69, 62, 43, 18, 
    67, 40, 35, 29, 22, 19, 16, 0, 11, 2, 14, 5, 6, 16, 11, 
    0, 0, 0, 0, 6, 10, 16, 21, 20, 10, 3, 0, 0, 0, 10, 
    4, 1, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 30, 9, 4, 
    0, 0, 0, 0, 0, 0, 2, 29, 28, 38, 35, 0, 0, 14, 16, 
    18, 0, 0, 0, 0, 0, 0, 20, 22, 0, 0, 16, 20, 14, 24, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 7, 26, 19, 19, 20, 24, 
    
    -- channel=72
    40, 38, 38, 38, 38, 38, 38, 40, 38, 38, 38, 38, 38, 38, 38, 
    40, 38, 38, 39, 38, 38, 37, 39, 37, 40, 13, 28, 39, 38, 38, 
    37, 37, 39, 39, 39, 40, 34, 39, 20, 28, 0, 12, 39, 38, 39, 
    29, 36, 36, 39, 40, 50, 17, 51, 32, 40, 33, 8, 36, 36, 38, 
    0, 0, 10, 35, 37, 50, 27, 41, 33, 38, 23, 11, 3, 0, 34, 
    35, 32, 32, 18, 22, 2, 0, 0, 5, 44, 41, 40, 52, 0, 29, 
    0, 0, 0, 16, 44, 37, 0, 0, 0, 29, 20, 13, 4, 10, 0, 
    0, 1, 10, 0, 27, 47, 27, 32, 10, 15, 18, 10, 6, 16, 4, 
    0, 36, 33, 22, 22, 31, 16, 32, 19, 6, 10, 11, 0, 0, 3, 
    0, 0, 0, 0, 0, 1, 13, 7, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 3, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 44, 42, 29, 4, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 22, 1, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    7, 8, 8, 8, 8, 9, 9, 8, 8, 9, 11, 9, 8, 8, 8, 
    8, 8, 8, 8, 8, 8, 8, 7, 8, 15, 29, 16, 7, 8, 8, 
    11, 10, 9, 7, 8, 9, 11, 11, 21, 19, 30, 32, 9, 9, 9, 
    12, 9, 10, 8, 9, 9, 21, 0, 0, 0, 0, 3, 11, 10, 10, 
    36, 42, 45, 10, 10, 0, 3, 5, 7, 17, 31, 37, 39, 42, 16, 
    0, 0, 0, 16, 33, 40, 67, 61, 43, 10, 0, 0, 0, 9, 13, 
    52, 48, 44, 22, 0, 0, 0, 0, 5, 21, 37, 45, 51, 37, 43, 
    15, 10, 0, 20, 9, 0, 0, 0, 19, 7, 0, 0, 0, 0, 4, 
    22, 0, 1, 4, 19, 23, 39, 33, 23, 32, 45, 39, 49, 39, 27, 
    43, 54, 52, 52, 46, 38, 24, 17, 23, 17, 22, 20, 18, 19, 17, 
    4, 21, 19, 35, 44, 52, 60, 58, 51, 39, 33, 24, 11, 3, 6, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 28, 16, 0, 2, 9, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 1, 14, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 13, 15, 20, 18, 18, 0, 7, 8, 5, 0, 0, 0, 0, 0, 
    0, 16, 17, 19, 18, 17, 16, 63, 61, 20, 0, 0, 0, 0, 0, 
    0, 3, 6, 7, 10, 9, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    91, 91, 91, 91, 91, 90, 91, 91, 91, 90, 91, 90, 90, 91, 91, 
    90, 90, 90, 90, 90, 90, 90, 90, 84, 44, 59, 87, 90, 90, 90, 
    86, 87, 91, 91, 92, 89, 87, 64, 32, 40, 37, 76, 89, 90, 91, 
    89, 90, 88, 91, 92, 69, 81, 85, 103, 105, 110, 97, 87, 89, 91, 
    0, 0, 75, 84, 88, 89, 93, 93, 100, 87, 39, 7, 0, 43, 89, 
    130, 137, 75, 38, 54, 0, 0, 9, 47, 84, 111, 124, 110, 108, 86, 
    0, 0, 20, 96, 64, 23, 26, 82, 104, 65, 31, 7, 19, 5, 31, 
    16, 94, 21, 36, 79, 143, 151, 50, 7, 22, 38, 59, 71, 96, 80, 
    122, 83, 125, 104, 81, 57, 46, 59, 79, 44, 57, 27, 6, 0, 11, 
    0, 0, 0, 0, 0, 12, 18, 27, 20, 26, 3, 9, 21, 20, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 46, 40, 
    0, 0, 14, 0, 0, 0, 87, 76, 52, 60, 81, 81, 31, 33, 57, 
    0, 0, 0, 0, 0, 0, 0, 48, 59, 31, 0, 0, 40, 44, 64, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 39, 29, 42, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 45, 28, 24, 37, 52, 66, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 41, 0, 0, 0, 
    0, 11, 16, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 
    0, 11, 2, 0, 0, 0, 13, 40, 69, 0, 0, 0, 0, 0, 10, 
    35, 39, 0, 48, 0, 0, 21, 0, 0, 0, 0, 0, 11, 7, 24, 
    159, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 12, 0, 1, 5, 6, 0, 0, 0, 0, 0, 0, 12, 9, 16, 
    0, 43, 0, 0, 0, 18, 43, 0, 10, 17, 28, 30, 4, 0, 22, 
    0, 19, 5, 0, 0, 5, 127, 0, 0, 0, 0, 0, 14, 16, 27, 
    0, 2, 7, 0, 2, 4, 64, 9, 0, 0, 24, 28, 0, 18, 19, 
    0, 0, 3, 1, 4, 6, 30, 13, 26, 40, 6, 0, 7, 11, 17, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 6, 0, 0, 2, 7, 
    0, 0, 10, 1, 0, 0, 39, 51, 47, 33, 23, 24, 13, 4, 1, 
    0, 0, 3, 1, 0, 0, 39, 108, 78, 53, 28, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 49, 30, 21, 4, 0, 0, 0, 0, 
    
    -- channel=78
    1, 1, 1, 1, 1, 1, 2, 2, 2, 1, 0, 2, 2, 1, 1, 
    1, 2, 2, 2, 2, 2, 2, 3, 2, 0, 11, 5, 1, 2, 2, 
    3, 3, 2, 2, 2, 1, 2, 0, 4, 0, 0, 10, 1, 2, 2, 
    0, 0, 1, 3, 2, 0, 9, 0, 0, 0, 0, 0, 0, 1, 1, 
    13, 18, 16, 5, 3, 0, 0, 0, 0, 0, 0, 3, 11, 19, 2, 
    0, 0, 0, 9, 11, 10, 19, 17, 12, 0, 0, 0, 0, 0, 0, 
    9, 19, 10, 3, 0, 0, 0, 0, 0, 0, 1, 8, 11, 6, 14, 
    0, 0, 0, 11, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 13, 6, 1, 0, 19, 11, 5, 7, 20, 24, 8, 2, 2, 
    0, 0, 4, 2, 1, 1, 28, 59, 59, 44, 17, 5, 7, 5, 3, 
    0, 0, 0, 0, 0, 0, 14, 37, 19, 8, 9, 10, 7, 3, 1, 
    
    -- channel=79
    29, 29, 29, 29, 28, 29, 29, 28, 26, 30, 32, 29, 29, 29, 29, 
    29, 29, 29, 29, 29, 28, 28, 28, 29, 37, 38, 29, 28, 28, 29, 
    30, 29, 28, 28, 28, 29, 32, 33, 47, 52, 39, 40, 28, 29, 29, 
    36, 34, 30, 28, 28, 30, 28, 35, 37, 39, 30, 23, 35, 33, 31, 
    47, 45, 37, 28, 28, 36, 23, 34, 32, 39, 50, 52, 47, 46, 34, 
    38, 30, 28, 29, 34, 49, 58, 56, 54, 47, 37, 32, 29, 16, 36, 
    54, 52, 44, 37, 42, 35, 31, 18, 12, 38, 46, 48, 51, 49, 46, 
    40, 11, 20, 16, 38, 27, 20, 30, 41, 40, 32, 26, 24, 28, 25, 
    0, 50, 32, 32, 43, 47, 50, 62, 51, 60, 64, 62, 62, 57, 51, 
    51, 70, 73, 75, 72, 71, 72, 58, 59, 56, 59, 59, 50, 45, 37, 
    20, 28, 33, 37, 39, 50, 67, 69, 67, 62, 57, 50, 43, 25, 20, 
    6, 10, 13, 3, 1, 5, 26, 13, 21, 20, 14, 10, 16, 16, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 23, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 14, 23, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    60, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 45, 13, 0, 0, 41, 37, 35, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 17, 9, 9, 0, 0, 0, 34, 51, 46, 25, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 28, 
    0, 19, 26, 29, 30, 30, 32, 29, 18, 16, 15, 17, 0, 0, 0, 
    47, 45, 45, 42, 38, 35, 29, 23, 22, 25, 18, 12, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 12, 5, 0, 0, 0, 0, 0, 
    1, 7, 20, 15, 4, 1, 0, 0, 0, 0, 0, 32, 0, 0, 0, 
    4, 0, 1, 3, 0, 0, 0, 0, 11, 26, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 4, 24, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 12, 11, 22, 27, 23, 7, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 27, 14, 5, 6, 60, 52, 45, 42, 49, 30, 0, 0, 0, 
    0, 3, 7, 5, 4, 4, 55, 104, 88, 36, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 25, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    51, 50, 50, 50, 49, 50, 50, 51, 48, 49, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 49, 50, 49, 51, 49, 56, 30, 42, 50, 50, 50, 
    47, 48, 49, 51, 50, 51, 45, 53, 33, 47, 14, 27, 50, 49, 50, 
    48, 51, 51, 49, 50, 65, 31, 64, 54, 66, 60, 32, 53, 51, 51, 
    0, 0, 32, 45, 47, 67, 45, 57, 49, 52, 41, 25, 13, 0, 50, 
    63, 59, 54, 26, 31, 11, 0, 6, 17, 65, 66, 67, 81, 25, 47, 
    0, 0, 12, 32, 75, 46, 18, 27, 21, 44, 29, 18, 15, 21, 0, 
    0, 39, 23, 0, 45, 74, 59, 54, 22, 30, 38, 38, 34, 48, 30, 
    0, 67, 58, 47, 41, 48, 34, 51, 39, 31, 35, 34, 16, 11, 21, 
    0, 4, 4, 9, 12, 21, 38, 30, 27, 28, 20, 25, 18, 16, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 26, 16, 
    0, 0, 23, 14, 0, 0, 16, 54, 36, 33, 32, 31, 18, 15, 15, 
    12, 0, 0, 0, 0, 0, 0, 13, 10, 2, 0, 0, 6, 13, 18, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 15, 11, 19, 
    36, 2, 0, 0, 0, 0, 0, 0, 0, 3, 12, 16, 16, 19, 24, 
    
    -- channel=84
    3, 4, 4, 4, 5, 4, 4, 4, 5, 4, 3, 4, 4, 4, 5, 
    4, 4, 4, 4, 5, 4, 5, 3, 2, 0, 7, 10, 4, 4, 5, 
    4, 5, 4, 4, 6, 2, 6, 0, 0, 0, 20, 14, 4, 5, 4, 
    6, 2, 6, 5, 4, 0, 17, 0, 0, 0, 4, 36, 2, 4, 5, 
    7, 19, 11, 6, 4, 0, 17, 0, 8, 0, 0, 0, 0, 25, 5, 
    0, 11, 10, 9, 0, 0, 0, 0, 5, 0, 0, 0, 0, 44, 8, 
    0, 17, 4, 6, 0, 0, 13, 28, 49, 2, 0, 0, 0, 0, 18, 
    23, 17, 12, 37, 0, 0, 19, 0, 0, 0, 0, 1, 13, 6, 25, 
    96, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 
    8, 7, 1, 2, 6, 6, 0, 0, 0, 0, 0, 0, 5, 7, 15, 
    0, 33, 0, 0, 3, 17, 7, 0, 2, 5, 16, 18, 10, 2, 21, 
    0, 23, 11, 0, 4, 10, 97, 5, 13, 7, 5, 3, 15, 19, 26, 
    0, 8, 11, 4, 8, 8, 69, 17, 0, 2, 18, 28, 12, 23, 22, 
    0, 9, 10, 9, 10, 10, 34, 9, 18, 38, 17, 11, 17, 20, 22, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    19, 5, 0, 7, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 
    25, 11, 0, 13, 5, 0, 0, 0, 1, 3, 1, 2, 1, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 6, 8, 
    8, 12, 12, 13, 13, 15, 13, 14, 10, 11, 10, 13, 11, 6, 11, 
    13, 26, 22, 24, 25, 29, 33, 13, 15, 16, 20, 20, 31, 15, 6, 
    17, 23, 27, 20, 20, 25, 59, 50, 62, 57, 46, 22, 7, 11, 0, 
    0, 24, 27, 25, 24, 24, 53, 100, 87, 47, 21, 21, 6, 0, 0, 
    0, 17, 18, 19, 21, 21, 27, 47, 24, 28, 13, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 10, 19, 34, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 18, 21, 19, 0, 
    0, 0, 0, 0, 0, 23, 50, 87, 41, 0, 0, 0, 0, 0, 0, 
    0, 34, 9, 12, 17, 25, 9, 0, 0, 24, 46, 50, 44, 38, 4, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    13, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 0, 
    0, 0, 0, 0, 0, 0, 52, 78, 68, 62, 57, 20, 0, 0, 12, 
    8, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 9, 22, 2, 6, 
    0, 2, 1, 1, 1, 1, 3, 0, 0, 13, 32, 4, 0, 3, 0, 
    1, 15, 14, 13, 14, 15, 19, 20, 31, 11, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 33, 25, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 62, 73, 94, 102, 92, 61, 43, 23, 21, 9, 0, 0, 0, 0, 
    28, 27, 0, 0, 36, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 68, 66, 50, 48, 49, 67, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 45, 49, 46, 47, 45, 63, 0, 15, 0, 0, 0, 0, 0, 0, 
    0, 13, 23, 28, 27, 25, 40, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 14, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 28, 17, 14, 0, 0, 
    0, 0, 11, 16, 0, 57, 3, 0, 0, 0, 0, 0, 6, 0, 0, 
    12, 0, 0, 0, 30, 48, 0, 0, 0, 13, 24, 24, 0, 20, 0, 
    0, 0, 9, 0, 0, 0, 0, 54, 9, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 11, 3, 4, 0, 20, 0, 27, 11, 8, 0, 
    11, 7, 5, 2, 0, 0, 5, 0, 2, 6, 12, 2, 0, 0, 0, 
    29, 0, 27, 18, 15, 7, 10, 10, 9, 13, 4, 0, 0, 0, 0, 
    15, 0, 4, 28, 20, 0, 0, 14, 0, 0, 0, 0, 17, 0, 0, 
    51, 6, 6, 19, 9, 8, 0, 0, 16, 37, 40, 0, 0, 0, 0, 
    66, 10, 8, 11, 8, 8, 0, 27, 66, 0, 0, 0, 0, 0, 0, 
    44, 9, 6, 4, 3, 2, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 20, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 24, 21, 21, 25, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 10, 13, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 32, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 16, 0, 
    8, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 48, 0, 
    0, 0, 0, 2, 0, 0, 7, 37, 53, 0, 0, 0, 0, 0, 0, 
    43, 36, 0, 37, 1, 0, 33, 0, 0, 0, 0, 0, 10, 17, 9, 
    136, 20, 5, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 15, 
    0, 41, 0, 0, 0, 9, 78, 0, 14, 20, 37, 32, 4, 0, 25, 
    0, 2, 3, 0, 0, 2, 111, 0, 0, 0, 0, 0, 11, 18, 26, 
    0, 2, 4, 0, 2, 4, 49, 21, 0, 0, 27, 26, 1, 14, 21, 
    0, 0, 5, 4, 7, 8, 16, 22, 25, 44, 6, 0, 10, 12, 17, 
    
    -- channel=92
    6, 6, 6, 6, 6, 7, 7, 7, 7, 5, 8, 7, 7, 6, 7, 
    6, 6, 6, 6, 6, 5, 5, 7, 2, 3, 16, 6, 5, 6, 5, 
    8, 6, 7, 6, 5, 5, 6, 0, 0, 20, 0, 22, 6, 6, 6, 
    1, 3, 5, 6, 6, 14, 7, 18, 9, 3, 0, 0, 7, 6, 7, 
    0, 0, 30, 7, 5, 30, 0, 16, 0, 0, 1, 1, 0, 11, 11, 
    14, 5, 0, 0, 13, 0, 19, 23, 29, 33, 12, 3, 9, 0, 3, 
    0, 0, 6, 28, 16, 0, 0, 0, 0, 0, 3, 8, 28, 9, 4, 
    13, 0, 0, 0, 28, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 17, 0, 0, 8, 4, 42, 12, 2, 28, 9, 9, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 27, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 38, 16, 6, 0, 16, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 14, 6, 22, 3, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 9, 3, 0, 0, 2, 1, 0, 0, 
    
    -- channel=93
    6, 4, 4, 4, 3, 4, 3, 6, 3, 4, 2, 4, 4, 4, 3, 
    6, 4, 4, 4, 3, 4, 3, 5, 6, 28, 0, 0, 5, 3, 3, 
    3, 3, 2, 5, 3, 6, 0, 18, 4, 15, 0, 0, 4, 3, 3, 
    0, 4, 2, 3, 4, 29, 0, 29, 6, 21, 11, 0, 3, 2, 2, 
    0, 0, 0, 1, 1, 22, 0, 11, 0, 10, 7, 0, 0, 0, 0, 
    15, 3, 4, 1, 0, 2, 0, 0, 0, 16, 16, 19, 45, 0, 0, 
    0, 0, 0, 0, 38, 66, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 27, 0, 31, 0, 5, 16, 5, 0, 0, 0, 
    0, 15, 10, 0, 0, 7, 0, 18, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 9, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 23, 29, 13, 0, 0, 44, 18, 10, 1, 1, 3, 0, 0, 
    43, 0, 0, 11, 6, 1, 0, 22, 25, 23, 11, 0, 0, 0, 0, 
    80, 4, 0, 6, 3, 2, 0, 33, 33, 4, 0, 0, 0, 0, 0, 
    63, 15, 6, 7, 6, 3, 0, 7, 2, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    42, 41, 41, 41, 40, 41, 41, 41, 40, 41, 42, 41, 40, 41, 40, 
    42, 41, 41, 41, 41, 41, 41, 41, 42, 52, 35, 36, 42, 41, 41, 
    40, 40, 41, 41, 41, 42, 41, 47, 49, 57, 25, 28, 42, 40, 41, 
    43, 45, 41, 40, 41, 50, 29, 56, 47, 56, 50, 27, 44, 42, 41, 
    40, 30, 23, 38, 41, 54, 32, 47, 41, 47, 46, 42, 38, 23, 39, 
    43, 34, 36, 35, 34, 36, 25, 27, 32, 57, 55, 49, 59, 14, 39, 
    40, 31, 35, 32, 57, 75, 41, 37, 17, 38, 38, 37, 32, 36, 27, 
    21, 18, 37, 11, 46, 52, 30, 45, 45, 57, 59, 49, 42, 44, 29, 
    0, 50, 38, 33, 36, 47, 38, 54, 38, 39, 40, 44, 36, 40, 46, 
    9, 47, 48, 53, 56, 59, 68, 60, 56, 61, 52, 56, 45, 37, 33, 
    33, 29, 40, 34, 27, 29, 42, 47, 48, 51, 49, 44, 41, 36, 25, 
    19, 0, 25, 26, 18, 11, 23, 58, 51, 47, 37, 27, 22, 31, 19, 
    24, 0, 9, 19, 12, 8, 0, 13, 9, 12, 16, 27, 19, 16, 14, 
    41, 8, 7, 13, 8, 8, 0, 1, 20, 24, 14, 4, 17, 13, 17, 
    41, 9, 7, 9, 9, 9, 0, 14, 11, 0, 8, 16, 14, 16, 19, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 48, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 39, 0, 0, 0, 
    16, 48, 54, 1, 0, 0, 11, 0, 0, 0, 0, 0, 0, 76, 5, 
    0, 4, 0, 0, 1, 0, 26, 27, 39, 0, 0, 0, 0, 57, 9, 
    13, 63, 30, 27, 0, 0, 23, 41, 58, 0, 0, 0, 13, 0, 53, 
    86, 19, 0, 69, 6, 0, 8, 0, 0, 0, 0, 0, 7, 2, 11, 
    174, 0, 0, 5, 7, 0, 0, 0, 0, 0, 3, 0, 6, 8, 3, 
    67, 12, 18, 14, 13, 6, 0, 0, 0, 0, 0, 0, 3, 9, 22, 
    0, 34, 2, 18, 31, 42, 29, 23, 10, 2, 7, 17, 28, 5, 24, 
    0, 60, 0, 0, 0, 20, 76, 0, 0, 0, 17, 6, 8, 6, 32, 
    0, 20, 19, 0, 0, 4, 171, 9, 0, 0, 0, 16, 13, 23, 37, 
    0, 0, 8, 0, 1, 2, 97, 26, 0, 13, 18, 20, 5, 27, 35, 
    0, 0, 0, 0, 0, 1, 36, 32, 13, 38, 2, 3, 16, 21, 29, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=99
    26, 25, 25, 25, 25, 25, 25, 26, 25, 27, 26, 25, 25, 25, 25, 
    27, 26, 26, 26, 26, 26, 25, 25, 27, 44, 22, 19, 26, 26, 26, 
    26, 25, 25, 26, 25, 27, 25, 37, 38, 42, 17, 13, 27, 25, 26, 
    23, 27, 26, 25, 25, 41, 17, 41, 30, 36, 27, 11, 28, 27, 27, 
    42, 26, 15, 24, 25, 33, 17, 28, 26, 37, 46, 47, 41, 11, 28, 
    20, 13, 26, 26, 27, 39, 29, 28, 23, 42, 34, 25, 35, 0, 26, 
    40, 22, 23, 11, 44, 57, 20, 9, 0, 33, 39, 40, 30, 38, 18, 
    0, 11, 31, 4, 29, 26, 10, 43, 37, 35, 34, 21, 15, 15, 16, 
    0, 25, 10, 5, 19, 37, 33, 40, 26, 32, 31, 40, 36, 41, 38, 
    9, 39, 39, 40, 40, 39, 46, 40, 35, 40, 39, 39, 27, 24, 20, 
    30, 21, 34, 33, 31, 30, 36, 35, 39, 37, 32, 25, 20, 20, 12, 
    11, 0, 11, 13, 5, 0, 0, 27, 20, 15, 8, 7, 12, 14, 0, 
    12, 0, 0, 3, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 2, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 10, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 8, 12, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 19, 5, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 56, 7, 0, 0, 0, 0, 0, 0, 0, 17, 45, 53, 35, 0, 
    0, 0, 0, 9, 12, 48, 70, 58, 36, 0, 0, 0, 0, 0, 0, 
    80, 76, 34, 0, 0, 16, 0, 0, 0, 0, 26, 50, 46, 42, 38, 
    26, 0, 4, 0, 0, 0, 0, 0, 34, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 13, 22, 0, 8, 16, 22, 44, 54, 41, 
    8, 72, 66, 67, 59, 47, 34, 21, 18, 24, 25, 32, 12, 11, 7, 
    45, 48, 52, 72, 81, 88, 88, 86, 74, 67, 52, 35, 11, 0, 0, 
    19, 3, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 11, 25, 21, 10, 5, 9, 22, 0, 3, 33, 29, 0, 0, 0, 
    0, 0, 3, 6, 3, 2, 0, 0, 17, 10, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=101
    56, 56, 56, 56, 56, 57, 56, 57, 56, 56, 57, 56, 56, 56, 56, 
    56, 56, 56, 56, 56, 56, 56, 56, 56, 54, 52, 55, 56, 56, 56, 
    58, 57, 57, 56, 57, 57, 56, 55, 50, 39, 45, 58, 56, 57, 57, 
    54, 55, 55, 57, 59, 55, 54, 45, 32, 23, 19, 40, 54, 55, 56, 
    33, 40, 56, 58, 58, 49, 50, 53, 52, 54, 53, 46, 46, 51, 54, 
    24, 30, 44, 54, 60, 59, 65, 65, 60, 44, 25, 22, 16, 36, 52, 
    35, 41, 47, 43, 37, 0, 0, 0, 31, 55, 60, 58, 57, 52, 53, 
    0, 9, 7, 37, 35, 20, 27, 37, 40, 29, 12, 7, 8, 15, 29, 
    12, 38, 34, 49, 58, 55, 59, 47, 38, 41, 45, 42, 41, 35, 27, 
    37, 43, 42, 42, 41, 36, 29, 19, 24, 16, 15, 8, 8, 10, 16, 
    0, 0, 0, 1, 6, 15, 22, 23, 18, 13, 7, 3, 0, 2, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 15, 16, 
    0, 0, 0, 0, 0, 0, 19, 52, 47, 45, 39, 23, 13, 14, 22, 
    0, 0, 0, 0, 0, 0, 0, 80, 79, 37, 9, 10, 10, 15, 27, 
    0, 0, 0, 0, 0, 0, 0, 15, 2, 2, 11, 7, 11, 17, 27, 
    
    -- channel=102
    17, 17, 17, 17, 17, 18, 17, 17, 15, 18, 20, 17, 17, 17, 17, 
    17, 17, 17, 17, 16, 16, 17, 15, 18, 36, 21, 14, 16, 16, 16, 
    19, 18, 16, 16, 16, 19, 19, 29, 39, 39, 37, 23, 17, 17, 17, 
    19, 20, 18, 16, 16, 25, 13, 20, 14, 13, 2, 6, 21, 20, 18, 
    38, 34, 20, 17, 17, 18, 11, 18, 18, 33, 56, 53, 47, 26, 20, 
    22, 14, 24, 28, 32, 68, 70, 63, 45, 27, 10, 7, 7, 1, 23, 
    53, 38, 35, 16, 34, 18, 0, 0, 0, 38, 55, 58, 54, 54, 36, 
    9, 0, 8, 2, 10, 0, 3, 36, 28, 13, 1, 0, 0, 0, 18, 
    0, 34, 15, 24, 38, 42, 49, 57, 48, 66, 63, 70, 68, 54, 34, 
    63, 68, 67, 66, 59, 53, 50, 35, 40, 38, 46, 40, 35, 34, 23, 
    13, 10, 24, 34, 40, 48, 63, 64, 60, 53, 44, 33, 17, 10, 10, 
    5, 6, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 20, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 5, 9, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 14, 0, 0, 
    0, 0, 0, 0, 1, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 3, 0, 0, 22, 11, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 9, 12, 0, 0, 0, 0, 11, 6, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 12, 24, 23, 19, 13, 9, 14, 7, 5, 5, 1, 0, 3, 1, 
    28, 6, 2, 13, 18, 16, 0, 0, 0, 0, 0, 0, 3, 6, 0, 
    37, 19, 16, 17, 18, 19, 0, 0, 0, 0, 7, 5, 9, 3, 0, 
    43, 29, 25, 24, 22, 22, 6, 0, 8, 9, 8, 13, 9, 6, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 28, 32, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 4, 0, 0, 0, 0, 0, 0, 
    77, 75, 12, 0, 0, 0, 0, 0, 0, 0, 25, 53, 53, 30, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 
    0, 51, 0, 0, 0, 67, 90, 4, 0, 0, 0, 0, 10, 31, 21, 
    45, 41, 65, 51, 7, 0, 0, 0, 21, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 25, 20, 1, 0, 48, 67, 35, 37, 49, 56, 12, 0, 7, 
    15, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 10, 8, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 31, 0, 0, 0, 
    0, 17, 13, 9, 10, 10, 0, 0, 33, 40, 9, 0, 2, 3, 1, 
    
    -- channel=106
    54, 54, 54, 54, 54, 54, 54, 55, 56, 53, 52, 54, 54, 54, 55, 
    53, 54, 54, 54, 53, 54, 54, 54, 53, 39, 34, 49, 54, 54, 54, 
    52, 53, 54, 54, 54, 54, 51, 48, 24, 10, 38, 44, 54, 54, 54, 
    45, 49, 53, 55, 55, 50, 49, 38, 36, 33, 37, 58, 49, 51, 53, 
    0, 2, 40, 53, 54, 44, 62, 48, 54, 46, 36, 19, 12, 23, 50, 
    48, 60, 64, 43, 42, 29, 21, 26, 32, 32, 31, 43, 39, 66, 50, 
    0, 0, 13, 34, 41, 0, 0, 11, 53, 50, 39, 27, 24, 29, 24, 
    0, 47, 20, 42, 24, 39, 71, 56, 15, 0, 0, 8, 21, 27, 47, 
    46, 45, 49, 62, 53, 39, 35, 15, 32, 29, 23, 21, 14, 5, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 
    0, 11, 11, 9, 1, 0, 4, 6, 0, 0, 11, 33, 42, 24, 39, 
    11, 7, 1, 0, 0, 3, 40, 49, 66, 63, 43, 17, 31, 43, 47, 
    4, 4, 5, 1, 2, 3, 36, 76, 60, 26, 39, 56, 38, 40, 44, 
    0, 16, 12, 8, 8, 8, 23, 26, 34, 63, 53, 34, 39, 43, 47, 
    
    -- channel=107
    4, 1, 1, 1, 0, 0, 0, 2, 0, 2, 0, 0, 1, 1, 0, 
    3, 1, 1, 1, 0, 1, 0, 1, 6, 30, 0, 0, 2, 1, 0, 
    0, 0, 0, 2, 0, 5, 0, 22, 4, 15, 0, 0, 2, 0, 0, 
    0, 3, 0, 0, 0, 29, 0, 32, 11, 31, 22, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 7, 0, 15, 10, 0, 0, 0, 0, 
    19, 7, 5, 0, 0, 0, 0, 0, 0, 14, 25, 28, 57, 0, 0, 
    0, 0, 0, 0, 42, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 34, 8, 45, 0, 7, 28, 15, 7, 6, 0, 
    0, 7, 8, 0, 0, 4, 0, 12, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 6, 0, 18, 1, 8, 0, 0, 0, 
    12, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    19, 0, 21, 39, 20, 0, 0, 77, 39, 26, 12, 11, 0, 0, 0, 
    62, 0, 0, 11, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    96, 9, 3, 8, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 26, 17, 15, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    20, 21, 21, 21, 21, 21, 21, 20, 20, 21, 23, 22, 21, 21, 21, 
    20, 21, 21, 21, 21, 21, 22, 20, 20, 19, 40, 29, 20, 21, 21, 
    21, 21, 21, 20, 21, 20, 24, 21, 29, 21, 54, 44, 22, 21, 22, 
    30, 26, 25, 20, 20, 14, 36, 7, 25, 20, 26, 51, 26, 26, 24, 
    53, 58, 52, 21, 22, 6, 30, 16, 29, 28, 40, 45, 45, 57, 31, 
    25, 33, 35, 25, 35, 36, 56, 52, 47, 21, 18, 19, 7, 62, 34, 
    57, 60, 47, 33, 17, 0, 41, 41, 57, 33, 36, 38, 40, 41, 54, 
    50, 57, 26, 54, 22, 8, 35, 30, 32, 20, 17, 23, 30, 27, 49, 
    95, 19, 22, 30, 38, 33, 44, 22, 41, 47, 51, 47, 57, 53, 40, 
    84, 54, 60, 58, 55, 48, 40, 43, 45, 36, 49, 38, 46, 48, 46, 
    37, 48, 42, 52, 58, 62, 62, 61, 56, 48, 49, 47, 47, 37, 39, 
    17, 47, 12, 9, 17, 30, 41, 13, 24, 26, 27, 30, 31, 18, 32, 
    0, 35, 18, 8, 16, 22, 77, 0, 0, 0, 0, 0, 12, 28, 42, 
    0, 18, 18, 15, 18, 19, 24, 0, 0, 0, 0, 23, 22, 36, 44, 
    0, 11, 17, 17, 16, 17, 24, 0, 0, 20, 17, 22, 29, 35, 44, 
    
    -- channel=109
    3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 4, 29, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 21, 13, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 24, 3, 12, 3, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 6, 0, 1, 0, 15, 19, 13, 9, 0, 0, 
    0, 0, 0, 11, 0, 29, 0, 0, 0, 4, 11, 6, 28, 0, 0, 
    3, 0, 0, 0, 16, 101, 0, 0, 0, 1, 13, 16, 0, 0, 0, 
    0, 0, 19, 0, 0, 18, 0, 31, 7, 12, 23, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 25, 0, 6, 0, 13, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 6, 8, 0, 26, 0, 13, 0, 0, 0, 
    21, 0, 14, 3, 0, 0, 0, 0, 0, 8, 1, 0, 0, 0, 0, 
    25, 0, 13, 28, 15, 0, 0, 33, 5, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 14, 10, 2, 0, 7, 11, 18, 14, 0, 0, 0, 0, 
    83, 3, 0, 5, 2, 1, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    68, 12, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 4, 1, 2, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 8, 8, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    28, 26, 26, 26, 25, 26, 26, 27, 24, 26, 27, 27, 26, 26, 25, 
    28, 26, 26, 26, 25, 26, 25, 28, 28, 56, 13, 11, 26, 25, 25, 
    30, 26, 25, 26, 23, 28, 25, 44, 47, 58, 2, 8, 27, 25, 25, 
    17, 27, 25, 25, 26, 50, 3, 50, 16, 19, 2, 0, 30, 27, 26, 
    24, 9, 2, 26, 25, 49, 2, 32, 14, 32, 50, 53, 44, 0, 23, 
    13, 0, 8, 33, 31, 64, 53, 48, 33, 47, 24, 10, 31, 0, 18, 
    35, 6, 17, 15, 48, 78, 0, 0, 0, 27, 50, 60, 48, 48, 10, 
    0, 0, 21, 0, 19, 22, 0, 35, 37, 34, 23, 0, 0, 0, 0, 
    0, 27, 19, 2, 15, 46, 34, 76, 29, 36, 37, 50, 41, 40, 33, 
    0, 38, 24, 28, 24, 25, 32, 15, 9, 27, 12, 28, 5, 6, 0, 
    6, 0, 1, 4, 3, 0, 13, 20, 25, 26, 16, 3, 0, 0, 0, 
    30, 0, 27, 22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    26, 0, 1, 21, 10, 0, 0, 14, 2, 14, 29, 17, 0, 0, 0, 
    80, 2, 0, 7, 2, 1, 0, 0, 28, 11, 0, 0, 9, 0, 0, 
    83, 7, 0, 2, 0, 0, 0, 0, 0, 0, 2, 17, 3, 0, 0, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 24, 41, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 44, 0, 0, 0, 0, 0, 0, 0, 0, 26, 43, 45, 32, 0, 
    0, 0, 0, 0, 0, 0, 14, 58, 39, 0, 0, 0, 0, 0, 0, 
    0, 58, 0, 0, 0, 60, 65, 0, 0, 0, 2, 28, 33, 43, 13, 
    78, 0, 36, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 1, 8, 0, 0, 66, 95, 65, 64, 68, 48, 0, 0, 8, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 2, 5, 
    8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 37, 19, 0, 0, 0, 
    0, 21, 17, 14, 16, 17, 14, 0, 39, 30, 0, 0, 0, 0, 0, 
    
    -- channel=113
    3, 4, 4, 4, 4, 3, 4, 3, 4, 3, 4, 2, 3, 4, 4, 
    2, 4, 4, 3, 4, 3, 4, 3, 0, 0, 0, 11, 3, 4, 4, 
    0, 1, 4, 4, 6, 1, 2, 0, 0, 0, 0, 5, 2, 3, 4, 
    13, 5, 4, 3, 4, 0, 12, 0, 30, 33, 47, 46, 1, 4, 4, 
    0, 0, 8, 0, 2, 0, 20, 5, 17, 0, 0, 0, 0, 0, 3, 
    49, 58, 6, 0, 0, 0, 0, 0, 0, 0, 33, 48, 36, 66, 6, 
    0, 0, 0, 21, 0, 0, 34, 72, 75, 0, 0, 0, 0, 0, 0, 
    35, 63, 0, 20, 13, 58, 77, 0, 0, 0, 8, 35, 44, 53, 37, 
    138, 11, 43, 31, 7, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 11, 6, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 29, 20, 
    0, 18, 3, 2, 1, 11, 96, 76, 66, 70, 79, 64, 9, 1, 33, 
    0, 0, 0, 0, 0, 3, 29, 0, 0, 0, 0, 0, 27, 24, 32, 
    0, 3, 2, 0, 2, 3, 22, 0, 0, 0, 43, 32, 5, 18, 20, 
    0, 11, 12, 10, 13, 15, 19, 7, 43, 43, 7, 0, 12, 18, 23, 
    
    -- channel=114
    56, 55, 55, 55, 55, 56, 55, 56, 55, 55, 57, 55, 55, 55, 55, 
    56, 55, 55, 55, 55, 55, 55, 55, 55, 58, 47, 52, 56, 55, 55, 
    56, 56, 55, 56, 56, 56, 55, 57, 55, 55, 39, 49, 55, 55, 56, 
    54, 56, 54, 56, 57, 58, 46, 57, 43, 44, 36, 35, 55, 55, 55, 
    37, 38, 44, 55, 56, 60, 46, 56, 51, 56, 56, 50, 47, 42, 52, 
    40, 37, 47, 51, 52, 57, 54, 55, 54, 56, 45, 40, 41, 23, 53, 
    39, 37, 45, 42, 52, 35, 10, 11, 22, 54, 57, 55, 53, 51, 45, 
    9, 6, 24, 21, 46, 39, 30, 45, 45, 44, 34, 26, 23, 30, 29, 
    0, 55, 43, 46, 54, 58, 56, 62, 46, 49, 50, 50, 44, 41, 40, 
    24, 50, 50, 53, 52, 52, 52, 41, 41, 38, 35, 34, 27, 23, 24, 
    1, 3, 11, 12, 12, 18, 33, 34, 33, 32, 26, 21, 18, 18, 19, 
    0, 0, 6, 0, 0, 0, 0, 5, 5, 6, 5, 14, 21, 24, 16, 
    0, 0, 0, 0, 0, 0, 0, 45, 41, 37, 31, 23, 13, 14, 18, 
    5, 0, 0, 0, 0, 0, 0, 43, 46, 25, 6, 3, 13, 13, 23, 
    6, 0, 0, 0, 0, 0, 0, 15, 2, 0, 8, 12, 12, 17, 24, 
    
    -- channel=115
    63, 63, 63, 63, 63, 63, 63, 62, 62, 65, 62, 63, 63, 63, 63, 
    62, 62, 62, 62, 61, 62, 61, 61, 63, 54, 36, 52, 62, 62, 62, 
    59, 59, 62, 62, 62, 64, 60, 63, 39, 36, 47, 47, 62, 62, 63, 
    61, 64, 62, 62, 62, 62, 50, 60, 67, 73, 72, 73, 65, 65, 64, 
    0, 0, 42, 57, 60, 59, 71, 63, 72, 72, 61, 35, 16, 18, 63, 
    95, 100, 78, 40, 48, 32, 23, 30, 39, 61, 69, 83, 80, 81, 64, 
    0, 0, 11, 52, 75, 26, 13, 29, 61, 64, 49, 32, 28, 36, 23, 
    0, 78, 25, 24, 37, 80, 109, 81, 19, 7, 16, 28, 42, 56, 74, 
    45, 74, 86, 87, 74, 60, 55, 53, 75, 68, 64, 60, 40, 22, 12, 
    57, 7, 10, 5, 9, 13, 19, 19, 22, 21, 20, 11, 24, 28, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 30, 33, 
    0, 2, 20, 15, 0, 0, 24, 50, 27, 25, 32, 51, 39, 18, 36, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 14, 40, 53, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 42, 35, 40, 53, 
    7, 9, 6, 2, 0, 1, 0, 0, 2, 37, 39, 32, 39, 50, 59, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 23, 29, 34, 33, 28, 22, 18, 12, 15, 8, 1, 0, 0, 0, 
    9, 0, 0, 1, 12, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 14, 28, 24, 16, 14, 17, 31, 22, 19, 27, 23, 0, 0, 0, 
    0, 12, 15, 17, 14, 13, 35, 85, 77, 42, 0, 0, 0, 0, 0, 
    0, 0, 1, 4, 6, 4, 10, 33, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 48, 14, 0, 0, 0, 
    3, 2, 0, 0, 0, 0, 5, 0, 37, 21, 33, 40, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 
    105, 110, 56, 6, 3, 0, 0, 0, 0, 0, 16, 57, 78, 91, 8, 
    0, 0, 0, 27, 38, 57, 94, 82, 62, 0, 0, 0, 0, 0, 6, 
    108, 128, 75, 12, 0, 0, 16, 0, 0, 2, 33, 56, 64, 53, 80, 
    54, 0, 5, 56, 21, 0, 0, 0, 57, 48, 11, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 11, 34, 4, 0, 0, 7, 6, 43, 67, 58, 
    32, 85, 86, 85, 77, 63, 38, 28, 30, 13, 31, 26, 12, 10, 17, 
    56, 76, 66, 91, 106, 117, 106, 97, 78, 66, 54, 38, 20, 0, 1, 
    1, 27, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 16, 41, 20, 3, 1, 87, 12, 0, 0, 35, 58, 0, 0, 0, 
    0, 0, 3, 2, 0, 0, 21, 19, 39, 40, 0, 0, 0, 6, 12, 
    0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 4, 1, 0, 4, 
    
    -- channel=118
    76, 75, 75, 75, 75, 75, 75, 76, 74, 76, 74, 76, 75, 75, 75, 
    75, 75, 75, 75, 74, 74, 74, 74, 74, 74, 47, 63, 75, 74, 75, 
    74, 74, 74, 75, 75, 76, 72, 77, 57, 49, 53, 55, 75, 75, 75, 
    68, 74, 76, 75, 75, 80, 56, 73, 62, 66, 59, 64, 76, 76, 76, 
    14, 14, 46, 72, 73, 74, 74, 75, 76, 79, 76, 55, 40, 29, 73, 
    79, 81, 86, 62, 59, 65, 49, 53, 55, 69, 63, 71, 70, 58, 74, 
    8, 0, 27, 46, 81, 30, 0, 4, 43, 80, 73, 60, 49, 57, 35, 
    0, 39, 32, 23, 42, 63, 81, 89, 35, 19, 18, 17, 27, 39, 60, 
    0, 79, 71, 81, 80, 77, 68, 66, 69, 71, 62, 67, 49, 36, 23, 
    47, 23, 22, 21, 21, 22, 29, 21, 23, 21, 21, 11, 14, 22, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 25, 
    0, 0, 7, 0, 0, 0, 0, 16, 0, 0, 4, 28, 37, 16, 23, 
    0, 0, 0, 0, 0, 0, 0, 25, 34, 30, 12, 0, 2, 27, 37, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 27, 28, 43, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 17, 30, 25, 29, 38, 48, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 12, 7, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 2, 2, 0, 0, 27, 84, 77, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 26, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    9, 7, 7, 7, 6, 7, 6, 8, 7, 8, 4, 7, 7, 7, 6, 
    9, 7, 7, 7, 6, 7, 6, 8, 11, 29, 0, 0, 8, 7, 6, 
    7, 6, 6, 8, 6, 10, 3, 23, 7, 6, 0, 0, 8, 6, 6, 
    0, 5, 4, 7, 7, 29, 0, 23, 3, 10, 3, 0, 5, 5, 5, 
    0, 0, 0, 5, 6, 15, 0, 9, 2, 10, 11, 2, 0, 0, 0, 
    3, 0, 0, 9, 0, 14, 0, 0, 0, 10, 7, 8, 30, 0, 0, 
    0, 0, 0, 0, 27, 59, 0, 0, 0, 3, 6, 5, 0, 0, 0, 
    0, 0, 6, 0, 0, 17, 0, 30, 0, 1, 9, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 9, 0, 13, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 13, 23, 10, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 13, 9, 5, 0, 9, 17, 24, 19, 0, 0, 0, 0, 
    74, 8, 3, 7, 6, 5, 0, 20, 43, 8, 1, 4, 7, 0, 0, 
    56, 20, 12, 10, 9, 7, 0, 0, 5, 0, 14, 9, 0, 0, 0, 
    
    -- channel=121
    102, 103, 103, 103, 103, 103, 103, 102, 102, 104, 104, 103, 103, 103, 103, 
    103, 103, 103, 103, 103, 103, 103, 102, 101, 100, 104, 105, 103, 103, 104, 
    103, 103, 104, 103, 103, 104, 104, 102, 100, 91, 100, 107, 104, 104, 105, 
    105, 104, 105, 103, 103, 101, 104, 96, 91, 89, 84, 107, 107, 106, 106, 
    97, 102, 112, 102, 104, 98, 101, 101, 104, 108, 110, 106, 101, 108, 110, 
    80, 84, 107, 94, 104, 101, 107, 108, 109, 105, 90, 84, 72, 98, 111, 
    89, 92, 99, 85, 95, 41, 56, 67, 97, 111, 108, 102, 100, 101, 105, 
    47, 70, 62, 91, 96, 72, 84, 94, 89, 77, 65, 61, 65, 73, 89, 
    56, 99, 72, 87, 105, 108, 114, 92, 90, 95, 98, 96, 95, 95, 87, 
    96, 96, 104, 103, 102, 100, 95, 85, 88, 73, 83, 69, 67, 67, 71, 
    31, 41, 45, 50, 56, 64, 73, 74, 72, 63, 58, 55, 60, 58, 62, 
    0, 21, 12, 0, 0, 0, 29, 27, 31, 32, 39, 50, 52, 49, 57, 
    0, 0, 2, 0, 0, 0, 57, 43, 33, 31, 28, 26, 29, 49, 70, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 45, 58, 82, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 38, 43, 51, 64, 84, 
    
    -- channel=122
    20, 20, 20, 20, 20, 21, 20, 21, 20, 21, 21, 20, 21, 20, 20, 
    22, 21, 21, 22, 21, 21, 21, 22, 24, 53, 36, 19, 21, 21, 21, 
    25, 24, 22, 21, 20, 24, 22, 40, 54, 44, 24, 26, 22, 21, 21, 
    15, 19, 20, 22, 22, 42, 18, 27, 0, 0, 0, 0, 22, 20, 21, 
    81, 62, 28, 26, 24, 27, 4, 18, 6, 18, 46, 69, 76, 37, 22, 
    0, 0, 17, 42, 46, 75, 81, 70, 47, 31, 0, 0, 0, 0, 20, 
    87, 76, 45, 0, 27, 23, 0, 0, 0, 30, 55, 71, 59, 72, 45, 
    0, 0, 21, 18, 19, 0, 0, 23, 65, 51, 20, 0, 0, 0, 0, 
    0, 9, 0, 0, 13, 42, 45, 30, 0, 14, 18, 34, 47, 65, 50, 
    24, 72, 72, 70, 63, 54, 49, 29, 30, 21, 32, 27, 5, 4, 8, 
    38, 34, 47, 58, 65, 69, 71, 66, 60, 54, 35, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 21, 14, 0, 0, 0, 35, 16, 31, 60, 45, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 55, 71, 27, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 2, 0, 0, 0, 
    
    -- channel=123
    22, 21, 21, 21, 21, 21, 21, 21, 21, 22, 23, 21, 21, 21, 21, 
    22, 22, 22, 22, 22, 22, 22, 21, 22, 32, 25, 21, 22, 21, 22, 
    23, 22, 21, 21, 21, 23, 23, 30, 37, 30, 30, 23, 22, 22, 22, 
    24, 25, 22, 21, 22, 23, 21, 20, 17, 16, 12, 21, 25, 24, 23, 
    48, 44, 21, 21, 23, 15, 16, 18, 23, 32, 44, 46, 45, 32, 24, 
    5, 5, 19, 29, 29, 50, 47, 43, 35, 24, 13, 7, 4, 13, 25, 
    51, 46, 35, 14, 18, 24, 9, 1, 14, 31, 41, 44, 36, 39, 38, 
    5, 0, 13, 17, 15, 0, 0, 29, 34, 27, 17, 7, 5, 3, 21, 
    0, 9, 1, 8, 26, 33, 38, 30, 24, 37, 34, 41, 43, 44, 34, 
    35, 55, 59, 60, 57, 52, 45, 39, 39, 36, 39, 32, 25, 22, 18, 
    17, 15, 29, 35, 37, 44, 53, 53, 46, 42, 34, 25, 17, 10, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=124
    49, 48, 48, 48, 49, 49, 49, 49, 48, 50, 50, 48, 48, 48, 48, 
    50, 49, 49, 49, 49, 49, 49, 48, 50, 61, 54, 49, 49, 49, 49, 
    51, 51, 49, 49, 49, 51, 50, 57, 65, 56, 54, 50, 49, 49, 49, 
    46, 48, 48, 49, 50, 54, 49, 48, 33, 28, 21, 39, 48, 48, 48, 
    82, 77, 50, 50, 51, 42, 39, 44, 45, 56, 67, 74, 79, 60, 49, 
    11, 11, 42, 60, 63, 81, 82, 76, 62, 46, 28, 17, 15, 26, 48, 
    86, 79, 66, 35, 38, 42, 23, 17, 30, 58, 72, 78, 69, 72, 67, 
    21, 11, 39, 48, 43, 7, 5, 48, 66, 55, 39, 24, 19, 16, 34, 
    1, 28, 10, 24, 47, 57, 66, 51, 41, 52, 51, 59, 64, 70, 61, 
    54, 84, 87, 87, 83, 74, 66, 57, 58, 53, 58, 50, 41, 37, 37, 
    46, 47, 60, 68, 73, 80, 86, 81, 73, 67, 56, 45, 34, 27, 28, 
    6, 11, 2, 1, 2, 9, 0, 0, 7, 7, 2, 14, 28, 31, 16, 
    0, 5, 18, 13, 0, 0, 41, 52, 45, 48, 52, 38, 14, 14, 20, 
    0, 0, 0, 0, 0, 0, 2, 27, 41, 19, 0, 0, 16, 20, 28, 
    1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 11, 16, 14, 19, 27, 
    
    -- channel=125
    28, 29, 29, 29, 28, 29, 29, 30, 30, 27, 25, 28, 29, 29, 29, 
    28, 28, 28, 28, 28, 28, 28, 29, 26, 19, 16, 26, 28, 28, 28, 
    28, 29, 29, 29, 29, 28, 26, 21, 9, 5, 6, 19, 28, 29, 28, 
    17, 20, 26, 30, 29, 29, 24, 25, 13, 9, 5, 9, 22, 24, 26, 
    0, 0, 17, 30, 28, 32, 27, 29, 21, 14, 7, 1, 0, 10, 23, 
    12, 14, 24, 23, 19, 13, 5, 9, 14, 17, 12, 14, 14, 9, 22, 
    0, 0, 4, 13, 19, 0, 0, 0, 7, 22, 15, 11, 14, 10, 6, 
    0, 0, 5, 17, 20, 18, 17, 14, 3, 0, 0, 0, 0, 5, 1, 
    0, 26, 13, 21, 15, 13, 8, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    5, 4, 13, 7, 4, 0, 0, 0, 0, 0, 0, 8, 18, 15, 18, 
    12, 1, 13, 13, 7, 6, 23, 78, 79, 66, 43, 30, 24, 22, 16, 
    15, 8, 8, 8, 8, 8, 19, 100, 83, 47, 35, 30, 24, 18, 17, 
    19, 16, 11, 9, 11, 9, 4, 42, 38, 40, 35, 22, 22, 19, 16, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 
    0, 1, 0, 21, 0, 39, 5, 14, 9, 0, 0, 0, 0, 0, 5, 
    27, 0, 5, 0, 0, 18, 4, 0, 0, 0, 3, 4, 5, 0, 2, 
    72, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    8, 8, 0, 0, 0, 11, 0, 1, 0, 6, 11, 0, 0, 0, 3, 
    0, 6, 0, 0, 6, 1, 0, 1, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 1, 1, 0, 39, 0, 0, 11, 16, 0, 0, 2, 0, 
    1, 2, 0, 1, 2, 2, 15, 0, 22, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 12, 0, 0, 0, 0, 
    36, 27, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 4, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 0, 0, 0, 0, 
    16, 35, 1, 0, 0, 41, 55, 69, 0, 0, 0, 0, 0, 0, 2, 
    21, 0, 19, 10, 23, 0, 0, 0, 25, 54, 54, 41, 32, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 4, 9, 16, 21, 27, 27, 12, 12, 5, 12, 0, 0, 0, 
    27, 37, 21, 14, 6, 4, 0, 0, 0, 7, 7, 10, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 33, 23, 31, 24, 12, 0, 0, 9, 1, 
    0, 0, 11, 8, 2, 0, 0, 0, 0, 0, 0, 40, 7, 0, 0, 
    0, 0, 1, 3, 0, 0, 0, 0, 7, 50, 14, 0, 0, 0, 0, 
    10, 2, 2, 4, 5, 6, 11, 45, 12, 0, 0, 1, 0, 0, 0, 
    
    -- channel=128
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 2, 0, 0, 3, 
    0, 0, 4, 0, 0, 0, 0, 0, 1, 0, 19, 10, 0, 0, 7, 
    0, 0, 12, 0, 1, 0, 0, 0, 6, 0, 32, 13, 0, 2, 9, 
    0, 9, 7, 17, 3, 7, 0, 0, 0, 0, 0, 0, 27, 3, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 19, 0, 0, 
    6, 0, 0, 10, 0, 0, 0, 0, 0, 0, 29, 28, 0, 25, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 24, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 13, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    
    -- channel=130
    0, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 
    0, 5, 10, 0, 0, 0, 0, 1, 4, 0, 52, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 45, 44, 59, 0, 0, 
    17, 19, 24, 30, 16, 16, 14, 0, 0, 2, 19, 16, 13, 0, 21, 
    40, 22, 0, 33, 26, 16, 12, 0, 11, 14, 36, 11, 0, 38, 0, 
    24, 12, 14, 44, 34, 12, 17, 13, 17, 15, 26, 3, 0, 0, 0, 
    11, 9, 10, 4, 3, 0, 0, 0, 0, 0, 32, 20, 0, 0, 27, 
    2, 8, 37, 16, 0, 0, 10, 15, 15, 0, 15, 0, 1, 0, 0, 
    14, 27, 7, 4, 19, 11, 0, 0, 9, 10, 3, 0, 0, 0, 19, 
    28, 10, 4, 0, 9, 26, 0, 10, 47, 14, 0, 4, 7, 14, 11, 
    51, 16, 0, 24, 33, 35, 0, 0, 21, 20, 9, 22, 19, 21, 20, 
    29, 2, 0, 7, 20, 31, 24, 16, 14, 24, 20, 24, 10, 26, 26, 
    30, 33, 30, 30, 22, 25, 31, 27, 40, 1, 25, 22, 24, 28, 23, 
    26, 32, 34, 35, 32, 26, 24, 17, 50, 0, 27, 24, 27, 31, 8, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 15, 24, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 1, 24, 22, 19, 24, 28, 11, 6, 4, 
    18, 15, 23, 24, 13, 8, 6, 4, 43, 40, 15, 59, 66, 38, 38, 
    58, 45, 47, 55, 61, 60, 52, 40, 15, 2, 5, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 25, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 21, 26, 10, 3, 0, 0, 
    15, 28, 10, 1, 11, 22, 14, 0, 0, 0, 0, 0, 1, 5, 23, 
    0, 0, 0, 4, 0, 0, 0, 22, 32, 3, 0, 13, 35, 41, 33, 
    3, 0, 2, 21, 36, 22, 7, 13, 2, 26, 41, 36, 27, 19, 17, 
    0, 4, 1, 1, 0, 0, 34, 17, 7, 12, 23, 16, 5, 9, 8, 
    21, 39, 43, 30, 25, 24, 11, 7, 24, 19, 8, 8, 12, 3, 0, 
    19, 22, 13, 10, 15, 18, 12, 8, 0, 0, 8, 4, 3, 0, 0, 
    2, 0, 0, 0, 0, 0, 1, 11, 9, 9, 2, 2, 0, 0, 8, 
    
    -- channel=132
    15, 27, 43, 37, 43, 42, 49, 43, 52, 51, 44, 54, 47, 52, 54, 
    14, 27, 44, 34, 45, 37, 41, 47, 50, 11, 36, 59, 44, 50, 53, 
    16, 24, 45, 36, 44, 38, 30, 27, 40, 0, 40, 51, 35, 43, 52, 
    13, 20, 31, 38, 35, 38, 29, 22, 0, 0, 0, 0, 20, 31, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 27, 0, 0, 
    0, 5, 0, 3, 16, 8, 12, 0, 0, 0, 29, 59, 0, 35, 0, 
    0, 0, 0, 5, 5, 5, 6, 8, 14, 14, 36, 27, 11, 0, 0, 
    9, 17, 37, 41, 35, 30, 25, 12, 13, 0, 3, 21, 20, 0, 14, 
    0, 0, 3, 18, 9, 1, 0, 0, 15, 14, 39, 25, 15, 8, 9, 
    0, 23, 23, 0, 2, 15, 18, 2, 7, 18, 18, 5, 0, 0, 0, 
    11, 4, 0, 0, 0, 8, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=133
    3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 0, 0, 
    5, 17, 11, 0, 25, 14, 9, 0, 0, 7, 29, 64, 23, 2, 1, 
    3, 0, 0, 0, 0, 4, 11, 25, 37, 29, 21, 0, 0, 0, 0, 
    24, 35, 60, 56, 32, 19, 13, 0, 0, 0, 0, 0, 0, 7, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 36, 3, 0, 0, 0, 
    0, 34, 21, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    13, 17, 21, 23, 23, 24, 28, 25, 29, 28, 26, 29, 28, 31, 27, 
    14, 16, 22, 24, 24, 25, 23, 18, 28, 26, 0, 26, 28, 27, 26, 
    15, 15, 23, 24, 31, 22, 23, 11, 8, 5, 2, 14, 20, 20, 25, 
    8, 8, 21, 8, 21, 19, 15, 29, 1, 0, 0, 0, 0, 9, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 37, 6, 0, 
    0, 5, 9, 0, 11, 8, 8, 0, 0, 0, 7, 48, 50, 0, 17, 
    6, 0, 0, 0, 0, 0, 5, 6, 21, 20, 35, 23, 0, 24, 0, 
    6, 10, 20, 39, 24, 21, 17, 19, 4, 6, 0, 0, 7, 0, 13, 
    0, 0, 0, 0, 6, 0, 0, 0, 9, 6, 36, 22, 6, 8, 4, 
    0, 10, 23, 4, 0, 10, 19, 14, 0, 1, 11, 8, 0, 0, 0, 
    0, 3, 2, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    29, 0, 23, 26, 31, 28, 37, 44, 35, 41, 40, 37, 33, 42, 29, 
    31, 4, 27, 30, 39, 31, 43, 45, 35, 60, 7, 37, 35, 47, 29, 
    37, 4, 29, 31, 47, 33, 52, 42, 34, 59, 15, 48, 45, 47, 34, 
    47, 7, 51, 43, 53, 38, 47, 50, 37, 2, 0, 0, 33, 65, 41, 
    28, 15, 21, 31, 36, 39, 29, 44, 14, 21, 9, 0, 22, 34, 14, 
    0, 0, 27, 0, 4, 3, 19, 19, 14, 11, 0, 20, 29, 39, 14, 
    12, 3, 2, 0, 0, 0, 0, 0, 0, 0, 8, 32, 36, 43, 15, 
    0, 0, 4, 13, 18, 19, 22, 28, 31, 44, 16, 21, 25, 0, 0, 
    20, 24, 0, 14, 28, 30, 18, 5, 8, 21, 16, 24, 21, 26, 46, 
    0, 0, 25, 18, 0, 10, 29, 46, 27, 25, 23, 39, 42, 30, 11, 
    9, 10, 18, 31, 36, 19, 29, 0, 0, 40, 38, 23, 21, 12, 24, 
    6, 7, 18, 0, 0, 17, 45, 25, 10, 11, 24, 9, 4, 5, 0, 
    21, 34, 36, 24, 14, 1, 0, 15, 21, 10, 3, 6, 10, 0, 0, 
    0, 0, 0, 2, 15, 13, 1, 2, 0, 17, 2, 1, 0, 0, 2, 
    1, 0, 0, 0, 0, 3, 8, 12, 0, 5, 1, 0, 0, 0, 14, 
    
    -- channel=136
    36, 0, 20, 28, 35, 33, 36, 47, 29, 38, 37, 36, 41, 43, 34, 
    37, 1, 18, 33, 34, 33, 34, 37, 30, 48, 0, 29, 42, 42, 33, 
    38, 0, 15, 36, 33, 32, 40, 13, 10, 66, 0, 10, 42, 35, 25, 
    32, 2, 17, 24, 33, 26, 36, 27, 7, 7, 0, 0, 0, 18, 6, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 32, 0, 
    0, 0, 6, 0, 1, 0, 0, 4, 0, 0, 0, 17, 48, 3, 10, 
    0, 0, 0, 0, 0, 11, 10, 14, 13, 12, 0, 15, 45, 0, 14, 
    1, 11, 5, 6, 12, 15, 17, 17, 8, 24, 0, 1, 17, 43, 17, 
    0, 0, 0, 1, 9, 5, 7, 13, 3, 35, 4, 12, 13, 14, 5, 
    10, 0, 0, 5, 6, 7, 10, 6, 0, 9, 12, 15, 2, 0, 0, 
    0, 2, 2, 2, 0, 0, 21, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=137
    17, 15, 25, 18, 22, 15, 16, 12, 14, 18, 11, 13, 6, 12, 9, 
    12, 13, 20, 13, 18, 10, 18, 19, 11, 12, 22, 15, 6, 15, 11, 
    10, 6, 16, 5, 11, 7, 12, 17, 23, 0, 41, 32, 14, 15, 14, 
    15, 11, 25, 22, 10, 10, 2, 11, 11, 10, 5, 19, 60, 30, 20, 
    32, 23, 21, 29, 30, 30, 26, 21, 16, 13, 12, 3, 0, 1, 12, 
    4, 0, 2, 0, 0, 0, 15, 13, 12, 6, 0, 0, 0, 10, 0, 
    11, 9, 3, 12, 12, 4, 0, 0, 0, 0, 8, 6, 0, 0, 0, 
    4, 0, 3, 5, 14, 15, 18, 20, 28, 17, 21, 11, 1, 0, 0, 
    30, 28, 28, 32, 30, 33, 24, 10, 6, 0, 0, 0, 4, 7, 7, 
    0, 18, 20, 19, 18, 14, 17, 25, 26, 16, 9, 15, 18, 14, 11, 
    36, 18, 25, 29, 38, 36, 13, 0, 11, 29, 25, 15, 13, 4, 7, 
    29, 21, 13, 4, 3, 24, 26, 18, 9, 9, 13, 5, 0, 2, 0, 
    31, 36, 33, 28, 21, 14, 10, 11, 14, 10, 4, 5, 0, 0, 0, 
    9, 12, 9, 10, 11, 10, 6, 3, 2, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 2, 10, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    75, 76, 93, 88, 96, 92, 93, 91, 91, 94, 81, 97, 95, 96, 98, 
    69, 70, 84, 83, 87, 80, 78, 84, 87, 43, 61, 93, 90, 88, 96, 
    65, 59, 77, 82, 77, 77, 64, 40, 61, 23, 44, 60, 73, 73, 84, 
    44, 56, 48, 60, 56, 68, 58, 53, 0, 0, 0, 0, 0, 33, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 18, 14, 62, 35, 28, 0, 
    31, 33, 24, 35, 56, 43, 40, 23, 24, 35, 78, 109, 57, 42, 10, 
    20, 16, 7, 29, 41, 61, 65, 76, 81, 72, 75, 49, 54, 0, 0, 
    58, 75, 94, 93, 84, 80, 76, 58, 46, 11, 13, 40, 49, 48, 88, 
    24, 1, 37, 59, 46, 31, 32, 48, 58, 72, 74, 54, 45, 43, 10, 
    49, 71, 55, 33, 56, 68, 59, 24, 19, 48, 51, 32, 0, 0, 0, 
    48, 48, 41, 20, 1, 32, 18, 0, 21, 8, 0, 0, 0, 0, 0, 
    25, 34, 17, 11, 31, 26, 3, 11, 5, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=140
    0, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 6, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    0, 11, 9, 0, 0, 0, 0, 0, 3, 0, 64, 2, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 37, 0, 1, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 10, 23, 0, 8, 
    13, 16, 0, 6, 1, 1, 0, 0, 0, 0, 34, 15, 0, 2, 0, 
    7, 0, 0, 25, 11, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 
    0, 0, 5, 11, 0, 0, 0, 0, 0, 0, 9, 5, 0, 0, 3, 
    0, 0, 19, 2, 0, 0, 0, 0, 4, 0, 19, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 1, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    0, 3, 2, 3, 2, 1, 0, 0, 33, 0, 0, 0, 0, 2, 0, 
    
    -- channel=141
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 2, 2, 
    0, 0, 2, 9, 6, 5, 0, 0, 0, 0, 0, 0, 18, 2, 5, 
    0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 14, 6, 0, 2, 3, 
    0, 0, 0, 0, 4, 4, 2, 9, 11, 0, 12, 12, 6, 10, 9, 
    0, 0, 9, 17, 16, 12, 8, 0, 5, 5, 0, 17, 35, 21, 25, 
    14, 13, 17, 25, 29, 28, 20, 2, 0, 0, 0, 0, 0, 9, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 5, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=143
    64, 50, 57, 54, 49, 41, 38, 39, 35, 36, 35, 32, 33, 35, 31, 
    53, 38, 43, 38, 36, 31, 32, 37, 32, 37, 29, 30, 29, 33, 26, 
    43, 29, 29, 25, 24, 25, 28, 30, 30, 45, 24, 37, 28, 25, 24, 
    35, 17, 19, 18, 15, 16, 24, 23, 37, 48, 29, 19, 34, 24, 14, 
    36, 25, 27, 22, 23, 25, 34, 50, 48, 44, 43, 19, 9, 7, 5, 
    34, 28, 35, 29, 31, 33, 50, 55, 43, 41, 25, 16, 0, 18, 17, 
    43, 34, 41, 39, 47, 51, 52, 49, 39, 36, 15, 15, 25, 4, 21, 
    51, 43, 48, 51, 58, 60, 61, 55, 56, 41, 23, 14, 19, 18, 0, 
    59, 62, 54, 64, 66, 68, 60, 48, 35, 36, 15, 20, 26, 20, 23, 
    54, 51, 61, 59, 58, 50, 48, 46, 47, 40, 32, 32, 33, 29, 21, 
    68, 63, 58, 60, 57, 58, 49, 38, 22, 39, 41, 38, 31, 28, 20, 
    52, 57, 57, 46, 42, 39, 55, 41, 31, 32, 33, 35, 23, 22, 17, 
    47, 55, 58, 47, 40, 35, 33, 30, 34, 33, 26, 22, 26, 19, 19, 
    24, 26, 26, 26, 27, 28, 28, 25, 25, 24, 23, 18, 20, 18, 15, 
    14, 13, 16, 17, 20, 21, 24, 20, 18, 27, 18, 17, 18, 18, 11, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 37, 64, 50, 69, 12, 0, 0, 
    29, 24, 38, 28, 32, 23, 25, 18, 0, 0, 0, 0, 0, 23, 31, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 13, 1, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 3, 0, 20, 0, 
    0, 6, 10, 0, 0, 0, 12, 12, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 1, 8, 0, 0, 0, 0, 0, 0, 0, 1, 21, 23, 
    0, 0, 0, 0, 0, 1, 15, 37, 9, 0, 9, 24, 9, 7, 0, 
    0, 1, 15, 25, 9, 0, 0, 0, 2, 12, 1, 15, 9, 6, 10, 
    0, 0, 0, 0, 12, 28, 11, 0, 0, 15, 5, 0, 6, 2, 0, 
    21, 20, 10, 0, 0, 1, 12, 12, 0, 0, 6, 2, 3, 0, 0, 
    0, 0, 2, 3, 0, 0, 0, 1, 0, 11, 0, 2, 0, 0, 4, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 3, 0, 1, 
    2, 0, 0, 9, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=147
    68, 21, 49, 50, 55, 46, 51, 64, 45, 52, 46, 49, 52, 59, 44, 
    63, 18, 40, 47, 52, 44, 48, 54, 43, 66, 4, 41, 49, 56, 38, 
    59, 10, 31, 47, 50, 43, 58, 25, 17, 82, 0, 21, 48, 47, 34, 
    45, 2, 23, 23, 38, 32, 47, 47, 21, 23, 1, 0, 0, 29, 4, 
    0, 0, 3, 0, 0, 0, 0, 30, 23, 27, 17, 17, 5, 46, 0, 
    16, 8, 38, 10, 40, 25, 28, 35, 23, 31, 11, 51, 67, 40, 25, 
    21, 15, 18, 4, 21, 42, 46, 50, 52, 50, 22, 27, 60, 1, 13, 
    35, 43, 44, 42, 45, 46, 49, 44, 35, 45, 5, 16, 28, 58, 51, 
    25, 18, 5, 31, 37, 32, 35, 42, 30, 62, 31, 30, 31, 31, 19, 
    38, 28, 36, 33, 33, 42, 40, 30, 10, 34, 32, 35, 20, 15, 0, 
    23, 37, 34, 31, 10, 16, 53, 23, 0, 18, 16, 18, 14, 9, 11, 
    6, 26, 50, 21, 23, 9, 32, 19, 9, 15, 11, 13, 13, 5, 7, 
    0, 9, 16, 7, 4, 5, 10, 11, 5, 8, 10, 0, 12, 2, 4, 
    0, 0, 0, 0, 1, 0, 1, 9, 0, 23, 5, 2, 3, 2, 4, 
    1, 0, 2, 2, 5, 6, 5, 9, 0, 23, 3, 0, 0, 1, 12, 
    
    -- channel=148
    0, 20, 2, 1, 0, 6, 3, 0, 9, 3, 5, 7, 4, 0, 12, 
    0, 24, 11, 3, 0, 6, 1, 0, 10, 0, 32, 12, 5, 0, 17, 
    0, 30, 18, 5, 3, 4, 0, 10, 19, 0, 50, 17, 0, 1, 17, 
    0, 33, 14, 11, 2, 10, 0, 0, 0, 0, 17, 34, 25, 2, 27, 
    0, 11, 1, 16, 5, 10, 3, 0, 0, 0, 0, 14, 34, 0, 24, 
    5, 18, 0, 12, 0, 6, 0, 0, 0, 0, 32, 11, 0, 0, 0, 
    3, 2, 0, 17, 6, 0, 0, 0, 0, 0, 34, 17, 0, 25, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 17, 15, 3, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 10, 0, 20, 9, 2, 1, 1, 
    0, 7, 0, 0, 0, 0, 0, 0, 5, 0, 4, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 2, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 21, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    4, 2, 0, 6, 2, 2, 2, 0, 11, 0, 0, 1, 0, 3, 3, 
    0, 6, 5, 7, 4, 4, 3, 0, 26, 0, 3, 0, 3, 5, 0, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 3, 0, 1, 0, 0, 0, 4, 6, 0, 22, 0, 0, 
    7, 4, 7, 8, 5, 0, 4, 0, 2, 0, 4, 10, 0, 8, 4, 
    12, 0, 2, 10, 0, 0, 0, 0, 0, 0, 4, 2, 0, 14, 0, 
    5, 4, 10, 14, 4, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 10, 
    0, 4, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    1, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 
    9, 0, 0, 0, 0, 6, 0, 4, 5, 0, 0, 1, 1, 8, 8, 
    11, 4, 1, 7, 4, 0, 0, 3, 6, 2, 0, 10, 9, 12, 13, 
    9, 4, 5, 8, 8, 7, 5, 1, 5, 10, 10, 12, 10, 14, 14, 
    14, 14, 10, 9, 7, 9, 9, 9, 15, 0, 16, 14, 14, 15, 15, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 25, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 16, 0, 
    14, 0, 0, 11, 19, 8, 0, 0, 0, 0, 13, 4, 14, 0, 0, 
    0, 0, 0, 8, 15, 17, 23, 26, 33, 24, 8, 0, 0, 0, 0, 
    1, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 66, 
    0, 0, 7, 0, 0, 0, 0, 15, 7, 3, 2, 0, 0, 0, 0, 
    29, 4, 0, 0, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 18, 23, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 0, 0, 0, 0, 0, 3, 6, 0, 0, 0, 0, 1, 0, 
    0, 3, 6, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=152
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 6, 2, 
    35, 32, 13, 2, 0, 3, 3, 0, 0, 0, 1, 4, 6, 2, 1, 
    9, 7, 3, 0, 0, 0, 0, 5, 5, 0, 7, 6, 7, 2, 24, 
    
    -- channel=153
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 10, 0, 0, 65, 0, 0, 1, 0, 0, 
    15, 0, 0, 0, 4, 0, 8, 20, 46, 9, 0, 16, 0, 0, 0, 
    4, 5, 7, 4, 4, 6, 0, 23, 0, 11, 0, 0, 0, 13, 10, 
    0, 0, 16, 0, 0, 1, 0, 11, 0, 0, 0, 0, 49, 0, 59, 
    0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 53, 36, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 38, 0, 0, 0, 23, 0, 
    10, 5, 0, 0, 7, 3, 0, 0, 0, 0, 0, 2, 0, 8, 14, 
    0, 0, 0, 7, 0, 0, 0, 21, 0, 0, 0, 19, 27, 27, 1, 
    0, 0, 0, 14, 7, 0, 26, 15, 0, 4, 18, 16, 15, 6, 25, 
    0, 0, 21, 0, 0, 0, 25, 6, 0, 3, 20, 1, 12, 10, 10, 
    0, 13, 15, 7, 6, 0, 0, 5, 15, 1, 3, 1, 18, 3, 4, 
    9, 0, 0, 0, 5, 4, 0, 4, 0, 34, 1, 10, 3, 1, 5, 
    4, 0, 0, 0, 0, 0, 6, 13, 0, 27, 6, 5, 3, 0, 38, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 
    19, 7, 0, 8, 12, 0, 0, 0, 0, 0, 34, 36, 0, 47, 0, 
    9, 0, 0, 15, 10, 0, 0, 0, 5, 9, 29, 0, 0, 0, 0, 
    2, 3, 22, 17, 6, 0, 0, 0, 0, 0, 2, 3, 0, 0, 22, 
    0, 0, 7, 2, 0, 0, 0, 0, 3, 0, 22, 0, 0, 0, 0, 
    0, 27, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 1, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 
    0, 2, 2, 2, 3, 1, 0, 0, 22, 0, 0, 0, 0, 4, 0, 
    
    -- channel=156
    13, 0, 3, 0, 6, 0, 6, 19, 2, 6, 5, 9, 0, 12, 0, 
    10, 0, 1, 0, 14, 0, 7, 24, 0, 5, 0, 6, 0, 15, 0, 
    14, 0, 0, 6, 12, 6, 16, 0, 0, 33, 0, 11, 12, 19, 1, 
    19, 0, 0, 18, 17, 10, 21, 8, 0, 8, 0, 0, 18, 21, 0, 
    5, 0, 0, 0, 0, 0, 0, 15, 9, 0, 0, 0, 0, 11, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 8, 0, 16, 0, 54, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 12, 
    0, 0, 6, 0, 0, 0, 0, 0, 7, 1, 0, 2, 2, 19, 7, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 29, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 2, 0, 0, 0, 4, 11, 0, 2, 1, 2, 0, 
    12, 0, 0, 1, 0, 14, 3, 0, 0, 0, 2, 6, 1, 3, 0, 
    0, 0, 3, 0, 0, 0, 18, 11, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=157
    20, 0, 0, 0, 0, 0, 0, 14, 0, 0, 4, 0, 8, 5, 0, 
    20, 0, 0, 3, 0, 3, 0, 0, 0, 37, 0, 0, 10, 5, 0, 
    22, 0, 0, 8, 0, 5, 17, 0, 0, 75, 0, 0, 12, 0, 0, 
    20, 0, 0, 0, 7, 0, 17, 20, 18, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 6, 6, 0, 0, 0, 24, 0, 
    0, 0, 19, 0, 3, 1, 0, 12, 0, 2, 0, 0, 63, 0, 44, 
    0, 0, 5, 0, 0, 6, 4, 11, 9, 7, 0, 0, 40, 8, 43, 
    0, 6, 0, 0, 0, 0, 0, 6, 0, 28, 0, 0, 7, 65, 20, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 30, 0, 4, 5, 12, 1, 
    11, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 13, 9, 14, 0, 
    0, 0, 0, 4, 0, 0, 27, 16, 0, 0, 0, 8, 7, 4, 10, 
    0, 0, 23, 1, 0, 0, 15, 5, 0, 0, 3, 2, 8, 3, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 14, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 2, 2, 0, 2, 
    1, 0, 0, 0, 0, 0, 0, 7, 0, 31, 0, 1, 0, 0, 26, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    68, 43, 50, 54, 51, 48, 44, 51, 39, 43, 44, 39, 46, 45, 41, 
    62, 36, 40, 47, 42, 42, 40, 43, 38, 56, 26, 35, 45, 43, 36, 
    54, 30, 29, 39, 34, 37, 43, 32, 28, 74, 2, 27, 42, 35, 30, 
    45, 22, 22, 24, 29, 26, 40, 35, 45, 62, 34, 24, 6, 22, 16, 
    33, 26, 32, 18, 25, 22, 32, 50, 47, 43, 37, 27, 11, 34, 15, 
    31, 27, 40, 32, 39, 40, 42, 54, 41, 42, 22, 25, 41, 21, 43, 
    36, 38, 45, 29, 44, 57, 59, 60, 52, 46, 16, 25, 51, 19, 44, 
    50, 49, 47, 46, 52, 55, 56, 53, 47, 50, 20, 22, 34, 61, 34, 
    48, 50, 41, 52, 58, 56, 53, 52, 39, 53, 22, 31, 37, 34, 28, 
    66, 41, 47, 55, 55, 48, 43, 39, 33, 38, 37, 41, 36, 38, 25, 
    46, 56, 52, 51, 38, 39, 57, 54, 19, 28, 38, 44, 33, 31, 24, 
    29, 50, 63, 52, 46, 25, 49, 37, 29, 35, 32, 34, 31, 25, 28, 
    25, 37, 45, 34, 34, 35, 36, 29, 27, 32, 30, 19, 33, 24, 24, 
    27, 27, 27, 22, 22, 22, 27, 29, 20, 34, 26, 24, 26, 22, 21, 
    21, 18, 20, 21, 23, 22, 23, 24, 6, 42, 22, 24, 22, 21, 27, 
    
    -- channel=160
    0, 26, 18, 0, 0, 0, 1, 0, 11, 0, 0, 4, 0, 0, 7, 
    0, 26, 24, 0, 2, 0, 0, 0, 7, 0, 52, 16, 0, 0, 11, 
    0, 24, 28, 0, 0, 0, 0, 12, 26, 0, 91, 39, 0, 0, 18, 
    0, 23, 13, 17, 0, 5, 0, 0, 0, 0, 17, 26, 92, 9, 32, 
    8, 16, 7, 33, 15, 21, 12, 0, 0, 0, 10, 14, 32, 0, 13, 
    21, 16, 0, 21, 0, 0, 0, 0, 0, 0, 47, 20, 0, 33, 0, 
    11, 0, 0, 39, 20, 0, 0, 0, 0, 0, 41, 11, 0, 0, 0, 
    0, 0, 5, 7, 3, 0, 0, 0, 2, 0, 39, 24, 0, 0, 0, 
    0, 3, 38, 18, 0, 0, 0, 0, 8, 0, 18, 0, 0, 0, 0, 
    0, 24, 9, 0, 3, 0, 0, 0, 19, 5, 0, 0, 0, 0, 4, 
    29, 0, 0, 0, 13, 31, 0, 0, 44, 13, 0, 0, 0, 0, 0, 
    55, 3, 0, 0, 5, 37, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    36, 1, 0, 2, 4, 6, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    5, 8, 4, 12, 4, 5, 5, 0, 26, 0, 0, 0, 0, 1, 0, 
    0, 5, 3, 4, 3, 1, 0, 0, 49, 0, 2, 0, 1, 7, 0, 
    
    -- channel=161
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=162
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=163
    55, 28, 37, 41, 38, 33, 31, 38, 26, 30, 32, 26, 31, 31, 23, 
    52, 24, 29, 37, 32, 31, 30, 29, 24, 53, 9, 19, 31, 30, 21, 
    46, 18, 20, 29, 27, 25, 35, 23, 18, 71, 0, 17, 34, 26, 17, 
    36, 10, 16, 13, 21, 17, 27, 29, 43, 42, 25, 25, 0, 19, 11, 
    23, 16, 18, 8, 12, 12, 16, 38, 32, 32, 25, 6, 1, 29, 5, 
    10, 8, 29, 9, 13, 15, 23, 38, 28, 28, 2, 4, 37, 0, 28, 
    23, 26, 28, 12, 24, 35, 36, 34, 29, 29, 7, 17, 28, 10, 37, 
    26, 23, 14, 20, 29, 36, 41, 45, 38, 51, 14, 5, 14, 35, 4, 
    37, 39, 25, 34, 45, 48, 49, 41, 25, 32, 3, 14, 20, 21, 17, 
    40, 16, 31, 44, 40, 35, 35, 38, 26, 26, 23, 30, 32, 32, 16, 
    32, 41, 41, 43, 35, 31, 53, 41, 8, 25, 35, 36, 27, 21, 19, 
    21, 40, 55, 36, 26, 17, 42, 29, 23, 27, 29, 29, 23, 19, 16, 
    19, 37, 42, 31, 35, 32, 23, 22, 25, 27, 23, 16, 23, 13, 10, 
    25, 23, 21, 16, 18, 20, 21, 24, 6, 28, 17, 14, 14, 11, 12, 
    10, 7, 12, 12, 13, 14, 17, 20, 0, 33, 11, 11, 11, 9, 20, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 6, 19, 4, 13, 0, 0, 0, 
    10, 6, 3, 9, 0, 0, 0, 0, 38, 51, 23, 52, 48, 16, 20, 
    53, 43, 39, 39, 46, 43, 42, 33, 22, 7, 13, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 
    0, 10, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 19, 23, 0, 0, 0, 0, 
    13, 38, 18, 7, 11, 27, 24, 5, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 11, 9, 0, 0, 12, 31, 1, 0, 3, 27, 37, 32, 
    18, 1, 6, 23, 32, 30, 13, 27, 4, 14, 37, 37, 26, 21, 15, 
    4, 14, 15, 18, 0, 0, 31, 22, 13, 15, 21, 26, 9, 15, 15, 
    17, 39, 46, 35, 36, 33, 18, 8, 23, 28, 14, 10, 19, 10, 5, 
    29, 32, 22, 14, 15, 21, 21, 15, 0, 0, 15, 9, 11, 3, 2, 
    8, 3, 2, 0, 0, 0, 5, 14, 11, 18, 7, 9, 6, 5, 12, 
    
    -- channel=165
    28, 27, 41, 44, 50, 50, 55, 53, 54, 60, 56, 57, 54, 57, 57, 
    30, 30, 44, 46, 51, 50, 56, 56, 54, 52, 49, 61, 57, 60, 59, 
    34, 30, 45, 45, 50, 49, 50, 50, 55, 34, 43, 61, 56, 56, 59, 
    41, 35, 55, 58, 55, 52, 45, 42, 30, 13, 5, 16, 51, 56, 56, 
    29, 23, 26, 36, 42, 45, 42, 31, 13, 5, 2, 2, 16, 25, 29, 
    0, 0, 3, 0, 6, 6, 16, 8, 4, 1, 0, 20, 11, 28, 4, 
    2, 0, 0, 5, 14, 10, 7, 0, 0, 0, 18, 38, 31, 29, 9, 
    4, 4, 12, 18, 25, 26, 26, 26, 29, 21, 23, 35, 35, 1, 0, 
    18, 17, 22, 31, 33, 29, 19, 12, 17, 13, 18, 28, 28, 26, 30, 
    0, 11, 20, 21, 15, 15, 22, 27, 25, 26, 29, 32, 26, 16, 8, 
    15, 13, 18, 19, 24, 23, 14, 0, 2, 25, 24, 12, 1, 0, 0, 
    8, 12, 5, 0, 0, 15, 19, 6, 0, 0, 0, 0, 0, 0, 0, 
    9, 15, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=166
    46, 30, 36, 36, 33, 27, 25, 26, 21, 25, 25, 18, 20, 22, 16, 
    37, 22, 26, 27, 23, 20, 23, 24, 19, 37, 10, 16, 19, 22, 13, 
    31, 18, 17, 15, 16, 15, 22, 25, 22, 41, 17, 30, 22, 17, 14, 
    31, 11, 22, 13, 13, 10, 17, 23, 37, 24, 12, 15, 24, 29, 14, 
    31, 21, 20, 22, 22, 25, 27, 43, 35, 36, 29, 3, 8, 2, 7, 
    12, 16, 28, 4, 8, 17, 37, 43, 30, 23, 0, 0, 1, 0, 16, 
    30, 22, 24, 17, 22, 23, 24, 17, 11, 14, 4, 10, 10, 20, 22, 
    29, 19, 23, 32, 38, 40, 43, 46, 45, 42, 11, 2, 9, 0, 0, 
    52, 50, 30, 43, 55, 56, 43, 24, 17, 16, 3, 12, 16, 17, 22, 
    21, 29, 47, 44, 31, 30, 37, 49, 38, 25, 20, 30, 35, 28, 15, 
    44, 43, 45, 53, 55, 40, 39, 20, 6, 38, 40, 31, 27, 20, 21, 
    33, 39, 42, 22, 16, 31, 53, 37, 22, 21, 32, 22, 15, 16, 8, 
    43, 55, 55, 44, 33, 21, 18, 26, 32, 23, 17, 17, 19, 10, 9, 
    17, 16, 17, 18, 23, 23, 17, 15, 6, 22, 13, 12, 10, 8, 9, 
    6, 4, 5, 5, 8, 12, 18, 16, 10, 19, 10, 8, 10, 8, 12, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=168
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 4, 11, 2, 0, 0, 
    2, 9, 9, 8, 2, 4, 0, 5, 6, 10, 11, 9, 6, 1, 22, 
    0, 1, 5, 0, 0, 2, 0, 9, 7, 6, 0, 0, 15, 0, 19, 
    6, 8, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 11, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 17, 1, 0, 0, 1, 3, 
    4, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 6, 14, 6, 
    0, 0, 0, 2, 2, 0, 7, 10, 1, 2, 8, 12, 8, 9, 15, 
    0, 0, 4, 2, 0, 0, 5, 6, 7, 6, 12, 9, 14, 12, 15, 
    0, 3, 8, 9, 10, 9, 8, 9, 16, 15, 12, 10, 14, 13, 12, 
    15, 14, 14, 13, 15, 15, 13, 13, 3, 21, 10, 12, 13, 13, 15, 
    
    -- channel=169
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 2, 0, 0, 
    4, 11, 8, 0, 24, 13, 4, 0, 0, 7, 25, 62, 29, 4, 0, 
    0, 0, 0, 0, 0, 2, 12, 25, 39, 32, 18, 0, 0, 0, 0, 
    20, 34, 55, 50, 26, 15, 10, 0, 0, 0, 0, 0, 0, 3, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 33, 1, 0, 0, 0, 
    0, 33, 12, 0, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=170
    11, 19, 29, 31, 37, 41, 48, 46, 51, 52, 49, 54, 50, 53, 52, 
    19, 27, 39, 40, 48, 47, 49, 47, 52, 41, 30, 56, 52, 55, 55, 
    28, 32, 48, 49, 58, 49, 49, 43, 45, 17, 39, 48, 49, 55, 58, 
    31, 37, 54, 51, 58, 56, 47, 48, 13, 0, 0, 0, 19, 50, 54, 
    0, 8, 4, 18, 16, 21, 12, 0, 0, 4, 1, 16, 50, 38, 26, 
    2, 12, 13, 6, 18, 13, 9, 0, 4, 4, 21, 58, 51, 40, 22, 
    6, 1, 0, 5, 2, 0, 2, 1, 12, 17, 47, 50, 28, 47, 0, 
    2, 9, 17, 25, 19, 17, 14, 16, 14, 15, 21, 37, 36, 9, 30, 
    0, 0, 0, 4, 6, 1, 0, 3, 22, 19, 47, 39, 28, 31, 34, 
    0, 8, 14, 3, 0, 12, 22, 21, 12, 21, 28, 27, 19, 4, 4, 
    0, 0, 2, 0, 4, 1, 3, 0, 8, 20, 9, 0, 0, 0, 7, 
    4, 0, 0, 0, 0, 18, 0, 3, 7, 1, 1, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 6, 0, 0, 0, 0, 1, 
    0, 1, 0, 0, 0, 3, 1, 0, 9, 0, 0, 0, 0, 0, 0, 
    
    -- channel=171
    28, 0, 0, 0, 0, 0, 0, 12, 0, 0, 1, 0, 9, 3, 0, 
    28, 0, 0, 7, 0, 4, 0, 0, 0, 43, 0, 0, 11, 0, 0, 
    26, 0, 0, 8, 0, 3, 15, 0, 0, 83, 0, 0, 10, 0, 0, 
    15, 0, 0, 0, 0, 0, 10, 22, 27, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 10, 14, 0, 0, 0, 27, 0, 
    0, 0, 26, 0, 7, 14, 2, 19, 4, 10, 0, 0, 83, 0, 61, 
    0, 11, 12, 0, 0, 16, 16, 24, 27, 21, 0, 0, 29, 17, 52, 
    9, 15, 1, 4, 0, 5, 9, 18, 0, 36, 0, 0, 5, 74, 28, 
    3, 0, 0, 0, 4, 0, 1, 8, 0, 33, 0, 7, 6, 14, 0, 
    27, 0, 0, 8, 0, 4, 6, 9, 0, 0, 1, 14, 10, 16, 0, 
    0, 6, 6, 9, 0, 0, 38, 28, 0, 0, 1, 12, 12, 9, 13, 
    0, 0, 36, 13, 3, 0, 15, 8, 0, 5, 12, 8, 17, 10, 16, 
    0, 0, 0, 0, 0, 0, 1, 4, 4, 1, 11, 0, 20, 6, 10, 
    1, 0, 0, 0, 0, 0, 0, 9, 0, 38, 5, 9, 9, 6, 10, 
    7, 2, 5, 4, 4, 7, 7, 14, 0, 43, 5, 7, 6, 0, 33, 
    
    -- channel=172
    38, 56, 54, 43, 40, 34, 32, 21, 34, 30, 24, 26, 21, 25, 25, 
    31, 49, 47, 32, 33, 26, 28, 26, 29, 17, 41, 29, 18, 22, 27, 
    23, 41, 41, 21, 25, 19, 18, 30, 37, 0, 71, 43, 20, 22, 27, 
    17, 34, 31, 20, 11, 17, 6, 20, 29, 14, 51, 53, 57, 27, 27, 
    33, 39, 30, 41, 28, 32, 30, 22, 31, 40, 45, 31, 39, 12, 30, 
    43, 42, 28, 34, 30, 33, 47, 37, 43, 36, 47, 29, 2, 15, 0, 
    51, 41, 29, 57, 48, 36, 40, 33, 37, 38, 53, 28, 0, 18, 0, 
    42, 35, 36, 49, 49, 48, 48, 48, 48, 31, 42, 25, 13, 0, 6, 
    55, 51, 61, 56, 53, 56, 53, 38, 40, 10, 34, 24, 24, 21, 20, 
    33, 57, 57, 51, 48, 48, 46, 45, 46, 36, 31, 26, 29, 22, 30, 
    64, 53, 54, 46, 61, 58, 33, 24, 57, 49, 37, 27, 31, 28, 31, 
    74, 53, 38, 39, 42, 66, 31, 37, 45, 36, 38, 34, 30, 34, 21, 
    66, 55, 43, 50, 52, 42, 34, 43, 43, 39, 33, 41, 24, 31, 28, 
    42, 40, 40, 44, 43, 42, 41, 37, 39, 30, 31, 31, 29, 32, 32, 
    28, 32, 34, 35, 35, 38, 40, 32, 53, 16, 32, 28, 33, 33, 19, 
    
    -- channel=173
    16, 0, 0, 0, 0, 2, 0, 4, 0, 0, 6, 0, 10, 0, 0, 
    18, 0, 0, 9, 0, 8, 0, 0, 0, 36, 0, 0, 15, 0, 0, 
    19, 4, 0, 9, 0, 5, 5, 0, 0, 73, 0, 0, 16, 0, 0, 
    18, 10, 0, 0, 0, 0, 5, 20, 38, 23, 0, 7, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 12, 16, 9, 0, 0, 0, 12, 7, 
    0, 0, 14, 0, 0, 3, 0, 16, 2, 1, 0, 0, 65, 0, 58, 
    0, 16, 10, 0, 0, 7, 0, 8, 3, 0, 0, 0, 21, 20, 80, 
    0, 0, 0, 0, 0, 0, 0, 15, 0, 36, 0, 0, 5, 70, 0, 
    7, 0, 0, 0, 5, 4, 3, 3, 0, 17, 0, 0, 4, 20, 0, 
    18, 0, 0, 4, 0, 0, 0, 13, 0, 0, 0, 15, 18, 26, 6, 
    0, 0, 4, 14, 0, 0, 29, 32, 0, 0, 11, 19, 19, 12, 11, 
    0, 0, 25, 13, 0, 0, 19, 15, 0, 4, 15, 7, 14, 10, 14, 
    0, 4, 8, 6, 3, 0, 4, 2, 7, 3, 12, 0, 18, 3, 5, 
    5, 2, 1, 0, 0, 0, 0, 7, 0, 26, 3, 7, 7, 0, 4, 
    3, 0, 0, 0, 0, 0, 1, 11, 0, 42, 0, 5, 1, 0, 24, 
    
    -- channel=174
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=175
    37, 0, 0, 13, 15, 19, 20, 38, 10, 22, 34, 19, 29, 25, 16, 
    40, 0, 0, 25, 20, 25, 23, 28, 15, 65, 0, 11, 34, 29, 14, 
    44, 1, 1, 30, 21, 29, 39, 21, 13, 110, 0, 17, 47, 29, 11, 
    52, 4, 17, 27, 36, 22, 45, 39, 53, 56, 0, 0, 0, 38, 21, 
    35, 22, 28, 11, 33, 26, 31, 56, 35, 22, 11, 0, 0, 38, 9, 
    0, 0, 30, 0, 0, 0, 3, 34, 17, 18, 0, 0, 50, 3, 45, 
    0, 14, 21, 0, 0, 12, 0, 7, 0, 0, 0, 11, 68, 18, 85, 
    2, 3, 0, 0, 0, 8, 16, 24, 22, 57, 6, 6, 25, 75, 0, 
    10, 27, 0, 0, 19, 28, 27, 23, 0, 45, 0, 11, 22, 30, 30, 
    15, 0, 0, 14, 10, 4, 14, 33, 27, 19, 15, 35, 45, 53, 23, 
    0, 7, 11, 33, 13, 12, 48, 38, 0, 13, 42, 48, 37, 32, 23, 
    0, 9, 41, 14, 0, 0, 55, 36, 9, 18, 30, 30, 17, 16, 23, 
    0, 25, 44, 24, 18, 15, 14, 12, 21, 23, 18, 5, 31, 9, 10, 
    4, 7, 9, 1, 11, 15, 10, 15, 0, 25, 14, 8, 12, 3, 5, 
    10, 0, 1, 0, 1, 3, 7, 21, 0, 49, 4, 7, 4, 2, 31, 
    
    -- channel=176
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    9, 4, 0, 2, 25, 11, 0, 0, 0, 0, 26, 40, 25, 0, 0, 
    0, 0, 0, 0, 0, 9, 17, 31, 47, 32, 16, 0, 0, 0, 0, 
    11, 29, 37, 27, 6, 0, 0, 0, 0, 0, 0, 0, 0, 15, 82, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 21, 0, 0, 0, 0, 
    12, 24, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=177
    7, 32, 28, 16, 15, 10, 8, 0, 13, 6, 0, 9, 5, 6, 13, 
    0, 24, 19, 4, 5, 1, 0, 0, 8, 0, 7, 10, 0, 0, 9, 
    0, 15, 13, 1, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 7, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 32, 13, 0, 0, 
    30, 27, 0, 23, 37, 25, 18, 0, 5, 12, 54, 55, 0, 12, 0, 
    17, 3, 0, 31, 24, 27, 36, 42, 51, 42, 43, 0, 0, 0, 0, 
    33, 38, 60, 54, 36, 27, 21, 5, 0, 0, 0, 2, 0, 0, 61, 
    5, 0, 18, 21, 2, 0, 0, 7, 23, 10, 38, 8, 0, 0, 0, 
    24, 56, 23, 0, 17, 28, 12, 0, 0, 3, 6, 0, 0, 0, 0, 
    20, 18, 9, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 
    29, 9, 0, 6, 28, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 
    0, 0, 0, 3, 0, 0, 0, 0, 27, 0, 0, 0, 1, 8, 4, 
    0, 8, 9, 11, 13, 11, 2, 0, 16, 0, 3, 3, 5, 9, 0, 
    
    -- channel=178
    52, 36, 49, 54, 56, 55, 56, 59, 52, 58, 58, 55, 57, 58, 56, 
    51, 34, 46, 52, 52, 52, 54, 56, 53, 59, 43, 54, 58, 59, 54, 
    50, 34, 42, 49, 47, 49, 52, 47, 47, 61, 23, 50, 55, 52, 51, 
    49, 32, 43, 47, 48, 46, 51, 41, 38, 40, 14, 16, 33, 47, 42, 
    32, 23, 31, 28, 36, 36, 39, 45, 31, 23, 19, 17, 15, 30, 22, 
    12, 11, 23, 14, 22, 23, 29, 34, 22, 20, 12, 25, 26, 29, 28, 
    18, 16, 24, 13, 28, 32, 32, 30, 22, 23, 17, 35, 51, 29, 25, 
    28, 26, 30, 33, 41, 43, 44, 41, 41, 39, 24, 31, 38, 33, 5, 
    35, 35, 31, 43, 48, 44, 38, 34, 30, 39, 22, 32, 35, 33, 34, 
    31, 24, 35, 38, 36, 33, 35, 37, 32, 35, 36, 39, 33, 29, 16, 
    31, 35, 36, 38, 32, 32, 37, 25, 6, 28, 32, 29, 17, 12, 6, 
    15, 31, 34, 21, 17, 18, 40, 22, 12, 17, 14, 10, 6, 1, 1, 
    16, 27, 31, 18, 12, 14, 14, 9, 10, 9, 4, 0, 7, 0, 0, 
    0, 2, 1, 0, 2, 2, 2, 2, 0, 6, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    
    -- channel=179
    65, 55, 68, 66, 68, 62, 66, 67, 65, 67, 58, 65, 65, 69, 61, 
    60, 49, 60, 61, 63, 57, 59, 59, 61, 60, 22, 59, 62, 64, 60, 
    56, 41, 54, 56, 62, 55, 58, 37, 43, 47, 30, 46, 55, 53, 56, 
    42, 32, 41, 33, 42, 45, 45, 62, 23, 0, 5, 0, 0, 37, 23, 
    0, 0, 0, 0, 0, 0, 4, 17, 24, 37, 25, 31, 46, 35, 7, 
    27, 34, 44, 23, 46, 44, 50, 34, 34, 38, 42, 74, 69, 23, 33, 
    36, 25, 15, 29, 29, 44, 48, 50, 62, 58, 58, 43, 29, 32, 7, 
    47, 54, 64, 79, 68, 67, 66, 63, 46, 38, 10, 23, 35, 28, 43, 
    38, 22, 23, 45, 52, 43, 38, 36, 45, 51, 60, 50, 37, 38, 25, 
    29, 54, 62, 42, 37, 55, 60, 50, 28, 41, 44, 39, 25, 6, 0, 
    41, 49, 47, 37, 31, 29, 40, 4, 17, 33, 21, 8, 13, 9, 12, 
    34, 36, 36, 12, 25, 40, 27, 30, 26, 16, 20, 10, 10, 9, 0, 
    28, 25, 15, 21, 11, 0, 8, 25, 19, 7, 10, 16, 6, 5, 8, 
    0, 0, 2, 10, 16, 12, 8, 7, 17, 30, 5, 7, 4, 9, 11, 
    5, 7, 10, 11, 15, 21, 20, 8, 11, 8, 6, 2, 8, 8, 0, 
    
    -- channel=180
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 15, 0, 0, 0, 
    3, 0, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 
    
    -- channel=181
    0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 5, 3, 0, 0, 0, 
    0, 7, 11, 0, 4, 1, 8, 11, 4, 0, 58, 11, 0, 3, 6, 
    0, 11, 15, 0, 2, 2, 0, 37, 38, 0, 62, 44, 7, 16, 15, 
    7, 14, 22, 32, 15, 14, 4, 0, 40, 68, 51, 99, 122, 40, 52, 
    76, 62, 69, 81, 81, 80, 71, 41, 13, 0, 10, 0, 0, 4, 53, 
    1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 3, 12, 17, 18, 0, 0, 0, 0, 0, 0, 11, 0, 1, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 3, 54, 29, 4, 0, 0, 
    7, 36, 44, 18, 8, 26, 29, 11, 0, 0, 0, 0, 3, 0, 23, 
    0, 0, 0, 9, 16, 0, 0, 6, 38, 12, 1, 3, 26, 38, 44, 
    24, 0, 1, 11, 40, 48, 1, 24, 32, 31, 41, 41, 23, 18, 9, 
    32, 16, 0, 17, 2, 14, 17, 4, 14, 22, 18, 23, 6, 9, 7, 
    31, 34, 38, 26, 39, 47, 23, 5, 19, 30, 9, 10, 6, 6, 0, 
    35, 41, 25, 18, 13, 21, 25, 15, 7, 0, 11, 4, 5, 0, 0, 
    3, 2, 2, 1, 0, 0, 0, 4, 34, 0, 3, 4, 1, 2, 0, 
    
    -- channel=182
    64, 46, 63, 70, 72, 71, 75, 79, 72, 78, 77, 75, 78, 80, 74, 
    64, 46, 62, 71, 71, 69, 70, 70, 71, 80, 34, 72, 78, 78, 71, 
    65, 45, 60, 69, 72, 66, 71, 55, 55, 71, 24, 62, 74, 69, 67, 
    59, 38, 58, 53, 66, 59, 64, 63, 39, 0, 2, 0, 3, 59, 50, 
    5, 5, 5, 9, 14, 18, 18, 33, 20, 27, 16, 15, 41, 38, 10, 
    4, 18, 33, 7, 25, 28, 33, 30, 24, 24, 21, 57, 67, 27, 37, 
    21, 15, 9, 8, 19, 30, 33, 32, 38, 40, 44, 53, 47, 48, 14, 
    30, 33, 38, 54, 54, 56, 57, 58, 47, 51, 16, 29, 42, 31, 16, 
    31, 25, 13, 37, 50, 45, 38, 33, 38, 47, 46, 48, 41, 41, 41, 
    15, 27, 48, 41, 27, 43, 53, 53, 32, 40, 43, 46, 36, 17, 1, 
    21, 37, 38, 37, 31, 24, 43, 7, 0, 33, 29, 14, 10, 3, 7, 
    14, 27, 32, 4, 6, 26, 36, 23, 14, 10, 14, 3, 0, 0, 0, 
    15, 24, 18, 13, 7, 0, 0, 11, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    
    -- channel=183
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=184
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 6, 0, 9, 4, 0, 
    6, 0, 0, 2, 0, 6, 2, 0, 0, 38, 0, 0, 14, 5, 0, 
    13, 0, 0, 10, 4, 10, 17, 0, 0, 64, 0, 0, 18, 4, 0, 
    17, 0, 0, 0, 14, 7, 16, 29, 28, 2, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 26, 5, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 28, 16, 54, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 11, 58, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 6, 5, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 11, 13, 15, 0, 
    0, 0, 0, 0, 0, 0, 17, 7, 0, 0, 2, 5, 9, 3, 10, 
    0, 0, 7, 0, 0, 0, 3, 3, 0, 0, 5, 0, 4, 3, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 1, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 4, 0, 22, 0, 0, 0, 0, 20, 
    
    -- channel=185
    107, 99, 120, 117, 118, 110, 113, 109, 111, 114, 108, 110, 106, 112, 106, 
    103, 92, 114, 106, 111, 101, 107, 109, 107, 103, 94, 109, 103, 111, 105, 
    97, 82, 103, 95, 103, 92, 97, 98, 100, 83, 93, 108, 100, 103, 102, 
    85, 69, 89, 86, 89, 87, 86, 78, 73, 63, 64, 71, 93, 91, 86, 
    62, 52, 59, 65, 63, 68, 70, 76, 61, 62, 59, 46, 57, 61, 50, 
    49, 49, 53, 46, 56, 57, 71, 69, 62, 59, 59, 69, 47, 67, 35, 
    65, 52, 52, 62, 81, 75, 81, 71, 70, 73, 77, 82, 61, 56, 22, 
    68, 63, 67, 82, 93, 98, 101, 96, 96, 80, 70, 67, 65, 26, 29, 
    84, 81, 89, 102, 104, 104, 99, 86, 81, 64, 63, 68, 69, 61, 68, 
    66, 76, 90, 93, 91, 89, 90, 88, 79, 82, 78, 75, 66, 52, 43, 
    89, 90, 91, 83, 90, 92, 80, 54, 59, 81, 71, 59, 45, 35, 31, 
    88, 86, 78, 59, 59, 83, 74, 52, 54, 55, 49, 41, 34, 27, 16, 
    73, 76, 71, 59, 60, 55, 45, 47, 45, 43, 34, 34, 25, 20, 15, 
    37, 35, 33, 35, 36, 36, 37, 35, 32, 33, 26, 22, 18, 19, 19, 
    14, 15, 20, 22, 25, 27, 30, 26, 36, 24, 20, 16, 18, 19, 10, 
    
    -- channel=186
    14, 0, 3, 11, 14, 13, 18, 26, 16, 21, 27, 19, 17, 22, 13, 
    21, 0, 11, 16, 23, 21, 29, 30, 18, 59, 21, 19, 23, 30, 16, 
    25, 0, 11, 17, 25, 22, 37, 43, 27, 76, 0, 34, 36, 36, 20, 
    40, 0, 33, 37, 41, 26, 37, 23, 69, 70, 34, 64, 49, 52, 42, 
    62, 42, 58, 58, 69, 65, 57, 60, 15, 6, 2, 0, 0, 44, 36, 
    0, 0, 4, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 17, 8, 
    0, 1, 15, 0, 3, 0, 0, 0, 0, 0, 0, 22, 32, 28, 39, 
    0, 0, 0, 0, 0, 0, 0, 7, 18, 44, 32, 19, 18, 7, 0, 
    8, 38, 12, 8, 19, 31, 29, 13, 0, 0, 0, 5, 15, 7, 40, 
    0, 0, 0, 21, 7, 0, 0, 25, 25, 16, 12, 26, 43, 51, 32, 
    3, 1, 7, 23, 33, 25, 35, 32, 0, 26, 49, 48, 23, 15, 16, 
    0, 11, 29, 11, 0, 0, 38, 11, 8, 18, 18, 20, 4, 5, 5, 
    5, 30, 40, 19, 29, 31, 8, 0, 16, 22, 0, 0, 13, 0, 0, 
    19, 17, 7, 0, 2, 9, 10, 6, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 11, 0, 0, 0, 0, 11, 
    
    -- channel=187
    38, 39, 38, 41, 37, 35, 29, 25, 26, 29, 29, 24, 27, 24, 26, 
    33, 32, 31, 32, 25, 27, 26, 22, 25, 33, 27, 22, 27, 23, 25, 
    26, 27, 22, 20, 16, 18, 18, 26, 27, 25, 25, 29, 24, 17, 21, 
    21, 21, 19, 14, 10, 11, 11, 14, 33, 25, 23, 37, 22, 16, 17, 
    23, 22, 18, 20, 18, 21, 24, 24, 20, 19, 17, 0, 2, 0, 14, 
    2, 6, 7, 2, 0, 10, 21, 26, 17, 8, 1, 0, 0, 0, 6, 
    16, 17, 14, 16, 24, 23, 23, 17, 11, 10, 9, 13, 0, 11, 10, 
    19, 10, 9, 21, 29, 33, 35, 38, 35, 29, 14, 5, 7, 0, 0, 
    40, 38, 36, 40, 48, 48, 40, 24, 19, 4, 0, 8, 12, 10, 7, 
    25, 21, 31, 40, 33, 27, 26, 33, 28, 17, 17, 20, 22, 17, 9, 
    33, 36, 38, 37, 40, 33, 28, 21, 17, 23, 27, 20, 11, 2, 0, 
    27, 35, 31, 23, 15, 24, 28, 16, 13, 13, 14, 5, 1, 0, 0, 
    26, 35, 31, 24, 22, 18, 10, 9, 12, 8, 1, 1, 0, 0, 0, 
    10, 9, 4, 3, 3, 4, 4, 2, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=188
    50, 49, 52, 57, 56, 56, 53, 51, 51, 55, 55, 50, 52, 51, 50, 
    50, 46, 51, 53, 51, 53, 55, 51, 50, 62, 56, 50, 54, 53, 53, 
    48, 47, 47, 46, 45, 47, 49, 58, 58, 57, 50, 57, 55, 51, 53, 
    50, 47, 53, 51, 47, 46, 43, 40, 62, 58, 47, 72, 60, 54, 56, 
    59, 49, 55, 57, 60, 61, 59, 55, 40, 34, 31, 17, 24, 37, 50, 
    17, 18, 24, 19, 12, 23, 34, 40, 30, 22, 12, 1, 18, 13, 29, 
    29, 31, 36, 29, 40, 32, 32, 22, 14, 18, 23, 43, 30, 48, 40, 
    26, 18, 13, 24, 36, 41, 44, 50, 51, 52, 43, 36, 37, 14, 0, 
    53, 55, 57, 54, 62, 62, 55, 40, 35, 21, 14, 32, 38, 35, 41, 
    36, 25, 38, 55, 47, 36, 39, 51, 47, 39, 40, 45, 48, 48, 39, 
    44, 45, 50, 52, 60, 51, 46, 43, 35, 45, 53, 49, 33, 25, 22, 
    40, 48, 45, 38, 27, 40, 50, 32, 30, 34, 33, 26, 21, 18, 14, 
    43, 54, 53, 42, 42, 42, 31, 26, 32, 30, 20, 20, 20, 14, 8, 
    34, 32, 24, 22, 22, 23, 24, 21, 9, 16, 17, 15, 12, 9, 10, 
    9, 7, 8, 8, 9, 8, 14, 16, 19, 20, 12, 13, 11, 9, 11, 
    
    -- channel=189
    0, 0, 0, 0, 6, 11, 19, 23, 20, 23, 26, 27, 23, 26, 25, 
    0, 0, 9, 13, 20, 20, 24, 27, 24, 19, 12, 28, 26, 30, 25, 
    12, 4, 20, 27, 33, 27, 29, 25, 20, 19, 3, 23, 27, 36, 30, 
    21, 10, 29, 36, 45, 38, 39, 22, 0, 0, 0, 0, 19, 35, 38, 
    1, 0, 3, 8, 15, 15, 7, 5, 0, 0, 0, 1, 17, 24, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 21, 48, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 26, 40, 25, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 25, 24, 16, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 16, 13, 15, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 11, 8, 4, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=190
    0, 28, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 1, 0, 9, 
    0, 43, 0, 0, 0, 0, 0, 0, 7, 0, 19, 0, 0, 0, 0, 
    0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 10, 
    0, 11, 0, 0, 0, 0, 2, 0, 6, 0, 0, 35, 4, 0, 11, 
    0, 22, 0, 17, 0, 4, 0, 0, 0, 0, 41, 0, 0, 0, 7, 
    0, 14, 0, 6, 0, 1, 0, 5, 0, 0, 9, 0, 0, 0, 40, 
    3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 5, 0, 
    9, 2, 0, 0, 1, 0, 0, 0, 11, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 3, 34, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 0, 0, 
    
    -- channel=191
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 58, 45, 42, 1, 0, 0, 
    13, 12, 26, 11, 15, 7, 17, 5, 0, 0, 0, 0, 0, 14, 13, 
    12, 0, 0, 23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 11, 16, 15, 11, 15, 8, 0, 0, 0, 3, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 0, 32, 20, 
    0, 1, 18, 0, 0, 0, 10, 18, 0, 0, 0, 0, 1, 0, 0, 
    31, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 
    0, 0, 0, 0, 0, 6, 1, 35, 14, 0, 0, 14, 0, 5, 0, 
    0, 2, 7, 28, 19, 0, 0, 0, 2, 7, 0, 16, 2, 0, 7, 
    0, 0, 0, 0, 3, 22, 8, 0, 0, 12, 0, 0, 1, 2, 2, 
    9, 12, 5, 0, 0, 0, 11, 7, 4, 0, 5, 0, 3, 0, 0, 
    0, 2, 5, 6, 1, 0, 0, 0, 0, 5, 0, 1, 0, 0, 0, 
    
    -- channel=192
    4, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 
    0, 0, 0, 0, 20, 19, 11, 21, 14, 13, 13, 16, 7, 0, 0, 
    2, 0, 0, 12, 19, 26, 22, 35, 22, 16, 23, 22, 11, 0, 0, 
    0, 0, 0, 30, 17, 19, 15, 24, 19, 13, 23, 17, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 16, 21, 2, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 12, 8, 0, 4, 1, 6, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 14, 13, 3, 0, 0, 0, 6, 7, 0, 
    6, 0, 0, 0, 4, 0, 14, 52, 9, 0, 19, 3, 42, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 3, 7, 23, 
    0, 2, 3, 4, 3, 13, 5, 12, 3, 5, 0, 4, 18, 4, 0, 
    
    -- channel=193
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 11, 25, 22, 23, 15, 22, 17, 13, 0, 0, 0, 
    0, 0, 0, 31, 13, 6, 14, 16, 11, 14, 12, 12, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 48, 27, 12, 25, 18, 25, 28, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 2, 4, 5, 4, 0, 0, 0, 0, 
    
    -- channel=194
    25, 3, 0, 0, 9, 3, 1, 7, 2, 5, 3, 2, 8, 0, 0, 
    22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 16, 0, 0, 
    2, 7, 0, 0, 1, 3, 5, 2, 0, 0, 6, 17, 0, 0, 0, 
    3, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 22, 27, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 42, 21, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 26, 40, 35, 8, 0, 2, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 27, 29, 18, 25, 31, 51, 19, 7, 0, 0, 
    17, 0, 0, 0, 0, 0, 41, 63, 0, 0, 19, 19, 60, 10, 6, 
    5, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    7, 1, 0, 0, 0, 0, 0, 4, 0, 0, 0, 4, 3, 0, 6, 
    15, 27, 23, 27, 23, 27, 27, 27, 23, 22, 27, 24, 24, 33, 54, 
    7, 22, 23, 25, 23, 30, 20, 28, 22, 23, 18, 20, 45, 36, 7, 
    
    -- channel=195
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 30, 26, 24, 26, 27, 25, 18, 0, 0, 0, 
    0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 4, 0, 0, 4, 3, 0, 0, 0, 0, 0, 
    0, 4, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 67, 12, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 58, 46, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 79, 77, 40, 8, 0, 0, 0, 0, 
    0, 0, 0, 12, 31, 17, 11, 0, 4, 38, 82, 100, 78, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 79, 86, 91, 94, 85, 60, 52, 62, 48, 43, 38, 32, 44, 44, 
    2, 0, 0, 2, 4, 7, 8, 19, 30, 36, 40, 43, 48, 48, 48, 
    22, 22, 22, 17, 15, 13, 10, 8, 7, 4, 3, 3, 2, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=196
    43, 41, 16, 17, 30, 29, 25, 28, 27, 27, 27, 26, 39, 47, 45, 
    37, 33, 27, 0, 11, 5, 0, 9, 7, 12, 10, 21, 44, 38, 41, 
    32, 29, 20, 21, 42, 58, 43, 60, 64, 60, 61, 59, 49, 40, 42, 
    30, 29, 12, 30, 29, 28, 32, 36, 24, 14, 26, 30, 40, 32, 35, 
    30, 29, 30, 21, 21, 17, 18, 23, 22, 18, 24, 43, 45, 35, 35, 
    37, 23, 13, 40, 41, 43, 47, 46, 43, 42, 44, 41, 34, 35, 37, 
    43, 13, 0, 0, 15, 37, 36, 36, 36, 33, 35, 34, 34, 32, 34, 
    48, 37, 41, 27, 0, 3, 37, 39, 32, 31, 35, 34, 35, 34, 35, 
    48, 42, 39, 37, 0, 0, 0, 0, 12, 27, 38, 35, 32, 31, 33, 
    49, 40, 40, 21, 0, 0, 0, 0, 0, 0, 0, 0, 18, 35, 37, 
    48, 39, 39, 19, 35, 8, 2, 51, 50, 11, 34, 6, 54, 41, 31, 
    16, 3, 0, 0, 0, 0, 14, 21, 0, 7, 13, 17, 14, 1, 6, 
    3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    
    -- channel=197
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 29, 18, 25, 37, 36, 33, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    2, 0, 0, 2, 28, 28, 27, 24, 26, 25, 23, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 68, 92, 38, 60, 93, 60, 86, 50, 47, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 9, 8, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 2, 8, 7, 6, 8, 6, 1, 10, 33, 0, 
    
    -- channel=198
    12, 13, 11, 12, 8, 11, 12, 9, 14, 12, 13, 10, 11, 26, 23, 
    14, 12, 6, 13, 8, 0, 0, 2, 3, 3, 5, 3, 15, 13, 19, 
    10, 13, 5, 2, 9, 18, 14, 13, 17, 24, 17, 26, 21, 19, 19, 
    15, 10, 5, 3, 6, 4, 7, 9, 6, 0, 3, 7, 13, 13, 15, 
    18, 13, 7, 14, 3, 3, 0, 4, 6, 0, 6, 2, 23, 17, 17, 
    18, 21, 6, 0, 27, 25, 27, 25, 25, 26, 25, 32, 13, 15, 18, 
    18, 8, 17, 0, 0, 0, 15, 17, 18, 20, 17, 16, 16, 14, 12, 
    20, 18, 9, 43, 37, 0, 0, 10, 15, 12, 15, 16, 17, 16, 16, 
    22, 21, 22, 11, 15, 0, 0, 0, 0, 0, 3, 16, 17, 15, 14, 
    21, 21, 18, 22, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 13, 
    16, 17, 19, 5, 7, 60, 17, 13, 55, 25, 43, 32, 31, 37, 17, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 1, 0, 0, 
    5, 0, 1, 4, 8, 2, 5, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 20, 21, 
    
    -- channel=199
    20, 26, 15, 15, 10, 16, 14, 9, 10, 8, 13, 13, 11, 29, 29, 
    18, 22, 25, 15, 22, 27, 28, 23, 30, 33, 30, 15, 28, 27, 27, 
    18, 21, 32, 15, 32, 26, 26, 20, 26, 35, 32, 28, 32, 31, 28, 
    17, 19, 27, 0, 6, 4, 7, 4, 0, 6, 5, 15, 0, 27, 23, 
    21, 18, 21, 33, 19, 17, 11, 14, 24, 21, 19, 14, 27, 26, 23, 
    28, 37, 38, 22, 22, 21, 22, 25, 25, 27, 25, 25, 23, 21, 18, 
    28, 3, 0, 17, 35, 28, 19, 22, 23, 27, 26, 29, 29, 29, 25, 
    29, 25, 31, 23, 8, 27, 39, 29, 25, 26, 25, 25, 25, 24, 22, 
    33, 30, 31, 33, 30, 10, 9, 32, 53, 48, 23, 22, 24, 25, 22, 
    34, 31, 30, 53, 35, 5, 9, 10, 6, 3, 9, 53, 57, 41, 25, 
    30, 28, 28, 24, 0, 0, 0, 0, 4, 0, 0, 0, 0, 6, 15, 
    63, 69, 70, 69, 67, 68, 66, 53, 44, 41, 46, 42, 39, 28, 33, 
    13, 14, 19, 25, 28, 26, 26, 26, 29, 28, 29, 27, 28, 29, 21, 
    0, 0, 2, 0, 5, 0, 1, 2, 7, 6, 4, 8, 6, 0, 0, 
    0, 4, 5, 5, 4, 0, 0, 0, 0, 0, 6, 9, 0, 16, 44, 
    
    -- channel=200
    0, 21, 39, 25, 14, 26, 28, 22, 27, 25, 26, 26, 22, 28, 27, 
    0, 13, 38, 60, 21, 30, 34, 27, 36, 31, 30, 17, 25, 30, 27, 
    0, 12, 40, 40, 46, 26, 38, 24, 32, 36, 30, 22, 14, 28, 28, 
    4, 13, 57, 35, 27, 28, 34, 26, 28, 43, 29, 36, 1, 26, 24, 
    18, 14, 27, 36, 14, 12, 15, 19, 16, 23, 14, 11, 25, 29, 24, 
    20, 20, 12, 27, 31, 29, 29, 34, 33, 30, 29, 23, 27, 29, 25, 
    18, 49, 39, 0, 0, 19, 29, 32, 33, 34, 28, 29, 27, 28, 24, 
    14, 32, 48, 72, 0, 0, 0, 29, 33, 32, 28, 29, 29, 30, 23, 
    17, 30, 35, 45, 74, 0, 0, 0, 0, 11, 20, 34, 30, 27, 24, 
    18, 30, 33, 42, 70, 0, 0, 0, 0, 0, 0, 0, 0, 11, 25, 
    12, 33, 31, 62, 55, 61, 8, 0, 41, 37, 22, 22, 0, 19, 16, 
    0, 0, 0, 0, 0, 3, 0, 0, 3, 4, 2, 7, 6, 6, 3, 
    0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=201
    15, 17, 0, 2, 7, 5, 0, 0, 0, 0, 0, 0, 2, 7, 9, 
    19, 23, 17, 0, 12, 16, 11, 16, 14, 17, 15, 10, 20, 13, 12, 
    20, 22, 23, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 17, 15, 
    15, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 
    12, 19, 17, 7, 13, 12, 10, 10, 15, 10, 8, 15, 10, 15, 16, 
    13, 20, 27, 24, 3, 6, 7, 7, 6, 6, 7, 11, 16, 12, 12, 
    14, 0, 0, 17, 61, 33, 15, 14, 13, 13, 16, 17, 17, 18, 19, 
    18, 13, 2, 0, 0, 48, 53, 22, 12, 14, 13, 13, 14, 13, 15, 
    18, 14, 12, 2, 0, 1, 11, 49, 62, 42, 23, 11, 13, 15, 16, 
    16, 12, 13, 22, 0, 0, 3, 0, 0, 5, 44, 70, 64, 38, 19, 
    17, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    49, 56, 57, 60, 61, 53, 47, 47, 41, 46, 37, 39, 31, 37, 41, 
    0, 7, 5, 7, 9, 10, 12, 19, 25, 29, 30, 34, 37, 36, 32, 
    0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=202
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=203
    67, 78, 71, 62, 68, 71, 70, 71, 74, 73, 73, 70, 83, 86, 85, 
    65, 72, 80, 46, 47, 42, 36, 47, 45, 46, 45, 56, 86, 80, 82, 
    62, 71, 68, 65, 71, 80, 66, 82, 85, 83, 86, 84, 72, 81, 84, 
    67, 73, 62, 76, 66, 68, 71, 66, 67, 58, 62, 66, 75, 75, 78, 
    76, 73, 80, 60, 52, 47, 56, 61, 54, 53, 53, 76, 83, 80, 80, 
    79, 61, 37, 90, 96, 97, 98, 98, 96, 92, 92, 85, 79, 82, 86, 
    80, 84, 50, 0, 10, 73, 86, 87, 88, 83, 81, 79, 76, 74, 75, 
    81, 88, 103, 114, 1, 0, 39, 81, 79, 77, 79, 80, 82, 80, 80, 
    81, 86, 86, 87, 32, 0, 0, 0, 0, 43, 75, 85, 79, 76, 79, 
    79, 81, 84, 60, 0, 0, 0, 9, 0, 0, 0, 0, 6, 55, 81, 
    76, 82, 82, 78, 137, 106, 66, 110, 123, 95, 110, 79, 97, 88, 72, 
    0, 0, 0, 0, 0, 0, 5, 10, 0, 23, 18, 34, 23, 16, 19, 
    25, 34, 31, 24, 20, 20, 19, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 
    0, 0, 0, 0, 0, 11, 8, 10, 8, 9, 0, 0, 13, 36, 0, 
    
    -- channel=204
    16, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    18, 0, 0, 0, 15, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 
    16, 0, 0, 0, 0, 5, 0, 11, 0, 0, 0, 10, 3, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 48, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 11, 31, 28, 2, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 3, 9, 2, 5, 0, 38, 10, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 13, 64, 0, 0, 3, 0, 68, 13, 6, 
    1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 2, 0, 5, 0, 6, 0, 0, 0, 0, 9, 28, 0, 
    
    -- channel=205
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 35, 27, 21, 29, 26, 24, 23, 20, 4, 0, 0, 
    0, 0, 0, 24, 27, 34, 33, 41, 31, 27, 25, 23, 8, 0, 0, 
    0, 0, 0, 43, 30, 23, 26, 35, 29, 31, 37, 33, 23, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 4, 0, 1, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 7, 8, 3, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 2, 0, 11, 24, 5, 0, 11, 0, 21, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 1, 3, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=206
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 9, 10, 8, 9, 11, 9, 7, 0, 0, 0, 
    0, 0, 0, 7, 11, 15, 12, 19, 13, 9, 10, 10, 1, 0, 0, 
    0, 0, 0, 11, 7, 0, 10, 8, 5, 7, 12, 6, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 15, 25, 19, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 10, 6, 9, 15, 25, 27, 18, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 9, 13, 15, 17, 9, 1, 3, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 11, 8, 10, 11, 10, 8, 8, 8, 7, 7, 5, 6, 7, 0, 
    6, 4, 4, 6, 7, 2, 0, 4, 1, 0, 1, 7, 5, 0, 0, 
    
    -- channel=207
    42, 53, 41, 28, 33, 35, 31, 30, 28, 29, 30, 31, 31, 33, 35, 
    47, 56, 52, 5, 0, 6, 4, 2, 5, 8, 9, 14, 36, 40, 39, 
    45, 55, 50, 3, 7, 0, 0, 0, 8, 9, 6, 6, 36, 41, 41, 
    44, 56, 40, 0, 4, 6, 0, 1, 0, 0, 0, 8, 6, 43, 44, 
    44, 52, 52, 44, 39, 38, 39, 35, 41, 39, 33, 40, 41, 46, 47, 
    44, 49, 54, 54, 44, 44, 43, 44, 44, 44, 42, 41, 46, 43, 44, 
    41, 43, 15, 19, 52, 52, 45, 45, 44, 44, 44, 46, 46, 46, 46, 
    41, 46, 44, 19, 2, 29, 49, 44, 42, 43, 41, 44, 45, 46, 48, 
    37, 40, 39, 40, 19, 2, 3, 25, 44, 47, 47, 43, 44, 45, 48, 
    34, 36, 39, 35, 33, 5, 5, 2, 0, 10, 22, 38, 48, 49, 46, 
    38, 38, 39, 42, 14, 0, 0, 0, 8, 1, 0, 0, 4, 21, 32, 
    47, 50, 50, 50, 50, 58, 50, 48, 58, 57, 56, 59, 57, 60, 58, 
    22, 27, 27, 25, 21, 24, 26, 28, 32, 30, 32, 31, 33, 33, 28, 
    4, 6, 7, 3, 0, 3, 2, 0, 1, 0, 0, 0, 0, 1, 2, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 22, 
    
    -- channel=208
    0, 0, 2, 0, 1, 2, 6, 3, 4, 7, 4, 6, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 6, 0, 0, 0, 1, 8, 16, 9, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 5, 1, 0, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 31, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 1, 25, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 11, 0, 0, 17, 55, 45, 8, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 18, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 16, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    27, 29, 26, 22, 21, 20, 14, 11, 8, 6, 4, 1, 3, 5, 0, 
    3, 3, 3, 1, 3, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    
    -- channel=209
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 21, 29, 26, 24, 24, 18, 17, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 20, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 1, 0, 4, 21, 31, 20, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 6, 9, 
    5, 12, 8, 6, 5, 4, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=211
    21, 46, 56, 41, 29, 45, 47, 39, 43, 42, 45, 42, 38, 46, 43, 
    22, 39, 59, 50, 9, 9, 13, 7, 16, 14, 14, 3, 35, 43, 40, 
    23, 38, 57, 26, 46, 27, 32, 18, 37, 44, 35, 25, 22, 44, 42, 
    29, 40, 73, 23, 21, 24, 35, 25, 20, 37, 21, 41, 0, 41, 39, 
    43, 40, 49, 57, 33, 32, 32, 35, 33, 39, 32, 27, 43, 46, 41, 
    46, 44, 27, 48, 55, 53, 50, 53, 54, 53, 51, 42, 46, 46, 43, 
    41, 70, 60, 0, 0, 32, 45, 48, 49, 50, 43, 45, 44, 43, 39, 
    38, 53, 70, 101, 12, 0, 1, 41, 47, 46, 43, 45, 47, 47, 42, 
    40, 48, 50, 61, 85, 2, 0, 0, 0, 19, 31, 48, 46, 44, 41, 
    40, 45, 46, 54, 73, 0, 0, 4, 0, 0, 0, 0, 0, 21, 38, 
    32, 46, 45, 82, 76, 91, 41, 18, 75, 54, 61, 49, 18, 37, 32, 
    0, 6, 1, 0, 0, 12, 6, 0, 11, 18, 15, 22, 19, 16, 14, 
    11, 21, 23, 20, 16, 15, 11, 1, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 1, 1, 
    0, 3, 5, 2, 4, 6, 12, 7, 13, 11, 8, 4, 0, 14, 19, 
    
    -- channel=212
    12, 0, 0, 4, 7, 0, 0, 4, 3, 4, 1, 2, 10, 5, 3, 
    11, 0, 0, 0, 20, 15, 8, 19, 12, 11, 8, 21, 1, 1, 3, 
    10, 0, 0, 4, 0, 5, 5, 10, 0, 0, 1, 14, 7, 0, 2, 
    7, 0, 0, 5, 6, 5, 0, 10, 8, 0, 6, 0, 29, 0, 2, 
    0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 1, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 3, 
    1, 0, 0, 31, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 23, 37, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 1, 0, 0, 0, 14, 37, 29, 9, 0, 2, 0, 0, 0, 0, 
    6, 3, 0, 0, 0, 12, 13, 10, 17, 15, 37, 13, 6, 1, 0, 
    9, 0, 1, 0, 0, 0, 13, 41, 0, 2, 3, 10, 42, 19, 9, 
    10, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 1, 0, 2, 9, 0, 0, 0, 3, 1, 0, 1, 
    12, 9, 4, 10, 7, 9, 9, 11, 5, 7, 10, 9, 9, 9, 21, 
    8, 8, 6, 11, 8, 12, 9, 15, 9, 11, 11, 10, 14, 20, 4, 
    
    -- channel=213
    8, 2, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    5, 0, 0, 23, 31, 31, 26, 29, 28, 27, 24, 22, 7, 0, 0, 
    3, 0, 0, 25, 34, 36, 39, 41, 33, 32, 30, 28, 18, 0, 0, 
    3, 0, 4, 34, 29, 27, 23, 35, 28, 27, 30, 27, 19, 0, 0, 
    1, 0, 0, 4, 3, 2, 0, 4, 3, 1, 5, 2, 6, 0, 0, 
    0, 0, 0, 0, 0, 1, 5, 5, 4, 2, 2, 4, 0, 0, 0, 
    0, 0, 0, 4, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 15, 9, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 17, 3, 6, 8, 5, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 16, 16, 18, 17, 6, 4, 0, 6, 6, 2, 
    4, 0, 0, 0, 0, 11, 13, 12, 12, 3, 12, 7, 13, 12, 0, 
    12, 5, 2, 3, 4, 0, 15, 22, 5, 1, 12, 7, 16, 7, 3, 
    14, 15, 15, 16, 16, 17, 22, 25, 15, 16, 17, 16, 16, 17, 15, 
    6, 9, 6, 6, 5, 8, 9, 9, 6, 9, 9, 11, 12, 9, 0, 
    10, 14, 13, 12, 10, 13, 12, 11, 10, 9, 10, 9, 8, 0, 0, 
    
    -- channel=214
    0, 0, 5, 6, 6, 10, 15, 14, 16, 18, 15, 12, 9, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 24, 16, 15, 14, 22, 24, 25, 26, 22, 19, 0, 0, 
    2, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 26, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 52, 58, 81, 62, 34, 53, 57, 72, 46, 20, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 9, 8, 8, 6, 8, 7, 7, 4, 4, 5, 0, 1, 9, 29, 
    2, 4, 3, 3, 4, 18, 14, 14, 16, 16, 3, 2, 15, 9, 0, 
    
    -- channel=215
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=216
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 22, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 47, 79, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    17, 17, 13, 10, 7, 10, 6, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=217
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 7, 3, 13, 0, 9, 6, 6, 0, 0, 0, 0, 
    0, 0, 0, 16, 11, 6, 15, 0, 4, 12, 4, 0, 0, 0, 0, 
    0, 0, 7, 4, 3, 0, 9, 1, 4, 12, 0, 3, 0, 0, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 99, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 90, 14, 0, 0, 10, 28, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 39, 0, 0, 0, 7, 0, 1, 0, 0, 0, 
    5, 20, 20, 18, 17, 18, 9, 0, 13, 1, 6, 0, 10, 6, 2, 
    3, 0, 7, 6, 6, 4, 6, 7, 16, 11, 13, 10, 10, 16, 14, 
    20, 8, 9, 2, 10, 6, 5, 3, 5, 8, 2, 4, 3, 0, 0, 
    16, 5, 4, 3, 3, 0, 4, 0, 1, 0, 9, 4, 0, 0, 33, 
    
    -- channel=218
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=219
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    17, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 5, 0, 8, 0, 0, 0, 0, 7, 0, 0, 
    10, 0, 0, 0, 0, 1, 0, 2, 0, 0, 7, 2, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    5, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 25, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 6, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 23, 77, 11, 0, 24, 3, 73, 11, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 29, 
    0, 0, 0, 0, 0, 8, 1, 7, 0, 2, 0, 0, 16, 24, 0, 
    
    -- channel=220
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 1, 2, 0, 2, 3, 6, 0, 6, 2, 0, 
    0, 0, 1, 1, 23, 6, 7, 3, 14, 11, 10, 0, 9, 3, 1, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 2, 0, 11, 0, 2, 0, 
    3, 0, 3, 3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    14, 0, 0, 33, 0, 2, 0, 4, 6, 4, 2, 0, 1, 0, 0, 
    10, 13, 0, 0, 19, 23, 0, 0, 2, 1, 0, 3, 0, 0, 0, 
    8, 6, 31, 39, 0, 0, 29, 15, 0, 3, 0, 2, 1, 0, 0, 
    9, 7, 4, 21, 7, 0, 0, 0, 24, 28, 12, 0, 0, 0, 0, 
    12, 2, 3, 0, 39, 0, 0, 3, 0, 0, 0, 5, 33, 28, 6, 
    7, 2, 1, 39, 23, 0, 0, 0, 11, 0, 1, 0, 0, 0, 0, 
    5, 10, 11, 11, 9, 39, 21, 1, 0, 12, 0, 13, 0, 0, 0, 
    0, 2, 0, 6, 5, 9, 4, 0, 6, 4, 6, 1, 5, 10, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    
    -- channel=221
    0, 0, 26, 10, 0, 6, 12, 3, 8, 5, 7, 7, 0, 1, 0, 
    0, 0, 12, 60, 0, 0, 8, 0, 8, 0, 3, 0, 0, 0, 0, 
    0, 0, 12, 34, 33, 15, 36, 10, 25, 30, 18, 11, 0, 0, 0, 
    0, 0, 36, 32, 12, 12, 28, 16, 11, 31, 8, 19, 0, 0, 0, 
    0, 0, 2, 28, 1, 2, 0, 1, 1, 9, 0, 0, 6, 0, 0, 
    0, 4, 0, 0, 10, 8, 5, 10, 13, 8, 5, 0, 0, 2, 0, 
    0, 35, 47, 0, 0, 0, 0, 3, 5, 8, 0, 2, 0, 0, 0, 
    0, 3, 23, 82, 30, 0, 0, 0, 6, 7, 1, 3, 2, 3, 0, 
    0, 0, 5, 19, 122, 0, 0, 0, 0, 0, 0, 5, 4, 1, 0, 
    0, 1, 2, 22, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 1, 47, 47, 93, 22, 0, 42, 50, 29, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 9, 7, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 3, 0, 0, 0, 1, 4, 0, 1, 0, 0, 0, 
    14, 4, 4, 1, 5, 0, 10, 1, 11, 8, 9, 3, 0, 0, 12, 
    
    -- channel=222
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=223
    30, 53, 62, 42, 40, 50, 49, 46, 47, 47, 47, 47, 42, 41, 44, 
    36, 49, 58, 53, 25, 23, 30, 21, 26, 25, 27, 26, 41, 49, 48, 
    36, 49, 53, 36, 41, 29, 31, 25, 35, 36, 32, 24, 35, 49, 48, 
    40, 50, 62, 48, 44, 48, 46, 45, 49, 54, 45, 50, 34, 50, 49, 
    47, 49, 55, 60, 48, 46, 47, 45, 48, 51, 44, 38, 52, 49, 52, 
    45, 48, 45, 50, 53, 51, 50, 53, 55, 51, 48, 46, 52, 52, 50, 
    40, 69, 59, 24, 22, 43, 52, 54, 54, 53, 49, 51, 50, 50, 50, 
    37, 52, 58, 64, 31, 6, 24, 47, 53, 53, 50, 51, 51, 53, 52, 
    34, 45, 48, 56, 79, 14, 6, 9, 19, 35, 44, 53, 53, 51, 51, 
    33, 43, 47, 48, 84, 16, 11, 14, 16, 24, 10, 14, 18, 34, 48, 
    32, 49, 48, 72, 61, 63, 38, 17, 44, 52, 37, 43, 13, 37, 44, 
    17, 33, 30, 28, 28, 41, 25, 23, 46, 44, 41, 45, 45, 52, 49, 
    25, 36, 35, 30, 24, 26, 25, 24, 33, 28, 29, 27, 28, 32, 29, 
    21, 22, 23, 18, 17, 17, 17, 15, 16, 15, 12, 12, 13, 15, 10, 
    17, 16, 17, 12, 14, 14, 17, 11, 16, 14, 12, 9, 13, 6, 15, 
    
    -- channel=224
    34, 5, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 8, 1, 0, 
    29, 14, 0, 0, 13, 17, 0, 19, 6, 10, 7, 30, 12, 0, 0, 
    29, 7, 0, 0, 0, 4, 0, 18, 3, 0, 0, 9, 26, 0, 1, 
    16, 9, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 26, 0, 2, 
    0, 8, 0, 0, 0, 1, 1, 4, 0, 0, 2, 32, 0, 0, 0, 
    2, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 
    11, 0, 0, 21, 70, 25, 2, 0, 0, 0, 0, 0, 0, 0, 2, 
    21, 0, 0, 0, 0, 79, 67, 7, 0, 0, 0, 0, 0, 0, 0, 
    21, 1, 0, 0, 0, 16, 42, 59, 53, 22, 22, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 10, 20, 10, 8, 4, 66, 54, 54, 30, 6, 
    28, 0, 0, 0, 0, 0, 0, 57, 0, 0, 0, 0, 61, 9, 7, 
    38, 10, 9, 13, 19, 0, 13, 39, 3, 0, 10, 3, 7, 8, 9, 
    2, 0, 0, 0, 0, 0, 3, 16, 0, 10, 9, 17, 17, 9, 14, 
    0, 8, 1, 7, 0, 2, 4, 7, 0, 0, 3, 1, 1, 7, 26, 
    0, 0, 0, 2, 0, 7, 0, 5, 0, 0, 0, 0, 21, 9, 0, 
    
    -- channel=225
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=226
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=227
    9, 25, 38, 23, 14, 23, 24, 19, 21, 21, 22, 21, 14, 17, 22, 
    19, 30, 37, 27, 8, 13, 19, 9, 14, 14, 14, 5, 19, 26, 25, 
    20, 34, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 26, 
    22, 32, 38, 0, 0, 0, 0, 0, 0, 6, 0, 3, 0, 31, 29, 
    30, 32, 31, 32, 20, 22, 23, 19, 23, 24, 18, 8, 20, 31, 31, 
    29, 37, 37, 26, 26, 23, 21, 23, 25, 26, 23, 26, 31, 30, 29, 
    24, 45, 46, 23, 13, 26, 29, 31, 32, 33, 30, 31, 32, 32, 29, 
    21, 33, 30, 36, 22, 3, 11, 28, 31, 31, 28, 30, 30, 31, 30, 
    21, 29, 31, 31, 63, 3, 7, 12, 17, 24, 22, 30, 32, 32, 31, 
    18, 26, 28, 40, 71, 1, 0, 0, 7, 23, 11, 19, 17, 22, 27, 
    15, 27, 29, 43, 10, 28, 0, 0, 7, 12, 0, 8, 0, 12, 22, 
    18, 31, 32, 31, 29, 33, 18, 14, 30, 25, 24, 22, 26, 29, 27, 
    10, 13, 15, 14, 13, 13, 12, 14, 27, 23, 25, 25, 27, 31, 26, 
    15, 14, 16, 10, 11, 9, 8, 8, 8, 7, 4, 3, 3, 0, 0, 
    5, 3, 2, 0, 3, 0, 3, 0, 4, 3, 3, 3, 0, 3, 37, 
    
    -- channel=228
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 20, 14, 17, 16, 18, 11, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 57, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 39, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 58, 63, 33, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 45, 10, 7, 0, 3, 37, 69, 80, 63, 27, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 60, 68, 72, 76, 68, 42, 41, 52, 42, 33, 30, 27, 40, 40, 
    0, 0, 0, 0, 0, 3, 4, 15, 30, 35, 40, 43, 48, 50, 51, 
    19, 25, 24, 18, 13, 12, 10, 8, 4, 3, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    
    -- channel=229
    40, 43, 30, 31, 38, 38, 36, 35, 34, 35, 37, 36, 39, 47, 48, 
    38, 41, 40, 40, 60, 57, 55, 58, 58, 59, 57, 54, 56, 51, 51, 
    36, 39, 41, 53, 54, 62, 56, 64, 61, 60, 60, 62, 57, 51, 53, 
    35, 38, 37, 65, 57, 54, 54, 61, 60, 58, 60, 56, 59, 49, 50, 
    37, 38, 37, 40, 38, 36, 34, 39, 42, 37, 38, 44, 52, 44, 48, 
    40, 42, 40, 40, 35, 37, 41, 44, 42, 38, 38, 45, 45, 45, 45, 
    44, 26, 7, 30, 55, 50, 48, 49, 47, 46, 47, 48, 47, 48, 51, 
    48, 46, 36, 11, 6, 41, 58, 53, 50, 49, 47, 46, 46, 45, 46, 
    48, 50, 49, 44, 5, 2, 16, 43, 58, 56, 50, 47, 46, 45, 47, 
    50, 52, 52, 54, 7, 0, 1, 4, 3, 9, 31, 52, 59, 53, 50, 
    52, 51, 51, 34, 9, 0, 0, 2, 7, 0, 0, 0, 14, 32, 45, 
    57, 59, 58, 58, 58, 49, 44, 51, 51, 47, 46, 47, 46, 49, 50, 
    16, 17, 14, 12, 10, 10, 12, 19, 20, 19, 20, 21, 23, 23, 21, 
    1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=230
    24, 34, 24, 15, 14, 15, 12, 10, 9, 8, 11, 12, 11, 21, 23, 
    31, 38, 31, 0, 0, 7, 6, 3, 9, 12, 12, 4, 25, 24, 24, 
    28, 37, 39, 4, 2, 0, 0, 0, 6, 11, 11, 15, 26, 26, 25, 
    28, 36, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 28, 
    28, 33, 33, 34, 26, 26, 23, 21, 30, 24, 19, 20, 29, 31, 31, 
    27, 44, 49, 31, 27, 26, 26, 27, 28, 29, 26, 28, 29, 25, 26, 
    23, 15, 0, 23, 44, 34, 26, 27, 27, 29, 29, 32, 32, 31, 30, 
    24, 28, 23, 1, 8, 32, 39, 27, 26, 27, 25, 28, 28, 28, 30, 
    23, 25, 25, 22, 23, 0, 4, 32, 48, 43, 29, 26, 28, 29, 30, 
    19, 22, 24, 37, 32, 2, 0, 0, 0, 7, 25, 50, 52, 39, 30, 
    20, 23, 24, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    56, 63, 64, 64, 64, 66, 61, 52, 56, 55, 54, 54, 52, 50, 51, 
    14, 17, 22, 23, 22, 23, 25, 30, 34, 34, 36, 35, 37, 37, 30, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 30, 
    
    -- channel=231
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=232
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 4, 2, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 25, 27, 7, 3, 19, 30, 18, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 1, 3, 7, 8, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 2, 7, 6, 5, 7, 11, 14, 13, 13, 13, 16, 20, 
    18, 13, 11, 11, 15, 13, 14, 15, 17, 16, 17, 18, 24, 14, 18, 
    
    -- channel=233
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 24, 14, 16, 26, 32, 25, 18, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 24, 24, 22, 20, 22, 21, 19, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 75, 99, 46, 64, 95, 66, 89, 57, 51, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 4, 9, 7, 8, 10, 5, 0, 5, 40, 0, 
    
    -- channel=234
    32, 24, 20, 29, 30, 29, 30, 30, 32, 31, 32, 30, 34, 43, 43, 
    27, 23, 21, 38, 50, 46, 45, 49, 48, 48, 47, 44, 40, 36, 38, 
    27, 21, 20, 42, 51, 59, 54, 60, 54, 56, 57, 58, 48, 38, 38, 
    28, 19, 23, 50, 43, 44, 45, 47, 45, 41, 46, 45, 48, 32, 32, 
    30, 23, 19, 24, 22, 21, 18, 25, 24, 20, 27, 28, 36, 31, 30, 
    35, 29, 19, 19, 33, 32, 35, 34, 33, 34, 35, 39, 29, 30, 32, 
    38, 17, 19, 19, 12, 25, 30, 32, 32, 33, 33, 32, 31, 31, 30, 
    40, 34, 29, 39, 34, 22, 27, 34, 33, 30, 33, 31, 31, 30, 29, 
    46, 41, 40, 34, 12, 25, 27, 16, 21, 29, 27, 31, 31, 30, 28, 
    49, 42, 39, 41, 0, 11, 17, 25, 26, 5, 1, 11, 22, 29, 31, 
    43, 37, 39, 23, 26, 39, 23, 40, 52, 28, 41, 30, 48, 45, 36, 
    30, 21, 18, 16, 15, 2, 21, 26, 3, 4, 12, 8, 13, 0, 3, 
    24, 16, 18, 20, 25, 21, 21, 20, 11, 11, 9, 9, 8, 7, 8, 
    11, 7, 6, 11, 13, 10, 11, 15, 15, 16, 16, 17, 17, 16, 23, 
    19, 16, 16, 19, 17, 19, 22, 24, 22, 22, 23, 23, 21, 33, 21, 
    
    -- channel=235
    0, 0, 34, 10, 0, 5, 13, 3, 12, 7, 8, 8, 0, 0, 0, 
    0, 0, 9, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 12, 10, 0, 12, 0, 1, 10, 0, 0, 0, 0, 0, 
    0, 0, 27, 11, 0, 0, 13, 0, 0, 15, 0, 3, 0, 0, 0, 
    0, 0, 4, 28, 0, 0, 0, 0, 0, 7, 0, 0, 3, 0, 0, 
    0, 8, 0, 0, 14, 10, 4, 8, 13, 10, 5, 1, 0, 2, 0, 
    0, 42, 68, 0, 0, 0, 0, 2, 4, 9, 0, 1, 0, 0, 0, 
    0, 3, 20, 89, 54, 0, 0, 0, 5, 4, 0, 3, 1, 4, 0, 
    0, 0, 4, 14, 143, 0, 0, 0, 0, 0, 0, 4, 4, 1, 0, 
    0, 0, 0, 25, 121, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 50, 119, 37, 0, 48, 71, 38, 59, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 8, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 6, 2, 0, 0, 4, 9, 2, 5, 3, 0, 0, 
    21, 8, 6, 4, 8, 3, 15, 5, 17, 15, 15, 8, 0, 0, 25, 
    
    -- channel=236
    40, 37, 20, 24, 26, 25, 19, 21, 20, 21, 21, 20, 24, 26, 27, 
    50, 47, 29, 0, 6, 3, 0, 5, 0, 4, 5, 8, 29, 25, 27, 
    49, 47, 35, 0, 0, 0, 0, 0, 0, 0, 0, 7, 27, 30, 29, 
    45, 45, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 31, 33, 
    37, 44, 34, 18, 29, 30, 30, 27, 28, 22, 27, 33, 27, 34, 35, 
    34, 39, 41, 33, 28, 28, 29, 24, 23, 28, 28, 37, 33, 30, 34, 
    35, 11, 13, 44, 55, 41, 31, 29, 28, 27, 31, 30, 33, 33, 34, 
    40, 31, 9, 0, 19, 64, 52, 30, 25, 25, 29, 29, 31, 30, 35, 
    40, 30, 27, 10, 0, 29, 47, 54, 49, 37, 34, 27, 29, 32, 34, 
    35, 26, 26, 25, 0, 20, 24, 17, 26, 32, 61, 58, 51, 39, 32, 
    34, 27, 27, 0, 0, 0, 4, 21, 0, 0, 5, 0, 40, 28, 32, 
    48, 44, 45, 46, 48, 27, 42, 54, 37, 38, 42, 36, 43, 40, 43, 
    22, 22, 22, 24, 27, 25, 30, 39, 34, 38, 38, 43, 42, 38, 39, 
    15, 24, 21, 23, 18, 19, 23, 23, 18, 18, 20, 19, 20, 20, 37, 
    6, 17, 17, 20, 16, 17, 14, 17, 12, 14, 16, 19, 24, 49, 43, 
    
    -- channel=237
    0, 0, 27, 4, 0, 0, 3, 0, 3, 0, 0, 1, 0, 0, 0, 
    0, 0, 7, 54, 0, 0, 9, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 31, 1, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 25, 0, 0, 12, 0, 5, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 4, 6, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 28, 54, 0, 0, 0, 0, 0, 1, 6, 0, 1, 0, 0, 0, 
    0, 0, 6, 61, 45, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 
    0, 0, 1, 4, 139, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 24, 128, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 28, 72, 0, 0, 8, 42, 0, 22, 0, 0, 0, 
    0, 0, 1, 0, 0, 11, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 1, 6, 2, 1, 3, 0, 0, 6, 0, 1, 0, 0, 3, 3, 
    21, 3, 6, 3, 9, 5, 3, 1, 3, 7, 1, 1, 1, 0, 0, 
    24, 4, 1, 0, 4, 0, 5, 0, 5, 5, 7, 4, 0, 0, 18, 
    
    -- channel=238
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 0, 8, 
    
    -- channel=239
    0, 9, 37, 9, 0, 14, 16, 8, 11, 8, 10, 13, 1, 8, 15, 
    0, 4, 34, 45, 0, 6, 20, 0, 13, 11, 14, 0, 6, 19, 14, 
    0, 5, 27, 30, 35, 4, 19, 0, 15, 15, 9, 0, 0, 20, 15, 
    0, 3, 56, 9, 4, 6, 22, 0, 3, 24, 2, 12, 0, 16, 13, 
    5, 2, 21, 38, 14, 14, 12, 8, 16, 27, 10, 0, 11, 15, 13, 
    9, 18, 31, 19, 13, 12, 8, 14, 18, 16, 13, 4, 17, 16, 8, 
    3, 42, 31, 0, 0, 16, 10, 14, 17, 21, 15, 21, 19, 19, 15, 
    0, 18, 44, 71, 1, 0, 2, 19, 20, 24, 16, 18, 17, 19, 11, 
    0, 16, 23, 39, 125, 0, 0, 0, 20, 28, 11, 16, 17, 18, 13, 
    0, 17, 21, 42, 153, 4, 1, 5, 0, 5, 0, 18, 25, 23, 12, 
    0, 18, 18, 63, 25, 36, 0, 0, 6, 14, 0, 0, 0, 0, 0, 
    16, 47, 52, 51, 47, 74, 41, 13, 38, 39, 26, 34, 20, 21, 23, 
    5, 12, 17, 19, 17, 19, 12, 3, 24, 17, 21, 14, 18, 25, 17, 
    17, 9, 15, 11, 18, 10, 8, 8, 15, 16, 9, 11, 10, 10, 0, 
    21, 10, 10, 6, 13, 0, 4, 0, 7, 4, 8, 13, 0, 0, 39, 
    
    -- channel=240
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 0, 5, 1, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 7, 4, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 6, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 87, 109, 86, 87, 86, 80, 102, 88, 64, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 11, 12, 12, 12, 15, 3, 0, 13, 34, 0, 
    
    -- channel=241
    32, 19, 6, 11, 20, 15, 14, 20, 19, 19, 18, 15, 26, 21, 14, 
    31, 18, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 16, 8, 11, 
    28, 18, 0, 0, 2, 25, 5, 24, 21, 18, 18, 17, 13, 10, 12, 
    29, 20, 0, 17, 19, 18, 13, 21, 18, 3, 16, 18, 36, 10, 11, 
    25, 22, 14, 0, 7, 6, 10, 12, 5, 0, 8, 26, 17, 12, 13, 
    21, 4, 0, 19, 29, 30, 31, 26, 25, 23, 24, 22, 12, 13, 19, 
    22, 14, 6, 0, 0, 4, 17, 16, 15, 11, 11, 8, 7, 6, 8, 
    24, 16, 16, 22, 0, 0, 0, 6, 7, 6, 11, 11, 13, 12, 16, 
    23, 12, 7, 3, 0, 2, 0, 0, 0, 0, 9, 14, 11, 10, 13, 
    21, 8, 7, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 11, 
    22, 8, 9, 0, 64, 51, 68, 102, 65, 50, 80, 60, 90, 38, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 8, 6, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 43, 
    0, 0, 1, 2, 0, 16, 12, 14, 11, 13, 5, 0, 23, 35, 0, 
    
    -- channel=242
    40, 51, 50, 40, 44, 46, 45, 44, 43, 44, 45, 45, 45, 49, 51, 
    39, 49, 57, 50, 42, 51, 49, 45, 52, 53, 51, 47, 57, 57, 53, 
    39, 47, 58, 56, 63, 57, 55, 58, 63, 62, 61, 52, 54, 54, 54, 
    41, 48, 61, 46, 49, 49, 53, 49, 49, 53, 47, 54, 39, 52, 54, 
    46, 47, 53, 57, 45, 44, 44, 47, 49, 49, 43, 50, 55, 53, 53, 
    48, 50, 50, 53, 50, 49, 51, 55, 53, 50, 49, 48, 55, 54, 52, 
    47, 52, 29, 27, 43, 52, 55, 57, 56, 55, 54, 55, 54, 55, 55, 
    46, 56, 58, 40, 16, 25, 46, 55, 57, 57, 53, 54, 54, 54, 53, 
    47, 54, 55, 60, 47, 4, 6, 28, 45, 52, 53, 56, 54, 53, 53, 
    48, 54, 56, 57, 54, 4, 5, 7, 5, 12, 18, 36, 45, 51, 54, 
    48, 55, 55, 61, 40, 20, 3, 8, 26, 21, 9, 8, 10, 35, 46, 
    45, 54, 51, 50, 49, 56, 43, 41, 56, 52, 51, 54, 51, 57, 54, 
    22, 28, 27, 22, 17, 19, 19, 21, 26, 24, 24, 23, 25, 27, 22, 
    11, 9, 10, 4, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=243
    54, 55, 52, 40, 41, 44, 45, 41, 47, 44, 45, 43, 47, 59, 60, 
    53, 57, 50, 5, 0, 0, 0, 1, 3, 8, 7, 11, 51, 50, 54, 
    49, 57, 46, 10, 28, 33, 19, 27, 38, 43, 44, 46, 46, 56, 55, 
    52, 54, 33, 0, 10, 11, 18, 7, 6, 0, 1, 13, 22, 49, 53, 
    59, 56, 54, 51, 38, 35, 35, 39, 39, 36, 38, 42, 56, 57, 56, 
    60, 59, 43, 51, 69, 67, 66, 65, 64, 67, 65, 64, 53, 54, 56, 
    59, 50, 41, 0, 1, 43, 52, 54, 56, 57, 54, 55, 54, 52, 51, 
    60, 60, 62, 82, 35, 0, 22, 50, 51, 48, 52, 54, 56, 55, 56, 
    60, 59, 59, 53, 45, 10, 0, 0, 4, 34, 41, 53, 53, 53, 54, 
    58, 54, 56, 58, 6, 0, 0, 10, 10, 0, 0, 0, 12, 38, 52, 
    55, 51, 54, 44, 52, 80, 31, 38, 82, 52, 65, 48, 51, 60, 45, 
    25, 17, 14, 10, 7, 7, 31, 30, 12, 22, 28, 29, 33, 14, 15, 
    30, 24, 29, 29, 32, 30, 29, 23, 13, 9, 7, 4, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 4, 7, 7, 8, 39, 
    9, 8, 7, 9, 7, 12, 15, 15, 17, 17, 16, 14, 19, 59, 36, 
    
    -- channel=244
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 5, 7, 7, 4, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 8, 0, 0, 0, 20, 23, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 6, 8, 
    7, 13, 11, 7, 5, 6, 5, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    14, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 0, 0, 20, 35, 32, 33, 27, 30, 32, 33, 9, 2, 0, 
    17, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 
    5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 13, 7, 8, 
    0, 4, 0, 0, 8, 11, 11, 5, 8, 7, 8, 15, 0, 0, 2, 
    0, 0, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    5, 0, 0, 69, 101, 29, 0, 0, 0, 0, 0, 0, 1, 4, 10, 
    10, 0, 0, 0, 0, 96, 77, 13, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 12, 61, 116, 98, 46, 22, 0, 0, 0, 2, 
    12, 2, 0, 0, 0, 24, 21, 4, 18, 69, 133, 128, 95, 41, 6, 
    19, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    76, 72, 82, 89, 96, 70, 38, 54, 66, 39, 39, 28, 31, 53, 54, 
    0, 0, 0, 0, 0, 0, 0, 16, 27, 38, 42, 51, 56, 54, 63, 
    32, 44, 40, 34, 25, 26, 22, 21, 14, 8, 9, 5, 6, 7, 0, 
    0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 
    
    -- channel=246
    38, 54, 57, 47, 38, 48, 48, 44, 48, 46, 48, 47, 48, 63, 63, 
    42, 53, 61, 50, 34, 36, 37, 34, 42, 42, 40, 34, 55, 60, 61, 
    38, 52, 67, 39, 45, 39, 43, 36, 47, 55, 51, 56, 49, 63, 62, 
    43, 50, 54, 22, 25, 28, 33, 27, 25, 26, 20, 31, 26, 57, 58, 
    50, 51, 55, 59, 40, 39, 37, 42, 44, 42, 40, 41, 61, 62, 59, 
    55, 64, 54, 47, 64, 62, 63, 64, 64, 65, 63, 64, 58, 60, 59, 
    55, 53, 43, 17, 14, 47, 58, 61, 63, 64, 61, 62, 61, 60, 57, 
    56, 63, 66, 74, 39, 6, 30, 56, 61, 59, 59, 60, 60, 60, 58, 
    58, 65, 68, 66, 64, 4, 2, 3, 24, 45, 48, 61, 60, 59, 58, 
    57, 65, 65, 74, 41, 0, 0, 4, 6, 0, 0, 8, 28, 47, 56, 
    51, 62, 63, 60, 40, 56, 5, 7, 59, 37, 33, 26, 23, 54, 49, 
    38, 45, 41, 37, 33, 33, 41, 37, 32, 34, 40, 39, 43, 31, 32, 
    21, 20, 24, 24, 24, 21, 22, 20, 18, 12, 12, 9, 8, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 3, 2, 4, 0, 0, 22, 37, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=248
    0, 0, 13, 2, 0, 0, 5, 0, 4, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 40, 0, 0, 8, 0, 4, 1, 2, 0, 0, 0, 0, 
    0, 0, 0, 20, 15, 8, 21, 2, 11, 14, 8, 6, 0, 0, 0, 
    0, 0, 11, 27, 8, 4, 19, 8, 10, 20, 5, 11, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 66, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 92, 0, 0, 4, 8, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 25, 77, 11, 0, 31, 35, 21, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 2, 1, 11, 6, 4, 3, 8, 12, 6, 9, 8, 5, 0, 
    24, 9, 8, 8, 11, 3, 13, 8, 15, 13, 15, 12, 0, 0, 23, 
    
    -- channel=249
    87, 99, 83, 81, 80, 85, 81, 80, 80, 82, 83, 82, 85, 92, 95, 
    96, 107, 98, 53, 72, 77, 72, 74, 75, 78, 77, 75, 97, 98, 99, 
    95, 105, 106, 45, 40, 35, 29, 35, 36, 43, 45, 51, 90, 99, 101, 
    93, 105, 78, 22, 47, 51, 37, 40, 51, 46, 49, 55, 69, 102, 103, 
    94, 103, 98, 83, 79, 79, 81, 81, 84, 78, 78, 88, 91, 103, 103, 
    99, 103, 99, 96, 90, 88, 90, 91, 89, 91, 90, 97, 100, 99, 102, 
    99, 83, 62, 81, 97, 101, 102, 103, 102, 100, 101, 100, 102, 102, 102, 
    104, 105, 89, 42, 42, 86, 100, 101, 100, 97, 97, 99, 100, 99, 102, 
    106, 105, 103, 94, 27, 31, 53, 83, 93, 95, 98, 100, 101, 101, 102, 
    102, 101, 102, 100, 30, 20, 23, 23, 32, 47, 71, 89, 94, 97, 100, 
    100, 100, 102, 82, 38, 13, 18, 37, 41, 23, 26, 23, 59, 77, 94, 
    94, 96, 94, 93, 92, 81, 74, 85, 92, 81, 88, 83, 90, 93, 94, 
    46, 50, 48, 46, 44, 43, 45, 55, 57, 57, 57, 60, 62, 60, 56, 
    26, 32, 31, 26, 23, 21, 22, 22, 20, 15, 15, 15, 15, 12, 27, 
    8, 14, 15, 15, 12, 14, 14, 14, 15, 14, 14, 12, 14, 43, 50, 
    
    -- channel=250
    1, 10, 12, 10, 12, 12, 13, 7, 7, 9, 10, 12, 1, 4, 9, 
    1, 12, 14, 46, 30, 50, 54, 42, 48, 46, 49, 33, 18, 20, 16, 
    3, 12, 22, 25, 18, 0, 10, 2, 0, 0, 0, 0, 20, 16, 16, 
    1, 10, 37, 10, 20, 17, 16, 16, 22, 38, 29, 24, 3, 20, 20, 
    5, 9, 10, 25, 17, 19, 15, 16, 20, 25, 18, 6, 7, 14, 14, 
    9, 16, 34, 10, 0, 0, 0, 0, 0, 0, 0, 3, 16, 14, 9, 
    10, 16, 9, 52, 49, 28, 14, 14, 12, 14, 15, 17, 19, 22, 21, 
    10, 14, 0, 0, 3, 41, 39, 25, 21, 22, 16, 15, 14, 15, 13, 
    11, 16, 18, 20, 24, 5, 35, 66, 62, 45, 23, 15, 17, 17, 15, 
    14, 21, 20, 37, 75, 12, 5, 0, 17, 59, 69, 80, 61, 35, 18, 
    16, 20, 19, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    58, 75, 80, 83, 84, 72, 40, 45, 68, 38, 45, 32, 45, 55, 50, 
    0, 3, 0, 0, 0, 0, 0, 13, 29, 30, 36, 37, 41, 46, 47, 
    26, 32, 29, 19, 19, 16, 11, 9, 8, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    
    -- channel=251
    17, 30, 26, 18, 20, 20, 17, 17, 17, 17, 18, 18, 17, 20, 24, 
    25, 38, 28, 6, 5, 15, 14, 14, 14, 15, 18, 18, 25, 27, 29, 
    26, 37, 30, 14, 0, 0, 0, 0, 0, 0, 0, 2, 24, 28, 30, 
    26, 35, 16, 0, 0, 2, 0, 0, 3, 0, 0, 0, 14, 30, 34, 
    25, 34, 32, 27, 24, 26, 25, 24, 28, 23, 20, 21, 27, 31, 35, 
    22, 36, 42, 24, 22, 21, 22, 23, 23, 22, 20, 29, 31, 29, 31, 
    20, 22, 12, 35, 38, 32, 31, 32, 31, 31, 31, 32, 32, 33, 34, 
    21, 31, 14, 0, 11, 32, 32, 29, 31, 29, 28, 29, 30, 30, 34, 
    20, 27, 28, 19, 7, 0, 11, 34, 36, 32, 30, 30, 32, 32, 34, 
    16, 25, 27, 31, 14, 0, 0, 0, 0, 15, 37, 41, 35, 30, 31, 
    18, 28, 28, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 27, 
    33, 46, 45, 45, 47, 37, 28, 34, 45, 38, 38, 34, 40, 46, 46, 
    1, 8, 7, 4, 3, 2, 5, 15, 20, 21, 22, 25, 27, 26, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    43, 47, 45, 42, 46, 41, 41, 40, 40, 41, 42, 43, 40, 42, 47, 
    48, 55, 48, 41, 58, 70, 68, 66, 68, 69, 66, 59, 57, 54, 52, 
    48, 54, 60, 47, 34, 32, 31, 35, 30, 31, 38, 42, 55, 51, 53, 
    47, 53, 41, 28, 37, 38, 30, 34, 42, 39, 37, 35, 48, 54, 56, 
    47, 52, 49, 50, 48, 49, 49, 50, 53, 49, 46, 47, 49, 52, 55, 
    46, 56, 64, 45, 38, 36, 39, 41, 40, 39, 38, 47, 53, 51, 52, 
    46, 41, 31, 74, 74, 57, 54, 55, 53, 53, 54, 54, 54, 56, 57, 
    48, 52, 33, 0, 35, 71, 64, 56, 56, 53, 51, 52, 51, 51, 54, 
    48, 52, 51, 44, 28, 18, 48, 79, 76, 65, 57, 53, 54, 54, 55, 
    47, 51, 53, 62, 46, 21, 17, 13, 25, 55, 82, 85, 73, 59, 55, 
    50, 52, 54, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 51, 
    74, 81, 83, 84, 86, 74, 57, 64, 80, 63, 66, 59, 66, 77, 73, 
    30, 32, 31, 27, 25, 26, 29, 42, 49, 51, 53, 57, 61, 61, 60, 
    34, 34, 33, 25, 20, 20, 18, 17, 13, 10, 8, 8, 8, 1, 0, 
    13, 9, 8, 7, 5, 3, 2, 0, 0, 0, 2, 1, 0, 0, 19, 
    
    -- channel=253
    4, 1, 0, 15, 9, 9, 13, 12, 12, 12, 13, 12, 13, 17, 16, 
    0, 0, 0, 41, 49, 49, 48, 50, 51, 47, 48, 42, 14, 13, 14, 
    0, 0, 1, 49, 44, 45, 54, 52, 44, 44, 42, 36, 26, 9, 12, 
    0, 0, 6, 40, 34, 31, 32, 35, 30, 36, 38, 37, 26, 9, 6, 
    2, 0, 0, 5, 4, 4, 2, 6, 6, 6, 10, 5, 12, 5, 4, 
    11, 3, 0, 4, 4, 4, 6, 8, 8, 7, 7, 5, 4, 7, 6, 
    12, 4, 1, 6, 7, 4, 6, 7, 9, 9, 8, 7, 6, 6, 5, 
    13, 9, 19, 23, 8, 5, 12, 11, 10, 10, 9, 8, 7, 5, 2, 
    17, 16, 15, 23, 15, 15, 8, 10, 16, 13, 9, 8, 8, 6, 4, 
    21, 19, 15, 15, 18, 13, 16, 21, 14, 3, 0, 9, 13, 12, 8, 
    18, 15, 15, 24, 24, 16, 10, 19, 27, 15, 18, 12, 15, 11, 11, 
    13, 8, 8, 7, 5, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 8, 7, 10, 11, 10, 8, 3, 4, 3, 2, 1, 1, 2, 2, 
    12, 11, 11, 13, 16, 13, 12, 14, 16, 15, 15, 15, 15, 12, 4, 
    19, 14, 15, 16, 17, 16, 18, 20, 20, 19, 19, 18, 12, 3, 10, 
    
    -- channel=254
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 32, 0, 0, 7, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 2, 0, 1, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 24, 0, 29, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    14, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 8, 0, 0, 
    
    -- channel=255
    0, 0, 9, 0, 8, 11, 13, 14, 13, 16, 11, 13, 8, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 23, 17, 19, 16, 19, 24, 28, 27, 21, 13, 0, 0, 
    0, 0, 0, 0, 2, 3, 9, 3, 0, 8, 6, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 4, 0, 0, 13, 33, 15, 0, 0, 0, 0, 
    0, 0, 0, 26, 21, 12, 48, 20, 0, 28, 11, 40, 1, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 18, 15, 16, 13, 15, 9, 7, 4, 5, 4, 0, 4, 15, 14, 
    4, 4, 4, 1, 5, 11, 2, 5, 8, 5, 0, 0, 20, 0, 0, 
    
    -- channel=256
    0, 0, 6, 0, 0, 38, 0, 14, 0, 4, 0, 49, 0, 22, 4, 
    0, 0, 0, 0, 0, 16, 0, 23, 0, 4, 0, 60, 0, 26, 0, 
    0, 4, 0, 0, 0, 40, 12, 0, 9, 0, 25, 51, 0, 0, 0, 
    0, 42, 0, 0, 11, 24, 0, 0, 33, 0, 29, 26, 0, 0, 0, 
    0, 46, 0, 0, 45, 1, 0, 40, 3, 17, 0, 16, 0, 0, 0, 
    0, 41, 0, 0, 14, 14, 0, 32, 0, 0, 0, 38, 0, 0, 0, 
    0, 24, 9, 0, 1, 28, 23, 16, 11, 22, 27, 24, 0, 1, 0, 
    0, 17, 7, 0, 30, 0, 39, 22, 29, 28, 14, 30, 0, 0, 0, 
    8, 3, 0, 0, 18, 18, 26, 22, 23, 21, 11, 18, 0, 0, 0, 
    0, 0, 0, 11, 1, 13, 33, 27, 17, 11, 17, 6, 0, 0, 23, 
    0, 26, 0, 18, 0, 5, 49, 16, 9, 1, 22, 13, 0, 5, 0, 
    29, 29, 0, 0, 0, 18, 34, 22, 10, 1, 32, 11, 1, 6, 0, 
    0, 33, 2, 0, 0, 8, 18, 0, 35, 22, 15, 8, 0, 8, 0, 
    0, 2, 50, 13, 0, 0, 0, 0, 29, 22, 23, 0, 0, 20, 28, 
    0, 3, 33, 46, 10, 0, 0, 0, 0, 18, 6, 10, 0, 12, 46, 
    
    -- channel=257
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 2, 6, 15, 2, 2, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 10, 3, 20, 24, 0, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 16, 5, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 3, 11, 0, 8, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 4, 5, 0, 6, 9, 0, 0, 
    0, 15, 3, 0, 0, 0, 0, 1, 0, 2, 11, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 9, 7, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    
    -- channel=258
    27, 17, 43, 39, 0, 68, 25, 41, 31, 40, 9, 73, 0, 65, 37, 
    26, 15, 25, 36, 0, 56, 42, 54, 27, 35, 10, 84, 0, 50, 15, 
    14, 33, 32, 21, 0, 67, 46, 17, 50, 5, 61, 77, 0, 30, 16, 
    20, 82, 10, 13, 36, 60, 18, 18, 72, 10, 62, 60, 10, 21, 0, 
    6, 83, 0, 8, 51, 30, 0, 64, 35, 43, 20, 52, 16, 21, 0, 
    0, 83, 27, 0, 57, 27, 0, 23, 9, 23, 16, 51, 0, 33, 0, 
    0, 62, 49, 8, 0, 9, 5, 16, 10, 8, 5, 13, 8, 34, 0, 
    12, 58, 36, 20, 11, 0, 30, 3, 0, 7, 1, 21, 0, 24, 0, 
    33, 29, 18, 29, 30, 0, 11, 0, 2, 12, 0, 1, 0, 0, 0, 
    15, 14, 14, 43, 32, 43, 0, 4, 0, 0, 0, 0, 0, 25, 56, 
    0, 55, 4, 54, 27, 15, 59, 0, 0, 0, 1, 2, 0, 25, 28, 
    38, 21, 0, 45, 18, 41, 24, 3, 0, 0, 7, 0, 0, 27, 32, 
    26, 59, 4, 1, 14, 41, 11, 0, 34, 0, 0, 0, 0, 39, 30, 
    7, 54, 85, 29, 0, 25, 37, 20, 39, 8, 3, 0, 0, 54, 60, 
    0, 26, 80, 74, 21, 4, 16, 36, 11, 13, 0, 11, 7, 50, 84, 
    
    -- channel=259
    0, 0, 0, 0, 4, 0, 0, 2, 10, 19, 8, 0, 0, 7, 0, 
    0, 0, 0, 0, 7, 8, 11, 0, 0, 0, 2, 0, 0, 0, 0, 
    32, 28, 1, 7, 8, 0, 0, 5, 13, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 24, 0, 0, 0, 0, 9, 0, 12, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 3, 24, 0, 0, 12, 
    13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 
    0, 0, 8, 1, 4, 1, 0, 0, 4, 6, 0, 0, 1, 0, 1, 
    5, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 21, 
    0, 0, 19, 15, 27, 0, 0, 0, 0, 0, 1, 0, 32, 30, 0, 
    3, 24, 16, 15, 9, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 3, 3, 0, 0, 0, 8, 3, 7, 
    47, 57, 0, 0, 0, 8, 15, 46, 43, 0, 0, 0, 2, 19, 17, 
    4, 58, 55, 0, 0, 0, 0, 0, 0, 7, 0, 11, 31, 12, 0, 
    13, 0, 30, 44, 7, 0, 0, 0, 19, 34, 49, 16, 0, 0, 0, 
    
    -- channel=260
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 36, 2, 1, 0, 
    0, 22, 0, 0, 0, 17, 0, 0, 0, 0, 18, 24, 5, 8, 0, 
    0, 37, 0, 0, 20, 5, 0, 9, 11, 18, 4, 9, 6, 7, 0, 
    0, 25, 14, 0, 12, 0, 0, 37, 4, 0, 0, 31, 0, 8, 0, 
    0, 14, 11, 6, 0, 13, 15, 4, 0, 13, 22, 16, 0, 12, 0, 
    0, 9, 8, 6, 36, 0, 22, 22, 31, 26, 9, 38, 5, 3, 0, 
    6, 10, 0, 0, 15, 24, 26, 27, 23, 16, 16, 21, 0, 0, 0, 
    1, 0, 0, 0, 0, 11, 32, 36, 27, 25, 17, 12, 0, 0, 10, 
    0, 7, 0, 12, 0, 0, 44, 31, 26, 8, 15, 11, 0, 4, 16, 
    25, 56, 0, 3, 0, 9, 32, 26, 23, 9, 31, 15, 0, 13, 0, 
    0, 28, 28, 8, 0, 19, 22, 0, 18, 25, 28, 6, 0, 0, 0, 
    0, 0, 23, 35, 9, 3, 1, 6, 23, 23, 26, 0, 0, 0, 6, 
    0, 0, 0, 34, 39, 24, 8, 3, 0, 9, 4, 1, 0, 0, 44, 
    
    -- channel=261
    16, 14, 25, 4, 0, 13, 8, 3, 0, 0, 0, 3, 0, 0, 1, 
    9, 20, 5, 5, 0, 0, 0, 1, 10, 9, 0, 6, 16, 43, 16, 
    0, 0, 0, 0, 0, 24, 35, 5, 0, 0, 0, 12, 13, 9, 9, 
    0, 28, 5, 0, 10, 35, 0, 0, 0, 11, 33, 2, 0, 7, 0, 
    4, 11, 22, 0, 22, 13, 0, 30, 30, 25, 4, 0, 0, 0, 0, 
    0, 0, 0, 35, 26, 0, 13, 46, 19, 0, 0, 23, 0, 0, 0, 
    17, 7, 0, 3, 0, 0, 14, 0, 0, 0, 14, 4, 0, 3, 0, 
    0, 0, 0, 0, 32, 0, 0, 3, 22, 23, 0, 5, 12, 0, 0, 
    18, 14, 0, 0, 0, 26, 9, 5, 2, 0, 0, 0, 0, 0, 5, 
    2, 0, 0, 0, 0, 0, 3, 14, 0, 2, 0, 0, 0, 0, 4, 
    0, 3, 2, 12, 0, 3, 0, 0, 1, 0, 0, 0, 0, 7, 27, 
    32, 81, 38, 2, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 0, 
    0, 0, 16, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 25, 7, 0, 10, 13, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 5, 32, 22, 0, 0, 0, 0, 0, 23, 24, 24, 
    
    -- channel=262
    8, 1, 24, 6, 0, 1, 12, 3, 19, 0, 1, 7, 15, 0, 0, 
    11, 18, 13, 9, 0, 6, 0, 5, 9, 21, 1, 19, 4, 35, 28, 
    2, 0, 0, 3, 0, 3, 32, 27, 0, 7, 0, 31, 25, 24, 12, 
    0, 15, 23, 0, 0, 47, 23, 0, 10, 0, 43, 45, 9, 22, 14, 
    8, 23, 17, 7, 14, 30, 4, 6, 38, 35, 33, 11, 23, 16, 0, 
    0, 15, 4, 17, 51, 8, 2, 46, 36, 23, 9, 40, 25, 10, 0, 
    8, 26, 16, 16, 18, 16, 15, 31, 2, 10, 12, 35, 13, 28, 0, 
    0, 11, 23, 9, 19, 20, 6, 11, 23, 31, 27, 10, 32, 19, 0, 
    10, 37, 12, 2, 6, 7, 30, 13, 31, 10, 5, 34, 0, 8, 0, 
    26, 0, 2, 3, 8, 0, 11, 29, 13, 27, 10, 16, 7, 5, 0, 
    5, 6, 12, 10, 24, 14, 10, 27, 22, 7, 10, 8, 14, 5, 50, 
    1, 79, 51, 38, 10, 7, 31, 14, 11, 9, 21, 19, 8, 28, 11, 
    14, 0, 29, 53, 31, 22, 17, 9, 0, 8, 24, 9, 17, 2, 20, 
    8, 3, 0, 18, 51, 44, 23, 1, 33, 17, 12, 13, 0, 5, 0, 
    3, 2, 19, 4, 20, 53, 49, 34, 14, 0, 4, 0, 7, 23, 63, 
    
    -- channel=263
    22, 0, 18, 15, 23, 0, 27, 9, 42, 26, 36, 0, 64, 8, 0, 
    11, 2, 27, 18, 13, 17, 13, 0, 33, 23, 38, 0, 44, 7, 35, 
    39, 23, 11, 17, 2, 0, 9, 40, 17, 27, 22, 0, 57, 22, 41, 
    19, 1, 23, 11, 0, 35, 56, 4, 1, 0, 25, 16, 59, 31, 69, 
    18, 28, 35, 22, 9, 39, 26, 0, 40, 22, 57, 24, 45, 33, 57, 
    18, 33, 36, 2, 26, 12, 19, 45, 37, 31, 30, 8, 53, 33, 50, 
    9, 21, 23, 40, 38, 27, 11, 18, 18, 27, 18, 19, 35, 31, 36, 
    15, 16, 14, 42, 30, 4, 19, 28, 27, 5, 8, 27, 33, 34, 24, 
    9, 23, 30, 31, 32, 23, 23, 27, 24, 19, 25, 25, 44, 45, 16, 
    35, 29, 22, 33, 32, 34, 22, 24, 25, 40, 18, 33, 32, 10, 0, 
    38, 16, 24, 22, 18, 14, 19, 36, 32, 34, 24, 25, 26, 3, 47, 
    0, 35, 30, 13, 38, 15, 37, 37, 26, 28, 28, 35, 40, 26, 35, 
    50, 51, 57, 41, 27, 39, 47, 64, 24, 24, 39, 23, 43, 5, 48, 
    41, 30, 48, 49, 48, 32, 33, 15, 3, 38, 27, 35, 40, 21, 2, 
    51, 19, 29, 55, 59, 44, 46, 32, 32, 47, 60, 19, 0, 2, 29, 
    
    -- channel=264
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 23, 
    0, 0, 24, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 42, 
    0, 0, 0, 29, 0, 0, 2, 0, 0, 0, 2, 0, 2, 0, 46, 
    0, 0, 0, 8, 13, 4, 5, 2, 2, 0, 5, 2, 0, 0, 36, 
    0, 0, 0, 0, 21, 0, 0, 8, 20, 18, 10, 0, 34, 0, 16, 
    0, 0, 0, 0, 0, 40, 0, 14, 16, 12, 12, 2, 19, 0, 9, 
    0, 0, 0, 0, 0, 0, 19, 16, 17, 28, 11, 17, 20, 0, 0, 
    10, 0, 0, 0, 0, 2, 0, 27, 24, 18, 14, 15, 9, 0, 0, 
    2, 10, 18, 0, 0, 0, 0, 18, 16, 29, 19, 15, 11, 0, 0, 
    0, 0, 19, 5, 0, 0, 2, 7, 0, 22, 12, 29, 13, 0, 0, 
    0, 0, 0, 0, 19, 0, 0, 1, 0, 5, 13, 19, 9, 0, 0, 
    2, 0, 0, 0, 1, 20, 1, 0, 0, 0, 0, 1, 4, 0, 0, 
    
    -- channel=265
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 32, 0, 0, 0, 8, 0, 0, 17, 0, 0, 0, 0, 0, 5, 
    0, 8, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 32, 0, 0, 0, 0, 0, 13, 15, 0, 0, 0, 0, 
    
    -- channel=266
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=267
    5, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 8, 
    15, 13, 0, 0, 0, 0, 0, 2, 0, 0, 0, 25, 22, 31, 5, 
    0, 0, 0, 0, 0, 15, 22, 0, 0, 0, 2, 30, 30, 18, 21, 
    0, 31, 0, 0, 6, 9, 0, 0, 5, 18, 15, 24, 13, 27, 0, 
    0, 25, 28, 0, 30, 12, 0, 37, 9, 30, 1, 0, 18, 23, 0, 
    0, 0, 32, 48, 14, 18, 31, 44, 26, 9, 3, 43, 8, 14, 0, 
    11, 8, 7, 32, 15, 23, 42, 21, 15, 24, 43, 39, 9, 23, 0, 
    0, 10, 26, 19, 62, 0, 27, 41, 52, 62, 40, 41, 48, 14, 0, 
    30, 26, 0, 0, 3, 83, 30, 41, 43, 33, 33, 36, 6, 0, 12, 
    13, 0, 0, 0, 0, 0, 64, 61, 47, 46, 38, 30, 9, 2, 27, 
    0, 15, 5, 12, 15, 32, 40, 55, 50, 21, 34, 31, 22, 29, 18, 
    79, 91, 41, 15, 0, 22, 39, 41, 43, 40, 54, 28, 8, 12, 2, 
    0, 0, 49, 37, 18, 13, 18, 0, 2, 55, 31, 35, 3, 0, 0, 
    0, 0, 0, 47, 41, 16, 2, 33, 34, 26, 46, 14, 0, 0, 32, 
    0, 0, 0, 0, 45, 59, 27, 13, 0, 0, 0, 9, 36, 23, 30, 
    
    -- channel=268
    0, 0, 17, 0, 0, 53, 0, 18, 0, 1, 0, 62, 0, 27, 3, 
    0, 0, 0, 0, 0, 34, 0, 36, 0, 13, 0, 81, 0, 42, 0, 
    0, 0, 0, 0, 0, 39, 19, 0, 2, 0, 10, 73, 0, 0, 0, 
    0, 47, 0, 0, 8, 40, 0, 0, 62, 0, 40, 51, 0, 0, 0, 
    0, 63, 0, 0, 40, 0, 0, 53, 0, 21, 0, 16, 0, 0, 0, 
    0, 67, 0, 0, 41, 0, 0, 17, 0, 0, 0, 58, 0, 0, 0, 
    0, 41, 25, 0, 0, 0, 0, 3, 0, 1, 0, 12, 0, 11, 0, 
    0, 25, 17, 0, 0, 0, 13, 1, 0, 0, 7, 11, 0, 0, 0, 
    2, 13, 0, 0, 21, 0, 18, 0, 0, 0, 0, 6, 0, 0, 0, 
    2, 0, 0, 16, 0, 31, 0, 3, 0, 0, 0, 0, 0, 0, 27, 
    0, 29, 0, 12, 17, 0, 54, 0, 0, 0, 0, 0, 0, 0, 11, 
    3, 15, 0, 23, 0, 21, 15, 0, 0, 0, 0, 0, 0, 17, 0, 
    13, 22, 0, 0, 0, 20, 0, 0, 17, 0, 0, 0, 0, 22, 0, 
    0, 43, 43, 0, 0, 0, 0, 0, 43, 1, 0, 0, 0, 49, 0, 
    0, 0, 79, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 
    
    -- channel=269
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 18, 10, 7, 16, 15, 4, 0, 0, 0, 
    0, 0, 0, 0, 26, 0, 28, 17, 22, 21, 8, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 17, 20, 19, 22, 14, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 15, 21, 15, 16, 13, 11, 6, 0, 0, 
    0, 1, 0, 0, 0, 0, 27, 11, 17, 8, 18, 18, 3, 0, 0, 
    0, 1, 0, 0, 0, 0, 16, 23, 13, 5, 25, 16, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 20, 18, 11, 5, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 21, 21, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 7, 0, 0, 3, 
    
    -- channel=270
    4, 0, 2, 0, 0, 11, 5, 11, 15, 23, 8, 19, 3, 20, 9, 
    2, 1, 3, 0, 0, 11, 14, 10, 10, 8, 9, 20, 6, 1, 1, 
    13, 22, 7, 0, 0, 9, 1, 2, 15, 3, 23, 17, 8, 7, 5, 
    3, 12, 0, 1, 5, 12, 17, 15, 14, 3, 10, 22, 17, 6, 0, 
    0, 17, 0, 2, 17, 10, 6, 11, 9, 15, 17, 33, 18, 8, 0, 
    1, 20, 11, 0, 8, 20, 11, 7, 12, 17, 19, 25, 19, 10, 0, 
    0, 8, 13, 7, 15, 31, 23, 17, 22, 26, 20, 16, 21, 11, 0, 
    7, 13, 8, 15, 18, 16, 34, 28, 24, 18, 17, 28, 6, 17, 0, 
    5, 3, 8, 15, 25, 14, 19, 25, 24, 31, 30, 21, 23, 17, 5, 
    4, 14, 11, 18, 23, 26, 22, 19, 22, 22, 23, 25, 16, 8, 12, 
    3, 19, 3, 9, 4, 14, 27, 18, 20, 22, 26, 25, 16, 7, 1, 
    3, 0, 6, 6, 7, 14, 21, 30, 23, 15, 22, 25, 30, 21, 10, 
    27, 50, 26, 17, 12, 15, 23, 32, 40, 21, 21, 21, 21, 24, 12, 
    6, 34, 62, 32, 18, 21, 28, 16, 12, 27, 28, 23, 22, 20, 18, 
    8, 12, 30, 58, 32, 16, 19, 25, 22, 32, 33, 33, 4, 1, 23, 
    
    -- channel=271
    3, 0, 0, 10, 13, 0, 0, 0, 0, 1, 6, 0, 2, 0, 0, 
    6, 0, 9, 11, 7, 0, 7, 0, 5, 0, 8, 0, 7, 0, 4, 
    2, 4, 8, 9, 4, 0, 0, 0, 14, 2, 2, 0, 7, 1, 7, 
    10, 0, 0, 0, 0, 0, 0, 8, 0, 4, 0, 0, 17, 8, 19, 
    5, 6, 15, 0, 0, 0, 3, 0, 0, 0, 0, 0, 3, 14, 25, 
    4, 6, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 16, 
    0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 18, 
    3, 5, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 
    3, 0, 12, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 
    5, 10, 4, 1, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    14, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 10, 0, 0, 0, 5, 0, 0, 1, 0, 0, 0, 0, 0, 7, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    6, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=272
    0, 0, 0, 0, 9, 0, 0, 0, 0, 2, 5, 0, 9, 6, 0, 
    0, 0, 0, 0, 8, 0, 9, 0, 0, 0, 2, 0, 8, 0, 0, 
    3, 6, 2, 0, 11, 0, 0, 0, 1, 16, 0, 0, 0, 0, 0, 
    11, 0, 0, 4, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 24, 
    5, 0, 0, 0, 0, 3, 0, 0, 0, 2, 7, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 0, 1, 0, 7, 
    8, 0, 0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 12, 0, 0, 5, 0, 4, 
    0, 9, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 6, 0, 4, 0, 
    8, 19, 7, 0, 0, 0, 0, 2, 0, 0, 0, 0, 24, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 15, 2, 4, 0, 
    
    -- channel=273
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 14, 21, 0, 0, 0, 0, 0, 0, 
    0, 22, 11, 0, 0, 0, 0, 0, 0, 3, 0, 0, 5, 0, 0, 
    0, 0, 14, 1, 0, 0, 0, 0, 0, 7, 18, 0, 0, 0, 0, 
    
    -- channel=274
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=275
    25, 11, 7, 8, 37, 0, 14, 0, 6, 0, 32, 0, 74, 0, 2, 
    21, 8, 17, 12, 28, 0, 2, 0, 22, 2, 35, 0, 83, 3, 31, 
    4, 0, 9, 5, 16, 0, 12, 14, 0, 16, 10, 0, 67, 21, 38, 
    30, 5, 24, 20, 0, 6, 25, 7, 0, 32, 13, 0, 52, 28, 64, 
    22, 0, 70, 13, 0, 23, 50, 0, 28, 13, 24, 0, 34, 26, 78, 
    17, 0, 31, 63, 14, 20, 10, 18, 29, 22, 27, 0, 33, 24, 83, 
    29, 0, 0, 43, 24, 11, 18, 14, 10, 9, 14, 9, 23, 15, 68, 
    18, 1, 8, 29, 52, 0, 8, 16, 28, 28, 13, 10, 45, 12, 43, 
    15, 14, 6, 13, 0, 50, 6, 21, 24, 19, 19, 7, 21, 0, 42, 
    15, 9, 12, 2, 23, 0, 19, 29, 20, 36, 16, 26, 40, 15, 0, 
    40, 2, 26, 13, 3, 31, 0, 33, 37, 24, 18, 25, 24, 7, 26, 
    31, 57, 59, 3, 37, 4, 19, 26, 20, 34, 30, 22, 20, 0, 21, 
    0, 0, 52, 43, 32, 6, 21, 11, 0, 29, 25, 30, 29, 0, 17, 
    41, 0, 0, 38, 54, 28, 20, 38, 0, 17, 22, 21, 22, 0, 20, 
    43, 20, 0, 0, 37, 54, 47, 35, 10, 0, 0, 11, 33, 30, 0, 
    
    -- channel=276
    0, 9, 17, 12, 0, 40, 8, 29, 19, 22, 0, 61, 0, 31, 17, 
    13, 22, 5, 11, 0, 32, 6, 41, 0, 27, 0, 71, 0, 38, 0, 
    10, 10, 11, 11, 0, 30, 27, 14, 19, 4, 5, 75, 0, 18, 0, 
    0, 33, 10, 0, 27, 33, 8, 0, 49, 0, 29, 63, 0, 13, 0, 
    3, 41, 0, 12, 39, 20, 0, 45, 12, 33, 14, 51, 4, 8, 0, 
    0, 45, 1, 0, 38, 31, 7, 23, 16, 24, 6, 64, 0, 9, 0, 
    0, 36, 37, 5, 14, 21, 15, 27, 19, 20, 18, 34, 2, 26, 0, 
    3, 29, 32, 9, 0, 33, 25, 20, 8, 21, 30, 21, 0, 12, 0, 
    17, 30, 20, 14, 41, 0, 34, 13, 20, 20, 11, 31, 0, 7, 0, 
    20, 9, 8, 20, 3, 39, 13, 17, 19, 3, 19, 8, 0, 7, 30, 
    0, 26, 1, 17, 36, 8, 44, 11, 3, 7, 13, 7, 0, 17, 15, 
    20, 19, 0, 42, 0, 35, 29, 13, 11, 1, 12, 11, 3, 27, 10, 
    32, 34, 0, 15, 12, 28, 21, 0, 31, 5, 15, 2, 0, 40, 16, 
    0, 59, 41, 11, 5, 22, 23, 0, 56, 17, 12, 7, 0, 37, 15, 
    0, 0, 74, 50, 7, 11, 13, 21, 26, 13, 12, 0, 0, 13, 70, 
    
    -- channel=277
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 12, 5, 11, 0, 11, 11, 3, 0, 0, 0, 
    0, 0, 0, 0, 6, 8, 10, 5, 15, 12, 8, 12, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 21, 13, 11, 4, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 9, 11, 7, 11, 3, 5, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 9, 6, 6, 10, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 6, 8, 1, 15, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 10, 10, 7, 18, 7, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 4, 4, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 0, 0, 
    
    -- channel=278
    6, 9, 8, 2, 0, 6, 0, 0, 0, 0, 0, 4, 0, 3, 17, 
    7, 8, 0, 0, 0, 0, 0, 14, 0, 0, 0, 9, 14, 13, 0, 
    0, 0, 6, 0, 0, 28, 21, 0, 0, 0, 10, 7, 2, 8, 1, 
    6, 33, 6, 7, 20, 7, 0, 0, 27, 10, 19, 14, 0, 0, 0, 
    0, 1, 9, 0, 0, 0, 9, 31, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 20, 13, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    6, 6, 0, 0, 0, 0, 13, 17, 7, 0, 0, 9, 0, 0, 0, 
    3, 7, 10, 0, 3, 3, 8, 0, 0, 28, 24, 0, 8, 0, 0, 
    7, 5, 0, 0, 0, 7, 0, 0, 11, 15, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 3, 0, 1, 18, 16, 
    0, 7, 2, 1, 9, 11, 7, 0, 0, 0, 0, 6, 3, 8, 0, 
    35, 21, 24, 18, 0, 9, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 9, 17, 0, 0, 0, 0, 1, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 9, 14, 13, 22, 20, 0, 0, 0, 0, 1, 23, 
    0, 13, 0, 0, 0, 10, 10, 22, 0, 0, 0, 0, 36, 41, 18, 
    
    -- channel=279
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=280
    0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 5, 35, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 14, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=281
    0, 8, 0, 0, 42, 0, 3, 0, 6, 0, 19, 0, 75, 0, 0, 
    0, 6, 10, 0, 42, 0, 0, 0, 0, 0, 17, 0, 34, 0, 13, 
    21, 0, 0, 14, 26, 0, 0, 26, 0, 50, 0, 0, 23, 0, 0, 
    18, 0, 29, 3, 0, 0, 21, 12, 0, 0, 0, 0, 2, 0, 64, 
    21, 0, 16, 39, 0, 0, 43, 0, 0, 0, 6, 0, 2, 0, 83, 
    39, 0, 0, 10, 0, 0, 10, 0, 0, 0, 5, 0, 19, 0, 82, 
    18, 0, 0, 0, 14, 0, 0, 8, 2, 0, 0, 0, 10, 0, 48, 
    5, 0, 0, 0, 0, 53, 0, 0, 0, 0, 14, 0, 24, 0, 67, 
    0, 0, 9, 0, 0, 0, 7, 0, 5, 0, 5, 5, 27, 21, 4, 
    5, 6, 14, 0, 0, 3, 0, 0, 2, 12, 0, 13, 32, 5, 0, 
    41, 0, 15, 0, 0, 0, 0, 3, 4, 23, 0, 4, 19, 0, 0, 
    0, 0, 26, 0, 1, 0, 0, 0, 1, 17, 0, 17, 22, 0, 0, 
    9, 0, 0, 11, 3, 0, 0, 57, 0, 0, 14, 17, 38, 0, 0, 
    29, 12, 0, 0, 14, 0, 0, 0, 0, 0, 0, 38, 64, 0, 0, 
    41, 0, 0, 0, 0, 0, 3, 0, 21, 0, 21, 0, 3, 0, 0, 
    
    -- channel=282
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=283
    5, 0, 21, 2, 0, 46, 0, 11, 0, 0, 0, 47, 0, 28, 0, 
    0, 0, 0, 2, 0, 27, 0, 20, 0, 6, 0, 63, 0, 43, 0, 
    0, 0, 0, 0, 0, 43, 24, 0, 9, 0, 31, 58, 0, 0, 0, 
    0, 61, 0, 0, 0, 44, 0, 0, 44, 0, 59, 24, 0, 0, 0, 
    0, 74, 0, 0, 29, 6, 0, 41, 18, 19, 0, 7, 0, 0, 0, 
    0, 69, 2, 0, 40, 3, 0, 31, 0, 0, 0, 28, 0, 3, 0, 
    0, 46, 20, 0, 0, 0, 0, 4, 0, 1, 1, 2, 0, 6, 0, 
    0, 28, 0, 0, 7, 0, 16, 5, 0, 7, 0, 21, 0, 0, 0, 
    8, 9, 0, 0, 12, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 38, 0, 4, 0, 0, 0, 0, 0, 0, 32, 
    0, 28, 0, 35, 0, 0, 64, 0, 0, 0, 0, 0, 0, 3, 10, 
    23, 41, 0, 10, 0, 23, 20, 2, 0, 0, 11, 0, 0, 0, 0, 
    0, 27, 0, 0, 0, 26, 2, 0, 11, 0, 7, 0, 0, 0, 0, 
    0, 0, 41, 3, 0, 0, 0, 0, 25, 5, 0, 0, 0, 17, 15, 
    0, 0, 53, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 77, 
    
    -- channel=284
    16, 0, 0, 0, 10, 0, 4, 0, 0, 4, 15, 0, 35, 0, 0, 
    0, 0, 1, 0, 1, 0, 11, 0, 22, 0, 25, 0, 63, 0, 8, 
    0, 22, 0, 0, 2, 2, 0, 0, 14, 0, 41, 0, 42, 0, 16, 
    16, 7, 0, 12, 0, 0, 0, 11, 0, 37, 0, 0, 51, 6, 23, 
    0, 5, 41, 0, 8, 5, 11, 0, 17, 0, 9, 0, 14, 5, 39, 
    0, 0, 32, 23, 0, 0, 6, 20, 0, 0, 9, 0, 10, 21, 42, 
    5, 0, 0, 16, 1, 8, 17, 0, 0, 5, 13, 0, 12, 0, 41, 
    2, 0, 0, 10, 56, 0, 11, 4, 30, 0, 0, 19, 6, 2, 3, 
    6, 0, 0, 7, 0, 59, 0, 16, 0, 0, 10, 0, 10, 4, 37, 
    0, 2, 0, 3, 30, 0, 23, 7, 0, 13, 0, 5, 30, 0, 0, 
    10, 14, 2, 17, 0, 18, 0, 9, 15, 0, 11, 14, 10, 2, 0, 
    20, 14, 13, 0, 26, 0, 6, 16, 6, 9, 16, 3, 15, 0, 11, 
    0, 33, 55, 2, 4, 6, 6, 0, 15, 26, 3, 10, 10, 0, 0, 
    16, 0, 34, 51, 10, 2, 4, 41, 0, 8, 20, 0, 20, 0, 42, 
    25, 29, 0, 21, 55, 14, 6, 4, 0, 15, 10, 40, 5, 4, 0, 
    
    -- channel=285
    8, 17, 0, 0, 48, 0, 4, 0, 0, 0, 25, 0, 87, 0, 0, 
    3, 7, 6, 0, 49, 0, 0, 0, 3, 0, 26, 0, 80, 0, 14, 
    0, 0, 0, 1, 37, 0, 0, 5, 0, 29, 0, 0, 45, 0, 7, 
    26, 0, 20, 17, 0, 0, 8, 24, 0, 27, 0, 0, 17, 0, 58, 
    23, 0, 52, 21, 0, 0, 62, 0, 0, 0, 0, 0, 6, 0, 95, 
    36, 0, 0, 60, 0, 0, 15, 0, 6, 1, 15, 0, 18, 0, 105, 
    34, 0, 0, 9, 21, 6, 15, 7, 5, 1, 3, 0, 12, 0, 80, 
    13, 0, 0, 0, 23, 29, 0, 6, 20, 20, 13, 0, 43, 0, 72, 
    0, 0, 0, 0, 0, 34, 0, 11, 14, 7, 14, 2, 19, 0, 40, 
    0, 0, 10, 0, 0, 0, 4, 7, 10, 24, 11, 21, 46, 5, 0, 
    42, 0, 21, 0, 0, 11, 0, 15, 20, 22, 8, 18, 26, 0, 0, 
    0, 6, 49, 0, 13, 0, 0, 6, 7, 31, 7, 20, 24, 0, 0, 
    0, 0, 14, 23, 15, 0, 0, 26, 0, 12, 12, 33, 37, 0, 0, 
    32, 0, 0, 0, 31, 5, 0, 21, 0, 1, 5, 32, 54, 0, 0, 
    41, 12, 0, 0, 0, 20, 16, 3, 8, 0, 0, 8, 34, 0, 0, 
    
    -- channel=286
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=287
    13, 15, 0, 5, 28, 0, 1, 0, 0, 0, 14, 0, 36, 0, 4, 
    14, 8, 9, 5, 27, 0, 5, 0, 7, 0, 16, 0, 45, 0, 12, 
    4, 0, 6, 12, 23, 0, 0, 0, 0, 14, 0, 0, 30, 4, 9, 
    23, 0, 14, 15, 5, 0, 0, 15, 0, 22, 0, 0, 20, 7, 35, 
    15, 0, 35, 13, 0, 0, 28, 0, 0, 0, 0, 0, 7, 12, 57, 
    22, 0, 13, 38, 0, 0, 12, 0, 0, 0, 6, 0, 10, 10, 55, 
    24, 0, 0, 12, 5, 0, 7, 2, 6, 0, 7, 0, 13, 0, 46, 
    15, 0, 0, 9, 13, 14, 0, 3, 10, 10, 7, 4, 25, 4, 41, 
    7, 0, 8, 8, 0, 24, 2, 13, 8, 10, 13, 1, 23, 12, 25, 
    4, 12, 10, 0, 6, 0, 10, 12, 15, 17, 13, 13, 31, 13, 0, 
    29, 0, 14, 2, 0, 7, 0, 17, 21, 23, 11, 15, 18, 12, 2, 
    12, 0, 17, 0, 16, 0, 0, 9, 19, 26, 9, 11, 11, 0, 8, 
    0, 0, 7, 0, 3, 0, 2, 14, 0, 18, 14, 23, 15, 0, 0, 
    16, 0, 0, 0, 3, 0, 0, 19, 0, 6, 10, 17, 33, 0, 0, 
    19, 3, 0, 0, 0, 2, 0, 0, 0, 0, 3, 21, 24, 12, 0, 
    
    -- channel=288
    0, 0, 9, 2, 0, 59, 0, 27, 1, 19, 0, 84, 0, 46, 1, 
    0, 0, 0, 1, 0, 39, 6, 34, 0, 10, 0, 103, 0, 35, 0, 
    0, 11, 0, 0, 0, 42, 11, 0, 32, 0, 29, 97, 0, 0, 0, 
    0, 60, 0, 0, 8, 33, 0, 0, 55, 0, 33, 56, 0, 0, 0, 
    0, 87, 0, 0, 51, 0, 0, 47, 0, 19, 0, 49, 0, 0, 0, 
    0, 90, 2, 0, 25, 17, 0, 27, 0, 0, 0, 61, 0, 11, 0, 
    0, 49, 42, 0, 0, 8, 0, 0, 0, 11, 6, 1, 0, 13, 0, 
    0, 41, 15, 0, 2, 0, 29, 0, 0, 0, 0, 39, 0, 0, 0, 
    8, 6, 0, 8, 40, 0, 21, 2, 0, 3, 0, 5, 0, 0, 0, 
    0, 0, 0, 24, 11, 56, 2, 6, 0, 0, 0, 0, 0, 0, 33, 
    0, 41, 0, 32, 0, 0, 77, 0, 0, 0, 0, 0, 0, 5, 0, 
    14, 0, 0, 17, 0, 28, 33, 6, 0, 0, 4, 0, 0, 19, 0, 
    21, 78, 0, 0, 0, 38, 16, 0, 60, 0, 3, 0, 0, 25, 0, 
    0, 47, 101, 6, 0, 0, 3, 0, 39, 14, 6, 0, 0, 36, 28, 
    0, 0, 81, 94, 2, 0, 0, 0, 0, 17, 10, 0, 0, 0, 82, 
    
    -- channel=289
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=290
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=291
    11, 11, 3, 17, 37, 0, 12, 1, 14, 10, 32, 0, 54, 0, 4, 
    15, 10, 20, 18, 33, 0, 12, 0, 16, 7, 31, 0, 45, 0, 23, 
    23, 13, 17, 20, 25, 0, 3, 20, 10, 32, 5, 0, 36, 17, 25, 
    28, 0, 23, 21, 0, 0, 34, 29, 0, 19, 0, 0, 31, 20, 53, 
    26, 0, 41, 15, 0, 15, 43, 0, 14, 2, 20, 4, 27, 21, 68, 
    31, 0, 24, 36, 3, 6, 1, 0, 20, 17, 21, 0, 32, 24, 62, 
    22, 0, 10, 29, 13, 0, 0, 1, 2, 0, 0, 0, 21, 18, 48, 
    25, 4, 12, 22, 0, 0, 0, 0, 0, 0, 0, 0, 19, 18, 52, 
    7, 14, 23, 22, 0, 7, 0, 0, 0, 0, 0, 0, 12, 18, 34, 
    18, 26, 27, 11, 16, 0, 0, 0, 0, 2, 0, 2, 17, 11, 0, 
    47, 0, 28, 5, 13, 17, 0, 4, 3, 6, 0, 0, 9, 6, 21, 
    2, 2, 35, 11, 29, 4, 0, 0, 1, 8, 0, 0, 7, 1, 33, 
    18, 0, 25, 31, 31, 2, 3, 10, 0, 0, 0, 4, 7, 0, 33, 
    32, 0, 0, 13, 35, 26, 15, 10, 0, 0, 0, 6, 25, 0, 18, 
    35, 13, 0, 0, 13, 30, 31, 26, 15, 0, 0, 3, 11, 13, 0, 
    
    -- channel=292
    0, 0, 0, 0, 4, 0, 0, 0, 0, 10, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 7, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 27, 0, 2, 14, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 11, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 3, 
    0, 18, 10, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 32, 0, 0, 0, 0, 0, 15, 29, 0, 0, 0, 0, 9, 0, 
    0, 26, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 7, 22, 16, 0, 0, 0, 
    
    -- channel=293
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 13, 9, 5, 9, 18, 16, 8, 0, 0, 0, 
    0, 0, 0, 2, 16, 3, 19, 25, 20, 12, 16, 32, 15, 0, 0, 
    0, 0, 0, 0, 19, 25, 21, 28, 25, 28, 26, 27, 27, 9, 0, 
    0, 0, 0, 0, 0, 23, 31, 31, 33, 33, 25, 24, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 35, 35, 32, 28, 23, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 38, 36, 24, 28, 28, 12, 4, 0, 
    7, 23, 1, 0, 0, 0, 18, 35, 35, 31, 33, 22, 13, 0, 0, 
    0, 0, 10, 2, 0, 0, 0, 0, 0, 34, 32, 25, 2, 0, 0, 
    0, 0, 0, 10, 11, 0, 0, 0, 0, 30, 34, 12, 0, 0, 0, 
    
    -- channel=294
    0, 0, 0, 4, 11, 0, 1, 0, 5, 2, 7, 0, 10, 0, 0, 
    0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 7, 0, 0, 0, 4, 
    16, 3, 1, 10, 0, 0, 0, 11, 5, 10, 0, 0, 5, 0, 7, 
    2, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 13, 2, 28, 
    5, 0, 5, 1, 0, 0, 0, 0, 0, 0, 3, 0, 2, 9, 27, 
    8, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 16, 
    0, 0, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 13, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 
    0, 0, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 4, 19, 0, 
    12, 11, 6, 4, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    18, 9, 0, 0, 0, 6, 0, 10, 0, 0, 0, 0, 0, 0, 16, 
    5, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    
    -- channel=295
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=296
    25, 39, 24, 30, 39, 18, 31, 28, 23, 27, 31, 17, 40, 16, 25, 
    32, 35, 36, 26, 43, 13, 26, 19, 35, 25, 36, 8, 51, 24, 29, 
    11, 21, 27, 24, 41, 28, 37, 29, 28, 24, 21, 17, 31, 28, 26, 
    37, 18, 25, 26, 38, 25, 34, 46, 5, 45, 20, 19, 28, 26, 20, 
    37, 7, 39, 27, 21, 34, 45, 25, 42, 33, 28, 38, 29, 20, 37, 
    37, 0, 31, 53, 17, 20, 29, 22, 30, 26, 31, 17, 33, 23, 47, 
    39, 12, 18, 26, 24, 16, 19, 8, 7, 9, 13, 6, 30, 21, 53, 
    30, 18, 14, 18, 19, 16, 0, 8, 21, 14, 3, 5, 10, 16, 42, 
    31, 23, 25, 25, 5, 13, 5, 10, 0, 0, 12, 2, 8, 20, 42, 
    16, 26, 24, 8, 21, 4, 8, 0, 5, 2, 5, 8, 17, 12, 28, 
    29, 15, 39, 28, 21, 22, 0, 4, 0, 2, 2, 7, 18, 31, 19, 
    38, 27, 53, 29, 33, 17, 0, 0, 3, 10, 0, 4, 19, 18, 38, 
    0, 9, 41, 48, 42, 20, 14, 1, 0, 7, 3, 10, 11, 24, 29, 
    22, 0, 3, 37, 50, 45, 32, 41, 9, 0, 1, 8, 24, 2, 46, 
    38, 34, 1, 12, 37, 47, 47, 36, 22, 2, 0, 22, 38, 36, 7, 
    
    -- channel=297
    19, 12, 27, 4, 0, 7, 12, 0, 0, 0, 0, 0, 12, 0, 3, 
    8, 16, 5, 5, 0, 0, 0, 0, 11, 7, 0, 0, 30, 43, 18, 
    0, 0, 0, 0, 0, 22, 39, 8, 0, 0, 0, 1, 24, 9, 19, 
    0, 29, 13, 0, 3, 35, 0, 0, 0, 9, 31, 1, 0, 7, 0, 
    5, 8, 25, 0, 13, 15, 0, 29, 31, 27, 8, 0, 0, 0, 0, 
    0, 0, 0, 40, 33, 0, 12, 38, 17, 0, 0, 12, 0, 0, 10, 
    16, 6, 0, 5, 0, 0, 13, 0, 0, 0, 6, 4, 0, 1, 11, 
    0, 0, 0, 0, 32, 0, 0, 6, 18, 27, 2, 0, 20, 0, 0, 
    14, 16, 0, 0, 0, 27, 4, 0, 1, 0, 0, 0, 0, 0, 4, 
    3, 0, 0, 0, 0, 0, 2, 11, 0, 2, 0, 0, 0, 0, 5, 
    0, 1, 5, 8, 4, 1, 0, 0, 0, 0, 0, 0, 1, 2, 23, 
    36, 85, 45, 6, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 15, 29, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 32, 10, 0, 15, 14, 0, 0, 0, 0, 0, 0, 
    1, 15, 0, 0, 2, 37, 25, 1, 0, 0, 0, 0, 30, 27, 27, 
    
    -- channel=298
    26, 16, 36, 18, 0, 30, 28, 28, 39, 28, 21, 41, 28, 23, 21, 
    27, 33, 24, 20, 0, 27, 10, 32, 30, 38, 20, 52, 23, 50, 37, 
    25, 18, 17, 17, 0, 30, 46, 38, 17, 17, 21, 57, 44, 39, 35, 
    8, 39, 33, 18, 15, 62, 39, 0, 41, 11, 61, 68, 40, 40, 23, 
    18, 49, 25, 25, 47, 46, 14, 39, 49, 60, 58, 42, 49, 36, 0, 
    13, 46, 31, 24, 61, 42, 40, 64, 54, 45, 37, 68, 46, 33, 5, 
    21, 45, 38, 39, 50, 60, 55, 61, 46, 54, 53, 65, 38, 47, 5, 
    19, 35, 42, 38, 55, 48, 55, 61, 63, 67, 63, 56, 56, 42, 0, 
    33, 47, 31, 29, 50, 46, 66, 56, 68, 57, 55, 67, 39, 35, 13, 
    42, 25, 20, 35, 31, 42, 55, 65, 58, 64, 53, 56, 37, 27, 28, 
    17, 38, 29, 33, 45, 35, 60, 65, 59, 50, 55, 52, 49, 33, 55, 
    35, 88, 58, 54, 27, 40, 66, 63, 54, 48, 64, 61, 52, 53, 30, 
    46, 46, 62, 68, 48, 50, 56, 52, 37, 53, 63, 52, 50, 34, 36, 
    26, 37, 45, 60, 68, 61, 55, 34, 60, 60, 57, 54, 22, 39, 23, 
    24, 24, 54, 61, 63, 69, 64, 56, 46, 48, 49, 28, 29, 37, 86, 
    
    -- channel=299
    16, 32, 1, 6, 65, 0, 17, 0, 4, 0, 41, 0, 105, 0, 5, 
    15, 29, 23, 6, 67, 0, 0, 0, 12, 0, 39, 0, 90, 0, 31, 
    14, 0, 8, 16, 52, 0, 8, 28, 0, 50, 0, 0, 54, 13, 21, 
    40, 0, 42, 29, 6, 0, 35, 36, 0, 34, 0, 0, 18, 9, 73, 
    44, 0, 66, 38, 0, 8, 81, 0, 12, 0, 16, 0, 17, 7, 111, 
    54, 0, 0, 84, 0, 3, 18, 0, 21, 11, 20, 0, 37, 0, 122, 
    52, 0, 0, 19, 23, 0, 9, 13, 5, 0, 0, 4, 17, 0, 94, 
    30, 0, 0, 3, 3, 43, 0, 0, 7, 18, 22, 0, 51, 0, 91, 
    0, 7, 7, 0, 0, 25, 0, 0, 10, 0, 4, 3, 15, 4, 54, 
    11, 10, 28, 0, 0, 0, 0, 0, 1, 16, 5, 16, 43, 18, 0, 
    57, 0, 43, 0, 13, 20, 0, 10, 10, 15, 0, 10, 28, 0, 3, 
    0, 16, 77, 6, 20, 0, 0, 0, 0, 28, 0, 11, 22, 0, 9, 
    0, 0, 18, 50, 44, 0, 0, 21, 0, 0, 0, 28, 35, 0, 11, 
    44, 0, 0, 0, 58, 31, 10, 30, 0, 0, 0, 32, 56, 0, 0, 
    55, 24, 0, 0, 0, 44, 43, 22, 22, 0, 0, 0, 53, 17, 0, 
    
    -- channel=300
    22, 13, 42, 45, 9, 57, 29, 44, 42, 42, 20, 63, 0, 44, 27, 
    25, 24, 28, 44, 4, 51, 30, 48, 27, 45, 17, 71, 0, 44, 29, 
    40, 39, 32, 35, 6, 42, 41, 39, 45, 23, 41, 64, 2, 38, 30, 
    15, 52, 23, 19, 20, 62, 41, 8, 62, 4, 46, 68, 16, 34, 8, 
    22, 75, 6, 16, 52, 35, 0, 45, 34, 44, 41, 49, 23, 34, 0, 
    8, 79, 37, 0, 55, 20, 0, 40, 29, 25, 10, 60, 19, 44, 0, 
    8, 57, 55, 29, 4, 0, 0, 5, 3, 5, 0, 16, 10, 51, 0, 
    23, 51, 50, 34, 0, 0, 10, 0, 0, 0, 0, 9, 0, 36, 0, 
    30, 45, 37, 38, 32, 0, 5, 0, 0, 0, 0, 11, 0, 23, 5, 
    43, 32, 31, 55, 32, 26, 3, 5, 0, 0, 0, 0, 0, 23, 40, 
    14, 48, 16, 41, 44, 27, 33, 0, 0, 0, 0, 0, 0, 19, 57, 
    16, 25, 2, 48, 27, 37, 28, 0, 0, 0, 1, 0, 0, 38, 47, 
    59, 53, 14, 21, 23, 47, 21, 0, 25, 0, 0, 0, 0, 39, 58, 
    19, 66, 73, 24, 14, 34, 33, 0, 36, 9, 2, 0, 0, 69, 38, 
    9, 22, 75, 72, 22, 19, 27, 34, 17, 15, 17, 0, 0, 22, 78, 
    
    -- channel=301
    0, 24, 0, 0, 47, 0, 4, 0, 0, 0, 28, 0, 75, 0, 2, 
    0, 29, 7, 0, 61, 0, 0, 0, 0, 0, 21, 0, 53, 0, 10, 
    20, 1, 3, 14, 56, 0, 0, 17, 0, 47, 0, 0, 24, 1, 3, 
    23, 0, 25, 25, 12, 0, 23, 40, 0, 29, 0, 0, 1, 0, 44, 
    39, 0, 43, 28, 0, 0, 58, 0, 0, 0, 3, 0, 1, 0, 82, 
    59, 0, 0, 65, 0, 0, 21, 0, 13, 4, 7, 0, 26, 0, 94, 
    49, 0, 0, 12, 23, 0, 8, 0, 7, 0, 0, 1, 11, 0, 76, 
    33, 0, 0, 0, 0, 45, 0, 0, 0, 2, 15, 0, 43, 0, 89, 
    0, 0, 10, 0, 0, 31, 0, 0, 3, 0, 5, 5, 18, 14, 52, 
    7, 17, 35, 0, 0, 0, 3, 0, 0, 7, 10, 10, 32, 10, 0, 
    49, 0, 34, 0, 6, 21, 0, 1, 8, 12, 2, 3, 19, 0, 0, 
    0, 0, 48, 0, 11, 0, 0, 0, 0, 26, 0, 9, 23, 0, 4, 
    0, 0, 11, 34, 30, 0, 0, 27, 0, 0, 0, 27, 28, 0, 9, 
    29, 0, 0, 0, 35, 17, 0, 12, 0, 0, 0, 34, 59, 0, 0, 
    38, 10, 0, 0, 0, 25, 21, 2, 24, 0, 0, 5, 38, 0, 0, 
    
    -- channel=302
    10, 16, 9, 17, 23, 6, 15, 12, 15, 20, 22, 8, 22, 15, 13, 
    13, 12, 21, 14, 21, 10, 19, 8, 18, 13, 22, 3, 24, 3, 13, 
    4, 16, 17, 8, 22, 12, 17, 14, 21, 18, 15, 6, 8, 16, 9, 
    25, 14, 8, 11, 15, 15, 31, 39, 1, 23, 6, 15, 11, 9, 10, 
    19, 1, 21, 7, 5, 22, 33, 9, 22, 15, 18, 31, 13, 5, 20, 
    15, 0, 10, 25, 13, 10, 0, 0, 14, 21, 17, 10, 17, 10, 22, 
    17, 3, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 23, 
    16, 10, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 27, 
    10, 6, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    1, 11, 17, 3, 17, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 
    18, 7, 17, 12, 3, 16, 0, 0, 0, 0, 0, 0, 0, 5, 4, 
    10, 0, 26, 16, 19, 0, 0, 0, 0, 0, 0, 0, 0, 2, 24, 
    0, 4, 22, 28, 27, 3, 0, 0, 0, 0, 0, 0, 0, 11, 23, 
    17, 9, 14, 25, 29, 32, 22, 22, 0, 0, 0, 0, 8, 4, 36, 
    18, 26, 3, 15, 18, 29, 36, 33, 10, 0, 0, 5, 17, 23, 2, 
    
    -- channel=303
    20, 28, 0, 13, 67, 0, 23, 3, 19, 23, 56, 0, 107, 0, 8, 
    20, 21, 29, 12, 70, 0, 23, 0, 36, 6, 59, 0, 103, 0, 32, 
    35, 34, 19, 23, 61, 0, 0, 24, 15, 47, 9, 0, 69, 18, 34, 
    53, 0, 23, 36, 6, 0, 49, 68, 0, 55, 0, 0, 61, 25, 84, 
    45, 0, 77, 31, 0, 23, 82, 0, 22, 3, 34, 16, 38, 28, 124, 
    65, 0, 37, 75, 0, 12, 31, 0, 32, 23, 40, 0, 57, 26, 126, 
    51, 0, 0, 46, 42, 23, 18, 2, 16, 14, 17, 0, 42, 9, 112, 
    46, 0, 0, 37, 33, 22, 1, 14, 31, 5, 0, 2, 43, 17, 104, 
    12, 0, 29, 33, 0, 57, 0, 24, 12, 14, 30, 3, 54, 44, 78, 
    16, 47, 42, 6, 38, 0, 27, 7, 17, 32, 21, 31, 59, 16, 0, 
    77, 0, 47, 2, 1, 40, 0, 25, 30, 33, 25, 26, 32, 12, 8, 
    9, 0, 60, 0, 50, 0, 0, 19, 22, 44, 10, 27, 50, 1, 42, 
    21, 16, 71, 50, 45, 0, 29, 59, 6, 27, 15, 43, 48, 1, 36, 
    56, 0, 1, 45, 64, 37, 31, 48, 0, 12, 22, 43, 89, 0, 28, 
    76, 37, 0, 0, 52, 55, 52, 31, 32, 23, 37, 55, 36, 4, 0, 
    
    -- channel=304
    12, 13, 22, 3, 0, 12, 1, 0, 0, 0, 0, 2, 0, 0, 16, 
    5, 20, 0, 2, 0, 0, 0, 15, 0, 2, 0, 9, 16, 39, 6, 
    0, 0, 0, 0, 0, 35, 40, 0, 0, 0, 0, 9, 4, 10, 8, 
    0, 43, 8, 2, 20, 26, 0, 0, 20, 13, 25, 15, 0, 0, 0, 
    0, 1, 20, 0, 17, 1, 0, 50, 10, 28, 0, 0, 0, 0, 0, 
    0, 0, 0, 48, 31, 0, 0, 7, 5, 0, 0, 21, 0, 0, 0, 
    17, 2, 0, 0, 0, 0, 12, 1, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 8, 0, 18, 0, 0, 0, 0, 30, 11, 0, 13, 0, 0, 
    14, 11, 0, 0, 0, 27, 0, 0, 2, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 11, 13, 
    0, 6, 3, 0, 8, 13, 0, 0, 0, 0, 0, 0, 0, 2, 6, 
    49, 66, 40, 14, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 12, 0, 19, 23, 0, 0, 0, 0, 3, 7, 
    0, 21, 0, 0, 0, 31, 21, 8, 0, 0, 0, 0, 44, 38, 27, 
    
    -- channel=305
    4, 3, 18, 1, 0, 29, 0, 4, 0, 0, 0, 34, 0, 1, 10, 
    3, 8, 0, 1, 0, 1, 0, 19, 0, 2, 0, 44, 0, 45, 0, 
    0, 0, 0, 0, 0, 37, 31, 0, 0, 0, 2, 45, 0, 3, 0, 
    0, 47, 0, 0, 21, 22, 0, 0, 30, 0, 31, 24, 0, 0, 0, 
    0, 33, 0, 0, 27, 0, 0, 52, 0, 20, 0, 0, 0, 0, 0, 
    0, 19, 0, 0, 26, 0, 0, 16, 0, 0, 0, 35, 0, 0, 0, 
    0, 22, 1, 0, 0, 0, 10, 1, 0, 0, 7, 7, 0, 3, 0, 
    0, 14, 10, 0, 12, 0, 3, 1, 1, 23, 8, 12, 0, 0, 0, 
    16, 9, 0, 0, 0, 6, 8, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 5, 21, 
    0, 18, 0, 12, 0, 0, 30, 0, 0, 0, 0, 0, 0, 13, 7, 
    42, 48, 0, 16, 0, 5, 2, 0, 0, 0, 7, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 30, 0, 0, 0, 0, 12, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 23, 44, 
    
    -- channel=306
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 16, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 22, 
    0, 0, 6, 0, 0, 0, 12, 0, 0, 0, 0, 0, 2, 2, 18, 
    0, 0, 0, 9, 7, 9, 6, 2, 9, 12, 15, 1, 6, 0, 18, 
    0, 0, 0, 9, 16, 14, 7, 18, 19, 12, 12, 23, 16, 0, 9, 
    0, 0, 1, 1, 13, 23, 16, 26, 17, 21, 24, 12, 36, 8, 0, 
    0, 0, 0, 0, 0, 18, 21, 23, 30, 30, 21, 22, 20, 0, 0, 
    7, 0, 0, 0, 0, 0, 10, 30, 32, 31, 22, 21, 12, 1, 0, 
    0, 0, 0, 0, 1, 0, 9, 28, 33, 30, 21, 23, 13, 0, 0, 
    0, 7, 4, 0, 0, 0, 16, 28, 19, 28, 30, 27, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 22, 24, 25, 19, 0, 0, 
    2, 0, 0, 0, 6, 0, 0, 0, 0, 17, 22, 17, 0, 0, 0, 
    
    -- channel=307
    35, 20, 47, 39, 20, 20, 41, 24, 43, 27, 37, 28, 50, 10, 26, 
    38, 39, 43, 40, 15, 15, 8, 27, 41, 45, 37, 36, 48, 53, 56, 
    28, 14, 32, 25, 7, 26, 59, 54, 24, 22, 22, 45, 64, 57, 57, 
    22, 44, 44, 25, 10, 67, 60, 0, 34, 21, 55, 68, 52, 55, 48, 
    37, 53, 60, 23, 40, 57, 32, 35, 62, 67, 67, 35, 59, 55, 30, 
    23, 40, 55, 58, 66, 28, 25, 67, 62, 42, 31, 62, 64, 46, 35, 
    35, 47, 40, 56, 31, 23, 22, 31, 13, 21, 24, 40, 36, 63, 35, 
    30, 40, 53, 49, 40, 14, 15, 25, 31, 35, 33, 22, 48, 49, 12, 
    42, 63, 38, 36, 28, 43, 26, 22, 34, 17, 16, 38, 11, 27, 36, 
    57, 28, 31, 37, 33, 0, 36, 40, 25, 40, 20, 29, 21, 27, 34, 
    31, 32, 47, 40, 56, 48, 24, 43, 35, 17, 20, 18, 28, 36, 74, 
    44, 96, 78, 66, 43, 39, 42, 25, 28, 25, 34, 24, 23, 44, 55, 
    34, 18, 68, 85, 67, 50, 39, 15, 0, 26, 26, 21, 23, 16, 62, 
    33, 8, 14, 61, 88, 74, 52, 44, 47, 24, 25, 22, 3, 38, 40, 
    39, 34, 19, 37, 63, 93, 85, 65, 30, 17, 11, 5, 38, 44, 70, 
    
    -- channel=308
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=309
    0, 0, 0, 0, 0, 17, 0, 12, 6, 33, 0, 30, 0, 35, 0, 
    0, 0, 0, 0, 0, 23, 26, 9, 0, 0, 0, 30, 0, 0, 0, 
    21, 40, 6, 4, 0, 0, 0, 0, 32, 0, 31, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 20, 0, 0, 8, 7, 0, 0, 
    0, 32, 0, 0, 8, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 
    0, 52, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 10, 33, 0, 0, 0, 0, 0, 8, 4, 0, 0, 6, 2, 0, 
    0, 20, 1, 9, 0, 0, 16, 0, 0, 0, 0, 16, 0, 14, 0, 
    0, 0, 18, 26, 32, 0, 0, 0, 0, 10, 2, 0, 19, 23, 0, 
    0, 26, 8, 30, 22, 54, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 20, 0, 8, 0, 0, 30, 0, 0, 3, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 4, 11, 6, 0, 0, 0, 0, 18, 13, 
    52, 100, 0, 0, 0, 16, 8, 25, 72, 0, 0, 0, 0, 44, 12, 
    0, 76, 120, 7, 0, 0, 8, 0, 0, 13, 4, 0, 8, 29, 20, 
    0, 0, 60, 93, 10, 0, 0, 0, 8, 37, 44, 30, 0, 0, 4, 
    
    -- channel=310
    14, 3, 10, 9, 12, 0, 17, 2, 26, 12, 24, 0, 49, 0, 0, 
    22, 18, 22, 14, 9, 0, 0, 0, 21, 20, 24, 1, 44, 15, 34, 
    20, 0, 9, 13, 0, 0, 16, 30, 5, 20, 0, 13, 57, 32, 39, 
    10, 0, 31, 8, 0, 26, 41, 0, 0, 8, 21, 30, 47, 40, 50, 
    22, 16, 45, 19, 1, 42, 32, 0, 38, 29, 45, 28, 47, 39, 41, 
    20, 10, 37, 38, 34, 25, 21, 44, 50, 39, 34, 27, 53, 32, 42, 
    20, 17, 26, 51, 42, 27, 21, 30, 18, 24, 24, 36, 37, 39, 39, 
    17, 13, 30, 41, 36, 27, 16, 31, 37, 33, 32, 24, 52, 31, 26, 
    20, 40, 32, 29, 32, 35, 34, 34, 38, 28, 30, 39, 30, 30, 17, 
    40, 25, 19, 15, 21, 17, 33, 40, 40, 47, 30, 37, 26, 9, 6, 
    36, 6, 28, 17, 33, 27, 20, 52, 43, 39, 29, 29, 29, 15, 47, 
    21, 67, 60, 30, 34, 25, 41, 40, 38, 40, 35, 37, 33, 21, 36, 
    33, 19, 63, 66, 42, 29, 45, 38, 6, 33, 43, 33, 32, 0, 40, 
    25, 1, 5, 52, 73, 48, 33, 21, 28, 34, 32, 38, 17, 0, 13, 
    33, 2, 2, 23, 55, 75, 64, 47, 31, 20, 27, 8, 18, 17, 37, 
    
    -- channel=311
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=312
    16, 26, 7, 7, 45, 0, 21, 0, 16, 7, 41, 0, 89, 0, 13, 
    12, 30, 22, 7, 49, 0, 6, 0, 21, 11, 37, 0, 75, 0, 30, 
    24, 11, 13, 14, 43, 0, 10, 29, 0, 45, 0, 0, 52, 18, 21, 
    32, 0, 32, 30, 9, 0, 43, 38, 0, 32, 0, 0, 29, 18, 59, 
    36, 0, 57, 28, 0, 20, 67, 0, 17, 13, 31, 0, 29, 14, 80, 
    49, 0, 3, 65, 5, 15, 28, 5, 35, 27, 31, 0, 46, 1, 91, 
    47, 0, 0, 25, 36, 24, 32, 26, 23, 17, 19, 26, 34, 7, 70, 
    32, 0, 8, 12, 28, 44, 8, 21, 31, 31, 31, 0, 58, 14, 73, 
    7, 10, 14, 5, 0, 48, 10, 20, 32, 23, 27, 26, 22, 23, 54, 
    17, 21, 36, 0, 18, 0, 21, 21, 18, 35, 27, 33, 53, 24, 0, 
    51, 0, 40, 0, 11, 35, 0, 24, 32, 27, 24, 29, 38, 5, 15, 
    0, 25, 71, 11, 27, 0, 5, 18, 19, 37, 17, 33, 42, 14, 15, 
    6, 0, 47, 60, 46, 0, 8, 43, 0, 21, 16, 42, 52, 2, 23, 
    45, 0, 0, 23, 65, 45, 24, 35, 0, 14, 21, 44, 65, 0, 0, 
    48, 33, 0, 0, 24, 57, 56, 35, 35, 4, 15, 24, 45, 10, 0, 
    
    -- channel=313
    24, 4, 23, 32, 12, 16, 21, 23, 38, 36, 30, 36, 24, 23, 18, 
    34, 16, 31, 37, 3, 18, 20, 22, 30, 32, 29, 42, 24, 26, 35, 
    37, 28, 32, 33, 0, 9, 22, 32, 38, 25, 35, 44, 52, 44, 49, 
    20, 32, 33, 18, 0, 40, 42, 7, 34, 9, 42, 50, 63, 54, 49, 
    22, 65, 36, 20, 23, 48, 20, 13, 38, 34, 48, 49, 59, 59, 30, 
    17, 67, 65, 15, 48, 34, 21, 47, 48, 46, 44, 41, 53, 63, 18, 
    12, 50, 66, 60, 37, 23, 14, 33, 33, 29, 24, 40, 49, 61, 21, 
    28, 47, 52, 62, 29, 12, 29, 31, 22, 21, 29, 42, 37, 58, 18, 
    36, 52, 54, 56, 53, 22, 35, 33, 34, 38, 33, 38, 44, 43, 13, 
    53, 45, 32, 50, 40, 55, 32, 41, 44, 42, 33, 35, 22, 25, 40, 
    40, 39, 29, 45, 47, 27, 56, 53, 45, 44, 35, 33, 28, 34, 60, 
    36, 51, 31, 46, 47, 51, 53, 51, 48, 37, 39, 32, 26, 40, 61, 
    63, 75, 58, 47, 37, 56, 50, 37, 44, 39, 46, 27, 21, 31, 60, 
    31, 40, 72, 62, 51, 40, 42, 20, 32, 45, 39, 30, 9, 36, 44, 
    27, 2, 43, 72, 65, 57, 51, 49, 36, 39, 41, 21, 7, 31, 66, 
    
    -- channel=314
    0, 0, 0, 0, 11, 0, 0, 0, 1, 4, 11, 0, 37, 0, 0, 
    0, 0, 0, 0, 5, 0, 6, 0, 0, 0, 13, 0, 21, 0, 0, 
    19, 8, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 15, 0, 0, 
    4, 0, 0, 0, 0, 0, 6, 27, 0, 0, 0, 0, 27, 0, 47, 
    0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 11, 1, 57, 
    10, 0, 1, 0, 0, 0, 0, 0, 0, 1, 11, 0, 19, 1, 39, 
    0, 0, 0, 0, 11, 10, 0, 3, 11, 5, 0, 0, 13, 0, 22, 
    0, 0, 0, 9, 0, 3, 5, 0, 0, 0, 0, 0, 2, 2, 40, 
    0, 0, 11, 13, 18, 0, 0, 9, 5, 18, 11, 3, 45, 27, 0, 
    0, 24, 6, 0, 14, 23, 3, 0, 9, 19, 6, 16, 28, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 17, 13, 28, 19, 15, 8, 0, 0, 
    0, 0, 0, 0, 4, 0, 4, 24, 20, 15, 5, 15, 19, 0, 0, 
    32, 36, 0, 0, 0, 0, 20, 61, 29, 11, 18, 19, 20, 0, 0, 
    16, 25, 34, 0, 0, 0, 0, 0, 0, 22, 8, 26, 54, 0, 0, 
    19, 0, 0, 21, 1, 0, 0, 0, 11, 33, 47, 28, 0, 0, 0, 
    
    -- channel=315
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=316
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 6, 2, 8, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 8, 1, 18, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 15, 
    10, 8, 6, 0, 0, 1, 10, 0, 0, 0, 0, 0, 9, 9, 2, 
    0, 0, 12, 6, 8, 5, 0, 8, 17, 12, 5, 8, 7, 4, 1, 
    4, 0, 6, 14, 0, 19, 6, 11, 0, 0, 17, 13, 11, 13, 12, 
    0, 0, 19, 13, 30, 1, 13, 13, 12, 19, 15, 20, 40, 28, 0, 
    13, 17, 10, 9, 0, 31, 15, 12, 22, 19, 17, 17, 9, 2, 0, 
    15, 0, 0, 0, 9, 0, 12, 24, 20, 30, 20, 14, 12, 3, 0, 
    0, 0, 0, 0, 0, 11, 11, 24, 30, 21, 12, 17, 11, 7, 2, 
    33, 27, 0, 0, 0, 3, 17, 40, 34, 16, 21, 18, 10, 14, 4, 
    1, 30, 16, 0, 0, 0, 0, 0, 0, 22, 17, 27, 21, 4, 0, 
    2, 0, 11, 10, 0, 0, 0, 0, 12, 29, 34, 12, 0, 0, 0, 
    
    -- channel=317
    20, 16, 14, 4, 9, 9, 16, 14, 21, 20, 18, 14, 37, 16, 13, 
    19, 16, 16, 7, 9, 12, 14, 9, 21, 15, 22, 14, 43, 19, 18, 
    8, 15, 10, 9, 8, 14, 18, 14, 13, 13, 21, 18, 42, 17, 20, 
    15, 16, 17, 14, 13, 25, 21, 16, 8, 21, 34, 18, 40, 22, 21, 
    11, 16, 21, 19, 18, 31, 29, 14, 32, 23, 31, 28, 37, 17, 20, 
    14, 15, 19, 17, 28, 37, 44, 37, 35, 40, 45, 25, 32, 18, 27, 
    16, 17, 19, 24, 47, 53, 55, 47, 46, 48, 47, 44, 44, 16, 26, 
    13, 15, 10, 20, 53, 41, 48, 56, 61, 56, 45, 50, 43, 26, 17, 
    20, 17, 17, 19, 28, 38, 52, 55, 51, 53, 58, 44, 45, 28, 14, 
    13, 18, 9, 12, 23, 40, 40, 47, 53, 53, 48, 51, 45, 17, 15, 
    18, 24, 20, 21, 11, 14, 44, 50, 48, 49, 48, 55, 49, 24, 18, 
    26, 50, 43, 17, 24, 18, 43, 58, 47, 46, 52, 56, 53, 31, 14, 
    16, 39, 54, 43, 25, 28, 37, 48, 38, 51, 58, 52, 50, 23, 11, 
    23, 12, 34, 53, 49, 33, 32, 34, 22, 51, 50, 50, 39, 7, 21, 
    25, 17, 21, 36, 54, 45, 41, 35, 34, 39, 42, 39, 26, 28, 35, 
    
    -- channel=318
    0, 18, 0, 0, 0, 16, 0, 21, 0, 6, 0, 46, 0, 0, 17, 
    0, 35, 0, 0, 4, 0, 0, 30, 0, 5, 0, 38, 0, 1, 0, 
    0, 16, 3, 0, 25, 10, 0, 0, 4, 0, 0, 40, 0, 0, 0, 
    0, 0, 0, 1, 54, 0, 0, 15, 1, 24, 0, 26, 0, 0, 0, 
    9, 0, 0, 0, 36, 0, 0, 42, 0, 3, 0, 36, 0, 0, 0, 
    15, 0, 0, 20, 0, 7, 18, 0, 0, 0, 0, 46, 0, 0, 0, 
    22, 0, 3, 0, 0, 0, 12, 0, 0, 0, 16, 8, 0, 0, 0, 
    14, 0, 18, 0, 0, 29, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    12, 0, 3, 0, 0, 22, 0, 0, 0, 0, 0, 6, 0, 0, 11, 
    0, 4, 11, 0, 0, 0, 22, 0, 0, 0, 14, 0, 0, 0, 18, 
    0, 0, 0, 0, 13, 20, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    37, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 41, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 18, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 7, 20, 0, 0, 
    
    -- channel=319
    0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 0, 13, 8, 
    9, 0, 0, 0, 0, 0, 12, 2, 0, 0, 0, 0, 11, 0, 0, 
    0, 2, 4, 0, 8, 13, 0, 0, 11, 0, 8, 0, 0, 0, 0, 
    12, 10, 0, 3, 20, 0, 0, 36, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 19, 0, 1, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 4, 
    7, 3, 0, 0, 0, 7, 10, 0, 0, 9, 0, 0, 0, 0, 18, 
    2, 0, 0, 4, 0, 0, 0, 0, 1, 14, 0, 0, 0, 0, 6, 
    0, 8, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 7, 4, 17, 
    3, 0, 0, 7, 0, 5, 0, 0, 0, 0, 3, 3, 0, 11, 0, 
    22, 0, 0, 0, 0, 7, 0, 0, 3, 0, 0, 0, 0, 0, 6, 
    0, 2, 0, 0, 1, 0, 0, 0, 7, 1, 0, 9, 0, 15, 0, 
    0, 0, 9, 0, 0, 0, 2, 22, 0, 0, 0, 0, 8, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 30, 20, 33, 0, 
    
    -- channel=320
    18, 50, 39, 50, 45, 44, 38, 42, 5, 23, 32, 24, 32, 37, 13, 
    36, 32, 46, 48, 49, 50, 44, 53, 18, 5, 39, 31, 43, 26, 29, 
    6, 49, 47, 49, 49, 48, 43, 54, 46, 21, 48, 26, 37, 36, 34, 
    21, 43, 43, 53, 45, 53, 42, 42, 50, 49, 40, 8, 30, 41, 36, 
    29, 46, 48, 48, 52, 39, 37, 44, 22, 58, 43, 0, 40, 31, 36, 
    96, 34, 51, 39, 36, 53, 0, 5, 23, 50, 17, 0, 36, 31, 39, 
    71, 65, 27, 28, 48, 24, 20, 17, 42, 32, 0, 0, 30, 35, 30, 
    21, 83, 23, 30, 53, 26, 34, 37, 22, 22, 0, 0, 41, 50, 0, 
    32, 79, 27, 2, 42, 47, 0, 28, 25, 1, 0, 3, 54, 62, 0, 
    28, 72, 23, 0, 61, 43, 0, 69, 0, 2, 19, 15, 52, 80, 0, 
    25, 58, 13, 0, 30, 7, 25, 46, 0, 4, 9, 32, 41, 74, 0, 
    34, 45, 32, 26, 12, 42, 43, 4, 0, 3, 1, 18, 50, 37, 37, 
    51, 44, 29, 41, 11, 30, 55, 17, 12, 13, 6, 24, 30, 32, 35, 
    26, 59, 20, 39, 9, 46, 54, 27, 35, 26, 37, 45, 33, 39, 19, 
    46, 52, 39, 47, 41, 44, 38, 38, 35, 39, 51, 50, 36, 28, 44, 
    
    -- channel=321
    23, 50, 38, 42, 40, 45, 40, 35, 31, 19, 22, 29, 25, 31, 23, 
    25, 27, 33, 39, 43, 45, 51, 47, 48, 32, 19, 24, 27, 34, 24, 
    33, 20, 36, 35, 39, 42, 49, 43, 40, 43, 45, 43, 37, 25, 31, 
    3, 24, 31, 34, 37, 41, 45, 40, 36, 35, 39, 46, 29, 34, 30, 
    6, 26, 32, 34, 37, 43, 30, 40, 45, 33, 29, 35, 20, 25, 26, 
    0, 31, 37, 36, 27, 15, 32, 16, 2, 26, 36, 15, 18, 23, 26, 
    37, 0, 24, 25, 16, 31, 0, 27, 40, 33, 28, 19, 16, 26, 29, 
    38, 13, 21, 11, 12, 17, 36, 19, 9, 9, 38, 19, 0, 26, 41, 
    45, 19, 22, 24, 10, 0, 41, 9, 3, 4, 0, 4, 7, 15, 36, 
    44, 23, 9, 45, 0, 9, 14, 32, 60, 11, 17, 37, 12, 9, 39, 
    48, 20, 9, 15, 35, 2, 0, 28, 4, 15, 8, 5, 28, 4, 14, 
    26, 45, 5, 33, 44, 40, 49, 40, 16, 8, 9, 9, 1, 22, 0, 
    42, 35, 37, 0, 34, 32, 34, 47, 34, 28, 27, 18, 29, 10, 31, 
    47, 20, 34, 27, 18, 36, 40, 43, 34, 39, 33, 43, 39, 44, 23, 
    33, 54, 37, 43, 35, 49, 44, 31, 37, 35, 41, 38, 41, 40, 34, 
    
    -- channel=322
    0, 3, 0, 0, 0, 0, 0, 3, 0, 10, 12, 8, 17, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 25, 6, 4, 0, 5, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 2, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 4, 
    1, 7, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 16, 3, 6, 
    78, 0, 13, 0, 0, 25, 0, 0, 0, 17, 0, 0, 26, 8, 13, 
    52, 20, 0, 0, 9, 0, 0, 0, 20, 2, 0, 0, 26, 17, 9, 
    0, 53, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 30, 25, 0, 
    0, 31, 0, 0, 20, 18, 0, 0, 0, 0, 0, 10, 51, 38, 0, 
    0, 44, 0, 0, 70, 0, 0, 13, 0, 1, 12, 1, 37, 56, 0, 
    0, 17, 0, 0, 38, 39, 20, 27, 0, 1, 20, 26, 20, 59, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 15, 30, 24, 40, 47, 21, 17, 
    0, 0, 0, 14, 0, 0, 7, 0, 0, 9, 15, 34, 34, 22, 31, 
    0, 12, 0, 0, 0, 8, 7, 0, 0, 0, 0, 3, 0, 1, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=323
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    9, 0, 0, 0, 1, 0, 3, 2, 7, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 11, 6, 11, 6, 6, 0, 
    17, 0, 0, 0, 7, 0, 0, 41, 25, 0, 5, 19, 6, 4, 1, 
    0, 17, 1, 0, 0, 0, 13, 0, 0, 0, 0, 1, 0, 0, 3, 
    0, 0, 3, 8, 0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 
    0, 0, 0, 14, 17, 15, 18, 44, 43, 61, 66, 17, 0, 0, 0, 
    0, 0, 0, 14, 56, 21, 26, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 5, 17, 11, 0, 50, 43, 34, 52, 16, 25, 10, 0, 10, 0, 
    9, 0, 2, 0, 0, 0, 0, 0, 7, 8, 6, 15, 11, 24, 13, 
    0, 0, 0, 25, 2, 5, 0, 0, 0, 0, 0, 0, 0, 2, 9, 
    4, 12, 8, 4, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=324
    7, 28, 15, 25, 17, 13, 5, 6, 0, 0, 0, 0, 0, 3, 0, 
    24, 18, 19, 21, 25, 24, 17, 19, 0, 0, 0, 0, 9, 0, 0, 
    6, 26, 24, 26, 30, 23, 19, 21, 25, 2, 17, 0, 2, 2, 5, 
    3, 24, 22, 32, 25, 27, 21, 18, 25, 22, 11, 0, 0, 2, 3, 
    10, 24, 28, 25, 29, 31, 26, 34, 3, 25, 22, 0, 2, 1, 4, 
    30, 16, 32, 31, 18, 55, 19, 5, 3, 28, 2, 0, 0, 0, 3, 
    27, 39, 28, 23, 33, 30, 4, 18, 37, 28, 0, 0, 0, 0, 0, 
    0, 49, 23, 23, 51, 35, 32, 42, 28, 28, 0, 0, 0, 24, 0, 
    11, 53, 32, 0, 30, 22, 2, 4, 5, 0, 0, 0, 0, 33, 0, 
    5, 46, 34, 0, 27, 34, 0, 57, 0, 0, 0, 0, 3, 55, 0, 
    12, 31, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 
    11, 22, 19, 12, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 14, 
    23, 21, 6, 23, 14, 12, 21, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 25, 6, 6, 0, 10, 24, 3, 8, 1, 1, 14, 3, 7, 0, 
    15, 27, 15, 25, 20, 19, 13, 13, 7, 3, 18, 23, 13, 4, 14, 
    
    -- channel=325
    16, 42, 1, 9, 2, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 
    1, 0, 0, 3, 6, 9, 8, 7, 4, 0, 0, 0, 6, 2, 0, 
    0, 0, 3, 0, 3, 0, 4, 0, 12, 32, 34, 15, 0, 0, 6, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 2, 0, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 1, 0, 13, 19, 0, 0, 3, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 7, 0, 0, 32, 47, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 12, 16, 4, 0, 6, 11, 0, 0, 28, 4, 
    8, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 
    0, 0, 0, 0, 0, 0, 0, 46, 4, 0, 6, 20, 5, 11, 16, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 2, 0, 32, 28, 44, 38, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 19, 3, 5, 24, 28, 25, 17, 17, 5, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 1, 14, 27, 29, 42, 36, 25, 6, 
    0, 17, 0, 15, 18, 10, 0, 0, 0, 0, 8, 8, 9, 7, 12, 
    
    -- channel=326
    3, 54, 15, 17, 13, 18, 8, 15, 1, 0, 0, 1, 0, 10, 0, 
    20, 16, 13, 19, 20, 18, 20, 20, 11, 1, 0, 0, 4, 7, 0, 
    24, 6, 21, 18, 20, 20, 17, 13, 14, 23, 28, 16, 4, 0, 6, 
    0, 23, 16, 20, 21, 18, 13, 16, 12, 10, 16, 9, 0, 0, 0, 
    9, 13, 20, 20, 16, 24, 5, 16, 18, 1, 9, 5, 0, 0, 0, 
    0, 22, 16, 24, 15, 12, 40, 5, 0, 7, 10, 0, 0, 0, 0, 
    40, 0, 22, 18, 11, 44, 0, 16, 34, 31, 6, 0, 0, 0, 0, 
    12, 14, 17, 10, 29, 21, 37, 25, 22, 20, 17, 0, 0, 12, 12, 
    6, 29, 17, 22, 15, 0, 17, 0, 0, 0, 0, 0, 0, 9, 3, 
    4, 19, 14, 15, 0, 23, 0, 21, 31, 0, 0, 8, 2, 14, 12, 
    13, 13, 9, 0, 15, 0, 0, 0, 0, 0, 0, 0, 10, 14, 0, 
    0, 22, 1, 9, 28, 16, 29, 8, 0, 0, 0, 0, 0, 10, 0, 
    13, 4, 21, 0, 16, 13, 0, 12, 11, 7, 1, 0, 11, 0, 0, 
    8, 0, 4, 14, 0, 1, 14, 4, 2, 18, 10, 28, 20, 27, 3, 
    0, 30, 0, 17, 15, 20, 13, 0, 9, 0, 10, 11, 13, 9, 7, 
    
    -- channel=327
    8, 18, 24, 27, 25, 23, 20, 9, 18, 7, 7, 1, 0, 7, 9, 
    30, 41, 15, 23, 27, 23, 25, 19, 14, 0, 6, 12, 16, 15, 2, 
    41, 31, 23, 27, 27, 28, 25, 19, 24, 2, 4, 8, 16, 14, 10, 
    14, 37, 28, 28, 34, 30, 32, 28, 29, 24, 6, 13, 9, 1, 10, 
    25, 24, 31, 23, 30, 35, 23, 18, 22, 24, 23, 42, 13, 19, 14, 
    0, 13, 19, 34, 33, 15, 41, 55, 40, 18, 27, 14, 15, 13, 11, 
    11, 21, 42, 35, 5, 45, 24, 5, 7, 15, 22, 2, 1, 8, 14, 
    12, 12, 39, 27, 26, 37, 29, 35, 37, 33, 34, 18, 0, 9, 13, 
    17, 13, 30, 31, 59, 2, 49, 49, 46, 54, 45, 0, 0, 13, 25, 
    13, 5, 35, 55, 43, 44, 36, 33, 31, 0, 0, 12, 0, 11, 43, 
    26, 14, 42, 29, 0, 6, 11, 24, 30, 7, 11, 9, 0, 16, 53, 
    15, 18, 20, 4, 12, 0, 6, 22, 0, 0, 2, 2, 0, 14, 32, 
    12, 15, 13, 31, 31, 33, 2, 8, 0, 0, 0, 0, 5, 0, 16, 
    26, 8, 32, 7, 27, 4, 15, 18, 1, 9, 0, 4, 1, 7, 25, 
    3, 14, 12, 12, 7, 21, 23, 24, 18, 4, 14, 15, 14, 18, 0, 
    
    -- channel=328
    33, 5, 15, 11, 20, 12, 12, 0, 11, 0, 0, 0, 0, 0, 5, 
    13, 24, 13, 19, 17, 21, 21, 13, 18, 0, 0, 0, 1, 7, 0, 
    22, 11, 15, 16, 17, 22, 27, 8, 15, 30, 1, 10, 0, 0, 1, 
    24, 11, 16, 12, 22, 23, 24, 15, 6, 21, 17, 14, 0, 0, 0, 
    0, 11, 20, 16, 22, 12, 19, 20, 20, 0, 7, 25, 0, 0, 0, 
    0, 25, 15, 18, 15, 0, 33, 0, 22, 0, 9, 10, 0, 0, 0, 
    0, 0, 28, 26, 7, 8, 27, 37, 11, 15, 25, 0, 0, 0, 0, 
    17, 0, 29, 8, 7, 38, 29, 15, 24, 29, 41, 0, 0, 0, 8, 
    20, 0, 27, 13, 6, 7, 35, 2, 3, 0, 12, 0, 0, 0, 38, 
    27, 0, 24, 51, 0, 0, 45, 13, 36, 0, 0, 0, 0, 0, 66, 
    29, 0, 18, 49, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 58, 
    22, 11, 4, 41, 19, 10, 10, 9, 0, 0, 0, 0, 0, 0, 6, 
    14, 19, 10, 0, 24, 17, 11, 22, 9, 0, 0, 0, 0, 0, 0, 
    18, 0, 27, 0, 15, 13, 6, 31, 10, 13, 14, 7, 14, 0, 5, 
    19, 15, 28, 15, 24, 25, 13, 12, 12, 13, 10, 12, 19, 20, 0, 
    
    -- channel=329
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 0, 1, 9, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=330
    0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 3, 3, 3, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 1, 6, 8, 4, 6, 1, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 6, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 14, 0, 0, 0, 
    0, 0, 0, 0, 5, 3, 5, 6, 11, 14, 10, 8, 4, 0, 0, 
    0, 0, 0, 0, 0, 8, 3, 5, 14, 15, 12, 9, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 7, 7, 5, 10, 6, 2, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 2, 2, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 2, 0, 0, 0, 1, 
    
    -- channel=331
    41, 48, 19, 27, 25, 15, 14, 16, 1, 0, 3, 6, 12, 12, 9, 
    34, 23, 29, 29, 28, 34, 25, 25, 14, 0, 0, 0, 18, 11, 10, 
    9, 27, 31, 27, 32, 26, 28, 19, 33, 52, 41, 21, 5, 6, 18, 
    28, 19, 25, 32, 28, 30, 22, 20, 15, 30, 28, 8, 0, 11, 11, 
    3, 34, 34, 30, 34, 25, 30, 50, 11, 13, 25, 0, 2, 0, 8, 
    23, 31, 44, 32, 11, 62, 37, 0, 7, 24, 2, 0, 0, 0, 6, 
    12, 35, 35, 33, 52, 28, 27, 69, 69, 54, 8, 0, 0, 3, 0, 
    14, 33, 35, 24, 62, 57, 53, 56, 46, 50, 29, 0, 0, 39, 0, 
    33, 52, 50, 9, 18, 33, 12, 0, 0, 0, 0, 0, 1, 35, 6, 
    22, 39, 51, 0, 0, 21, 7, 67, 7, 0, 6, 0, 0, 51, 22, 
    29, 26, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 21, 
    21, 35, 23, 71, 22, 52, 43, 0, 0, 0, 0, 0, 0, 0, 17, 
    37, 33, 23, 9, 37, 13, 38, 33, 26, 14, 0, 5, 0, 0, 0, 
    14, 21, 18, 17, 0, 32, 29, 27, 35, 32, 41, 48, 43, 31, 0, 
    37, 46, 37, 44, 51, 35, 19, 12, 15, 22, 29, 34, 32, 20, 33, 
    
    -- channel=332
    0, 26, 0, 4, 0, 0, 0, 9, 0, 1, 2, 0, 8, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 16, 5, 7, 0, 1, 
    0, 3, 0, 0, 0, 0, 0, 10, 0, 0, 22, 0, 6, 0, 2, 
    0, 2, 0, 7, 0, 0, 0, 0, 6, 0, 0, 0, 0, 17, 5, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 16, 2, 0, 11, 0, 1, 
    73, 0, 15, 0, 0, 21, 0, 0, 0, 15, 0, 0, 18, 2, 10, 
    94, 20, 0, 0, 11, 11, 0, 0, 21, 9, 0, 0, 15, 8, 4, 
    0, 74, 0, 0, 20, 0, 0, 6, 0, 0, 0, 0, 18, 15, 0, 
    0, 54, 0, 0, 7, 8, 0, 0, 0, 0, 0, 0, 52, 38, 0, 
    0, 69, 0, 0, 57, 11, 0, 18, 0, 0, 0, 0, 42, 63, 0, 
    0, 41, 0, 0, 38, 18, 0, 33, 0, 0, 0, 0, 28, 78, 0, 
    0, 15, 0, 0, 0, 7, 15, 0, 0, 1, 0, 21, 31, 41, 0, 
    9, 0, 8, 7, 0, 0, 7, 0, 0, 0, 0, 13, 34, 3, 38, 
    0, 26, 0, 12, 0, 7, 23, 0, 0, 0, 0, 14, 0, 18, 0, 
    0, 20, 0, 10, 0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 15, 
    
    -- channel=333
    27, 37, 45, 52, 50, 50, 48, 42, 20, 23, 33, 29, 30, 35, 22, 
    35, 36, 46, 49, 56, 53, 51, 60, 41, 14, 34, 34, 42, 35, 31, 
    24, 44, 45, 52, 52, 53, 55, 52, 54, 29, 43, 32, 41, 40, 37, 
    16, 37, 46, 52, 47, 58, 54, 48, 54, 55, 44, 30, 40, 42, 39, 
    30, 43, 45, 47, 52, 49, 44, 49, 33, 59, 44, 15, 35, 35, 40, 
    54, 38, 49, 43, 40, 44, 12, 15, 27, 47, 32, 9, 31, 32, 39, 
    37, 47, 31, 36, 36, 27, 24, 31, 34, 23, 12, 10, 22, 32, 34, 
    29, 57, 32, 29, 38, 29, 35, 36, 20, 26, 7, 2, 22, 44, 11, 
    46, 54, 32, 9, 41, 36, 24, 32, 34, 18, 7, 12, 28, 45, 0, 
    50, 55, 25, 0, 44, 31, 25, 67, 20, 16, 18, 21, 32, 53, 0, 
    46, 48, 22, 5, 21, 17, 37, 49, 23, 10, 12, 32, 30, 51, 5, 
    48, 49, 36, 27, 25, 39, 37, 25, 6, 7, 4, 9, 34, 29, 42, 
    56, 55, 32, 40, 17, 38, 58, 34, 18, 13, 7, 14, 23, 26, 29, 
    46, 55, 38, 36, 35, 47, 56, 48, 40, 32, 34, 39, 31, 34, 34, 
    57, 56, 52, 51, 42, 53, 49, 50, 46, 46, 53, 54, 45, 41, 43, 
    
    -- channel=334
    33, 28, 47, 49, 50, 49, 46, 39, 27, 26, 26, 22, 22, 24, 20, 
    46, 50, 50, 49, 53, 53, 51, 51, 38, 22, 28, 28, 28, 27, 26, 
    39, 51, 51, 56, 56, 57, 56, 59, 50, 20, 21, 24, 32, 34, 28, 
    38, 44, 53, 56, 54, 62, 57, 55, 56, 51, 44, 35, 33, 32, 32, 
    40, 45, 51, 55, 59, 59, 48, 42, 39, 57, 50, 34, 34, 33, 33, 
    54, 40, 49, 52, 57, 50, 19, 37, 43, 42, 36, 28, 29, 31, 32, 
    28, 55, 41, 44, 43, 36, 38, 18, 15, 19, 20, 15, 20, 28, 30, 
    23, 46, 39, 42, 40, 35, 37, 35, 26, 27, 14, 13, 21, 25, 16, 
    33, 38, 34, 32, 47, 50, 38, 52, 49, 45, 37, 22, 23, 35, 10, 
    37, 43, 31, 17, 53, 41, 36, 37, 20, 27, 13, 7, 23, 37, 0, 
    35, 42, 34, 18, 15, 40, 45, 52, 45, 21, 22, 25, 20, 43, 15, 
    41, 34, 38, 17, 11, 9, 14, 22, 18, 14, 9, 18, 31, 35, 40, 
    42, 39, 31, 48, 34, 36, 36, 18, 4, 1, 0, 2, 16, 27, 33, 
    38, 46, 35, 37, 36, 32, 37, 33, 25, 13, 14, 13, 13, 19, 24, 
    37, 32, 37, 33, 29, 32, 43, 43, 38, 35, 37, 39, 33, 33, 30, 
    
    -- channel=335
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=336
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 4, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 2, 0, 0, 0, 
    2, 10, 0, 0, 4, 0, 0, 0, 0, 0, 4, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 7, 10, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 0, 7, 4, 9, 34, 21, 0, 0, 8, 
    10, 0, 0, 20, 0, 0, 11, 0, 1, 21, 2, 0, 0, 0, 7, 
    0, 0, 2, 31, 20, 45, 30, 21, 20, 5, 9, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 10, 27, 14, 6, 10, 5, 0, 1, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 12, 
    2, 0, 0, 2, 7, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=337
    9, 11, 35, 33, 37, 42, 38, 35, 17, 23, 24, 20, 19, 21, 13, 
    16, 26, 34, 35, 37, 34, 40, 44, 26, 15, 30, 29, 30, 25, 22, 
    14, 24, 30, 38, 33, 41, 37, 44, 32, 3, 14, 21, 36, 33, 24, 
    15, 29, 33, 33, 37, 46, 44, 40, 43, 42, 34, 18, 33, 28, 29, 
    29, 22, 30, 35, 35, 29, 23, 12, 27, 47, 31, 11, 28, 30, 30, 
    42, 26, 18, 25, 36, 0, 0, 17, 28, 25, 24, 18, 27, 28, 31, 
    25, 31, 15, 15, 8, 9, 20, 0, 0, 0, 5, 6, 18, 23, 29, 
    27, 31, 14, 19, 4, 1, 15, 5, 0, 0, 0, 4, 22, 8, 9, 
    24, 26, 3, 11, 22, 29, 13, 48, 38, 42, 40, 20, 23, 18, 0, 
    34, 25, 0, 0, 45, 27, 27, 14, 21, 21, 5, 9, 28, 15, 0, 
    28, 35, 15, 7, 21, 42, 46, 62, 34, 21, 24, 26, 22, 35, 0, 
    41, 28, 19, 0, 18, 9, 17, 25, 10, 9, 7, 21, 33, 42, 23, 
    36, 37, 25, 30, 0, 33, 30, 11, 2, 0, 0, 1, 17, 26, 29, 
    31, 44, 29, 35, 24, 27, 38, 31, 17, 13, 15, 10, 9, 16, 25, 
    33, 28, 32, 27, 20, 34, 38, 40, 39, 36, 36, 34, 28, 28, 21, 
    
    -- channel=338
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=339
    25, 12, 5, 4, 10, 2, 2, 0, 10, 0, 0, 3, 0, 0, 6, 
    8, 19, 0, 10, 9, 9, 6, 3, 13, 0, 0, 0, 0, 6, 0, 
    24, 13, 6, 4, 6, 8, 14, 0, 3, 28, 8, 4, 0, 0, 0, 
    8, 12, 7, 2, 8, 2, 6, 0, 0, 6, 1, 10, 0, 0, 0, 
    0, 9, 11, 3, 10, 1, 13, 17, 12, 0, 0, 24, 0, 0, 0, 
    0, 19, 14, 9, 3, 0, 43, 0, 15, 0, 6, 6, 0, 0, 0, 
    0, 0, 22, 23, 1, 12, 18, 47, 31, 20, 27, 6, 0, 0, 0, 
    9, 0, 24, 1, 9, 37, 15, 14, 24, 34, 48, 6, 0, 13, 10, 
    8, 0, 25, 1, 19, 0, 28, 0, 0, 0, 8, 0, 0, 0, 42, 
    14, 0, 27, 53, 0, 0, 31, 23, 25, 0, 3, 9, 0, 0, 83, 
    16, 0, 18, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 
    2, 0, 5, 43, 19, 13, 7, 12, 0, 0, 0, 0, 0, 0, 12, 
    0, 5, 0, 0, 15, 11, 5, 19, 14, 9, 8, 2, 0, 0, 0, 
    7, 0, 14, 0, 18, 8, 0, 17, 5, 14, 13, 13, 16, 1, 14, 
    8, 8, 11, 2, 12, 18, 0, 1, 1, 0, 0, 2, 8, 14, 0, 
    
    -- channel=340
    2, 43, 25, 25, 19, 27, 19, 33, 2, 22, 15, 14, 21, 30, 3, 
    26, 13, 32, 26, 25, 26, 24, 27, 2, 22, 24, 20, 19, 11, 19, 
    7, 21, 32, 30, 28, 28, 19, 39, 19, 6, 31, 19, 21, 16, 19, 
    14, 28, 27, 33, 30, 29, 23, 25, 32, 22, 27, 9, 13, 27, 21, 
    24, 28, 27, 33, 29, 23, 15, 16, 21, 33, 28, 0, 23, 18, 17, 
    66, 22, 31, 27, 25, 34, 3, 14, 0, 27, 12, 0, 24, 19, 23, 
    77, 37, 15, 10, 36, 32, 8, 0, 22, 26, 0, 0, 24, 21, 19, 
    13, 61, 9, 25, 36, 11, 28, 20, 14, 5, 0, 0, 29, 19, 9, 
    11, 51, 13, 21, 12, 38, 2, 19, 13, 12, 0, 0, 50, 36, 0, 
    4, 59, 9, 0, 40, 33, 0, 14, 1, 6, 9, 4, 42, 48, 0, 
    7, 47, 7, 0, 41, 29, 9, 35, 0, 9, 13, 6, 35, 65, 0, 
    13, 26, 15, 0, 12, 19, 29, 0, 7, 10, 3, 26, 32, 53, 0, 
    28, 16, 31, 24, 10, 8, 17, 1, 4, 9, 8, 17, 34, 23, 37, 
    11, 38, 3, 37, 0, 21, 33, 0, 16, 13, 14, 23, 16, 31, 0, 
    13, 31, 11, 26, 19, 19, 22, 12, 18, 19, 24, 24, 18, 8, 30, 
    
    -- channel=341
    16, 30, 35, 36, 34, 37, 33, 35, 22, 31, 35, 31, 29, 37, 28, 
    16, 19, 29, 33, 35, 33, 39, 42, 30, 26, 35, 37, 42, 37, 33, 
    16, 18, 27, 29, 30, 31, 32, 36, 36, 26, 40, 41, 45, 38, 37, 
    7, 26, 25, 28, 28, 34, 36, 34, 37, 36, 33, 27, 38, 38, 38, 
    22, 21, 25, 27, 24, 34, 28, 29, 29, 40, 29, 18, 34, 38, 38, 
    21, 26, 19, 25, 21, 16, 16, 22, 20, 37, 30, 16, 34, 33, 38, 
    42, 21, 19, 18, 14, 20, 6, 17, 24, 23, 19, 21, 28, 31, 37, 
    37, 38, 18, 19, 18, 12, 26, 24, 15, 15, 10, 21, 29, 34, 29, 
    41, 44, 17, 14, 18, 11, 16, 27, 21, 22, 13, 18, 30, 33, 10, 
    43, 37, 13, 6, 33, 30, 18, 45, 38, 23, 24, 37, 39, 36, 5, 
    42, 40, 16, 8, 32, 16, 25, 46, 20, 28, 26, 33, 39, 42, 2, 
    42, 44, 23, 12, 42, 41, 48, 41, 16, 18, 23, 27, 31, 38, 21, 
    44, 45, 29, 23, 17, 45, 44, 36, 31, 29, 24, 24, 35, 28, 33, 
    42, 43, 35, 34, 21, 36, 49, 39, 36, 38, 36, 42, 35, 39, 40, 
    41, 49, 40, 45, 38, 47, 43, 43, 43, 41, 46, 45, 40, 37, 38, 
    
    -- channel=342
    12, 13, 0, 0, 3, 3, 0, 5, 2, 0, 2, 13, 21, 3, 0, 
    0, 0, 4, 7, 4, 6, 1, 4, 15, 9, 2, 0, 0, 0, 4, 
    0, 6, 4, 0, 3, 3, 8, 3, 0, 22, 14, 1, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 4, 13, 2, 
    0, 5, 0, 8, 5, 0, 3, 17, 4, 0, 0, 0, 0, 0, 0, 
    12, 19, 24, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 15, 0, 0, 28, 33, 18, 0, 3, 6, 7, 0, 
    6, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 3, 10, 9, 2, 
    9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 6, 7, 
    0, 0, 0, 0, 36, 1, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 4, 0, 27, 0, 11, 3, 0, 15, 6, 0, 0, 6, 0, 0, 
    1, 3, 10, 0, 0, 0, 14, 10, 13, 21, 25, 26, 3, 15, 10, 
    0, 0, 0, 0, 0, 18, 2, 2, 11, 1, 11, 12, 14, 7, 0, 
    16, 9, 3, 1, 7, 4, 0, 0, 0, 6, 2, 2, 2, 2, 7, 
    
    -- channel=343
    11, 9, 21, 18, 25, 29, 28, 21, 10, 0, 0, 0, 0, 0, 0, 
    10, 17, 24, 25, 26, 29, 32, 28, 22, 3, 0, 3, 0, 0, 1, 
    8, 11, 22, 28, 23, 35, 30, 37, 25, 0, 2, 3, 5, 5, 0, 
    8, 14, 22, 24, 29, 36, 33, 29, 25, 26, 23, 12, 3, 4, 2, 
    7, 10, 20, 26, 31, 19, 1, 0, 16, 22, 18, 2, 0, 2, 0, 
    5, 11, 15, 16, 28, 0, 0, 1, 0, 0, 4, 3, 0, 2, 1, 
    1, 4, 3, 0, 3, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 6, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 6, 0, 7, 7, 19, 7, 12, 7, 0, 0, 0, 0, 
    7, 2, 0, 0, 1, 0, 6, 0, 8, 0, 0, 0, 0, 0, 0, 
    4, 7, 0, 0, 0, 14, 4, 20, 8, 0, 0, 0, 0, 0, 0, 
    11, 2, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    9, 7, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    4, 8, 9, 8, 2, 2, 6, 8, 0, 0, 0, 0, 0, 0, 0, 
    7, 1, 7, 5, 0, 8, 15, 10, 11, 10, 9, 8, 7, 6, 0, 
    
    -- channel=344
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 27, 13, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 10, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 27, 77, 28, 19, 6, 24, 41, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 38, 41, 33, 58, 17, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=345
    18, 6, 17, 8, 12, 18, 17, 7, 35, 11, 4, 11, 0, 4, 20, 
    5, 15, 5, 10, 10, 10, 24, 9, 33, 33, 0, 10, 0, 20, 7, 
    45, 0, 8, 7, 7, 16, 19, 13, 8, 17, 0, 27, 18, 7, 8, 
    7, 8, 9, 2, 15, 10, 24, 20, 9, 6, 18, 42, 13, 2, 9, 
    9, 0, 5, 7, 5, 22, 8, 0, 41, 0, 8, 59, 0, 13, 6, 
    0, 16, 0, 14, 23, 0, 43, 41, 9, 0, 36, 45, 0, 9, 1, 
    0, 0, 19, 12, 0, 20, 5, 0, 0, 4, 48, 33, 0, 1, 13, 
    30, 0, 18, 9, 0, 9, 20, 0, 8, 3, 54, 41, 0, 0, 55, 
    20, 0, 8, 49, 0, 0, 59, 18, 7, 44, 58, 13, 0, 0, 69, 
    29, 0, 0, 106, 0, 0, 41, 0, 79, 24, 0, 24, 0, 0, 80, 
    35, 0, 18, 73, 6, 19, 0, 12, 43, 29, 17, 0, 0, 0, 50, 
    17, 12, 0, 0, 43, 0, 11, 52, 27, 10, 16, 7, 0, 14, 0, 
    6, 10, 22, 0, 34, 26, 0, 33, 21, 12, 16, 0, 8, 0, 9, 
    33, 0, 36, 8, 24, 0, 2, 28, 4, 18, 1, 0, 7, 9, 22, 
    0, 9, 12, 8, 5, 19, 25, 17, 21, 11, 5, 3, 19, 26, 0, 
    
    -- channel=346
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=347
    0, 25, 0, 7, 0, 2, 0, 5, 0, 0, 6, 0, 9, 17, 0, 
    0, 0, 0, 6, 9, 5, 0, 7, 0, 0, 17, 7, 14, 0, 2, 
    0, 16, 0, 3, 3, 0, 0, 7, 1, 0, 32, 0, 6, 4, 2, 
    0, 13, 0, 8, 0, 0, 0, 0, 6, 3, 0, 0, 0, 13, 5, 
    0, 12, 1, 0, 5, 0, 0, 6, 0, 16, 0, 0, 12, 2, 5, 
    60, 0, 22, 0, 0, 27, 0, 0, 0, 20, 0, 0, 21, 1, 11, 
    70, 18, 0, 0, 7, 2, 0, 0, 39, 10, 0, 0, 13, 10, 5, 
    0, 68, 0, 0, 20, 0, 0, 15, 0, 0, 0, 0, 18, 35, 0, 
    0, 52, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 39, 46, 0, 
    0, 57, 0, 0, 79, 0, 0, 54, 0, 0, 0, 3, 37, 74, 0, 
    0, 27, 0, 0, 8, 0, 0, 21, 0, 0, 0, 16, 19, 69, 0, 
    0, 7, 7, 0, 0, 19, 20, 0, 0, 0, 0, 8, 31, 10, 17, 
    3, 8, 0, 18, 0, 0, 18, 0, 0, 0, 0, 21, 25, 0, 23, 
    0, 19, 0, 0, 0, 15, 27, 0, 5, 0, 9, 28, 6, 16, 4, 
    13, 18, 0, 11, 0, 13, 0, 0, 0, 0, 13, 16, 0, 0, 12, 
    
    -- channel=348
    28, 0, 7, 14, 19, 4, 16, 0, 7, 0, 7, 0, 0, 0, 10, 
    7, 25, 5, 11, 15, 13, 10, 15, 18, 0, 0, 0, 11, 5, 0, 
    4, 26, 2, 11, 12, 11, 16, 0, 27, 19, 0, 0, 0, 10, 3, 
    10, 7, 11, 10, 8, 13, 12, 7, 6, 21, 0, 0, 9, 0, 0, 
    7, 9, 13, 3, 14, 8, 16, 15, 0, 6, 3, 20, 7, 4, 8, 
    4, 0, 3, 5, 3, 17, 1, 0, 45, 8, 0, 6, 0, 2, 1, 
    0, 21, 12, 20, 0, 0, 27, 40, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 18, 2, 8, 23, 0, 16, 10, 26, 14, 0, 0, 20, 0, 
    10, 0, 12, 0, 34, 0, 0, 8, 22, 0, 36, 10, 0, 5, 12, 
    12, 0, 18, 10, 19, 0, 37, 51, 0, 0, 1, 1, 0, 6, 42, 
    8, 0, 12, 52, 0, 0, 17, 0, 34, 0, 0, 28, 0, 0, 67, 
    15, 0, 19, 27, 0, 10, 0, 3, 0, 0, 0, 0, 1, 0, 63, 
    1, 15, 0, 20, 3, 20, 19, 10, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 29, 5, 0, 20, 8, 3, 12, 5, 5, 0, 27, 
    22, 0, 16, 0, 9, 6, 0, 19, 4, 3, 7, 9, 3, 11, 0, 
    
    -- channel=349
    56, 15, 28, 21, 31, 27, 30, 12, 39, 10, 12, 21, 12, 3, 31, 
    17, 32, 23, 25, 26, 29, 38, 27, 49, 23, 0, 10, 10, 27, 15, 
    45, 8, 22, 21, 22, 31, 41, 17, 30, 53, 14, 34, 16, 13, 18, 
    28, 14, 22, 14, 25, 27, 34, 27, 15, 27, 30, 48, 22, 7, 14, 
    13, 9, 22, 19, 23, 25, 29, 26, 43, 3, 12, 63, 2, 13, 14, 
    0, 34, 11, 24, 26, 0, 52, 11, 32, 2, 31, 47, 0, 12, 7, 
    0, 0, 27, 30, 3, 10, 27, 48, 13, 16, 57, 38, 1, 9, 13, 
    34, 0, 31, 10, 0, 35, 32, 3, 16, 25, 71, 37, 0, 5, 47, 
    34, 0, 25, 33, 0, 0, 55, 0, 0, 9, 48, 18, 0, 0, 83, 
    45, 0, 15, 105, 0, 0, 63, 2, 70, 23, 20, 27, 0, 0, 111, 
    44, 0, 15, 102, 0, 0, 6, 0, 39, 18, 1, 2, 0, 0, 81, 
    32, 14, 3, 52, 52, 25, 22, 46, 22, 5, 10, 0, 0, 0, 0, 
    19, 22, 15, 0, 46, 36, 16, 51, 39, 26, 26, 5, 0, 6, 0, 
    32, 0, 41, 6, 37, 18, 6, 48, 23, 34, 28, 18, 32, 15, 29, 
    23, 17, 35, 20, 30, 32, 23, 26, 26, 24, 18, 17, 31, 39, 9, 
    
    -- channel=350
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=351
    18, 0, 0, 0, 0, 0, 0, 0, 9, 0, 4, 6, 4, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 1, 0, 6, 5, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 3, 0, 2, 1, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 2, 
    0, 0, 0, 0, 0, 0, 4, 3, 3, 0, 0, 18, 0, 0, 1, 
    0, 5, 0, 0, 0, 0, 17, 2, 10, 0, 8, 26, 0, 0, 0, 
    0, 0, 3, 3, 0, 0, 11, 24, 6, 5, 26, 22, 0, 0, 0, 
    8, 0, 8, 1, 0, 11, 0, 1, 11, 15, 30, 18, 0, 0, 16, 
    8, 0, 10, 7, 0, 0, 13, 0, 0, 3, 31, 15, 0, 0, 38, 
    16, 0, 12, 41, 0, 0, 28, 0, 19, 15, 14, 10, 0, 0, 56, 
    11, 0, 11, 56, 0, 0, 7, 0, 26, 10, 4, 6, 0, 0, 49, 
    11, 0, 8, 18, 12, 2, 0, 18, 15, 8, 11, 0, 0, 0, 11, 
    0, 8, 0, 0, 5, 4, 5, 19, 15, 13, 14, 4, 0, 4, 0, 
    7, 0, 13, 0, 15, 0, 0, 15, 7, 8, 6, 0, 5, 0, 12, 
    10, 0, 11, 0, 7, 3, 0, 5, 2, 5, 0, 0, 4, 8, 0, 
    
    -- channel=352
    0, 10, 0, 3, 0, 0, 0, 8, 0, 8, 7, 0, 5, 20, 0, 
    0, 0, 1, 0, 1, 0, 0, 3, 0, 0, 26, 11, 15, 0, 2, 
    0, 14, 1, 4, 2, 0, 0, 9, 0, 0, 16, 0, 5, 7, 2, 
    0, 11, 1, 12, 0, 0, 0, 0, 13, 0, 0, 0, 0, 15, 7, 
    10, 14, 0, 2, 2, 0, 0, 0, 0, 30, 2, 0, 21, 7, 9, 
    119, 0, 10, 0, 0, 35, 0, 0, 0, 28, 0, 0, 28, 6, 18, 
    89, 51, 0, 0, 15, 1, 0, 0, 7, 0, 0, 0, 18, 10, 7, 
    0, 96, 0, 5, 32, 0, 0, 11, 0, 0, 0, 0, 36, 25, 0, 
    0, 71, 0, 0, 27, 35, 0, 8, 11, 0, 0, 0, 64, 56, 0, 
    0, 79, 0, 0, 115, 28, 0, 37, 0, 0, 0, 0, 56, 89, 0, 
    0, 51, 0, 0, 22, 28, 19, 43, 0, 0, 7, 21, 26, 107, 0, 
    0, 5, 15, 0, 0, 0, 3, 0, 0, 0, 0, 25, 54, 44, 18, 
    10, 3, 0, 38, 0, 0, 15, 0, 0, 0, 0, 10, 32, 15, 28, 
    0, 43, 0, 12, 0, 7, 30, 0, 0, 0, 0, 5, 0, 6, 0, 
    5, 14, 0, 5, 0, 0, 0, 0, 0, 0, 10, 12, 0, 0, 14, 
    
    -- channel=353
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=354
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=355
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 17, 
    0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=356
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 18, 30, 55, 19, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 8, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 31, 34, 5, 38, 10, 14, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 5, 6, 4, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=357
    12, 9, 27, 33, 28, 26, 23, 17, 7, 4, 9, 3, 1, 13, 10, 
    33, 30, 27, 28, 32, 30, 29, 29, 13, 0, 8, 15, 20, 17, 11, 
    27, 27, 30, 35, 36, 33, 32, 32, 32, 3, 7, 14, 23, 22, 18, 
    21, 25, 32, 36, 38, 41, 42, 35, 38, 34, 23, 18, 15, 17, 21, 
    23, 29, 33, 33, 36, 44, 37, 34, 26, 42, 38, 20, 15, 19, 20, 
    19, 22, 33, 39, 33, 37, 26, 40, 28, 30, 31, 7, 7, 12, 18, 
    12, 42, 39, 35, 27, 38, 27, 15, 12, 20, 16, 0, 0, 6, 15, 
    13, 35, 40, 34, 39, 37, 37, 45, 36, 32, 19, 3, 0, 10, 6, 
    33, 37, 41, 30, 44, 37, 46, 46, 45, 43, 21, 0, 0, 24, 7, 
    33, 40, 43, 19, 33, 46, 34, 37, 20, 3, 0, 0, 0, 30, 6, 
    42, 42, 39, 4, 0, 9, 21, 42, 30, 2, 0, 2, 4, 36, 19, 
    40, 40, 29, 12, 2, 2, 7, 7, 0, 0, 0, 0, 3, 22, 29, 
    41, 42, 30, 36, 31, 31, 32, 15, 0, 0, 0, 0, 0, 0, 19, 
    41, 44, 39, 28, 23, 20, 36, 33, 18, 10, 1, 4, 0, 8, 12, 
    33, 38, 38, 36, 27, 34, 39, 40, 31, 29, 31, 33, 30, 23, 21, 
    
    -- channel=358
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=359
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=360
    37, 11, 12, 2, 10, 6, 11, 8, 15, 11, 6, 7, 7, 0, 13, 
    5, 13, 13, 7, 7, 10, 12, 6, 18, 14, 1, 5, 2, 5, 9, 
    10, 5, 8, 7, 6, 9, 9, 5, 17, 27, 10, 12, 0, 4, 4, 
    20, 7, 7, 5, 5, 6, 5, 7, 2, 8, 12, 13, 6, 0, 1, 
    10, 1, 6, 6, 6, 8, 6, 3, 4, 0, 2, 19, 4, 4, 2, 
    0, 9, 0, 7, 9, 13, 11, 0, 14, 0, 0, 19, 3, 6, 0, 
    0, 0, 5, 6, 10, 0, 15, 21, 7, 5, 15, 16, 6, 6, 2, 
    7, 0, 4, 9, 0, 14, 10, 0, 6, 9, 15, 17, 11, 9, 14, 
    4, 0, 4, 7, 0, 0, 0, 0, 0, 0, 13, 13, 0, 0, 20, 
    2, 0, 0, 11, 0, 0, 16, 1, 9, 12, 15, 11, 1, 0, 27, 
    0, 0, 0, 38, 0, 0, 0, 0, 12, 11, 4, 11, 1, 0, 23, 
    5, 0, 4, 22, 28, 16, 9, 10, 11, 12, 14, 2, 0, 0, 7, 
    0, 0, 0, 4, 18, 7, 0, 15, 23, 22, 20, 18, 1, 8, 0, 
    0, 0, 2, 0, 7, 0, 0, 3, 9, 12, 18, 13, 19, 7, 15, 
    1, 0, 0, 0, 8, 0, 0, 1, 0, 1, 0, 1, 4, 7, 4, 
    
    -- channel=361
    19, 45, 1, 9, 5, 1, 0, 0, 0, 0, 0, 1, 1, 3, 0, 
    0, 0, 0, 5, 7, 12, 10, 8, 7, 0, 0, 0, 5, 1, 0, 
    0, 0, 3, 0, 3, 0, 7, 0, 14, 37, 36, 13, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 1, 3, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 3, 0, 13, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 4, 0, 0, 34, 53, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 13, 16, 4, 0, 5, 18, 0, 0, 28, 6, 
    11, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 
    0, 0, 0, 0, 0, 0, 0, 43, 8, 0, 6, 23, 0, 9, 28, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 5, 
    0, 2, 0, 44, 29, 46, 39, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 20, 0, 7, 28, 30, 27, 21, 20, 3, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 2, 15, 27, 31, 45, 38, 28, 2, 
    0, 17, 1, 14, 17, 14, 0, 0, 0, 0, 8, 7, 9, 7, 11, 
    
    -- channel=362
    57, 96, 79, 83, 80, 82, 73, 70, 49, 41, 42, 43, 40, 54, 38, 
    82, 79, 79, 86, 88, 88, 88, 86, 65, 40, 41, 46, 56, 54, 45, 
    73, 73, 87, 87, 90, 91, 87, 89, 82, 64, 73, 61, 58, 51, 55, 
    52, 81, 83, 91, 91, 94, 87, 85, 82, 80, 77, 59, 47, 54, 54, 
    60, 77, 86, 89, 91, 93, 69, 75, 72, 77, 77, 51, 48, 52, 52, 
    43, 76, 86, 88, 83, 76, 70, 60, 47, 66, 62, 21, 42, 47, 51, 
    84, 68, 80, 75, 73, 87, 56, 56, 71, 71, 44, 23, 35, 47, 48, 
    57, 79, 73, 69, 84, 77, 90, 80, 69, 65, 51, 28, 32, 58, 46, 
    64, 86, 73, 67, 73, 59, 72, 64, 58, 51, 10, 9, 39, 64, 33, 
    61, 81, 66, 42, 41, 76, 41, 79, 67, 21, 20, 38, 46, 72, 33, 
    70, 74, 61, 10, 43, 18, 21, 59, 20, 25, 19, 23, 51, 71, 33, 
    58, 77, 56, 57, 61, 56, 69, 45, 9, 6, 8, 17, 28, 57, 41, 
    76, 69, 70, 61, 67, 64, 58, 55, 40, 30, 21, 23, 43, 27, 53, 
    66, 62, 63, 66, 43, 58, 74, 61, 55, 56, 53, 66, 59, 67, 46, 
    58, 84, 63, 74, 68, 77, 75, 62, 65, 57, 70, 72, 69, 62, 61, 
    
    -- channel=363
    44, 9, 7, 0, 8, 7, 9, 0, 33, 0, 0, 13, 3, 0, 21, 
    1, 13, 4, 5, 1, 7, 17, 1, 36, 26, 0, 0, 0, 12, 1, 
    35, 0, 4, 0, 0, 8, 18, 0, 5, 49, 0, 24, 0, 0, 1, 
    21, 0, 1, 0, 4, 0, 7, 6, 0, 0, 16, 41, 4, 0, 0, 
    0, 0, 1, 1, 0, 4, 6, 6, 32, 0, 0, 55, 0, 0, 0, 
    0, 21, 0, 5, 7, 0, 48, 0, 9, 0, 17, 43, 0, 0, 0, 
    0, 0, 11, 12, 0, 2, 9, 37, 6, 14, 52, 36, 0, 0, 0, 
    26, 0, 13, 0, 0, 16, 19, 0, 4, 9, 70, 37, 0, 0, 48, 
    13, 0, 8, 32, 0, 0, 42, 0, 0, 0, 32, 13, 0, 0, 88, 
    24, 0, 0, 111, 0, 0, 40, 0, 69, 16, 13, 22, 0, 0, 116, 
    22, 0, 1, 92, 2, 0, 0, 0, 16, 16, 0, 0, 0, 0, 70, 
    3, 0, 0, 44, 45, 10, 11, 37, 27, 5, 8, 0, 0, 0, 0, 
    0, 0, 10, 0, 38, 14, 0, 39, 38, 30, 33, 7, 0, 0, 0, 
    12, 0, 19, 0, 13, 0, 0, 25, 7, 21, 16, 6, 24, 7, 7, 
    0, 0, 8, 0, 12, 8, 1, 0, 5, 3, 0, 0, 12, 20, 0, 
    
    -- channel=364
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 5, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 24, 7, 0, 
    0, 9, 0, 0, 30, 4, 0, 0, 0, 0, 0, 0, 14, 16, 0, 
    0, 0, 0, 0, 20, 14, 0, 0, 0, 0, 8, 0, 2, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 24, 11, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=365
    37, 0, 5, 0, 3, 3, 9, 0, 30, 3, 0, 9, 0, 0, 23, 
    10, 11, 8, 0, 0, 2, 15, 0, 28, 26, 0, 0, 0, 9, 2, 
    29, 0, 6, 0, 0, 5, 13, 0, 3, 36, 0, 22, 0, 0, 1, 
    31, 0, 1, 0, 4, 6, 9, 12, 0, 0, 15, 38, 0, 0, 0, 
    2, 0, 0, 2, 0, 6, 5, 0, 29, 0, 4, 53, 0, 0, 0, 
    0, 11, 0, 3, 12, 0, 31, 2, 19, 0, 18, 45, 0, 0, 0, 
    0, 0, 5, 9, 0, 0, 21, 20, 0, 0, 48, 37, 0, 0, 0, 
    19, 0, 12, 0, 0, 9, 20, 0, 0, 0, 60, 41, 0, 0, 40, 
    11, 0, 3, 47, 0, 0, 46, 0, 0, 14, 46, 19, 0, 0, 82, 
    18, 0, 0, 109, 0, 0, 46, 0, 54, 24, 11, 8, 0, 0, 87, 
    19, 0, 1, 82, 0, 0, 0, 0, 37, 26, 1, 0, 0, 0, 49, 
    10, 0, 0, 32, 29, 2, 0, 25, 29, 5, 5, 0, 0, 0, 0, 
    1, 0, 15, 0, 47, 13, 0, 30, 29, 15, 18, 0, 0, 4, 0, 
    10, 0, 21, 10, 16, 0, 0, 25, 3, 14, 7, 0, 12, 0, 0, 
    0, 0, 10, 0, 11, 0, 4, 0, 6, 8, 0, 0, 10, 14, 0, 
    
    -- channel=366
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=367
    52, 0, 21, 12, 24, 13, 20, 0, 34, 9, 6, 7, 0, 0, 27, 
    23, 43, 17, 16, 14, 18, 23, 9, 31, 9, 0, 4, 1, 15, 5, 
    46, 16, 16, 18, 17, 23, 28, 8, 19, 28, 0, 13, 3, 10, 5, 
    49, 16, 22, 12, 22, 23, 27, 25, 12, 20, 16, 32, 13, 0, 3, 
    26, 9, 22, 15, 22, 23, 30, 12, 29, 1, 15, 70, 2, 10, 8, 
    0, 22, 0, 21, 36, 0, 44, 29, 67, 0, 25, 59, 0, 9, 0, 
    0, 3, 33, 36, 4, 1, 50, 35, 0, 0, 53, 35, 0, 0, 5, 
    17, 0, 38, 21, 0, 40, 22, 3, 25, 32, 63, 41, 0, 0, 29, 
    14, 0, 25, 39, 11, 9, 54, 27, 30, 43, 94, 31, 0, 0, 80, 
    27, 0, 26, 107, 0, 11, 82, 0, 41, 29, 11, 6, 0, 0, 106, 
    25, 0, 32, 114, 0, 0, 29, 0, 74, 25, 13, 11, 0, 0, 100, 
    28, 0, 14, 35, 21, 0, 0, 33, 20, 5, 13, 0, 0, 0, 26, 
    2, 8, 0, 16, 49, 35, 0, 21, 15, 2, 0, 0, 0, 6, 0, 
    17, 0, 37, 0, 44, 0, 0, 32, 3, 7, 5, 0, 5, 0, 24, 
    5, 0, 20, 0, 13, 5, 10, 22, 14, 11, 0, 0, 12, 24, 0, 
    
    -- channel=368
    10, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 26, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 10, 0, 0, 35, 51, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 0, 0, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 13, 10, 0, 1, 10, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 42, 6, 35, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 15, 25, 29, 28, 29, 1, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 10, 13, 23, 32, 30, 19, 0, 
    0, 10, 0, 1, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    
    -- channel=369
    0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 30, 2, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 9, 0, 0, 22, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 13, 0, 0, 19, 44, 18, 0, 0, 6, 1, 0, 
    0, 30, 0, 0, 14, 0, 0, 5, 0, 0, 0, 0, 6, 25, 0, 
    0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 21, 0, 
    0, 34, 0, 0, 0, 0, 0, 31, 0, 0, 10, 5, 20, 38, 0, 
    0, 8, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 17, 23, 0, 
    0, 6, 0, 14, 0, 35, 23, 0, 0, 0, 0, 0, 7, 0, 0, 
    6, 0, 0, 0, 0, 0, 14, 4, 14, 20, 18, 27, 13, 1, 0, 
    0, 1, 0, 0, 0, 9, 10, 0, 14, 12, 18, 31, 20, 19, 0, 
    7, 19, 0, 11, 10, 2, 0, 0, 0, 0, 5, 6, 0, 0, 18, 
    
    -- channel=370
    18, 0, 16, 14, 14, 10, 10, 2, 10, 3, 6, 3, 2, 4, 13, 
    15, 18, 11, 15, 15, 14, 13, 10, 9, 1, 1, 11, 12, 13, 10, 
    22, 12, 12, 15, 17, 16, 17, 13, 13, 7, 1, 12, 13, 15, 11, 
    22, 14, 16, 15, 19, 17, 24, 16, 16, 19, 14, 13, 11, 7, 13, 
    14, 13, 16, 14, 17, 19, 25, 19, 18, 17, 18, 22, 5, 12, 13, 
    0, 18, 15, 19, 18, 13, 28, 30, 25, 15, 20, 19, 1, 5, 9, 
    0, 17, 29, 24, 13, 15, 27, 22, 9, 14, 24, 10, 0, 0, 9, 
    15, 4, 30, 24, 16, 34, 22, 27, 30, 30, 28, 11, 0, 4, 14, 
    23, 10, 31, 21, 18, 24, 36, 24, 25, 27, 32, 2, 0, 5, 24, 
    28, 8, 36, 30, 14, 20, 43, 21, 24, 11, 3, 0, 0, 3, 35, 
    31, 14, 31, 35, 0, 4, 17, 15, 31, 0, 0, 4, 0, 2, 41, 
    34, 19, 23, 17, 12, 4, 6, 14, 0, 0, 0, 0, 0, 1, 23, 
    22, 30, 14, 27, 24, 23, 21, 16, 2, 0, 0, 0, 0, 1, 3, 
    28, 23, 33, 10, 24, 12, 20, 26, 15, 11, 5, 1, 4, 0, 17, 
    25, 19, 30, 21, 21, 24, 23, 28, 19, 21, 16, 20, 21, 19, 10, 
    
    -- channel=371
    2, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 10, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 4, 6, 0, 3, 0, 0, 0, 0, 20, 13, 3, 0, 0, 0, 
    2, 11, 2, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 7, 5, 0, 9, 0, 10, 1, 0, 0, 7, 0, 0, 0, 
    0, 7, 7, 11, 0, 22, 42, 5, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 20, 16, 11, 35, 0, 28, 36, 35, 7, 0, 0, 0, 0, 
    2, 0, 16, 6, 31, 23, 24, 28, 29, 27, 27, 2, 0, 10, 5, 
    0, 14, 20, 15, 22, 0, 10, 0, 0, 0, 0, 0, 0, 9, 15, 
    0, 3, 26, 21, 0, 18, 0, 14, 15, 0, 0, 4, 0, 14, 35, 
    0, 0, 14, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 5, 0, 19, 9, 7, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 21, 4, 0, 1, 9, 8, 4, 3, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 17, 13, 13, 0, 
    0, 7, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=372
    2, 0, 10, 9, 11, 14, 16, 11, 11, 13, 16, 14, 15, 10, 14, 
    0, 0, 8, 8, 8, 9, 14, 16, 15, 14, 18, 19, 13, 15, 16, 
    0, 0, 3, 7, 4, 10, 12, 16, 8, 0, 0, 13, 21, 20, 12, 
    2, 0, 4, 2, 4, 12, 16, 13, 13, 14, 12, 14, 23, 19, 17, 
    4, 0, 0, 3, 5, 2, 6, 0, 13, 19, 8, 8, 14, 16, 16, 
    12, 3, 0, 0, 6, 0, 0, 1, 11, 5, 12, 24, 13, 16, 17, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 7, 15, 12, 13, 18, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 11, 
    16, 0, 0, 0, 0, 4, 4, 16, 10, 17, 35, 26, 9, 0, 6, 
    24, 0, 0, 9, 9, 0, 21, 0, 13, 24, 15, 10, 10, 0, 0, 
    17, 7, 0, 25, 12, 35, 39, 36, 37, 21, 22, 21, 9, 0, 0, 
    26, 10, 0, 0, 7, 3, 4, 20, 23, 18, 14, 18, 22, 18, 5, 
    17, 18, 8, 4, 0, 14, 20, 12, 5, 4, 7, 4, 7, 23, 14, 
    20, 23, 17, 13, 15, 14, 16, 22, 11, 7, 7, 0, 1, 2, 13, 
    22, 9, 21, 11, 7, 14, 19, 24, 21, 25, 17, 14, 14, 16, 10, 
    
    -- channel=373
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 7, 1, 0, 
    71, 0, 0, 0, 0, 2, 0, 22, 9, 1, 0, 3, 11, 1, 3, 
    2, 37, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 7, 0, 0, 33, 40, 0, 48, 47, 52, 49, 20, 17, 13, 0, 
    0, 26, 0, 0, 101, 15, 0, 0, 0, 14, 0, 0, 10, 23, 0, 
    0, 24, 16, 0, 0, 76, 56, 61, 40, 6, 25, 18, 0, 50, 0, 
    1, 0, 17, 0, 0, 0, 0, 0, 5, 12, 4, 22, 35, 29, 37, 
    0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 25, 
    0, 25, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=374
    22, 30, 17, 16, 16, 15, 8, 7, 7, 0, 0, 0, 0, 0, 1, 
    28, 30, 16, 20, 19, 19, 18, 12, 6, 0, 0, 0, 3, 6, 0, 
    35, 18, 23, 21, 22, 23, 20, 11, 16, 19, 11, 9, 2, 0, 4, 
    20, 30, 23, 21, 29, 22, 22, 16, 15, 17, 13, 10, 0, 0, 0, 
    18, 20, 27, 23, 24, 22, 17, 19, 22, 4, 13, 23, 0, 1, 0, 
    0, 25, 20, 31, 25, 17, 54, 28, 16, 7, 15, 0, 0, 0, 0, 
    6, 10, 42, 33, 17, 49, 25, 23, 26, 33, 23, 0, 0, 0, 0, 
    11, 3, 38, 26, 34, 48, 44, 37, 45, 41, 39, 5, 0, 5, 14, 
    12, 13, 37, 34, 31, 9, 43, 18, 15, 18, 1, 0, 0, 4, 24, 
    10, 3, 39, 42, 0, 33, 24, 20, 36, 0, 0, 0, 0, 4, 46, 
    22, 8, 32, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 40, 
    9, 16, 13, 27, 23, 5, 14, 5, 0, 0, 0, 0, 0, 0, 2, 
    11, 11, 19, 10, 34, 18, 0, 13, 3, 0, 0, 0, 0, 0, 0, 
    13, 0, 22, 8, 9, 4, 10, 13, 3, 14, 6, 12, 12, 11, 7, 
    1, 18, 11, 15, 17, 21, 12, 7, 9, 0, 7, 10, 14, 12, 2, 
    
    -- channel=375
    3, 0, 20, 21, 23, 28, 24, 17, 11, 10, 11, 11, 10, 8, 6, 
    5, 12, 20, 19, 21, 24, 29, 27, 21, 15, 14, 14, 9, 12, 11, 
    9, 9, 17, 22, 19, 26, 28, 33, 19, 0, 1, 12, 22, 16, 10, 
    4, 8, 17, 17, 21, 28, 31, 27, 27, 22, 20, 21, 19, 19, 16, 
    4, 7, 14, 19, 22, 20, 16, 9, 26, 30, 19, 15, 15, 14, 14, 
    7, 9, 12, 14, 23, 0, 0, 7, 9, 9, 20, 19, 12, 16, 15, 
    6, 2, 0, 3, 0, 0, 0, 0, 0, 0, 5, 6, 7, 13, 17, 
    14, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 3, 0, 0, 13, 
    16, 0, 0, 7, 0, 2, 17, 21, 10, 19, 23, 13, 4, 0, 4, 
    23, 1, 0, 15, 2, 0, 15, 0, 21, 13, 4, 6, 4, 0, 0, 
    19, 8, 0, 9, 14, 31, 29, 43, 29, 16, 15, 8, 9, 0, 0, 
    20, 14, 0, 0, 2, 0, 3, 16, 15, 8, 3, 14, 14, 22, 0, 
    21, 16, 14, 1, 5, 15, 16, 8, 0, 0, 0, 0, 7, 14, 22, 
    24, 21, 16, 15, 9, 14, 16, 21, 6, 1, 0, 0, 0, 5, 2, 
    16, 13, 18, 12, 4, 17, 24, 23, 22, 23, 19, 16, 16, 17, 9, 
    
    -- channel=376
    61, 39, 44, 40, 47, 46, 48, 33, 50, 21, 19, 31, 18, 14, 36, 
    44, 53, 44, 42, 45, 47, 57, 46, 65, 38, 7, 16, 17, 35, 22, 
    63, 26, 46, 44, 45, 52, 60, 40, 49, 64, 21, 43, 23, 22, 28, 
    44, 30, 44, 39, 48, 52, 52, 54, 37, 42, 48, 62, 29, 18, 23, 
    31, 29, 43, 45, 45, 54, 43, 40, 57, 23, 39, 76, 13, 23, 22, 
    0, 48, 30, 47, 52, 14, 59, 23, 44, 16, 46, 52, 5, 24, 16, 
    0, 3, 42, 48, 28, 35, 39, 52, 16, 27, 60, 43, 8, 19, 21, 
    41, 0, 45, 28, 16, 42, 53, 20, 26, 32, 73, 45, 0, 10, 51, 
    40, 0, 35, 58, 13, 10, 67, 22, 22, 32, 51, 24, 0, 0, 84, 
    49, 0, 26, 113, 0, 19, 60, 7, 75, 33, 19, 29, 0, 0, 98, 
    50, 0, 29, 85, 14, 0, 12, 0, 45, 33, 10, 1, 11, 0, 70, 
    34, 29, 16, 51, 51, 26, 26, 50, 33, 11, 14, 0, 0, 5, 4, 
    34, 27, 37, 5, 63, 44, 18, 51, 42, 28, 25, 7, 3, 16, 0, 
    42, 4, 46, 32, 44, 22, 13, 53, 29, 37, 30, 23, 36, 26, 28, 
    23, 28, 38, 28, 38, 33, 37, 31, 37, 30, 27, 26, 40, 45, 22, 
    
    -- channel=377
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 6, 1, 0, 12, 21, 26, 0, 0, 0, 0, 0, 0, 0, 
    17, 15, 21, 11, 4, 35, 20, 1, 15, 17, 0, 0, 0, 0, 0, 
    0, 23, 20, 17, 29, 25, 7, 35, 40, 33, 7, 0, 0, 0, 0, 
    0, 19, 22, 9, 44, 23, 13, 24, 25, 25, 6, 0, 0, 18, 0, 
    0, 23, 36, 0, 39, 25, 3, 9, 0, 0, 0, 0, 0, 28, 6, 
    0, 16, 37, 0, 0, 11, 0, 8, 0, 0, 0, 0, 0, 32, 25, 
    0, 4, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 24, 
    0, 0, 9, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 1, 1, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=378
    0, 0, 12, 3, 12, 10, 9, 0, 15, 2, 3, 0, 0, 0, 4, 
    3, 21, 4, 8, 9, 3, 7, 3, 10, 0, 3, 5, 2, 8, 0, 
    25, 12, 4, 12, 9, 14, 13, 6, 3, 0, 0, 0, 11, 11, 0, 
    20, 15, 14, 7, 15, 18, 22, 14, 14, 15, 6, 9, 12, 0, 6, 
    17, 4, 10, 13, 12, 18, 14, 0, 14, 18, 10, 33, 4, 11, 9, 
    0, 15, 0, 13, 26, 0, 9, 36, 39, 4, 22, 36, 3, 7, 7, 
    0, 13, 24, 21, 0, 12, 30, 0, 0, 0, 22, 8, 0, 0, 10, 
    13, 0, 25, 18, 0, 9, 1, 10, 16, 15, 14, 10, 0, 0, 5, 
    6, 0, 11, 20, 39, 25, 37, 58, 51, 66, 86, 20, 0, 0, 21, 
    24, 0, 16, 56, 34, 22, 52, 0, 27, 20, 0, 0, 0, 0, 31, 
    19, 6, 39, 59, 0, 47, 44, 50, 58, 11, 17, 8, 0, 0, 48, 
    27, 7, 18, 0, 0, 0, 0, 27, 6, 0, 0, 3, 0, 11, 34, 
    2, 21, 10, 26, 0, 22, 0, 0, 0, 0, 0, 0, 0, 1, 16, 
    26, 14, 29, 8, 29, 1, 6, 20, 0, 0, 0, 0, 0, 0, 16, 
    10, 0, 13, 0, 0, 9, 18, 24, 16, 10, 2, 4, 4, 11, 0, 
    
    -- channel=379
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=380
    0, 0, 0, 0, 0, 0, 0, 2, 9, 5, 3, 0, 1, 5, 8, 
    5, 1, 0, 0, 0, 0, 0, 0, 0, 6, 5, 9, 5, 6, 6, 
    8, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 11, 9, 4, 
    16, 2, 2, 0, 6, 1, 6, 2, 3, 1, 2, 4, 4, 5, 9, 
    8, 2, 1, 3, 0, 2, 2, 0, 7, 8, 9, 10, 4, 8, 7, 
    3, 2, 0, 3, 5, 0, 9, 35, 11, 2, 14, 18, 2, 4, 7, 
    5, 13, 14, 7, 0, 17, 19, 0, 0, 3, 13, 8, 1, 0, 8, 
    10, 8, 16, 16, 5, 7, 5, 18, 21, 12, 11, 13, 1, 0, 9, 
    9, 6, 13, 23, 20, 25, 27, 39, 34, 45, 39, 12, 1, 4, 12, 
    11, 13, 22, 24, 24, 22, 24, 0, 16, 16, 0, 0, 0, 1, 8, 
    16, 22, 32, 14, 6, 38, 23, 36, 28, 11, 15, 0, 0, 16, 16, 
    19, 16, 14, 0, 0, 0, 0, 9, 8, 3, 0, 7, 4, 24, 13, 
    9, 15, 21, 16, 6, 7, 3, 0, 0, 0, 0, 0, 0, 5, 25, 
    20, 20, 20, 18, 11, 3, 11, 10, 2, 0, 0, 0, 0, 0, 3, 
    9, 7, 12, 8, 3, 8, 16, 15, 11, 12, 4, 4, 6, 3, 2, 
    
    -- channel=381
    83, 76, 87, 87, 92, 90, 90, 76, 63, 45, 51, 49, 48, 51, 49, 
    77, 86, 87, 92, 98, 97, 98, 96, 86, 44, 46, 56, 62, 61, 55, 
    77, 80, 87, 95, 95, 102, 100, 94, 100, 73, 71, 64, 62, 64, 60, 
    63, 81, 89, 93, 96, 103, 101, 92, 91, 96, 85, 69, 61, 58, 60, 
    67, 77, 89, 91, 99, 94, 77, 77, 74, 84, 80, 66, 53, 59, 60, 
    45, 79, 85, 89, 89, 76, 60, 59, 61, 66, 65, 48, 46, 54, 57, 
    42, 70, 80, 77, 72, 71, 72, 64, 58, 54, 55, 38, 35, 52, 53, 
    62, 64, 76, 73, 68, 81, 84, 74, 64, 66, 56, 35, 35, 60, 49, 
    78, 66, 72, 60, 62, 64, 75, 68, 65, 56, 49, 30, 29, 56, 44, 
    79, 66, 61, 52, 55, 58, 74, 87, 72, 41, 33, 42, 40, 61, 49, 
    80, 67, 59, 63, 21, 28, 44, 57, 56, 30, 24, 42, 42, 57, 61, 
    80, 71, 66, 67, 73, 64, 64, 57, 22, 18, 16, 12, 35, 45, 67, 
    78, 84, 62, 74, 64, 67, 71, 71, 47, 33, 26, 26, 33, 36, 42, 
    71, 69, 79, 59, 68, 66, 75, 80, 66, 63, 63, 65, 62, 59, 66, 
    80, 76, 80, 78, 72, 84, 79, 79, 74, 70, 76, 80, 77, 74, 64, 
    
    -- channel=382
    18, 0, 0, 0, 0, 0, 0, 7, 0, 9, 0, 1, 7, 0, 7, 
    12, 0, 18, 0, 0, 0, 0, 0, 0, 14, 0, 1, 0, 0, 9, 
    0, 0, 8, 0, 0, 0, 0, 10, 1, 8, 0, 9, 0, 0, 3, 
    32, 0, 0, 2, 0, 5, 0, 8, 0, 0, 12, 0, 0, 4, 0, 
    9, 0, 0, 4, 0, 0, 3, 0, 0, 1, 17, 0, 4, 0, 0, 
    64, 0, 0, 0, 1, 13, 0, 0, 1, 0, 0, 1, 0, 2, 0, 
    0, 26, 0, 0, 33, 0, 10, 0, 0, 0, 0, 9, 4, 0, 0, 
    0, 3, 0, 4, 6, 0, 13, 0, 0, 0, 0, 6, 22, 0, 0, 
    0, 4, 0, 21, 0, 33, 0, 0, 0, 0, 0, 5, 29, 0, 0, 
    0, 5, 0, 0, 0, 4, 0, 0, 0, 15, 18, 0, 13, 0, 0, 
    0, 13, 0, 0, 3, 0, 2, 0, 1, 17, 0, 0, 13, 0, 0, 
    9, 0, 0, 13, 0, 12, 1, 0, 13, 5, 0, 0, 16, 16, 0, 
    14, 0, 6, 0, 29, 0, 3, 0, 6, 4, 0, 0, 0, 31, 0, 
    0, 19, 0, 28, 0, 0, 0, 0, 7, 0, 6, 0, 5, 3, 0, 
    0, 0, 4, 4, 14, 0, 0, 0, 0, 11, 0, 0, 1, 0, 20, 
    
    -- channel=383
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 11, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 4, 1, 2, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 7, 3, 0, 
    0, 0, 0, 4, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 
    28, 20, 4, 0, 5, 7, 0, 0, 0, 2, 0, 20, 0, 0, 0, 
    0, 4, 0, 0, 12, 0, 5, 13, 0, 0, 1, 7, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 11, 18, 2, 0, 0, 
    13, 0, 0, 0, 0, 0, 3, 0, 0, 18, 9, 0, 0, 0, 0, 
    0, 0, 0, 22, 14, 23, 21, 8, 9, 2, 0, 4, 0, 0, 0, 
    6, 0, 7, 0, 0, 0, 0, 3, 21, 9, 2, 6, 15, 0, 9, 
    0, 7, 0, 0, 0, 0, 10, 0, 0, 3, 3, 5, 0, 26, 1, 
    0, 4, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    
    -- channel=384
    120, 104, 115, 105, 95, 89, 94, 76, 75, 52, 55, 49, 0, 39, 52, 
    103, 88, 87, 86, 82, 75, 80, 68, 67, 64, 67, 9, 0, 65, 58, 
    67, 65, 74, 71, 72, 70, 73, 70, 68, 72, 23, 0, 29, 65, 48, 
    66, 72, 71, 69, 76, 76, 81, 75, 70, 55, 0, 34, 60, 57, 56, 
    72, 74, 73, 71, 79, 72, 65, 71, 79, 22, 0, 28, 50, 54, 56, 
    74, 73, 70, 69, 75, 76, 41, 14, 0, 0, 31, 0, 30, 42, 50, 
    73, 71, 63, 71, 47, 9, 0, 0, 0, 75, 27, 0, 0, 16, 40, 
    72, 68, 68, 31, 1, 25, 0, 49, 59, 40, 0, 0, 0, 18, 57, 
    69, 73, 0, 4, 0, 7, 50, 49, 0, 0, 0, 0, 47, 45, 22, 
    82, 89, 0, 7, 0, 16, 73, 2, 0, 0, 8, 0, 5, 0, 0, 
    81, 0, 0, 0, 0, 40, 61, 0, 0, 0, 0, 46, 0, 0, 0, 
    42, 0, 0, 0, 18, 21, 61, 0, 0, 8, 0, 38, 7, 0, 11, 
    34, 5, 4, 0, 42, 17, 24, 0, 0, 28, 0, 0, 18, 0, 21, 
    33, 6, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 12, 
    30, 1, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 4, 6, 13, 
    
    -- channel=385
    117, 112, 109, 108, 105, 99, 94, 91, 87, 53, 63, 59, 42, 4, 56, 
    104, 104, 102, 101, 94, 87, 85, 81, 77, 71, 60, 64, 12, 31, 67, 
    76, 73, 79, 84, 79, 79, 81, 77, 76, 71, 57, 0, 31, 56, 69, 
    70, 77, 78, 78, 80, 81, 81, 83, 79, 72, 22, 0, 45, 63, 66, 
    75, 81, 80, 80, 78, 78, 58, 57, 58, 85, 26, 21, 56, 65, 65, 
    80, 82, 80, 78, 68, 49, 47, 22, 0, 0, 0, 51, 0, 44, 61, 
    82, 81, 82, 64, 64, 5, 0, 0, 0, 0, 0, 13, 31, 1, 30, 
    79, 80, 55, 63, 13, 4, 0, 0, 39, 46, 0, 0, 0, 0, 22, 
    80, 61, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 31, 5, 
    62, 57, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 
    55, 0, 0, 7, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    53, 0, 0, 3, 0, 1, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 4, 0, 0, 2, 0, 17, 10, 0, 0, 7, 
    39, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 7, 
    33, 13, 0, 19, 2, 3, 6, 6, 7, 0, 0, 0, 7, 6, 3, 
    
    -- channel=386
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 1, 28, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 8, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 6, 0, 0, 0, 6, 0, 47, 0, 0, 
    0, 0, 0, 0, 4, 5, 13, 15, 38, 107, 56, 0, 2, 37, 7, 
    0, 0, 7, 0, 0, 23, 8, 61, 68, 36, 0, 0, 0, 37, 52, 
    0, 5, 3, 33, 0, 47, 77, 41, 0, 0, 0, 0, 47, 33, 14, 
    5, 48, 0, 35, 0, 44, 90, 24, 0, 0, 7, 0, 0, 0, 0, 
    19, 9, 0, 5, 15, 71, 92, 12, 0, 0, 50, 103, 0, 0, 0, 
    13, 19, 30, 0, 47, 60, 78, 0, 0, 35, 16, 74, 29, 0, 21, 
    18, 28, 43, 0, 76, 37, 53, 6, 0, 53, 0, 18, 64, 0, 35, 
    12, 20, 14, 0, 35, 28, 23, 16, 0, 56, 12, 2, 48, 23, 35, 
    9, 14, 41, 21, 32, 34, 30, 28, 28, 53, 4, 7, 32, 33, 40, 
    
    -- channel=387
    0, 0, 11, 20, 19, 18, 17, 15, 13, 24, 6, 0, 19, 24, 0, 
    13, 7, 15, 18, 17, 14, 11, 9, 4, 0, 0, 0, 2, 0, 0, 
    32, 30, 18, 11, 5, 0, 0, 0, 0, 0, 2, 18, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 13, 0, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 16, 67, 76, 0, 0, 35, 0, 0, 
    0, 0, 0, 0, 0, 40, 46, 56, 31, 0, 0, 0, 0, 31, 13, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 45, 8, 0, 0, 
    0, 0, 0, 25, 22, 19, 0, 0, 11, 10, 0, 8, 0, 0, 0, 
    0, 0, 0, 1, 16, 13, 0, 0, 4, 66, 80, 0, 0, 0, 24, 
    4, 75, 24, 1, 11, 0, 0, 0, 35, 62, 40, 69, 29, 43, 67, 
    2, 2, 0, 0, 0, 0, 0, 0, 15, 0, 0, 22, 16, 22, 5, 
    3, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 37, 40, 7, 
    0, 7, 40, 57, 73, 112, 124, 128, 87, 5, 11, 5, 25, 20, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 32, 15, 0, 0, 0, 
    
    -- channel=388
    43, 38, 44, 38, 32, 27, 29, 18, 17, 0, 0, 1, 0, 0, 0, 
    43, 37, 27, 25, 22, 17, 17, 12, 9, 3, 16, 0, 0, 0, 0, 
    19, 6, 11, 11, 11, 10, 9, 10, 9, 13, 24, 0, 0, 6, 0, 
    1, 6, 8, 7, 11, 13, 20, 20, 20, 19, 0, 0, 0, 0, 0, 
    6, 8, 9, 8, 15, 25, 27, 28, 44, 22, 0, 0, 6, 0, 0, 
    8, 10, 9, 8, 20, 47, 76, 70, 47, 23, 67, 0, 0, 0, 0, 
    11, 9, 5, 14, 33, 0, 0, 0, 0, 24, 68, 0, 0, 0, 0, 
    10, 9, 33, 25, 0, 1, 0, 19, 67, 97, 46, 0, 0, 0, 30, 
    8, 25, 0, 0, 0, 0, 21, 98, 51, 40, 3, 0, 10, 45, 47, 
    26, 102, 0, 0, 0, 0, 49, 40, 30, 0, 34, 49, 58, 23, 0, 
    41, 5, 0, 0, 0, 3, 50, 31, 0, 0, 0, 28, 0, 0, 0, 
    5, 0, 0, 0, 0, 10, 56, 35, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 3, 0, 30, 32, 49, 19, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=389
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 8, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 15, 1, 14, 20, 5, 
    0, 0, 0, 2, 3, 3, 9, 13, 13, 12, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 2, 12, 7, 7, 26, 39, 29, 30, 5, 0, 0, 
    1, 1, 0, 0, 4, 26, 76, 65, 3, 0, 77, 17, 0, 9, 0, 
    1, 0, 0, 3, 17, 0, 0, 0, 0, 0, 16, 48, 10, 0, 0, 
    0, 0, 20, 28, 0, 4, 6, 60, 120, 120, 5, 0, 3, 10, 55, 
    0, 11, 0, 0, 0, 0, 0, 67, 0, 0, 0, 0, 23, 79, 44, 
    12, 79, 24, 0, 0, 0, 8, 0, 0, 0, 0, 74, 75, 12, 0, 
    3, 0, 0, 0, 0, 27, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 16, 15, 5, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 50, 61, 25, 0, 0, 16, 23, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 2, 5, 33, 21, 21, 14, 6, 2, 0, 0, 0, 3, 5, 8, 
    
    -- channel=390
    46, 27, 18, 12, 6, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 
    1, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 16, 0, 0, 11, 4, 
    0, 0, 0, 0, 0, 0, 0, 8, 8, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 5, 0, 4, 25, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 33, 43, 29, 0, 18, 42, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 39, 0, 21, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 43, 120, 34, 1, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 67, 42, 5, 27, 0, 0, 35, 41, 
    0, 30, 22, 0, 0, 0, 7, 20, 5, 22, 0, 11, 62, 23, 12, 
    2, 0, 0, 0, 0, 0, 35, 16, 23, 0, 0, 0, 1, 0, 0, 
    2, 0, 0, 0, 0, 19, 5, 27, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 10, 30, 55, 6, 0, 0, 1, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=391
    25, 31, 42, 39, 39, 31, 32, 27, 19, 22, 13, 6, 27, 2, 4, 
    27, 28, 31, 23, 22, 18, 19, 15, 12, 10, 0, 13, 0, 0, 4, 
    33, 20, 12, 12, 8, 5, 6, 7, 7, 2, 31, 16, 0, 6, 15, 
    2, 1, 3, 3, 3, 3, 2, 5, 7, 9, 27, 0, 1, 8, 7, 
    1, 1, 2, 4, 2, 16, 23, 3, 0, 0, 0, 0, 15, 11, 6, 
    0, 1, 3, 5, 0, 0, 33, 81, 102, 80, 28, 8, 2, 20, 5, 
    1, 2, 8, 0, 20, 32, 20, 0, 0, 0, 37, 30, 0, 21, 9, 
    1, 2, 0, 12, 14, 0, 6, 0, 0, 3, 30, 93, 12, 0, 0, 
    3, 0, 2, 4, 34, 0, 0, 53, 59, 36, 49, 0, 0, 0, 30, 
    0, 0, 28, 0, 1, 0, 0, 39, 25, 85, 62, 20, 20, 25, 48, 
    0, 72, 33, 12, 0, 0, 0, 28, 82, 0, 0, 16, 45, 51, 36, 
    0, 0, 31, 9, 0, 6, 0, 32, 66, 0, 0, 0, 16, 42, 0, 
    0, 0, 23, 0, 0, 0, 2, 11, 41, 0, 0, 0, 35, 13, 0, 
    0, 10, 44, 22, 36, 47, 51, 50, 39, 1, 3, 0, 8, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 28, 0, 0, 0, 0, 
    
    -- channel=392
    45, 40, 37, 35, 35, 27, 23, 23, 7, 16, 6, 0, 0, 0, 5, 
    29, 33, 34, 26, 20, 17, 16, 14, 10, 10, 1, 0, 0, 0, 11, 
    11, 17, 16, 15, 11, 15, 16, 13, 12, 8, 0, 0, 0, 4, 13, 
    10, 12, 15, 16, 15, 18, 20, 22, 16, 0, 0, 0, 13, 12, 9, 
    14, 16, 16, 16, 14, 10, 11, 14, 22, 31, 9, 0, 8, 6, 4, 
    16, 17, 17, 14, 2, 0, 0, 0, 0, 0, 37, 53, 0, 23, 4, 
    16, 18, 17, 4, 0, 0, 0, 0, 0, 0, 0, 119, 0, 0, 0, 
    17, 17, 0, 0, 1, 0, 0, 11, 8, 0, 33, 68, 30, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 22, 34, 60, 75, 0, 0, 8, 
    0, 0, 53, 0, 0, 0, 0, 6, 21, 11, 0, 67, 9, 17, 17, 
    0, 0, 43, 0, 0, 0, 0, 14, 40, 14, 0, 0, 26, 16, 19, 
    0, 0, 0, 7, 0, 0, 0, 22, 91, 0, 0, 0, 0, 39, 0, 
    0, 0, 0, 10, 0, 8, 0, 20, 84, 0, 14, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=393
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 39, 35, 10, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 4, 11, 0, 15, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 31, 22, 22, 8, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 6, 27, 22, 21, 40, 62, 0, 0, 1, 17, 
    0, 25, 19, 0, 0, 0, 2, 16, 32, 2, 17, 76, 25, 30, 0, 
    0, 0, 15, 0, 0, 9, 31, 12, 0, 0, 0, 13, 36, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 11, 0, 0, 0, 0, 44, 0, 0, 
    0, 3, 27, 28, 46, 64, 71, 70, 35, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 0, 0, 0, 0, 
    
    -- channel=394
    54, 57, 58, 63, 64, 63, 59, 60, 60, 43, 50, 40, 21, 17, 42, 
    61, 59, 62, 71, 69, 65, 61, 59, 57, 54, 36, 34, 22, 18, 48, 
    51, 58, 64, 66, 62, 60, 58, 55, 52, 47, 16, 0, 12, 22, 44, 
    58, 61, 59, 60, 59, 58, 53, 46, 41, 33, 14, 7, 32, 43, 52, 
    57, 63, 63, 62, 57, 46, 25, 23, 1, 0, 0, 0, 24, 49, 49, 
    61, 63, 61, 60, 47, 10, 0, 0, 0, 0, 0, 0, 0, 15, 47, 
    62, 62, 61, 49, 24, 0, 0, 0, 5, 0, 0, 0, 0, 0, 26, 
    61, 59, 33, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 41, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    32, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 14, 12, 
    19, 4, 0, 0, 0, 0, 0, 1, 6, 0, 0, 9, 13, 11, 5, 
    
    -- channel=395
    47, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 12, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 9, 3, 
    0, 0, 0, 0, 0, 4, 4, 5, 7, 12, 8, 0, 7, 17, 1, 
    0, 4, 7, 7, 10, 14, 24, 26, 23, 16, 0, 0, 9, 0, 0, 
    7, 8, 8, 8, 13, 19, 14, 26, 71, 68, 32, 6, 0, 0, 0, 
    11, 11, 8, 5, 15, 63, 82, 47, 0, 0, 132, 0, 0, 7, 0, 
    11, 10, 4, 10, 22, 0, 0, 0, 0, 51, 76, 81, 0, 0, 0, 
    10, 10, 31, 26, 0, 11, 5, 107, 164, 149, 94, 0, 14, 0, 73, 
    9, 25, 0, 0, 0, 0, 39, 110, 68, 78, 49, 1, 54, 107, 68, 
    27, 130, 14, 0, 0, 0, 49, 57, 74, 0, 20, 134, 94, 56, 7, 
    29, 0, 13, 0, 0, 33, 70, 65, 0, 0, 0, 0, 27, 0, 0, 
    0, 12, 20, 0, 5, 11, 82, 77, 0, 0, 0, 0, 39, 0, 0, 
    0, 2, 14, 16, 71, 99, 78, 69, 7, 19, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=396
    19, 3, 9, 2, 0, 0, 6, 0, 9, 0, 0, 0, 0, 8, 0, 
    4, 0, 0, 0, 0, 0, 6, 0, 4, 2, 9, 0, 0, 33, 0, 
    0, 0, 0, 1, 7, 6, 8, 7, 7, 9, 22, 0, 0, 24, 0, 
    7, 11, 9, 6, 11, 9, 10, 9, 10, 12, 0, 25, 10, 2, 0, 
    11, 11, 9, 7, 13, 15, 6, 4, 12, 0, 0, 15, 0, 0, 3, 
    10, 9, 7, 6, 17, 32, 35, 1, 0, 0, 0, 0, 25, 0, 3, 
    11, 8, 1, 10, 38, 3, 0, 0, 0, 94, 59, 0, 1, 3, 0, 
    9, 4, 19, 9, 0, 16, 0, 8, 61, 95, 0, 0, 0, 17, 31, 
    7, 17, 7, 5, 0, 15, 70, 69, 0, 0, 0, 0, 20, 60, 18, 
    21, 83, 0, 20, 0, 37, 108, 12, 0, 0, 0, 0, 16, 0, 0, 
    80, 4, 0, 0, 0, 40, 127, 0, 0, 0, 41, 81, 0, 0, 0, 
    33, 8, 0, 0, 17, 58, 88, 0, 0, 5, 0, 94, 0, 0, 0, 
    25, 12, 5, 0, 58, 19, 67, 0, 0, 31, 0, 19, 43, 0, 14, 
    16, 21, 0, 0, 27, 0, 0, 0, 0, 39, 0, 0, 15, 0, 11, 
    6, 0, 0, 0, 2, 3, 1, 0, 0, 44, 0, 0, 3, 6, 15, 
    
    -- channel=397
    131, 126, 135, 131, 127, 118, 117, 106, 102, 72, 77, 68, 20, 33, 62, 
    130, 118, 116, 119, 113, 102, 102, 94, 89, 81, 79, 40, 9, 44, 72, 
    93, 96, 100, 98, 95, 92, 93, 88, 86, 85, 43, 6, 28, 61, 69, 
    86, 90, 90, 88, 93, 94, 96, 91, 84, 72, 1, 15, 61, 72, 76, 
    87, 93, 92, 91, 95, 88, 76, 83, 82, 47, 0, 13, 59, 72, 73, 
    92, 93, 91, 89, 92, 74, 36, 7, 0, 0, 11, 0, 17, 45, 66, 
    94, 92, 88, 88, 58, 20, 0, 0, 11, 25, 12, 0, 0, 21, 42, 
    92, 91, 78, 42, 6, 15, 1, 22, 24, 9, 0, 0, 0, 9, 35, 
    92, 88, 18, 7, 0, 0, 6, 18, 0, 0, 0, 0, 42, 16, 7, 
    97, 70, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 0, 0, 0, 0, 14, 6, 0, 0, 0, 0, 25, 0, 0, 0, 
    65, 0, 0, 0, 3, 3, 9, 0, 0, 4, 0, 2, 0, 0, 5, 
    47, 3, 1, 0, 11, 0, 1, 0, 0, 9, 0, 0, 10, 0, 13, 
    41, 11, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 4, 
    36, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=398
    97, 111, 123, 128, 123, 113, 110, 101, 91, 74, 65, 57, 29, 33, 41, 
    121, 108, 105, 105, 97, 87, 84, 80, 72, 62, 62, 34, 8, 20, 46, 
    90, 86, 84, 77, 73, 66, 66, 65, 62, 61, 41, 18, 13, 33, 50, 
    62, 61, 61, 61, 62, 63, 61, 61, 60, 57, 17, 11, 33, 54, 55, 
    54, 60, 61, 61, 63, 63, 62, 59, 50, 21, 0, 7, 45, 52, 54, 
    58, 60, 61, 61, 62, 45, 22, 16, 27, 23, 0, 0, 32, 30, 47, 
    62, 60, 59, 59, 43, 30, 19, 13, 18, 11, 0, 0, 0, 25, 35, 
    61, 61, 55, 27, 15, 11, 0, 0, 0, 0, 0, 0, 0, 2, 3, 
    59, 57, 23, 16, 0, 12, 7, 0, 0, 0, 0, 0, 1, 0, 0, 
    60, 26, 0, 0, 0, 2, 6, 0, 0, 0, 19, 0, 0, 0, 0, 
    52, 20, 0, 0, 0, 0, 0, 0, 0, 5, 9, 28, 0, 0, 5, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 5, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 10, 
    20, 2, 0, 0, 7, 19, 24, 24, 10, 3, 0, 0, 6, 4, 3, 
    19, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 1, 
    
    -- channel=399
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 23, 55, 37, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 13, 5, 2, 37, 33, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 44, 54, 10, 0, 0, 
    0, 0, 0, 18, 22, 8, 11, 27, 44, 51, 40, 11, 0, 0, 19, 
    0, 0, 22, 12, 10, 3, 15, 47, 49, 47, 69, 34, 20, 33, 23, 
    0, 44, 51, 11, 3, 6, 6, 48, 43, 36, 3, 53, 54, 40, 33, 
    0, 6, 41, 15, 4, 18, 29, 47, 52, 7, 8, 4, 45, 35, 0, 
    0, 15, 41, 18, 12, 23, 22, 44, 42, 16, 10, 0, 32, 27, 0, 
    0, 4, 31, 29, 31, 45, 50, 51, 53, 12, 25, 4, 8, 5, 0, 
    0, 0, 12, 6, 10, 9, 5, 3, 0, 5, 19, 6, 0, 0, 0, 
    
    -- channel=400
    0, 0, 0, 5, 9, 9, 7, 8, 7, 22, 9, 2, 4, 8, 0, 
    10, 3, 8, 11, 9, 7, 6, 6, 3, 0, 6, 2, 8, 0, 0, 
    6, 20, 12, 6, 5, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 8, 0, 3, 4, 
    0, 0, 0, 0, 0, 0, 0, 4, 15, 13, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 13, 4, 0, 0, 
    0, 0, 0, 3, 0, 10, 51, 66, 44, 10, 0, 13, 2, 9, 4, 
    0, 0, 0, 0, 14, 0, 2, 12, 0, 0, 0, 0, 1, 0, 0, 
    0, 4, 16, 13, 7, 21, 0, 0, 0, 0, 18, 66, 5, 0, 0, 
    3, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 2, 14, 0, 0, 0, 10, 71, 43, 2, 0, 6, 47, 
    0, 8, 0, 10, 0, 0, 0, 0, 30, 5, 5, 0, 2, 25, 6, 
    1, 0, 0, 16, 0, 0, 0, 6, 27, 0, 0, 0, 0, 31, 3, 
    0, 0, 0, 0, 5, 33, 38, 44, 39, 0, 25, 12, 22, 18, 0, 
    0, 9, 18, 0, 0, 0, 0, 3, 5, 0, 0, 13, 0, 0, 0, 
    
    -- channel=401
    124, 127, 138, 138, 132, 122, 120, 107, 101, 96, 81, 56, 19, 42, 60, 
    125, 108, 120, 118, 110, 101, 101, 90, 85, 79, 61, 27, 13, 46, 67, 
    98, 104, 99, 95, 91, 85, 87, 81, 77, 75, 7, 3, 21, 50, 62, 
    84, 85, 84, 82, 86, 86, 80, 73, 66, 51, 10, 32, 65, 76, 74, 
    82, 88, 88, 86, 86, 67, 63, 62, 33, 0, 0, 7, 49, 69, 69, 
    87, 86, 84, 84, 75, 24, 0, 0, 0, 0, 0, 0, 19, 38, 65, 
    86, 86, 82, 74, 19, 34, 17, 27, 24, 0, 0, 0, 0, 19, 46, 
    87, 83, 44, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    85, 60, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 23, 0, 0, 0, 0, 0, 0, 0, 14, 22, 7, 0, 0, 25, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 4, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 21, 
    30, 1, 0, 0, 23, 37, 37, 38, 10, 2, 0, 0, 25, 3, 6, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 2, 0, 0, 0, 
    
    -- channel=402
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=403
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 32, 30, 6, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 15, 0, 10, 78, 57, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 32, 147, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 18, 46, 52, 35, 53, 93, 41, 0, 34, 
    0, 0, 0, 0, 23, 0, 0, 33, 40, 46, 84, 62, 10, 6, 37, 
    0, 0, 67, 0, 12, 0, 0, 37, 40, 27, 2, 84, 45, 43, 34, 
    0, 0, 66, 16, 0, 0, 0, 42, 70, 9, 0, 0, 45, 32, 26, 
    0, 0, 45, 32, 0, 0, 0, 46, 116, 4, 10, 0, 21, 64, 0, 
    0, 0, 28, 32, 3, 51, 19, 42, 107, 0, 41, 0, 0, 34, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 22, 9, 0, 0, 0, 
    0, 0, 11, 26, 4, 8, 7, 4, 1, 0, 2, 0, 0, 0, 0, 
    
    -- channel=404
    57, 50, 51, 52, 41, 41, 42, 32, 40, 22, 24, 19, 0, 22, 19, 
    44, 39, 37, 35, 31, 29, 31, 27, 29, 25, 26, 10, 0, 41, 20, 
    31, 23, 27, 25, 29, 28, 28, 29, 28, 32, 13, 0, 17, 33, 17, 
    27, 30, 30, 27, 32, 30, 27, 28, 30, 29, 0, 37, 30, 26, 19, 
    29, 30, 30, 27, 32, 25, 25, 23, 27, 1, 0, 32, 13, 20, 24, 
    30, 28, 28, 26, 31, 28, 20, 9, 11, 0, 0, 0, 28, 0, 22, 
    30, 28, 20, 26, 27, 19, 0, 0, 0, 73, 27, 0, 24, 2, 12, 
    30, 24, 24, 16, 0, 20, 0, 4, 35, 63, 4, 0, 0, 22, 14, 
    27, 25, 18, 5, 0, 19, 63, 31, 7, 0, 0, 0, 10, 41, 15, 
    32, 35, 0, 18, 0, 31, 83, 5, 0, 0, 0, 0, 12, 0, 0, 
    64, 10, 0, 0, 0, 24, 93, 0, 0, 0, 42, 42, 0, 0, 0, 
    26, 17, 0, 0, 15, 32, 58, 0, 0, 5, 0, 80, 0, 0, 5, 
    22, 8, 0, 0, 34, 8, 44, 0, 0, 20, 0, 28, 17, 0, 18, 
    20, 13, 0, 0, 27, 10, 5, 1, 0, 24, 0, 0, 15, 0, 14, 
    12, 0, 0, 0, 6, 4, 5, 3, 3, 35, 0, 0, 8, 10, 16, 
    
    -- channel=405
    91, 87, 86, 83, 81, 80, 79, 74, 78, 60, 60, 59, 43, 33, 57, 
    85, 79, 86, 88, 86, 81, 80, 74, 73, 68, 65, 47, 24, 48, 68, 
    75, 76, 78, 82, 79, 78, 78, 73, 72, 72, 51, 21, 37, 57, 65, 
    73, 78, 80, 78, 80, 81, 81, 73, 68, 63, 28, 22, 51, 64, 66, 
    80, 83, 83, 81, 82, 74, 66, 65, 54, 35, 10, 32, 58, 65, 67, 
    83, 84, 81, 79, 79, 56, 36, 36, 33, 16, 3, 2, 24, 50, 64, 
    84, 83, 80, 76, 58, 43, 6, 0, 10, 16, 16, 0, 18, 30, 49, 
    83, 81, 68, 55, 25, 24, 21, 7, 12, 20, 0, 0, 9, 29, 25, 
    83, 75, 37, 11, 13, 13, 8, 22, 2, 0, 0, 0, 43, 25, 29, 
    82, 48, 4, 19, 7, 23, 25, 4, 0, 0, 1, 0, 22, 5, 0, 
    73, 38, 0, 15, 9, 22, 20, 0, 0, 0, 10, 8, 0, 0, 1, 
    70, 8, 10, 8, 19, 26, 8, 0, 0, 16, 11, 34, 0, 0, 11, 
    57, 23, 16, 0, 17, 9, 13, 0, 0, 23, 11, 20, 22, 0, 30, 
    52, 33, 19, 5, 19, 6, 0, 0, 0, 26, 8, 9, 26, 5, 28, 
    48, 31, 8, 10, 17, 16, 17, 19, 18, 31, 18, 10, 22, 22, 22, 
    
    -- channel=406
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 4, 13, 5, 
    0, 0, 0, 0, 0, 3, 3, 5, 4, 7, 0, 0, 10, 7, 0, 
    4, 3, 3, 3, 4, 6, 12, 15, 10, 0, 0, 11, 6, 1, 1, 
    3, 2, 2, 1, 2, 0, 0, 14, 62, 69, 31, 1, 1, 0, 1, 
    4, 2, 3, 2, 9, 38, 0, 0, 0, 0, 8, 11, 0, 0, 1, 
    3, 3, 0, 6, 0, 0, 0, 8, 15, 50, 4, 19, 10, 0, 0, 
    1, 3, 8, 1, 6, 0, 3, 97, 114, 33, 0, 0, 0, 10, 48, 
    0, 14, 10, 0, 0, 1, 18, 0, 0, 0, 2, 34, 49, 44, 0, 
    14, 41, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 3, 37, 32, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 16, 3, 0, 17, 2, 12, 0, 0, 15, 9, 0, 0, 0, 9, 
    0, 0, 1, 23, 48, 52, 28, 12, 0, 7, 20, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 4, 1, 
    0, 13, 39, 29, 12, 17, 17, 16, 14, 0, 0, 0, 5, 5, 6, 
    
    -- channel=407
    119, 119, 127, 130, 121, 107, 102, 92, 76, 70, 60, 33, 0, 1, 34, 
    108, 96, 98, 92, 81, 71, 71, 65, 58, 55, 29, 12, 0, 8, 36, 
    65, 67, 64, 61, 59, 53, 56, 56, 53, 49, 0, 0, 0, 22, 36, 
    49, 51, 50, 52, 54, 54, 46, 49, 46, 31, 0, 0, 37, 47, 46, 
    45, 52, 52, 51, 50, 40, 26, 25, 1, 0, 0, 0, 10, 38, 38, 
    50, 50, 50, 50, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    50, 50, 48, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    50, 47, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=408
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 14, 35, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 51, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 1, 
    0, 0, 0, 0, 0, 9, 23, 86, 53, 0, 0, 0, 22, 28, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 27, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 38, 0, 0, 0, 0, 46, 92, 0, 0, 0, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 21, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 4, 19, 43, 
    0, 0, 14, 45, 84, 100, 99, 100, 35, 3, 0, 28, 80, 53, 40, 
    0, 0, 0, 0, 0, 0, 0, 10, 22, 50, 17, 36, 36, 35, 24, 
    
    -- channel=409
    28, 43, 35, 41, 44, 42, 34, 42, 35, 39, 27, 20, 62, 0, 22, 
    34, 40, 50, 44, 40, 38, 33, 34, 30, 28, 4, 58, 18, 0, 25, 
    42, 40, 31, 38, 29, 27, 29, 25, 24, 16, 29, 20, 12, 3, 35, 
    21, 24, 26, 29, 23, 24, 15, 22, 22, 26, 73, 0, 3, 28, 28, 
    22, 27, 28, 29, 20, 24, 16, 6, 0, 31, 29, 10, 25, 30, 24, 
    24, 29, 30, 30, 10, 0, 0, 32, 39, 12, 0, 132, 0, 18, 27, 
    28, 30, 37, 11, 17, 33, 31, 37, 0, 0, 0, 72, 61, 5, 14, 
    27, 31, 0, 33, 26, 0, 15, 0, 0, 0, 0, 132, 15, 0, 0, 
    31, 1, 56, 0, 54, 0, 0, 0, 6, 0, 40, 73, 0, 0, 0, 
    0, 0, 110, 0, 44, 0, 0, 0, 0, 80, 0, 0, 7, 8, 47, 
    0, 48, 19, 32, 11, 0, 0, 0, 90, 25, 19, 0, 26, 40, 74, 
    21, 0, 0, 58, 0, 0, 0, 0, 127, 0, 17, 0, 0, 100, 0, 
    12, 0, 0, 23, 0, 0, 0, 0, 107, 0, 27, 23, 0, 61, 0, 
    11, 8, 26, 19, 13, 18, 19, 23, 31, 0, 22, 44, 16, 3, 2, 
    12, 16, 0, 13, 2, 0, 6, 8, 11, 0, 23, 15, 6, 4, 0, 
    
    -- channel=410
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 15, 3, 
    
    -- channel=411
    30, 6, 15, 1, 0, 0, 6, 0, 0, 0, 0, 3, 0, 11, 4, 
    5, 0, 0, 0, 0, 0, 6, 0, 3, 4, 17, 0, 0, 39, 7, 
    0, 0, 0, 0, 6, 6, 9, 9, 10, 15, 9, 0, 4, 36, 0, 
    8, 11, 9, 7, 13, 13, 18, 16, 14, 4, 0, 15, 16, 3, 2, 
    15, 11, 9, 7, 16, 16, 14, 16, 29, 0, 0, 14, 3, 4, 6, 
    13, 9, 7, 7, 19, 43, 47, 0, 0, 0, 27, 0, 23, 0, 4, 
    10, 8, 2, 16, 22, 0, 0, 0, 0, 73, 83, 0, 0, 18, 0, 
    8, 4, 26, 0, 0, 12, 0, 41, 95, 79, 0, 0, 0, 13, 58, 
    5, 19, 0, 2, 0, 2, 55, 89, 0, 0, 0, 0, 52, 50, 42, 
    26, 89, 0, 10, 0, 21, 71, 24, 0, 0, 0, 0, 18, 0, 0, 
    39, 1, 0, 0, 0, 47, 87, 5, 0, 0, 0, 81, 0, 0, 0, 
    15, 0, 26, 0, 19, 53, 72, 0, 0, 4, 0, 50, 8, 0, 0, 
    11, 9, 36, 0, 67, 40, 58, 0, 0, 41, 0, 0, 48, 0, 12, 
    11, 13, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 11, 0, 9, 
    11, 0, 6, 0, 6, 8, 4, 0, 0, 36, 0, 0, 5, 6, 15, 
    
    -- channel=412
    17, 15, 21, 15, 18, 12, 14, 14, 0, 7, 13, 6, 0, 11, 7, 
    16, 11, 8, 8, 11, 8, 9, 9, 5, 11, 8, 0, 12, 0, 5, 
    7, 10, 9, 8, 6, 6, 6, 8, 7, 5, 0, 28, 0, 0, 9, 
    5, 2, 2, 3, 4, 6, 14, 7, 6, 0, 3, 0, 4, 0, 12, 
    2, 1, 1, 5, 5, 9, 14, 16, 7, 0, 0, 0, 7, 7, 4, 
    3, 2, 3, 5, 4, 6, 1, 8, 3, 65, 91, 0, 0, 22, 0, 
    1, 2, 5, 9, 0, 0, 0, 0, 8, 0, 0, 83, 0, 11, 7, 
    1, 4, 11, 0, 2, 0, 16, 25, 0, 0, 0, 32, 45, 0, 17, 
    1, 9, 0, 2, 6, 0, 0, 7, 0, 19, 16, 6, 7, 0, 0, 
    5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 63, 68, 0, 0, 0, 
    0, 0, 74, 0, 0, 0, 0, 3, 0, 20, 0, 15, 13, 0, 23, 
    0, 0, 43, 0, 0, 0, 0, 0, 52, 0, 0, 0, 36, 9, 8, 
    0, 0, 22, 0, 0, 0, 0, 0, 37, 0, 0, 0, 5, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 70, 0, 11, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 11, 0, 0, 0, 
    
    -- channel=413
    49, 54, 48, 50, 56, 50, 42, 52, 35, 28, 35, 25, 27, 3, 35, 
    47, 54, 59, 51, 47, 44, 40, 42, 37, 36, 21, 39, 28, 1, 38, 
    37, 44, 41, 44, 37, 39, 40, 37, 37, 31, 0, 36, 31, 19, 43, 
    35, 35, 37, 39, 37, 38, 36, 39, 38, 26, 42, 0, 25, 32, 39, 
    36, 38, 37, 39, 33, 28, 24, 28, 24, 58, 47, 13, 38, 38, 33, 
    37, 39, 40, 38, 21, 0, 0, 12, 0, 0, 8, 122, 0, 49, 33, 
    38, 40, 43, 25, 0, 0, 8, 15, 0, 0, 0, 163, 33, 0, 26, 
    38, 41, 9, 27, 24, 0, 23, 6, 0, 0, 1, 112, 59, 0, 0, 
    40, 16, 17, 0, 37, 0, 0, 0, 0, 0, 53, 115, 0, 0, 0, 
    15, 0, 114, 0, 42, 0, 0, 0, 0, 18, 0, 57, 13, 12, 26, 
    0, 0, 61, 23, 16, 0, 0, 0, 58, 38, 0, 0, 22, 20, 62, 
    0, 0, 0, 57, 0, 0, 0, 0, 144, 0, 18, 0, 0, 92, 8, 
    0, 0, 0, 49, 0, 2, 0, 0, 136, 0, 45, 0, 0, 72, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 38, 0, 25, 35, 0, 9, 0, 
    14, 13, 6, 26, 5, 6, 9, 11, 11, 0, 9, 23, 3, 1, 0, 
    
    -- channel=414
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=415
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 31, 45, 1, 3, 0, 0, 
    0, 0, 0, 0, 0, 4, 4, 7, 1, 36, 37, 58, 0, 11, 0, 
    0, 0, 0, 0, 0, 10, 35, 36, 22, 0, 21, 106, 20, 9, 7, 
    0, 0, 0, 11, 33, 9, 36, 35, 27, 0, 47, 86, 38, 11, 9, 
    0, 0, 18, 23, 37, 8, 0, 1, 37, 51, 66, 88, 27, 14, 23, 
    0, 0, 77, 18, 36, 0, 0, 38, 47, 41, 31, 64, 36, 44, 37, 
    0, 22, 70, 28, 23, 9, 0, 45, 58, 62, 3, 0, 56, 44, 57, 
    0, 21, 38, 47, 12, 3, 0, 47, 105, 18, 28, 0, 35, 71, 15, 
    4, 20, 31, 54, 14, 40, 18, 51, 99, 13, 42, 10, 2, 60, 2, 
    4, 11, 17, 21, 0, 14, 17, 22, 58, 1, 44, 32, 7, 21, 6, 
    9, 27, 34, 30, 22, 23, 22, 21, 19, 0, 21, 27, 9, 8, 5, 
    
    -- channel=416
    15, 2, 14, 5, 0, 0, 8, 0, 10, 0, 0, 4, 0, 32, 0, 
    8, 0, 0, 0, 1, 0, 7, 0, 3, 0, 17, 0, 0, 46, 0, 
    6, 0, 6, 0, 8, 5, 5, 4, 4, 13, 3, 0, 0, 29, 0, 
    10, 11, 9, 3, 10, 8, 9, 0, 2, 4, 0, 44, 18, 3, 0, 
    13, 9, 9, 4, 17, 7, 14, 11, 15, 0, 0, 17, 0, 0, 4, 
    12, 7, 4, 3, 26, 32, 20, 0, 13, 1, 0, 0, 56, 0, 1, 
    8, 6, 0, 20, 20, 17, 0, 0, 5, 135, 71, 0, 0, 30, 6, 
    9, 1, 26, 0, 0, 23, 0, 14, 28, 54, 0, 0, 0, 25, 38, 
    5, 25, 0, 20, 0, 32, 102, 81, 3, 0, 0, 0, 29, 28, 25, 
    36, 66, 0, 23, 0, 44, 153, 27, 2, 0, 57, 0, 0, 0, 0, 
    75, 34, 0, 0, 0, 53, 130, 9, 0, 0, 36, 160, 0, 0, 0, 
    26, 3, 0, 0, 24, 59, 120, 0, 0, 10, 0, 112, 27, 0, 0, 
    20, 16, 23, 0, 63, 6, 60, 0, 0, 50, 0, 1, 75, 0, 22, 
    11, 20, 10, 0, 53, 43, 38, 27, 0, 61, 0, 0, 24, 0, 14, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 1, 4, 16, 
    
    -- channel=417
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=418
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=419
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 45, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 26, 32, 12, 0, 1, 76, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 33, 80, 26, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 0, 28, 35, 62, 59, 0, 0, 0, 
    0, 0, 51, 1, 25, 0, 0, 25, 32, 50, 15, 18, 0, 23, 36, 
    0, 7, 59, 21, 7, 0, 0, 31, 74, 53, 13, 0, 49, 48, 55, 
    0, 3, 24, 32, 0, 0, 0, 33, 96, 2, 10, 0, 21, 66, 0, 
    0, 0, 17, 26, 0, 10, 4, 36, 85, 0, 22, 2, 3, 49, 0, 
    0, 0, 23, 25, 18, 32, 35, 40, 52, 0, 25, 18, 7, 9, 0, 
    0, 0, 5, 9, 2, 3, 6, 6, 4, 0, 15, 13, 0, 0, 0, 
    
    -- channel=420
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 59, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 26, 48, 63, 42, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 26, 0, 0, 
    0, 0, 0, 22, 19, 20, 0, 0, 0, 7, 0, 30, 0, 0, 0, 
    0, 0, 0, 4, 23, 8, 0, 0, 0, 32, 68, 0, 0, 0, 7, 
    0, 46, 44, 4, 21, 0, 0, 0, 20, 89, 35, 58, 27, 32, 76, 
    0, 9, 0, 5, 0, 0, 0, 0, 22, 0, 0, 11, 22, 26, 14, 
    0, 2, 0, 0, 0, 0, 0, 0, 11, 0, 0, 1, 26, 53, 5, 
    0, 1, 29, 58, 64, 102, 114, 120, 100, 11, 22, 9, 25, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 32, 27, 0, 0, 0, 
    
    -- channel=421
    62, 71, 76, 77, 75, 69, 66, 60, 58, 41, 35, 31, 20, 2, 15, 
    80, 73, 70, 73, 69, 60, 55, 50, 44, 36, 32, 23, 0, 0, 25, 
    64, 61, 58, 56, 48, 45, 43, 39, 37, 35, 45, 4, 0, 10, 29, 
    38, 41, 42, 41, 42, 45, 47, 41, 39, 40, 9, 0, 9, 28, 31, 
    37, 44, 45, 46, 47, 52, 46, 46, 35, 29, 0, 0, 28, 33, 30, 
    42, 46, 45, 45, 45, 40, 48, 57, 66, 51, 19, 0, 2, 19, 26, 
    46, 47, 47, 41, 51, 34, 18, 0, 0, 0, 42, 0, 0, 2, 14, 
    47, 47, 44, 39, 14, 7, 0, 0, 0, 21, 43, 30, 0, 0, 0, 
    48, 44, 23, 10, 0, 0, 0, 47, 58, 56, 43, 0, 1, 4, 22, 
    44, 58, 0, 0, 0, 0, 12, 42, 43, 53, 59, 29, 26, 25, 30, 
    61, 51, 6, 0, 0, 0, 3, 34, 37, 0, 0, 45, 36, 26, 0, 
    41, 0, 1, 0, 0, 0, 22, 37, 0, 0, 0, 2, 25, 0, 0, 
    24, 0, 2, 0, 0, 0, 20, 33, 0, 0, 0, 0, 17, 0, 0, 
    11, 7, 5, 0, 8, 25, 32, 33, 4, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=422
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 30, 60, 64, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 18, 9, 0, 0, 18, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 74, 9, 0, 0, 
    0, 0, 0, 9, 26, 0, 0, 19, 43, 32, 31, 0, 0, 0, 6, 
    0, 0, 25, 4, 8, 0, 0, 32, 33, 76, 60, 10, 11, 23, 34, 
    0, 60, 38, 12, 0, 0, 0, 30, 64, 21, 9, 32, 51, 48, 36, 
    0, 0, 23, 12, 0, 10, 2, 34, 52, 0, 0, 4, 25, 39, 0, 
    0, 5, 21, 0, 0, 0, 4, 23, 38, 0, 0, 0, 29, 25, 0, 
    0, 6, 42, 39, 48, 60, 66, 67, 50, 3, 11, 4, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 25, 0, 0, 0, 0, 
    
    -- channel=423
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=424
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 2, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 19, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 22, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 14, 18, 29, 6, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 14, 0, 1, 
    0, 0, 0, 0, 4, 6, 20, 26, 23, 0, 0, 17, 22, 18, 4, 
    0, 0, 0, 1, 13, 4, 13, 0, 0, 0, 0, 28, 7, 2, 2, 
    0, 0, 31, 1, 23, 5, 0, 0, 0, 0, 3, 29, 2, 0, 0, 
    0, 0, 18, 6, 22, 14, 0, 0, 0, 17, 0, 0, 0, 0, 19, 
    0, 1, 1, 26, 19, 0, 0, 0, 33, 6, 16, 0, 0, 19, 17, 
    0, 1, 0, 31, 10, 10, 0, 0, 33, 10, 17, 2, 0, 31, 7, 
    0, 0, 0, 9, 0, 0, 0, 0, 18, 0, 11, 17, 0, 19, 14, 
    3, 9, 18, 18, 21, 19, 18, 17, 18, 0, 5, 24, 20, 19, 18, 
    
    -- channel=425
    27, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 10, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 8, 0, 21, 23, 6, 
    0, 0, 0, 0, 3, 2, 10, 15, 16, 8, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 10, 3, 2, 27, 54, 36, 24, 8, 0, 0, 
    0, 0, 0, 0, 0, 24, 74, 52, 0, 0, 76, 26, 0, 14, 0, 
    0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 19, 58, 9, 0, 0, 
    0, 0, 10, 27, 0, 1, 2, 65, 135, 120, 6, 0, 2, 0, 61, 
    0, 0, 0, 0, 0, 0, 0, 62, 0, 0, 0, 0, 26, 82, 41, 
    0, 83, 27, 0, 0, 0, 0, 0, 0, 0, 0, 68, 72, 10, 0, 
    0, 0, 0, 0, 0, 23, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 12, 12, 0, 3, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 9, 49, 67, 25, 0, 2, 10, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 7, 39, 20, 22, 16, 8, 4, 0, 0, 0, 3, 3, 6, 
    
    -- channel=426
    164, 154, 153, 148, 136, 125, 122, 110, 100, 75, 76, 66, 38, 18, 60, 
    134, 125, 120, 112, 103, 95, 96, 89, 83, 82, 73, 52, 8, 47, 68, 
    94, 81, 83, 85, 83, 81, 85, 84, 85, 83, 68, 9, 34, 73, 72, 
    70, 78, 80, 81, 84, 87, 89, 93, 90, 85, 16, 10, 62, 74, 69, 
    76, 81, 81, 82, 85, 91, 83, 80, 77, 67, 14, 38, 60, 66, 67, 
    82, 82, 81, 81, 79, 69, 78, 73, 60, 14, 37, 28, 11, 47, 58, 
    83, 81, 81, 72, 73, 36, 0, 0, 0, 11, 56, 0, 17, 11, 34, 
    80, 81, 69, 64, 19, 28, 14, 12, 51, 97, 42, 7, 0, 12, 35, 
    80, 71, 40, 0, 3, 3, 7, 79, 52, 30, 33, 0, 24, 47, 52, 
    75, 86, 8, 6, 0, 10, 31, 36, 24, 32, 8, 28, 54, 31, 29, 
    79, 27, 0, 6, 0, 7, 43, 28, 23, 0, 8, 4, 12, 9, 0, 
    57, 5, 5, 0, 3, 25, 31, 33, 0, 5, 0, 27, 4, 0, 0, 
    36, 10, 8, 0, 18, 26, 52, 20, 0, 11, 8, 14, 15, 0, 13, 
    37, 22, 10, 0, 5, 0, 0, 0, 0, 16, 0, 0, 1, 0, 8, 
    36, 14, 0, 4, 0, 1, 3, 1, 1, 13, 2, 0, 4, 5, 9, 
    
    -- channel=427
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 22, 0, 6, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 30, 25, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 21, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 45, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 60, 10, 8, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 166, 0, 22, 4, 
    0, 0, 2, 0, 0, 0, 5, 22, 0, 0, 0, 171, 58, 0, 0, 
    0, 0, 0, 13, 24, 0, 23, 11, 12, 0, 7, 116, 56, 0, 0, 
    0, 0, 24, 0, 40, 0, 0, 0, 0, 0, 56, 127, 0, 0, 0, 
    0, 0, 143, 0, 51, 0, 0, 0, 0, 24, 0, 51, 21, 17, 34, 
    0, 0, 61, 32, 22, 0, 0, 0, 72, 43, 0, 0, 23, 27, 62, 
    0, 0, 0, 70, 0, 0, 0, 5, 157, 0, 26, 0, 0, 104, 5, 
    0, 0, 0, 65, 0, 14, 0, 5, 156, 0, 60, 13, 0, 80, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 24, 45, 0, 11, 0, 
    0, 15, 16, 42, 16, 15, 21, 20, 19, 0, 5, 27, 8, 6, 0, 
    
    -- channel=428
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 31, 13, 20, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 11, 17, 15, 19, 55, 60, 0, 13, 8, 0, 
    0, 0, 0, 0, 0, 14, 0, 2, 3, 65, 36, 0, 0, 14, 8, 
    0, 0, 0, 19, 11, 35, 44, 70, 42, 30, 14, 0, 0, 23, 25, 
    0, 0, 0, 38, 2, 42, 88, 51, 39, 44, 40, 0, 27, 29, 27, 
    0, 38, 0, 26, 9, 35, 90, 44, 31, 0, 64, 88, 30, 33, 0, 
    0, 25, 32, 0, 25, 64, 84, 39, 0, 27, 11, 80, 42, 0, 8, 
    0, 27, 42, 0, 45, 30, 69, 36, 0, 36, 2, 36, 68, 0, 19, 
    0, 23, 49, 39, 77, 68, 68, 62, 0, 56, 8, 8, 39, 12, 20, 
    0, 0, 14, 16, 25, 25, 24, 20, 17, 44, 27, 6, 19, 20, 24, 
    
    -- channel=429
    0, 9, 0, 4, 7, 6, 0, 12, 0, 0, 8, 1, 19, 0, 8, 
    0, 8, 10, 6, 2, 4, 0, 5, 2, 5, 0, 24, 25, 0, 5, 
    1, 8, 3, 4, 0, 1, 0, 0, 1, 0, 0, 27, 9, 0, 9, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 2, 36, 0, 2, 3, 6, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 25, 40, 2, 2, 4, 1, 
    0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 154, 0, 14, 3, 
    0, 3, 7, 0, 0, 0, 13, 42, 0, 0, 0, 148, 51, 0, 2, 
    1, 5, 0, 6, 12, 0, 9, 0, 0, 0, 0, 102, 68, 0, 0, 
    4, 0, 21, 0, 30, 0, 0, 0, 0, 0, 42, 140, 0, 0, 0, 
    0, 0, 123, 0, 57, 0, 0, 0, 0, 40, 0, 41, 0, 3, 35, 
    0, 0, 63, 25, 32, 0, 0, 0, 62, 76, 0, 0, 31, 35, 75, 
    0, 18, 0, 60, 0, 0, 0, 0, 128, 0, 17, 0, 0, 91, 16, 
    0, 0, 0, 63, 0, 0, 0, 4, 140, 0, 39, 22, 0, 94, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 49, 0, 18, 44, 0, 23, 0, 
    0, 10, 1, 20, 3, 0, 6, 9, 9, 0, 13, 35, 1, 0, 0, 
    
    -- channel=430
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 1, 0, 0, 0, 4, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 4, 0, 2, 1, 1, 0, 1, 0, 0, 6, 4, 4, 3, 
    
    -- channel=431
    0, 16, 17, 23, 29, 23, 17, 26, 2, 26, 10, 4, 26, 12, 6, 
    18, 20, 26, 18, 15, 14, 9, 14, 6, 7, 0, 8, 23, 0, 3, 
    22, 26, 15, 11, 3, 1, 1, 0, 0, 0, 0, 59, 7, 0, 11, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 6, 9, 
    0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 28, 2, 20, 10, 3, 
    0, 0, 0, 0, 0, 0, 0, 27, 38, 78, 25, 90, 0, 36, 5, 
    0, 0, 4, 0, 0, 8, 34, 45, 16, 0, 0, 169, 1, 14, 22, 
    0, 1, 0, 0, 30, 0, 27, 0, 0, 0, 10, 144, 80, 0, 0, 
    0, 0, 0, 5, 54, 0, 0, 0, 23, 34, 66, 127, 0, 0, 0, 
    0, 0, 106, 0, 54, 0, 0, 0, 18, 57, 49, 79, 0, 16, 43, 
    0, 10, 114, 22, 30, 0, 0, 7, 78, 101, 0, 0, 60, 58, 116, 
    0, 0, 13, 61, 0, 0, 0, 16, 174, 0, 16, 0, 10, 109, 18, 
    0, 0, 0, 51, 0, 0, 0, 15, 156, 0, 31, 0, 0, 113, 0, 
    0, 0, 11, 38, 0, 24, 35, 45, 118, 0, 39, 34, 0, 30, 0, 
    0, 5, 0, 4, 0, 0, 0, 2, 5, 0, 34, 45, 0, 0, 0, 
    
    -- channel=432
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 13, 0, 
    0, 0, 0, 0, 0, 0, 5, 11, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 59, 79, 43, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 39, 0, 0, 0, 52, 26, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 49, 15, 0, 0, 
    0, 0, 6, 15, 0, 0, 0, 116, 172, 109, 0, 0, 0, 6, 77, 
    0, 2, 0, 0, 0, 0, 5, 20, 0, 0, 0, 0, 45, 95, 9, 
    1, 85, 7, 0, 0, 0, 0, 0, 0, 0, 0, 46, 44, 0, 0, 
    0, 0, 0, 0, 0, 45, 41, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 5, 9, 0, 0, 9, 4, 0, 0, 0, 0, 
    0, 0, 0, 25, 70, 78, 29, 0, 0, 9, 31, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 31, 49, 23, 27, 22, 15, 10, 0, 0, 0, 4, 5, 8, 
    
    -- channel=433
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 0, 7, 16, 0, 
    0, 0, 0, 0, 0, 0, 7, 6, 5, 2, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 6, 45, 41, 25, 19, 0, 0, 0, 
    0, 0, 0, 0, 11, 47, 54, 0, 0, 0, 52, 0, 0, 0, 0, 
    0, 0, 0, 5, 21, 0, 0, 0, 0, 81, 53, 0, 7, 0, 0, 
    0, 0, 25, 16, 0, 16, 1, 91, 149, 127, 18, 0, 0, 25, 68, 
    0, 20, 1, 0, 0, 0, 58, 69, 0, 0, 0, 0, 58, 98, 36, 
    25, 105, 0, 13, 0, 14, 73, 12, 8, 0, 0, 25, 56, 12, 0, 
    36, 0, 0, 0, 0, 60, 101, 13, 0, 0, 0, 16, 0, 0, 0, 
    9, 19, 10, 0, 32, 43, 71, 12, 0, 17, 2, 25, 7, 0, 1, 
    10, 17, 15, 4, 88, 77, 68, 13, 0, 38, 9, 5, 0, 0, 0, 
    11, 11, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 5, 
    8, 10, 27, 30, 22, 24, 18, 13, 6, 6, 0, 0, 7, 7, 15, 
    
    -- channel=434
    14, 23, 22, 24, 25, 24, 21, 22, 16, 26, 8, 10, 13, 5, 6, 
    29, 28, 30, 30, 29, 26, 22, 21, 16, 13, 14, 8, 0, 0, 12, 
    29, 30, 28, 27, 21, 21, 20, 15, 14, 12, 18, 21, 0, 3, 15, 
    18, 19, 21, 20, 18, 20, 21, 17, 16, 13, 19, 0, 2, 14, 14, 
    18, 21, 22, 22, 22, 22, 23, 23, 19, 19, 14, 0, 18, 13, 14, 
    21, 23, 23, 21, 20, 20, 32, 43, 44, 57, 32, 18, 6, 18, 13, 
    23, 24, 23, 20, 19, 22, 24, 13, 1, 0, 36, 60, 0, 14, 12, 
    24, 24, 24, 20, 21, 4, 13, 0, 0, 1, 52, 73, 17, 0, 3, 
    25, 21, 14, 16, 16, 0, 0, 25, 54, 60, 57, 48, 12, 0, 30, 
    21, 17, 39, 0, 5, 0, 0, 43, 50, 55, 60, 56, 30, 38, 36, 
    8, 43, 42, 1, 0, 0, 0, 43, 49, 31, 0, 22, 51, 40, 34, 
    7, 3, 21, 12, 0, 0, 7, 47, 64, 0, 0, 0, 31, 37, 0, 
    4, 7, 17, 12, 0, 12, 14, 44, 55, 0, 11, 0, 7, 26, 0, 
    2, 4, 10, 7, 1, 20, 25, 29, 38, 0, 18, 0, 0, 0, 0, 
    9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    
    -- channel=435
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 19, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 49, 63, 49, 9, 80, 45, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 56, 13, 0, 0, 
    0, 0, 0, 6, 0, 2, 11, 29, 72, 128, 76, 35, 8, 0, 26, 
    0, 0, 0, 0, 5, 0, 0, 97, 74, 50, 55, 0, 0, 51, 58, 
    0, 48, 47, 3, 0, 0, 25, 57, 53, 45, 9, 74, 84, 54, 37, 
    0, 0, 15, 12, 0, 13, 48, 56, 54, 0, 0, 0, 41, 28, 0, 
    0, 5, 29, 5, 5, 35, 43, 67, 28, 4, 0, 3, 21, 10, 0, 
    0, 8, 27, 10, 38, 63, 71, 49, 31, 11, 28, 8, 6, 0, 0, 
    0, 2, 12, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 1, 24, 12, 13, 10, 3, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=436
    59, 67, 73, 75, 76, 73, 71, 69, 66, 64, 56, 44, 21, 37, 47, 
    75, 67, 77, 81, 78, 72, 70, 65, 62, 55, 43, 27, 23, 29, 52, 
    65, 77, 76, 73, 68, 65, 65, 58, 55, 53, 2, 16, 19, 29, 47, 
    65, 65, 64, 63, 63, 63, 57, 50, 45, 34, 20, 25, 42, 52, 57, 
    63, 67, 67, 65, 64, 47, 38, 41, 22, 1, 0, 5, 40, 53, 53, 
    65, 67, 66, 64, 55, 18, 0, 0, 0, 0, 0, 0, 19, 33, 52, 
    66, 67, 64, 57, 14, 19, 21, 40, 31, 0, 0, 0, 3, 22, 43, 
    67, 65, 36, 11, 12, 0, 0, 0, 0, 0, 0, 0, 9, 6, 0, 
    67, 48, 15, 7, 4, 7, 0, 0, 0, 0, 0, 35, 7, 0, 0, 
    57, 0, 0, 0, 17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 1, 17, 0, 0, 0, 0, 36, 17, 0, 0, 0, 34, 
    38, 0, 0, 7, 0, 0, 0, 0, 0, 0, 4, 0, 0, 7, 18, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 24, 20, 
    30, 2, 0, 7, 7, 22, 23, 27, 31, 0, 10, 14, 20, 21, 12, 
    23, 9, 0, 0, 0, 0, 0, 4, 8, 7, 7, 18, 9, 8, 3, 
    
    -- channel=437
    0, 0, 0, 0, 2, 2, 6, 0, 6, 28, 5, 0, 1, 26, 0, 
    2, 0, 0, 2, 4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 60, 0, 0, 49, 0, 0, 
    0, 0, 0, 0, 0, 44, 70, 71, 64, 61, 8, 0, 0, 39, 1, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 1, 41, 41, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 27, 51, 21, 12, 27, 97, 0, 0, 0, 0, 
    29, 87, 0, 0, 6, 0, 7, 7, 0, 67, 72, 159, 13, 23, 43, 
    26, 11, 3, 0, 0, 5, 38, 0, 0, 0, 0, 64, 45, 0, 6, 
    18, 14, 15, 0, 0, 0, 0, 6, 0, 5, 0, 0, 81, 1, 12, 
    0, 17, 40, 45, 92, 140, 152, 153, 79, 36, 17, 0, 48, 22, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 19, 5, 0, 0, 0, 
    
    -- channel=438
    10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 31, 64, 62, 38, 48, 52, 0, 1, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 55, 67, 4, 0, 0, 
    0, 0, 0, 3, 0, 0, 3, 0, 17, 77, 75, 82, 6, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 67, 83, 65, 77, 11, 0, 12, 50, 
    0, 4, 55, 0, 0, 0, 0, 55, 55, 77, 31, 59, 62, 52, 49, 
    0, 28, 19, 4, 0, 0, 3, 54, 75, 0, 0, 0, 54, 42, 8, 
    0, 0, 13, 8, 0, 3, 8, 67, 67, 0, 0, 0, 10, 37, 0, 
    0, 0, 11, 0, 0, 30, 46, 49, 56, 0, 13, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=439
    94, 106, 118, 122, 120, 112, 108, 100, 91, 77, 68, 49, 27, 28, 49, 
    116, 106, 112, 112, 104, 94, 92, 84, 78, 68, 50, 39, 6, 23, 55, 
    89, 94, 92, 88, 81, 75, 76, 70, 66, 61, 13, 0, 14, 32, 53, 
    73, 72, 71, 71, 72, 72, 67, 65, 59, 47, 10, 7, 39, 58, 63, 
    67, 73, 74, 72, 71, 61, 48, 48, 29, 16, 0, 1, 49, 64, 59, 
    70, 73, 73, 72, 59, 20, 0, 0, 0, 0, 0, 0, 7, 35, 57, 
    73, 73, 72, 60, 27, 10, 1, 17, 9, 0, 0, 0, 0, 8, 41, 
    73, 72, 37, 21, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    73, 47, 19, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=440
    78, 89, 84, 92, 93, 83, 73, 80, 62, 43, 53, 39, 45, 1, 39, 
    81, 84, 82, 75, 67, 62, 56, 60, 52, 52, 35, 55, 28, 0, 42, 
    60, 58, 53, 55, 48, 48, 48, 49, 48, 43, 25, 29, 26, 20, 49, 
    40, 42, 44, 47, 45, 45, 44, 51, 49, 47, 49, 0, 28, 42, 46, 
    37, 43, 44, 46, 40, 42, 36, 38, 34, 63, 44, 13, 37, 45, 40, 
    41, 44, 46, 45, 33, 8, 5, 21, 9, 0, 0, 115, 0, 39, 38, 
    44, 45, 50, 33, 18, 10, 13, 15, 0, 0, 0, 125, 39, 0, 21, 
    43, 47, 19, 37, 21, 0, 19, 0, 0, 0, 0, 78, 50, 0, 0, 
    44, 28, 38, 0, 29, 0, 0, 0, 0, 0, 43, 86, 0, 0, 0, 
    26, 0, 99, 0, 36, 0, 0, 0, 0, 20, 0, 40, 6, 3, 26, 
    0, 0, 44, 19, 18, 0, 0, 0, 51, 29, 0, 0, 15, 16, 48, 
    14, 4, 0, 41, 0, 0, 0, 0, 100, 0, 12, 0, 0, 66, 8, 
    8, 0, 0, 37, 0, 0, 0, 0, 102, 0, 32, 10, 0, 56, 0, 
    14, 0, 0, 3, 0, 0, 0, 0, 21, 0, 12, 31, 0, 11, 0, 
    14, 18, 0, 20, 3, 2, 6, 7, 9, 0, 12, 23, 5, 5, 0, 
    
    -- channel=441
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 27, 53, 62, 60, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 42, 24, 16, 30, 117, 20, 0, 1, 0, 
    0, 0, 0, 0, 4, 6, 16, 3, 22, 77, 109, 76, 0, 0, 2, 
    0, 0, 0, 23, 24, 16, 30, 103, 110, 112, 100, 8, 1, 19, 64, 
    0, 8, 11, 25, 1, 12, 49, 111, 104, 106, 98, 38, 58, 73, 68, 
    0, 77, 42, 19, 0, 6, 63, 103, 97, 27, 44, 103, 89, 78, 27, 
    0, 15, 59, 8, 0, 48, 83, 102, 51, 11, 8, 45, 75, 37, 0, 
    0, 24, 62, 5, 30, 54, 94, 98, 37, 25, 14, 9, 70, 6, 0, 
    0, 21, 55, 30, 61, 77, 81, 80, 35, 34, 26, 0, 19, 0, 0, 
    0, 0, 8, 3, 2, 3, 4, 0, 0, 23, 18, 0, 0, 0, 0, 
    
    -- channel=442
    6, 29, 40, 45, 50, 43, 41, 38, 32, 55, 26, 16, 25, 7, 8, 
    41, 32, 45, 44, 41, 34, 31, 28, 22, 15, 6, 9, 3, 0, 9, 
    44, 53, 35, 31, 23, 17, 18, 13, 10, 6, 1, 12, 0, 0, 14, 
    20, 13, 13, 13, 11, 13, 8, 5, 1, 4, 39, 0, 3, 22, 19, 
    10, 13, 15, 16, 13, 9, 15, 14, 0, 0, 0, 0, 15, 15, 13, 
    13, 14, 15, 17, 10, 0, 0, 0, 39, 66, 0, 4, 5, 15, 13, 
    13, 15, 21, 12, 0, 46, 72, 67, 42, 0, 0, 20, 0, 27, 13, 
    15, 18, 0, 0, 22, 0, 4, 0, 0, 0, 8, 84, 10, 0, 0, 
    18, 4, 7, 15, 34, 8, 0, 0, 27, 37, 56, 55, 0, 0, 0, 
    2, 0, 14, 0, 15, 0, 0, 24, 17, 66, 63, 0, 0, 1, 37, 
    0, 78, 48, 5, 0, 0, 0, 14, 76, 80, 34, 35, 46, 54, 95, 
    13, 0, 11, 13, 0, 0, 0, 6, 89, 0, 0, 0, 21, 62, 0, 
    1, 0, 9, 0, 0, 0, 0, 13, 54, 0, 0, 0, 31, 49, 0, 
    0, 0, 35, 29, 49, 97, 107, 114, 93, 0, 28, 3, 27, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 7, 0, 0, 0, 
    
    -- channel=443
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 12, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 33, 33, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 27, 33, 56, 32, 0, 0, 14, 22, 
    0, 28, 8, 0, 0, 0, 5, 27, 42, 21, 20, 29, 37, 32, 13, 
    0, 0, 0, 0, 0, 0, 13, 30, 15, 0, 0, 11, 15, 13, 0, 
    0, 0, 0, 0, 0, 0, 14, 31, 12, 0, 0, 0, 9, 3, 0, 
    0, 0, 14, 16, 29, 46, 50, 52, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=444
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 16, 3, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 6, 7, 0, 0, 
    8, 12, 4, 4, 1, 1, 0, 0, 0, 0, 16, 5, 0, 0, 0, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 29, 10, 0, 4, 0, 
    0, 2, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 3, 3, 0, 0, 0, 16, 49, 52, 0, 15, 13, 0, 0, 
    2, 4, 5, 0, 12, 41, 56, 53, 30, 11, 35, 4, 4, 13, 0, 
    5, 4, 0, 3, 23, 6, 7, 0, 0, 0, 49, 64, 12, 0, 0, 
    7, 0, 24, 27, 23, 16, 11, 13, 55, 60, 54, 38, 0, 0, 13, 
    0, 0, 22, 18, 16, 14, 16, 50, 55, 84, 67, 4, 8, 34, 53, 
    23, 73, 35, 16, 6, 0, 13, 45, 71, 58, 53, 63, 60, 63, 52, 
    19, 25, 17, 13, 0, 11, 28, 46, 43, 3, 8, 37, 42, 39, 2, 
    15, 20, 20, 3, 0, 0, 24, 49, 34, 1, 5, 17, 42, 32, 1, 
    7, 24, 43, 42, 61, 87, 94, 97, 55, 18, 24, 10, 24, 9, 0, 
    4, 9, 0, 0, 0, 0, 0, 0, 0, 21, 23, 7, 0, 0, 0, 
    
    -- channel=445
    186, 183, 189, 188, 180, 164, 159, 149, 130, 109, 108, 90, 39, 38, 84, 
    173, 162, 158, 151, 141, 129, 128, 121, 112, 109, 93, 67, 33, 46, 91, 
    122, 120, 119, 119, 115, 111, 114, 113, 111, 108, 57, 28, 49, 78, 95, 
    101, 107, 107, 108, 112, 114, 113, 114, 112, 96, 36, 18, 80, 96, 99, 
    102, 109, 109, 110, 111, 108, 95, 99, 86, 64, 20, 23, 71, 92, 92, 
    108, 109, 108, 108, 100, 77, 54, 44, 31, 32, 20, 10, 20, 58, 82, 
    110, 109, 107, 97, 66, 34, 11, 0, 9, 0, 18, 20, 3, 22, 49, 
    108, 108, 86, 55, 24, 22, 21, 9, 24, 13, 8, 26, 12, 13, 22, 
    106, 93, 31, 11, 12, 2, 0, 21, 14, 13, 16, 20, 34, 12, 24, 
    102, 52, 8, 0, 4, 0, 0, 7, 0, 5, 15, 14, 12, 6, 8, 
    71, 26, 0, 0, 2, 0, 0, 3, 0, 0, 0, 2, 0, 0, 12, 
    69, 0, 5, 4, 1, 0, 0, 3, 17, 2, 5, 0, 0, 7, 12, 
    51, 6, 1, 0, 0, 0, 0, 0, 8, 4, 4, 0, 3, 1, 15, 
    47, 20, 2, 0, 0, 0, 0, 0, 5, 0, 7, 5, 4, 2, 8, 
    45, 16, 0, 0, 0, 0, 0, 1, 4, 3, 4, 4, 7, 7, 8, 
    
    -- channel=446
    0, 5, 0, 7, 0, 4, 0, 4, 5, 0, 0, 1, 0, 20, 2, 
    9, 8, 2, 6, 2, 5, 0, 3, 4, 4, 6, 0, 5, 11, 0, 
    1, 2, 10, 4, 5, 6, 1, 2, 2, 11, 0, 17, 9, 0, 0, 
    5, 8, 7, 7, 7, 3, 2, 0, 3, 8, 0, 35, 6, 0, 0, 
    3, 7, 8, 5, 9, 0, 0, 2, 16, 0, 5, 21, 0, 1, 2, 
    6, 8, 6, 3, 10, 13, 0, 0, 0, 0, 0, 22, 21, 0, 2, 
    7, 8, 0, 10, 0, 0, 0, 3, 0, 87, 0, 0, 22, 0, 8, 
    11, 6, 15, 2, 0, 19, 0, 26, 14, 0, 0, 0, 23, 21, 0, 
    7, 16, 0, 4, 0, 8, 87, 0, 0, 0, 0, 37, 0, 44, 0, 
    28, 0, 0, 6, 13, 20, 82, 0, 0, 0, 0, 25, 0, 0, 0, 
    54, 0, 0, 0, 28, 20, 58, 0, 0, 36, 0, 0, 0, 0, 0, 
    0, 47, 0, 0, 21, 0, 41, 0, 0, 1, 0, 34, 0, 0, 32, 
    9, 0, 0, 36, 19, 0, 0, 0, 0, 3, 0, 26, 0, 14, 1, 
    3, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 2, 
    0, 0, 6, 0, 6, 1, 0, 0, 0, 0, 0, 19, 0, 2, 6, 
    
    -- channel=447
    0, 0, 0, 0, 2, 3, 2, 4, 2, 17, 5, 4, 0, 10, 0, 
    14, 2, 3, 6, 6, 5, 3, 4, 2, 0, 20, 0, 5, 0, 0, 
    0, 13, 9, 6, 4, 2, 1, 0, 0, 3, 0, 8, 3, 0, 0, 
    6, 0, 0, 0, 0, 0, 3, 3, 0, 0, 4, 8, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 23, 60, 34, 12, 0, 7, 2, 0, 
    0, 0, 0, 0, 13, 36, 0, 0, 0, 0, 0, 0, 10, 3, 0, 
    0, 0, 0, 13, 0, 1, 26, 41, 31, 58, 0, 7, 0, 4, 7, 
    0, 1, 15, 0, 22, 0, 16, 74, 41, 0, 0, 0, 0, 17, 14, 
    0, 25, 10, 16, 0, 20, 32, 0, 0, 5, 0, 56, 44, 0, 0, 
    28, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 12, 31, 0, 0, 0, 62, 12, 4, 0, 0, 21, 
    1, 9, 0, 3, 14, 0, 2, 0, 1, 8, 3, 0, 7, 0, 7, 
    6, 0, 2, 30, 24, 17, 0, 10, 0, 8, 2, 0, 0, 13, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 20, 0, 10, 12, 1, 
    0, 19, 39, 2, 5, 8, 5, 7, 7, 0, 0, 11, 1, 1, 2, 
    
    -- channel=448
    0, 0, 7, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 6, 3, 
    0, 0, 3, 4, 6, 13, 8, 3, 0, 7, 8, 12, 13, 14, 9, 
    0, 0, 0, 15, 8, 15, 16, 20, 18, 14, 11, 10, 5, 3, 2, 
    0, 5, 0, 8, 14, 17, 22, 25, 19, 11, 14, 1, 8, 6, 14, 
    23, 22, 0, 0, 9, 33, 19, 10, 20, 19, 20, 12, 20, 22, 23, 
    11, 2, 0, 0, 18, 34, 0, 6, 19, 20, 15, 20, 24, 25, 14, 
    0, 0, 0, 0, 7, 25, 3, 16, 17, 10, 12, 24, 13, 17, 0, 
    8, 12, 0, 6, 0, 30, 11, 25, 16, 1, 9, 13, 11, 12, 13, 
    16, 27, 22, 0, 13, 0, 29, 8, 11, 3, 8, 6, 16, 6, 5, 
    26, 16, 0, 0, 6, 0, 26, 1, 10, 8, 9, 0, 8, 0, 22, 
    0, 0, 0, 0, 0, 0, 4, 11, 15, 8, 8, 5, 8, 24, 14, 
    0, 0, 0, 0, 0, 8, 23, 0, 18, 17, 14, 9, 6, 36, 12, 
    0, 0, 3, 8, 0, 9, 21, 2, 17, 28, 4, 4, 10, 26, 30, 
    7, 10, 3, 2, 18, 22, 18, 10, 13, 11, 7, 5, 3, 25, 30, 
    1, 8, 20, 21, 36, 30, 17, 21, 25, 22, 22, 17, 17, 30, 27, 
    
    -- channel=449
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 11, 14, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 7, 4, 3, 2, 
    0, 0, 6, 7, 0, 0, 0, 1, 3, 0, 0, 0, 4, 6, 9, 
    2, 6, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 15, 18, 
    0, 0, 0, 18, 8, 0, 0, 0, 0, 0, 0, 0, 4, 6, 5, 
    0, 0, 0, 0, 20, 16, 7, 0, 0, 0, 0, 0, 0, 2, 10, 
    0, 0, 0, 25, 0, 28, 0, 3, 0, 0, 0, 0, 0, 5, 12, 
    6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 35, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 12, 14, 27, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 9, 26, 13, 
    0, 0, 0, 0, 0, 9, 8, 5, 0, 0, 0, 0, 3, 18, 22, 
    1, 0, 6, 20, 21, 15, 14, 16, 22, 17, 8, 3, 9, 27, 28, 
    
    -- channel=450
    19, 17, 26, 14, 21, 27, 15, 19, 17, 20, 19, 18, 23, 29, 25, 
    20, 17, 25, 20, 20, 33, 21, 23, 21, 25, 26, 25, 22, 17, 12, 
    22, 22, 9, 27, 32, 39, 42, 42, 33, 16, 13, 11, 9, 7, 8, 
    25, 28, 12, 30, 46, 49, 47, 40, 34, 37, 23, 11, 16, 9, 12, 
    31, 21, 0, 0, 39, 53, 32, 21, 36, 35, 40, 28, 20, 6, 6, 
    9, 4, 0, 0, 37, 61, 28, 27, 40, 33, 34, 49, 30, 6, 0, 
    9, 7, 4, 0, 33, 40, 19, 38, 42, 27, 30, 48, 24, 20, 2, 
    18, 14, 0, 0, 0, 43, 16, 37, 39, 20, 28, 39, 41, 32, 15, 
    17, 25, 13, 0, 0, 0, 23, 10, 44, 30, 31, 33, 48, 19, 0, 
    5, 0, 0, 0, 16, 0, 30, 5, 42, 37, 30, 25, 41, 12, 12, 
    0, 0, 0, 27, 26, 21, 32, 29, 35, 32, 27, 32, 34, 18, 0, 
    0, 0, 0, 0, 4, 49, 52, 7, 58, 53, 37, 25, 16, 27, 0, 
    11, 14, 19, 13, 0, 0, 32, 19, 39, 55, 25, 22, 10, 18, 18, 
    23, 15, 5, 4, 18, 19, 21, 23, 24, 37, 39, 30, 21, 13, 17, 
    3, 9, 18, 11, 22, 18, 8, 7, 12, 19, 28, 23, 13, 14, 11, 
    
    -- channel=451
    0, 2, 0, 7, 8, 0, 0, 3, 0, 0, 4, 3, 0, 0, 0, 
    0, 0, 1, 9, 5, 18, 8, 0, 2, 0, 0, 0, 0, 0, 0, 
    4, 3, 16, 15, 9, 5, 9, 3, 0, 0, 0, 0, 0, 5, 8, 
    0, 0, 0, 0, 4, 0, 0, 0, 3, 14, 4, 3, 0, 0, 0, 
    0, 0, 0, 2, 5, 0, 0, 0, 2, 2, 10, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 3, 6, 4, 0, 0, 
    11, 9, 0, 0, 9, 31, 15, 2, 0, 0, 2, 6, 10, 15, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 2, 11, 22, 
    0, 0, 26, 23, 22, 9, 5, 3, 0, 2, 0, 1, 8, 9, 1, 
    0, 13, 39, 39, 39, 42, 29, 30, 7, 12, 11, 2, 2, 0, 0, 
    81, 69, 27, 5, 2, 14, 0, 0, 10, 5, 0, 0, 3, 4, 0, 
    30, 21, 8, 0, 0, 0, 9, 1, 0, 0, 0, 6, 0, 1, 1, 
    1, 0, 16, 30, 18, 0, 0, 6, 11, 24, 33, 13, 13, 10, 8, 
    21, 28, 13, 2, 2, 0, 3, 7, 0, 0, 8, 19, 12, 6, 6, 
    
    -- channel=452
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 33, 3, 0, 0, 9, 9, 0, 0, 0, 0, 0, 1, 0, 1, 
    28, 21, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 3, 7, 0, 
    11, 8, 8, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 1, 0, 
    13, 20, 14, 17, 0, 3, 0, 2, 10, 0, 0, 0, 0, 0, 0, 
    29, 42, 53, 19, 36, 1, 15, 0, 1, 0, 0, 0, 0, 0, 0, 
    77, 79, 40, 9, 14, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 3, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=453
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 27, 29, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 26, 18, 11, 3, 0, 0, 
    0, 0, 8, 3, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 4, 
    39, 54, 40, 5, 0, 10, 23, 8, 0, 0, 0, 0, 1, 10, 16, 
    14, 0, 0, 6, 14, 13, 0, 0, 3, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 
    0, 3, 1, 13, 50, 27, 14, 5, 5, 4, 1, 0, 0, 0, 0, 
    10, 17, 47, 37, 30, 21, 13, 9, 0, 0, 5, 2, 0, 0, 0, 
    64, 48, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 7, 
    0, 0, 0, 7, 0, 0, 1, 0, 0, 0, 8, 5, 0, 0, 4, 
    0, 0, 0, 0, 17, 26, 0, 0, 7, 6, 13, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=454
    2, 1, 0, 2, 4, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 3, 0, 14, 12, 9, 15, 0, 0, 1, 4, 10, 14, 10, 
    0, 0, 0, 0, 2, 14, 18, 12, 14, 22, 17, 14, 7, 0, 0, 
    0, 1, 0, 15, 7, 14, 17, 24, 26, 6, 12, 7, 0, 0, 1, 
    20, 35, 42, 5, 17, 14, 32, 30, 23, 27, 21, 13, 10, 10, 14, 
    29, 22, 0, 7, 12, 31, 23, 15, 20, 24, 28, 17, 10, 7, 7, 
    8, 5, 0, 18, 8, 7, 16, 20, 24, 23, 22, 24, 14, 0, 0, 
    12, 16, 25, 0, 36, 26, 26, 26, 29, 25, 22, 27, 11, 4, 0, 
    24, 24, 30, 57, 30, 40, 10, 35, 23, 19, 24, 26, 19, 13, 0, 
    57, 67, 46, 14, 15, 10, 18, 22, 27, 21, 26, 27, 21, 0, 0, 
    33, 30, 0, 0, 4, 0, 9, 0, 23, 22, 19, 16, 15, 3, 7, 
    0, 0, 0, 11, 9, 3, 6, 21, 0, 7, 20, 23, 12, 5, 2, 
    0, 0, 0, 4, 4, 25, 20, 1, 23, 22, 32, 20, 14, 12, 0, 
    0, 9, 10, 0, 0, 0, 13, 10, 12, 14, 0, 8, 8, 0, 4, 
    3, 0, 0, 0, 0, 5, 8, 0, 2, 2, 7, 0, 0, 0, 0, 
    
    -- channel=455
    16, 16, 11, 20, 25, 21, 16, 14, 13, 15, 10, 8, 4, 0, 0, 
    16, 16, 18, 2, 36, 37, 36, 21, 8, 6, 0, 0, 0, 2, 5, 
    15, 16, 26, 18, 29, 31, 35, 27, 11, 17, 19, 20, 17, 20, 16, 
    12, 8, 0, 6, 26, 23, 24, 38, 31, 27, 29, 23, 8, 10, 9, 
    0, 6, 53, 13, 32, 35, 39, 39, 41, 36, 36, 32, 12, 9, 13, 
    27, 32, 49, 3, 17, 20, 38, 41, 39, 40, 43, 31, 19, 20, 21, 
    31, 27, 24, 4, 26, 45, 51, 38, 35, 38, 45, 33, 33, 27, 24, 
    17, 16, 37, 28, 19, 0, 33, 36, 43, 45, 42, 38, 35, 12, 4, 
    20, 4, 0, 12, 49, 41, 36, 38, 39, 42, 40, 43, 33, 28, 28, 
    18, 45, 71, 85, 52, 69, 33, 40, 38, 39, 43, 46, 34, 16, 4, 
    45, 64, 31, 36, 45, 51, 42, 38, 45, 45, 44, 37, 26, 14, 8, 
    80, 42, 26, 44, 28, 28, 22, 17, 25, 24, 33, 39, 23, 18, 14, 
    24, 25, 11, 18, 35, 34, 37, 26, 30, 26, 44, 44, 31, 16, 20, 
    10, 19, 35, 30, 7, 15, 12, 31, 29, 33, 44, 37, 38, 17, 16, 
    32, 22, 10, 8, 5, 22, 22, 16, 12, 16, 19, 26, 21, 11, 14, 
    
    -- channel=456
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    5, 6, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 
    1, 5, 17, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 6, 12, 10, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 15, 40, 31, 29, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 35, 26, 58, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 48, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 13, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=457
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 15, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=458
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 4, 0, 0, 0, 4, 0, 0, 0, 0, 6, 11, 
    
    -- channel=459
    4, 0, 6, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 22, 23, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 29, 19, 16, 6, 0, 0, 
    0, 6, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 4, 
    63, 78, 38, 0, 0, 0, 5, 0, 0, 0, 0, 0, 15, 24, 22, 
    52, 41, 20, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 18, 11, 
    24, 27, 39, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 51, 37, 40, 47, 26, 2, 0, 0, 0, 0, 0, 0, 0, 11, 
    56, 83, 121, 79, 67, 38, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    137, 121, 48, 40, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 19, 5, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 6, 15, 14, 5, 0, 0, 0, 0, 7, 0, 0, 0, 2, 
    5, 9, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=460
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 1, 0, 0, 7, 0, 0, 0, 0, 0, 1, 3, 4, 0, 
    0, 0, 0, 4, 0, 0, 1, 2, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 1, 5, 7, 4, 5, 0, 0, 0, 0, 0, 
    14, 14, 0, 0, 6, 15, 0, 0, 0, 1, 6, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 5, 8, 0, 0, 
    0, 0, 0, 0, 22, 15, 0, 0, 1, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 9, 3, 0, 0, 0, 0, 0, 0, 
    3, 7, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 5, 0, 0, 
    17, 7, 0, 0, 0, 0, 12, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 11, 0, 14, 6, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 9, 20, 0, 0, 0, 8, 0, 
    0, 3, 0, 0, 0, 0, 3, 0, 0, 14, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 17, 8, 0, 0, 0, 1, 11, 0, 0, 3, 0, 
    
    -- channel=461
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 2, 2, 3, 
    0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 8, 3, 9, 
    3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 17, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 24, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 17, 6, 
    0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 7, 11, 
    2, 11, 10, 0, 6, 0, 13, 0, 0, 0, 0, 0, 0, 0, 15, 
    6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 21, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 28, 18, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 24, 29, 
    0, 1, 0, 5, 16, 19, 4, 2, 0, 0, 0, 0, 0, 25, 27, 
    0, 9, 20, 22, 29, 25, 12, 19, 23, 18, 10, 11, 16, 30, 31, 
    
    -- channel=462
    2, 2, 6, 4, 15, 22, 9, 5, 2, 4, 3, 2, 2, 2, 0, 
    2, 2, 6, 10, 21, 35, 31, 22, 10, 6, 5, 2, 0, 0, 0, 
    4, 4, 6, 20, 30, 39, 46, 48, 27, 6, 9, 10, 11, 10, 12, 
    5, 5, 0, 12, 38, 40, 44, 50, 50, 37, 25, 21, 12, 8, 13, 
    0, 0, 0, 13, 34, 38, 34, 41, 54, 52, 49, 39, 20, 16, 19, 
    4, 7, 3, 6, 26, 31, 35, 43, 47, 51, 55, 52, 36, 29, 24, 
    10, 10, 6, 0, 21, 42, 40, 44, 41, 40, 49, 52, 43, 33, 22, 
    8, 6, 7, 13, 0, 11, 27, 45, 42, 35, 45, 50, 44, 27, 14, 
    8, 8, 0, 0, 16, 8, 29, 36, 43, 37, 41, 46, 43, 30, 28, 
    0, 0, 6, 13, 30, 24, 31, 39, 41, 37, 40, 43, 43, 31, 27, 
    4, 4, 11, 35, 41, 47, 45, 46, 44, 41, 43, 45, 40, 30, 21, 
    22, 24, 12, 11, 20, 43, 35, 17, 43, 44, 36, 36, 37, 37, 25, 
    14, 13, 12, 11, 8, 13, 36, 28, 30, 37, 27, 36, 39, 36, 36, 
    12, 11, 19, 27, 31, 25, 22, 30, 35, 39, 42, 39, 43, 39, 37, 
    18, 27, 31, 29, 31, 30, 29, 33, 33, 31, 32, 36, 38, 38, 36, 
    
    -- channel=463
    9, 7, 5, 6, 0, 0, 0, 1, 3, 1, 2, 1, 0, 0, 0, 
    9, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 9, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 13, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 3, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 12, 22, 24, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 29, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 36, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=464
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 11, 0, 4, 7, 1, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 
    0, 0, 48, 45, 7, 14, 6, 3, 0, 0, 1, 6, 0, 0, 0, 
    12, 46, 7, 0, 18, 10, 0, 11, 16, 5, 0, 0, 1, 0, 0, 
    11, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 8, 16, 0, 0, 0, 0, 3, 6, 7, 3, 2, 0, 
    0, 12, 15, 3, 0, 0, 0, 5, 1, 0, 2, 6, 9, 1, 2, 
    
    -- channel=465
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 8, 5, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 6, 12, 1, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 5, 0, 1, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 9, 10, 5, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 2, 3, 10, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 13, 23, 
    0, 0, 0, 3, 0, 9, 2, 7, 0, 0, 0, 0, 0, 6, 16, 
    0, 3, 0, 0, 0, 1, 0, 0, 3, 0, 0, 0, 10, 22, 10, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 1, 24, 17, 
    0, 0, 4, 24, 28, 7, 5, 7, 9, 11, 4, 0, 6, 29, 30, 
    11, 29, 28, 23, 28, 19, 12, 28, 28, 20, 25, 27, 28, 33, 32, 
    
    -- channel=466
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=467
    12, 11, 4, 10, 6, 10, 10, 8, 10, 7, 4, 3, 2, 0, 4, 
    12, 16, 8, 0, 10, 0, 9, 5, 2, 9, 10, 12, 13, 13, 14, 
    8, 12, 7, 0, 1, 0, 0, 0, 0, 18, 17, 15, 7, 8, 5, 
    8, 12, 34, 0, 0, 2, 0, 0, 0, 0, 6, 12, 8, 12, 10, 
    26, 34, 66, 7, 0, 0, 16, 11, 0, 0, 0, 5, 11, 14, 11, 
    27, 26, 73, 5, 10, 0, 6, 13, 7, 3, 0, 0, 0, 8, 9, 
    20, 22, 37, 56, 0, 0, 13, 5, 6, 12, 7, 0, 2, 0, 5, 
    23, 26, 33, 28, 66, 1, 22, 0, 4, 21, 10, 0, 4, 0, 11, 
    27, 34, 65, 41, 58, 53, 25, 7, 0, 18, 13, 8, 0, 0, 3, 
    57, 54, 35, 80, 16, 61, 0, 15, 1, 12, 15, 12, 0, 10, 0, 
    53, 61, 40, 15, 0, 2, 0, 0, 0, 4, 8, 10, 0, 15, 4, 
    22, 19, 29, 31, 22, 0, 1, 13, 0, 0, 9, 20, 4, 0, 17, 
    9, 8, 12, 13, 26, 15, 0, 14, 0, 0, 24, 15, 19, 0, 1, 
    8, 8, 6, 0, 0, 7, 0, 6, 0, 0, 0, 10, 11, 0, 0, 
    3, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=468
    8, 8, 15, 7, 15, 13, 12, 6, 6, 7, 7, 5, 6, 11, 7, 
    7, 4, 11, 21, 13, 31, 12, 19, 12, 8, 13, 12, 14, 14, 9, 
    9, 5, 5, 18, 18, 29, 33, 35, 30, 15, 13, 11, 12, 6, 6, 
    10, 11, 0, 31, 26, 30, 36, 39, 39, 28, 19, 12, 10, 8, 11, 
    19, 19, 0, 10, 33, 31, 24, 28, 33, 38, 38, 21, 20, 15, 17, 
    16, 11, 0, 18, 17, 46, 27, 20, 29, 34, 33, 39, 36, 16, 11, 
    9, 7, 0, 0, 30, 34, 13, 29, 29, 25, 24, 48, 27, 16, 2, 
    13, 15, 7, 0, 0, 46, 18, 37, 30, 16, 24, 36, 22, 24, 13, 
    19, 20, 4, 27, 0, 0, 7, 27, 33, 19, 24, 26, 35, 30, 8, 
    23, 19, 12, 0, 19, 0, 33, 14, 33, 27, 25, 22, 36, 15, 12, 
    6, 0, 0, 0, 25, 7, 28, 25, 29, 30, 22, 22, 34, 13, 15, 
    0, 0, 0, 0, 4, 32, 30, 15, 31, 35, 26, 19, 28, 32, 1, 
    4, 8, 8, 14, 0, 16, 29, 6, 31, 44, 16, 22, 14, 31, 14, 
    13, 17, 14, 11, 18, 10, 26, 21, 28, 40, 20, 20, 21, 22, 30, 
    12, 11, 15, 17, 32, 19, 19, 17, 23, 21, 33, 27, 16, 26, 18, 
    
    -- channel=469
    0, 0, 6, 4, 0, 0, 0, 4, 5, 5, 8, 9, 11, 15, 13, 
    0, 0, 6, 0, 0, 0, 0, 0, 6, 7, 8, 9, 14, 19, 18, 
    0, 1, 5, 0, 0, 0, 0, 0, 0, 9, 8, 10, 13, 15, 15, 
    1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 12, 15, 
    2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 17, 19, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 19, 
    0, 0, 0, 2, 0, 3, 2, 0, 0, 0, 0, 0, 0, 22, 21, 
    1, 5, 6, 10, 13, 11, 7, 0, 0, 0, 0, 0, 0, 20, 27, 
    13, 15, 15, 21, 31, 23, 10, 18, 23, 15, 11, 6, 10, 28, 32, 
    
    -- channel=470
    0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 1, 6, 13, 
    0, 0, 0, 0, 0, 0, 0, 6, 4, 7, 18, 21, 15, 9, 5, 
    0, 0, 0, 0, 0, 1, 0, 9, 7, 4, 0, 0, 0, 0, 0, 
    1, 8, 31, 8, 6, 17, 15, 0, 4, 0, 0, 2, 4, 3, 4, 
    31, 20, 0, 0, 0, 0, 1, 0, 2, 4, 1, 0, 7, 10, 4, 
    0, 0, 0, 0, 13, 16, 1, 0, 4, 0, 1, 4, 3, 0, 0, 
    0, 0, 1, 27, 0, 0, 0, 1, 5, 3, 0, 0, 0, 0, 0, 
    6, 9, 0, 0, 18, 35, 7, 0, 0, 0, 0, 2, 2, 9, 12, 
    6, 27, 46, 25, 0, 9, 0, 0, 0, 0, 3, 2, 1, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 5, 4, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 7, 5, 7, 3, 
    0, 0, 0, 0, 4, 0, 8, 8, 9, 10, 3, 4, 1, 0, 7, 
    0, 0, 6, 0, 0, 0, 0, 4, 0, 1, 0, 0, 2, 3, 0, 
    6, 0, 0, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    
    -- channel=471
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 18, 29, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 15, 16, 23, 32, 27, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 23, 33, 33, 28, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 11, 16, 18, 33, 35, 20, 3, 0, 0, 
    0, 0, 0, 0, 4, 5, 12, 20, 6, 14, 29, 28, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 21, 3, 6, 25, 27, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 7, 5, 16, 23, 12, 0, 4, 
    0, 0, 0, 0, 0, 0, 3, 17, 9, 6, 13, 23, 16, 5, 2, 
    0, 0, 0, 3, 6, 19, 10, 17, 14, 12, 17, 23, 16, 0, 2, 
    0, 0, 0, 0, 1, 19, 0, 0, 16, 11, 0, 8, 19, 7, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 7, 0, 0, 8, 6, 14, 2, 
    0, 0, 0, 3, 7, 0, 3, 13, 18, 15, 9, 10, 13, 16, 15, 
    0, 5, 11, 9, 8, 2, 5, 15, 19, 14, 20, 22, 20, 17, 12, 
    
    -- channel=472
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 2, 3, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 8, 0, 0, 0, 2, 21, 1, 0, 0, 0, 0, 
    0, 17, 8, 0, 0, 0, 0, 0, 0, 0, 14, 14, 4, 7, 1, 
    
    -- channel=473
    0, 4, 0, 8, 0, 0, 12, 1, 6, 6, 7, 10, 6, 0, 2, 
    0, 4, 0, 0, 7, 0, 0, 3, 7, 0, 0, 0, 0, 0, 6, 
    1, 0, 25, 0, 2, 0, 0, 0, 0, 0, 0, 4, 9, 13, 15, 
    0, 0, 3, 19, 0, 0, 0, 0, 0, 0, 0, 11, 0, 9, 5, 
    0, 0, 41, 23, 0, 0, 0, 11, 0, 0, 0, 0, 0, 2, 5, 
    0, 0, 33, 34, 0, 0, 9, 0, 0, 0, 2, 0, 0, 2, 15, 
    0, 0, 0, 39, 14, 0, 1, 0, 0, 2, 5, 0, 0, 3, 24, 
    0, 0, 11, 0, 31, 0, 8, 0, 0, 4, 4, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 34, 0, 19, 0, 0, 0, 3, 0, 7, 29, 
    0, 0, 37, 32, 4, 31, 0, 13, 0, 0, 0, 8, 0, 14, 10, 
    0, 24, 78, 13, 4, 10, 0, 0, 0, 0, 1, 0, 0, 0, 30, 
    40, 16, 2, 13, 31, 0, 0, 29, 0, 0, 0, 0, 14, 0, 21, 
    5, 3, 0, 0, 10, 11, 0, 0, 0, 0, 0, 5, 7, 11, 0, 
    0, 0, 16, 21, 1, 0, 6, 9, 1, 0, 0, 0, 11, 8, 9, 
    21, 17, 3, 11, 0, 2, 10, 11, 12, 6, 3, 4, 7, 10, 15, 
    
    -- channel=474
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=475
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 1, 0, 0, 3, 0, 0, 0, 0, 2, 7, 11, 11, 2, 
    0, 0, 0, 0, 0, 0, 2, 4, 10, 8, 2, 1, 0, 0, 0, 
    0, 1, 0, 3, 0, 5, 7, 11, 0, 7, 0, 0, 0, 0, 0, 
    26, 28, 0, 0, 1, 28, 7, 0, 1, 0, 6, 0, 7, 2, 3, 
    6, 0, 0, 0, 3, 39, 0, 0, 4, 0, 0, 8, 11, 0, 0, 
    0, 0, 0, 0, 12, 10, 0, 0, 10, 0, 0, 9, 0, 1, 0, 
    0, 4, 0, 0, 0, 30, 0, 9, 9, 0, 0, 0, 4, 1, 0, 
    8, 18, 19, 0, 0, 0, 15, 0, 4, 0, 0, 0, 12, 0, 0, 
    31, 12, 0, 0, 0, 0, 14, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 23, 0, 10, 7, 5, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 9, 22, 0, 0, 0, 3, 11, 
    0, 1, 0, 0, 0, 7, 0, 1, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 11, 12, 0, 0, 0, 2, 6, 0, 0, 1, 0, 
    
    -- channel=476
    0, 0, 0, 0, 2, 15, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 10, 1, 30, 7, 0, 4, 0, 0, 0, 0, 0, 
    0, 4, 0, 8, 9, 8, 6, 10, 12, 5, 4, 4, 0, 1, 2, 
    0, 1, 12, 0, 8, 5, 1, 4, 0, 10, 15, 6, 5, 0, 5, 
    0, 0, 18, 0, 0, 23, 15, 2, 12, 7, 9, 22, 9, 5, 3, 
    0, 0, 51, 0, 16, 0, 0, 19, 14, 6, 8, 7, 0, 9, 2, 
    1, 4, 22, 3, 0, 8, 28, 15, 12, 7, 15, 0, 4, 8, 3, 
    4, 2, 0, 35, 32, 0, 1, 2, 14, 17, 13, 1, 18, 0, 4, 
    2, 4, 19, 0, 52, 9, 37, 0, 6, 17, 14, 11, 6, 0, 6, 
    0, 0, 0, 77, 6, 65, 0, 16, 6, 11, 14, 12, 0, 1, 5, 
    6, 12, 0, 11, 1, 29, 5, 13, 12, 8, 15, 13, 0, 21, 0, 
    14, 19, 25, 23, 0, 0, 14, 0, 0, 4, 9, 13, 0, 2, 14, 
    3, 3, 4, 1, 26, 0, 0, 26, 0, 1, 15, 9, 22, 0, 22, 
    1, 0, 0, 4, 4, 17, 0, 1, 0, 0, 17, 14, 4, 7, 0, 
    0, 4, 6, 0, 0, 7, 1, 6, 0, 1, 0, 0, 8, 0, 2, 
    
    -- channel=477
    0, 3, 0, 2, 0, 0, 9, 2, 7, 4, 5, 7, 6, 1, 10, 
    0, 6, 0, 0, 1, 0, 2, 5, 5, 4, 9, 9, 9, 10, 15, 
    0, 1, 11, 0, 0, 0, 0, 0, 0, 4, 9, 10, 9, 11, 14, 
    0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 15, 14, 
    0, 1, 53, 26, 0, 0, 0, 14, 0, 0, 0, 0, 7, 17, 16, 
    0, 0, 60, 29, 1, 0, 0, 6, 0, 3, 0, 0, 0, 12, 18, 
    0, 1, 14, 74, 0, 0, 5, 0, 0, 8, 7, 0, 3, 0, 19, 
    0, 0, 12, 14, 73, 0, 17, 0, 0, 11, 8, 0, 0, 2, 13, 
    0, 0, 18, 37, 24, 49, 1, 13, 0, 3, 5, 6, 0, 6, 25, 
    1, 3, 10, 59, 0, 50, 0, 20, 0, 0, 0, 10, 0, 27, 19, 
    3, 24, 71, 0, 0, 0, 0, 0, 0, 0, 2, 6, 3, 18, 31, 
    7, 5, 20, 20, 29, 0, 0, 26, 0, 0, 0, 13, 20, 0, 41, 
    0, 0, 0, 2, 22, 16, 0, 12, 0, 0, 1, 7, 29, 8, 6, 
    0, 0, 6, 12, 3, 7, 4, 7, 0, 0, 0, 0, 16, 16, 0, 
    10, 10, 9, 16, 0, 0, 12, 21, 13, 8, 0, 0, 16, 13, 13, 
    
    -- channel=478
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=479
    15, 15, 10, 16, 3, 0, 8, 13, 14, 11, 12, 14, 12, 10, 14, 
    15, 17, 10, 9, 0, 0, 0, 0, 7, 12, 10, 10, 9, 10, 13, 
    13, 14, 12, 0, 0, 0, 0, 0, 0, 3, 7, 7, 9, 13, 13, 
    11, 12, 27, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 14, 8, 
    14, 13, 27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 
    16, 19, 49, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 
    21, 23, 30, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    17, 18, 19, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    14, 20, 35, 21, 16, 16, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    24, 24, 29, 46, 4, 26, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    40, 45, 56, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    34, 41, 31, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    19, 15, 18, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 4, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=480
    0, 0, 12, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 5, 1, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 3, 6, 10, 18, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 5, 2, 4, 9, 5, 21, 8, 0, 0, 0, 0, 
    9, 5, 0, 0, 4, 32, 0, 0, 0, 2, 16, 5, 8, 0, 0, 
    6, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 21, 24, 0, 0, 
    2, 0, 0, 0, 6, 35, 0, 2, 7, 0, 0, 23, 4, 12, 0, 
    7, 6, 0, 0, 0, 17, 0, 9, 10, 0, 0, 0, 7, 9, 0, 
    12, 19, 0, 0, 0, 0, 2, 0, 10, 0, 0, 0, 16, 3, 0, 
    8, 2, 0, 0, 8, 0, 18, 0, 6, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 5, 0, 6, 5, 3, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 26, 0, 17, 18, 2, 0, 0, 28, 0, 
    0, 1, 0, 0, 0, 0, 17, 0, 8, 36, 0, 0, 0, 8, 10, 
    2, 3, 0, 0, 7, 1, 0, 0, 0, 20, 15, 0, 0, 1, 14, 
    0, 0, 1, 0, 21, 11, 0, 0, 0, 0, 12, 7, 0, 7, 1, 
    
    -- channel=481
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=482
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=483
    12, 13, 5, 11, 9, 7, 12, 10, 9, 9, 9, 10, 6, 1, 2, 
    12, 14, 7, 6, 8, 0, 8, 7, 5, 4, 1, 0, 0, 0, 0, 
    12, 12, 13, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 
    9, 7, 14, 0, 1, 0, 0, 0, 0, 0, 3, 6, 0, 2, 0, 
    0, 0, 26, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 14, 41, 7, 0, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 
    15, 16, 19, 30, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 8, 15, 5, 22, 0, 2, 0, 0, 10, 1, 0, 0, 0, 0, 
    6, 2, 6, 14, 12, 18, 0, 0, 0, 10, 3, 1, 0, 0, 0, 
    0, 8, 27, 51, 13, 29, 0, 8, 2, 7, 4, 7, 0, 0, 0, 
    26, 39, 61, 29, 13, 18, 0, 0, 1, 3, 5, 5, 0, 0, 0, 
    48, 44, 22, 16, 21, 0, 0, 9, 0, 0, 0, 4, 0, 0, 0, 
    21, 17, 13, 5, 7, 1, 0, 7, 0, 0, 9, 8, 0, 0, 0, 
    6, 2, 7, 6, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=484
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 39, 23, 15, 22, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    61, 63, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 12, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    6, 18, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=485
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    19, 22, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 13, 
    22, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 9, 
    11, 15, 19, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 19, 17, 7, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    34, 52, 60, 37, 14, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 62, 17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 35, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    9, 5, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 
    0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    
    -- channel=486
    4, 4, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 37, 32, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 30, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 32, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=487
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=488
    16, 16, 12, 12, 17, 27, 23, 20, 18, 17, 19, 20, 20, 18, 21, 
    16, 17, 11, 21, 24, 29, 39, 36, 25, 20, 22, 22, 24, 20, 19, 
    16, 17, 14, 17, 34, 40, 40, 43, 39, 23, 22, 18, 15, 12, 13, 
    18, 18, 24, 21, 41, 41, 41, 42, 36, 29, 26, 25, 14, 14, 18, 
    20, 20, 19, 38, 38, 36, 42, 46, 45, 44, 39, 39, 21, 16, 17, 
    7, 5, 25, 31, 38, 29, 39, 46, 42, 45, 45, 42, 22, 11, 10, 
    3, 4, 16, 27, 9, 23, 41, 46, 40, 42, 46, 43, 30, 10, 10, 
    10, 8, 6, 32, 42, 19, 31, 38, 40, 45, 49, 45, 38, 25, 17, 
    9, 7, 16, 17, 22, 15, 20, 40, 39, 44, 48, 51, 44, 28, 12, 
    6, 0, 0, 19, 18, 29, 22, 43, 41, 43, 45, 53, 44, 28, 12, 
    0, 0, 16, 7, 18, 34, 29, 32, 38, 41, 39, 47, 41, 26, 17, 
    0, 0, 12, 24, 29, 37, 35, 27, 24, 38, 36, 42, 36, 14, 20, 
    6, 9, 10, 12, 28, 29, 23, 37, 37, 40, 35, 42, 40, 14, 16, 
    14, 12, 13, 12, 12, 15, 23, 24, 29, 21, 26, 39, 35, 20, 8, 
    11, 10, 13, 15, 10, 9, 16, 20, 17, 18, 17, 18, 22, 14, 9, 
    
    -- channel=489
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 29, 30, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 25, 18, 13, 2, 0, 0, 
    0, 0, 14, 0, 0, 1, 6, 4, 0, 0, 0, 0, 0, 0, 4, 
    42, 56, 49, 0, 0, 8, 23, 9, 2, 0, 0, 0, 4, 12, 17, 
    12, 0, 4, 0, 15, 14, 0, 0, 6, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 5, 6, 2, 0, 0, 0, 0, 
    0, 4, 3, 8, 52, 29, 17, 4, 5, 6, 3, 0, 0, 0, 3, 
    8, 15, 53, 45, 34, 29, 13, 7, 0, 0, 7, 5, 0, 0, 0, 
    67, 46, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 
    0, 0, 0, 2, 0, 0, 6, 0, 0, 0, 8, 9, 0, 0, 7, 
    0, 0, 0, 0, 16, 23, 0, 0, 4, 5, 15, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=490
    22, 21, 24, 25, 37, 38, 34, 24, 20, 20, 16, 13, 11, 13, 11, 
    21, 21, 26, 22, 45, 52, 48, 46, 27, 22, 25, 28, 31, 34, 31, 
    20, 19, 21, 29, 42, 55, 61, 60, 52, 48, 42, 43, 35, 29, 25, 
    22, 23, 17, 41, 45, 53, 60, 70, 70, 52, 51, 42, 31, 30, 34, 
    40, 51, 52, 33, 49, 56, 66, 68, 72, 73, 70, 56, 48, 49, 53, 
    51, 47, 23, 29, 41, 66, 58, 57, 65, 70, 74, 62, 58, 55, 49, 
    36, 34, 30, 29, 42, 49, 55, 62, 65, 63, 67, 69, 59, 47, 30, 
    39, 45, 51, 38, 46, 55, 59, 69, 68, 60, 64, 68, 54, 42, 35, 
    50, 53, 55, 70, 61, 62, 56, 70, 63, 56, 63, 64, 59, 50, 40, 
    75, 82, 68, 45, 56, 46, 63, 62, 63, 59, 64, 64, 57, 36, 36, 
    61, 57, 21, 25, 45, 45, 55, 46, 64, 62, 61, 57, 52, 47, 46, 
    32, 7, 16, 35, 37, 41, 45, 45, 44, 51, 59, 58, 52, 57, 46, 
    19, 25, 24, 37, 37, 49, 55, 40, 57, 60, 61, 58, 57, 59, 49, 
    27, 40, 43, 35, 32, 42, 48, 48, 50, 51, 42, 47, 50, 49, 54, 
    36, 31, 33, 41, 48, 52, 50, 44, 49, 47, 48, 45, 41, 50, 48, 
    
    -- channel=491
    6, 10, 0, 5, 0, 4, 20, 7, 13, 10, 11, 14, 12, 6, 16, 
    7, 13, 0, 5, 8, 0, 6, 17, 13, 8, 15, 15, 15, 14, 18, 
    5, 6, 18, 0, 8, 4, 2, 0, 0, 9, 11, 12, 9, 10, 12, 
    5, 5, 41, 13, 2, 8, 5, 0, 3, 0, 0, 20, 6, 16, 12, 
    5, 7, 62, 40, 4, 0, 9, 28, 6, 6, 0, 3, 4, 13, 12, 
    0, 1, 59, 47, 9, 0, 18, 19, 5, 12, 12, 0, 0, 2, 11, 
    0, 1, 12, 94, 0, 0, 12, 5, 0, 21, 17, 0, 6, 0, 14, 
    0, 0, 15, 4, 83, 4, 28, 0, 0, 25, 21, 10, 0, 4, 12, 
    0, 0, 19, 68, 18, 60, 0, 28, 0, 16, 19, 22, 0, 10, 15, 
    3, 3, 9, 53, 0, 42, 0, 33, 0, 7, 14, 28, 6, 29, 6, 
    0, 22, 91, 4, 0, 2, 0, 0, 0, 4, 10, 21, 14, 8, 26, 
    2, 2, 19, 19, 48, 0, 0, 44, 0, 0, 2, 24, 25, 0, 36, 
    1, 0, 2, 3, 20, 24, 0, 19, 0, 0, 14, 19, 30, 3, 0, 
    2, 1, 6, 7, 0, 0, 10, 8, 2, 0, 0, 11, 20, 5, 0, 
    8, 3, 0, 8, 0, 0, 11, 13, 6, 4, 0, 0, 9, 0, 0, 
    
    -- channel=492
    27, 26, 29, 25, 28, 19, 17, 19, 20, 23, 20, 20, 19, 20, 14, 
    27, 24, 28, 22, 24, 30, 17, 15, 12, 17, 11, 10, 10, 11, 8, 
    28, 25, 21, 33, 21, 21, 21, 15, 10, 14, 13, 10, 9, 9, 7, 
    25, 24, 0, 24, 27, 19, 15, 12, 13, 18, 20, 3, 5, 6, 2, 
    18, 19, 3, 4, 28, 32, 18, 8, 9, 15, 19, 7, 1, 0, 0, 
    24, 24, 0, 3, 18, 37, 21, 15, 13, 9, 10, 18, 4, 0, 0, 
    25, 21, 8, 0, 27, 40, 19, 18, 18, 11, 9, 23, 6, 2, 0, 
    24, 19, 17, 0, 0, 19, 6, 18, 24, 15, 11, 18, 14, 7, 0, 
    22, 16, 0, 3, 4, 0, 8, 7, 28, 20, 15, 13, 21, 10, 0, 
    17, 23, 24, 0, 22, 0, 20, 2, 28, 26, 19, 13, 21, 0, 0, 
    22, 16, 0, 19, 34, 17, 23, 15, 26, 23, 15, 11, 9, 0, 0, 
    33, 20, 7, 11, 10, 27, 21, 7, 32, 25, 19, 10, 0, 0, 0, 
    24, 27, 17, 16, 0, 12, 26, 6, 29, 35, 24, 17, 0, 0, 0, 
    17, 19, 16, 5, 0, 0, 6, 10, 16, 33, 32, 21, 2, 0, 0, 
    12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 10, 6, 0, 0, 0, 
    
    -- channel=493
    2, 7, 0, 3, 0, 0, 13, 4, 8, 4, 8, 10, 7, 0, 8, 
    2, 7, 0, 12, 2, 0, 3, 7, 10, 0, 4, 2, 0, 0, 7, 
    2, 1, 15, 0, 4, 0, 0, 0, 0, 0, 1, 2, 7, 7, 11, 
    0, 0, 23, 9, 0, 0, 0, 0, 0, 0, 0, 14, 2, 10, 7, 
    0, 0, 30, 49, 0, 0, 0, 20, 0, 0, 0, 0, 0, 7, 5, 
    0, 0, 34, 55, 0, 0, 10, 16, 0, 4, 4, 0, 0, 0, 9, 
    0, 2, 2, 87, 0, 0, 12, 0, 0, 12, 7, 0, 1, 0, 15, 
    0, 0, 8, 3, 55, 0, 13, 0, 0, 15, 13, 3, 0, 0, 6, 
    0, 0, 0, 56, 0, 43, 0, 23, 0, 7, 10, 9, 0, 8, 19, 
    0, 0, 16, 53, 0, 19, 0, 34, 0, 0, 4, 18, 0, 25, 6, 
    0, 20, 113, 5, 6, 6, 6, 1, 0, 0, 7, 13, 6, 0, 19, 
    26, 22, 38, 11, 42, 0, 0, 40, 0, 0, 0, 10, 20, 0, 31, 
    12, 3, 2, 2, 15, 18, 0, 13, 0, 0, 0, 10, 22, 1, 0, 
    0, 0, 7, 15, 4, 0, 7, 1, 5, 0, 0, 9, 11, 6, 0, 
    11, 11, 4, 9, 0, 0, 12, 14, 7, 1, 0, 0, 10, 2, 1, 
    
    -- channel=494
    0, 0, 0, 0, 1, 13, 4, 0, 1, 1, 2, 2, 4, 2, 4, 
    0, 0, 0, 2, 10, 17, 22, 19, 7, 3, 5, 2, 0, 0, 0, 
    0, 1, 0, 7, 24, 34, 38, 37, 19, 0, 0, 0, 0, 0, 0, 
    2, 3, 6, 8, 39, 43, 41, 37, 31, 16, 7, 7, 0, 0, 0, 
    0, 0, 0, 17, 33, 30, 31, 38, 41, 39, 31, 25, 2, 0, 0, 
    0, 0, 2, 12, 30, 23, 31, 42, 41, 43, 44, 41, 10, 0, 0, 
    0, 0, 0, 7, 3, 19, 34, 40, 34, 36, 42, 40, 21, 0, 0, 
    0, 0, 0, 0, 10, 6, 21, 30, 33, 36, 43, 45, 34, 14, 0, 
    0, 0, 0, 0, 0, 0, 4, 25, 36, 38, 42, 47, 39, 17, 0, 
    0, 0, 0, 0, 0, 7, 4, 30, 38, 38, 38, 47, 43, 21, 0, 
    0, 0, 0, 8, 18, 24, 29, 29, 33, 35, 34, 46, 38, 9, 0, 
    0, 0, 0, 5, 23, 43, 30, 19, 31, 39, 29, 36, 26, 0, 0, 
    0, 0, 0, 0, 0, 9, 13, 24, 26, 33, 25, 30, 28, 1, 0, 
    0, 0, 0, 0, 0, 0, 10, 16, 23, 23, 25, 37, 31, 7, 0, 
    0, 0, 2, 0, 0, 0, 2, 5, 3, 7, 11, 13, 13, 0, 0, 
    
    -- channel=495
    17, 20, 5, 20, 23, 24, 20, 18, 19, 17, 17, 19, 14, 4, 8, 
    17, 22, 9, 19, 31, 20, 42, 23, 15, 15, 7, 2, 0, 0, 7, 
    17, 20, 27, 21, 36, 28, 29, 23, 3, 7, 16, 15, 16, 22, 24, 
    14, 10, 31, 2, 30, 24, 22, 24, 20, 11, 23, 31, 12, 18, 16, 
    0, 0, 49, 55, 19, 13, 29, 47, 34, 28, 21, 29, 9, 12, 11, 
    7, 18, 88, 41, 25, 0, 37, 55, 33, 39, 36, 20, 5, 16, 21, 
    23, 26, 37, 70, 0, 20, 57, 36, 23, 43, 45, 15, 28, 15, 34, 
    13, 8, 25, 45, 66, 0, 35, 21, 23, 53, 50, 31, 28, 11, 11, 
    6, 0, 8, 20, 47, 48, 28, 41, 23, 49, 46, 44, 18, 20, 36, 
    0, 0, 42, 123, 36, 87, 14, 61, 23, 36, 42, 54, 25, 39, 13, 
    28, 55, 118, 51, 40, 65, 36, 43, 31, 36, 47, 48, 24, 21, 15, 
    81, 75, 63, 51, 60, 28, 5, 39, 15, 20, 25, 44, 32, 0, 40, 
    34, 28, 22, 15, 42, 31, 15, 44, 17, 5, 34, 49, 49, 4, 15, 
    15, 10, 25, 36, 19, 15, 12, 22, 23, 11, 34, 48, 43, 22, 0, 
    28, 31, 20, 16, 0, 5, 22, 29, 13, 11, 4, 18, 33, 11, 10, 
    
    -- channel=496
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 26, 28, 24, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 7, 3, 0, 0, 0, 
    0, 1, 27, 4, 0, 12, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 50, 21, 0, 0, 0, 16, 6, 0, 0, 0, 0, 0, 9, 9, 
    0, 0, 0, 4, 19, 18, 0, 0, 6, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 43, 46, 15, 1, 0, 0, 0, 0, 0, 0, 5, 
    4, 23, 61, 48, 15, 22, 4, 1, 0, 0, 6, 3, 0, 0, 0, 
    55, 17, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 8, 2, 
    0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 7, 7, 0, 0, 5, 
    0, 0, 0, 0, 0, 6, 0, 0, 1, 5, 5, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=497
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 20, 23, 22, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 16, 5, 2, 0, 0, 0, 
    0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    45, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 6, 
    12, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 13, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    15, 33, 52, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=498
    2, 1, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 7, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 
    0, 5, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 
    19, 23, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 
    23, 24, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 
    14, 18, 21, 25, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 21, 30, 15, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    34, 44, 53, 47, 14, 24, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    58, 61, 40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    52, 44, 26, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    15, 10, 10, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    2, 1, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=499
    26, 24, 21, 19, 22, 28, 27, 19, 20, 17, 12, 9, 6, 5, 6, 
    25, 24, 22, 8, 27, 26, 30, 30, 17, 13, 15, 19, 24, 26, 22, 
    21, 20, 15, 10, 18, 27, 25, 26, 33, 42, 32, 28, 20, 12, 4, 
    21, 22, 18, 12, 24, 30, 29, 28, 29, 20, 30, 23, 12, 12, 9, 
    44, 60, 67, 16, 32, 36, 51, 39, 33, 33, 30, 31, 19, 14, 17, 
    51, 46, 37, 15, 30, 42, 42, 37, 38, 33, 36, 30, 17, 11, 11, 
    33, 30, 31, 39, 14, 21, 35, 37, 43, 39, 33, 36, 29, 9, 3, 
    37, 41, 46, 25, 52, 31, 38, 35, 50, 47, 38, 39, 30, 14, 9, 
    47, 49, 64, 76, 62, 59, 28, 41, 45, 44, 44, 42, 36, 25, 0, 
    88, 94, 64, 58, 36, 37, 26, 37, 47, 46, 47, 46, 37, 6, 0, 
    69, 64, 18, 0, 22, 13, 30, 11, 40, 42, 33, 35, 28, 12, 0, 
    29, 0, 15, 33, 28, 18, 32, 30, 13, 28, 42, 40, 16, 2, 6, 
    11, 17, 12, 22, 27, 39, 23, 24, 36, 44, 58, 41, 26, 3, 0, 
    13, 23, 19, 0, 0, 4, 15, 16, 20, 23, 18, 32, 22, 0, 0, 
    10, 0, 0, 0, 0, 3, 11, 0, 0, 0, 3, 0, 0, 0, 0, 
    
    -- channel=500
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 
    0, 0, 0, 6, 14, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 
    0, 14, 15, 13, 12, 0, 0, 11, 10, 2, 0, 0, 7, 16, 18, 
    
    -- channel=501
    0, 0, 7, 6, 11, 5, 0, 3, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 5, 11, 1, 23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 4, 4, 21, 13, 9, 15, 12, 0, 0, 0, 0, 0, 0, 2, 
    1, 0, 0, 0, 13, 1, 0, 1, 10, 29, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 12, 0, 0, 2, 6, 19, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 19, 6, 0, 0, 
    15, 13, 0, 0, 10, 41, 8, 5, 1, 0, 0, 13, 5, 19, 10, 
    1, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 3, 13, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 10, 0, 9, 
    0, 0, 1, 0, 28, 0, 14, 0, 9, 3, 0, 0, 6, 0, 0, 
    0, 0, 8, 65, 45, 52, 26, 30, 12, 9, 9, 0, 0, 0, 0, 
    72, 84, 14, 0, 0, 22, 8, 0, 36, 20, 0, 0, 0, 10, 0, 
    35, 27, 19, 0, 0, 0, 17, 0, 0, 9, 0, 0, 0, 0, 7, 
    9, 0, 7, 24, 29, 1, 0, 1, 8, 29, 50, 11, 0, 3, 11, 
    9, 27, 19, 0, 4, 6, 0, 0, 0, 0, 11, 19, 8, 2, 4, 
    
    -- channel=502
    14, 13, 9, 14, 14, 14, 15, 5, 7, 5, 0, 0, 0, 0, 0, 
    13, 13, 10, 2, 18, 15, 17, 13, 1, 0, 0, 0, 5, 8, 8, 
    9, 9, 12, 0, 6, 9, 12, 11, 8, 20, 21, 19, 14, 10, 3, 
    7, 7, 4, 0, 4, 7, 9, 17, 16, 7, 17, 17, 4, 8, 4, 
    20, 36, 58, 11, 11, 12, 29, 28, 19, 18, 14, 17, 12, 12, 14, 
    45, 45, 47, 13, 10, 15, 28, 22, 19, 22, 20, 13, 12, 14, 14, 
    36, 34, 34, 31, 6, 14, 28, 21, 20, 24, 21, 15, 18, 6, 8, 
    32, 35, 47, 32, 43, 9, 29, 21, 28, 33, 24, 18, 13, 5, 4, 
    41, 41, 53, 69, 56, 51, 22, 33, 23, 29, 26, 24, 15, 19, 7, 
    75, 92, 89, 76, 46, 49, 23, 30, 25, 28, 30, 29, 18, 6, 0, 
    83, 87, 54, 15, 22, 17, 17, 13, 26, 28, 25, 21, 16, 5, 2, 
    62, 28, 23, 34, 23, 5, 9, 16, 0, 9, 21, 29, 14, 1, 8, 
    16, 19, 10, 18, 24, 28, 17, 11, 13, 18, 37, 31, 20, 2, 0, 
    8, 16, 21, 10, 0, 0, 6, 15, 12, 13, 12, 21, 20, 0, 0, 
    15, 0, 0, 0, 0, 2, 9, 1, 0, 0, 1, 4, 1, 0, 0, 
    
    -- channel=503
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 
    0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 1, 17, 16, 
    0, 8, 12, 14, 14, 3, 3, 15, 16, 9, 7, 8, 14, 23, 22, 
    
    -- channel=504
    9, 12, 1, 10, 13, 21, 24, 12, 15, 13, 13, 14, 12, 7, 13, 
    9, 14, 7, 10, 26, 18, 32, 31, 19, 12, 17, 16, 15, 14, 19, 
    9, 9, 19, 12, 29, 34, 37, 35, 21, 18, 21, 21, 19, 19, 21, 
    10, 8, 31, 22, 31, 37, 39, 40, 42, 16, 19, 31, 17, 20, 22, 
    4, 7, 52, 50, 31, 12, 38, 58, 48, 46, 32, 33, 19, 26, 28, 
    8, 11, 49, 48, 30, 8, 41, 51, 43, 52, 55, 31, 21, 27, 31, 
    8, 10, 13, 82, 14, 8, 48, 40, 33, 50, 54, 33, 37, 18, 29, 
    6, 7, 22, 15, 74, 13, 47, 35, 32, 51, 54, 49, 32, 22, 21, 
    7, 3, 15, 55, 35, 65, 21, 56, 30, 43, 51, 54, 29, 32, 37, 
    5, 11, 22, 67, 11, 54, 12, 63, 34, 36, 45, 59, 40, 45, 27, 
    8, 27, 83, 17, 27, 33, 36, 31, 35, 38, 45, 53, 42, 31, 38, 
    23, 13, 31, 32, 55, 31, 13, 55, 19, 25, 32, 49, 49, 13, 52, 
    12, 11, 8, 14, 31, 39, 19, 39, 25, 14, 37, 42, 57, 32, 20, 
    10, 13, 23, 28, 19, 20, 31, 32, 35, 24, 16, 40, 45, 35, 22, 
    23, 24, 23, 30, 17, 18, 35, 37, 35, 31, 24, 28, 38, 30, 30, 
    
    -- channel=505
    34, 30, 32, 34, 30, 23, 23, 23, 21, 20, 16, 12, 7, 5, 1, 
    33, 29, 30, 20, 22, 22, 16, 12, 12, 14, 8, 7, 6, 8, 8, 
    31, 29, 25, 14, 10, 3, 5, 3, 6, 20, 19, 20, 17, 17, 12, 
    26, 25, 8, 5, 4, 0, 0, 0, 2, 20, 24, 16, 15, 14, 5, 
    31, 39, 38, 0, 5, 16, 13, 0, 0, 0, 9, 9, 12, 8, 4, 
    58, 63, 48, 0, 5, 21, 22, 7, 3, 0, 0, 6, 9, 8, 8, 
    60, 59, 54, 3, 20, 27, 18, 11, 13, 5, 0, 4, 4, 11, 11, 
    54, 54, 56, 37, 4, 11, 12, 9, 21, 16, 2, 0, 8, 7, 8, 
    57, 60, 60, 43, 47, 26, 25, 8, 23, 21, 8, 2, 9, 8, 1, 
    78, 93, 101, 71, 62, 41, 30, 9, 22, 24, 17, 6, 6, 0, 0, 
    110, 106, 51, 56, 37, 29, 16, 13, 21, 21, 15, 6, 1, 0, 0, 
    99, 80, 42, 36, 14, 6, 15, 1, 15, 13, 15, 11, 0, 1, 0, 
    49, 45, 38, 32, 22, 10, 19, 7, 12, 20, 30, 19, 0, 0, 0, 
    28, 28, 27, 17, 6, 5, 2, 12, 8, 20, 33, 18, 2, 0, 0, 
    20, 10, 0, 0, 0, 4, 1, 0, 0, 0, 3, 7, 0, 0, 0, 
    
    -- channel=506
    0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 12, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 
    18, 18, 12, 0, 0, 7, 6, 0, 0, 0, 0, 0, 4, 15, 22, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 35, 54, 30, 43, 1, 0, 0, 0, 0, 0, 0, 11, 3, 
    24, 44, 74, 60, 25, 41, 11, 11, 0, 0, 6, 0, 0, 0, 0, 
    95, 92, 19, 13, 11, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 
    27, 24, 15, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 4, 
    2, 0, 14, 32, 20, 0, 0, 0, 0, 6, 22, 3, 8, 8, 6, 
    18, 30, 17, 3, 0, 3, 0, 10, 1, 0, 0, 13, 15, 4, 8, 
    
    -- channel=507
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 29, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 26, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=508
    10, 11, 12, 16, 8, 0, 6, 9, 6, 5, 7, 6, 2, 0, 0, 
    10, 8, 9, 11, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    11, 9, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 11, 
    5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 25, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 
    30, 30, 19, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 
    17, 16, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    12, 9, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    5, 24, 58, 31, 22, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    51, 58, 55, 33, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    78, 70, 27, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 25, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 9, 14, 19, 13, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 
    16, 17, 6, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=509
    13, 13, 15, 19, 26, 33, 26, 20, 16, 16, 15, 13, 13, 13, 14, 
    13, 14, 17, 18, 37, 42, 45, 39, 25, 22, 24, 25, 26, 26, 25, 
    13, 15, 18, 23, 39, 48, 55, 58, 46, 32, 32, 34, 30, 27, 28, 
    16, 16, 21, 30, 40, 47, 54, 66, 61, 49, 40, 39, 32, 30, 37, 
    24, 28, 34, 31, 38, 47, 52, 58, 67, 65, 61, 53, 46, 49, 51, 
    29, 28, 35, 26, 38, 45, 46, 51, 59, 66, 68, 57, 54, 55, 49, 
    22, 24, 30, 24, 33, 41, 53, 57, 54, 53, 65, 57, 50, 46, 35, 
    25, 29, 32, 44, 44, 36, 52, 60, 54, 51, 59, 57, 51, 41, 39, 
    31, 34, 41, 31, 49, 44, 54, 58, 49, 48, 55, 58, 52, 44, 49, 
    37, 38, 37, 44, 44, 59, 50, 58, 50, 48, 55, 58, 49, 44, 50, 
    31, 33, 22, 35, 36, 50, 43, 52, 54, 51, 56, 56, 51, 55, 53, 
    20, 16, 22, 36, 32, 42, 43, 32, 41, 45, 48, 53, 57, 59, 53, 
    19, 19, 23, 30, 43, 38, 46, 44, 42, 43, 44, 48, 58, 59, 60, 
    25, 31, 37, 42, 44, 49, 44, 52, 49, 40, 43, 44, 52, 61, 57, 
    35, 41, 48, 51, 52, 55, 49, 57, 59, 54, 51, 54, 56, 59, 58, 
    
    -- channel=510
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 1, 3, 3, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 35, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 6, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 3, 0, 30, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 1, 1, 
    0, 0, 22, 0, 0, 0, 1, 10, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 21, 0, 0, 4, 0, 5, 0, 2, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 6, 0, 10, 0, 4, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 2, 12, 0, 0, 4, 2, 0, 0, 0, 0, 3, 0, 
    
    -- channel=511
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 6, 
    0, 0, 0, 8, 0, 0, 0, 0, 1, 6, 9, 3, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 22, 0, 5, 11, 5, 0, 0, 0, 0, 1, 3, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 7, 0, 0, 0, 1, 0, 0, 3, 0, 0, 0, 
    0, 0, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 1, 11, 1, 
    0, 18, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 
    0, 0, 27, 28, 0, 5, 0, 0, 0, 0, 0, 5, 0, 1, 0, 
    0, 29, 0, 0, 10, 7, 2, 7, 15, 11, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 12, 0, 2, 0, 0, 0, 0, 2, 0, 1, 0, 
    0, 0, 9, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=512
    2, 79, 58, 12, 21, 34, 27, 30, 11, 0, 78, 39, 34, 33, 30, 
    3, 44, 70, 22, 17, 1, 24, 31, 9, 0, 88, 23, 20, 25, 25, 
    4, 17, 94, 22, 28, 0, 0, 16, 3, 28, 33, 18, 10, 16, 15, 
    0, 58, 59, 0, 37, 0, 0, 0, 15, 45, 13, 38, 8, 0, 21, 
    0, 33, 12, 0, 39, 7, 0, 0, 15, 32, 29, 34, 6, 0, 18, 
    6, 12, 3, 0, 22, 0, 0, 0, 15, 28, 23, 37, 4, 0, 3, 
    3, 11, 0, 29, 0, 13, 0, 21, 0, 16, 22, 41, 6, 0, 0, 
    0, 13, 0, 59, 0, 3, 0, 0, 27, 6, 4, 14, 37, 0, 13, 
    0, 11, 18, 30, 10, 10, 0, 0, 32, 6, 14, 6, 26, 1, 39, 
    0, 6, 15, 7, 5, 0, 6, 1, 0, 26, 0, 25, 29, 9, 21, 
    2, 0, 26, 9, 9, 0, 22, 7, 0, 0, 23, 24, 18, 1, 8, 
    3, 0, 30, 6, 0, 0, 24, 11, 0, 0, 37, 9, 22, 3, 7, 
    0, 0, 23, 4, 0, 19, 26, 7, 0, 0, 28, 8, 5, 16, 10, 
    0, 0, 21, 12, 0, 30, 3, 9, 0, 10, 21, 13, 1, 31, 20, 
    0, 4, 5, 25, 0, 0, 0, 16, 0, 30, 17, 18, 13, 19, 18, 
    
    -- channel=513
    4, 0, 6, 14, 9, 6, 15, 11, 15, 38, 0, 16, 20, 17, 19, 
    5, 0, 0, 0, 0, 11, 0, 0, 8, 6, 2, 0, 9, 11, 13, 
    7, 4, 0, 19, 0, 5, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    52, 12, 32, 9, 0, 0, 15, 18, 5, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 12, 0, 0, 4, 3, 0, 0, 2, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 4, 2, 0, 6, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 9, 4, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 5, 1, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 22, 4, 0, 1, 0, 4, 1, 3, 0, 1, 
    0, 0, 0, 0, 0, 2, 0, 0, 6, 0, 0, 3, 1, 11, 0, 
    
    -- channel=514
    25, 81, 20, 0, 0, 9, 0, 6, 0, 0, 70, 3, 0, 0, 0, 
    25, 54, 53, 11, 1, 0, 3, 2, 0, 0, 71, 0, 0, 0, 0, 
    23, 33, 92, 12, 20, 0, 4, 21, 0, 19, 30, 15, 0, 0, 0, 
    0, 62, 46, 0, 34, 0, 0, 0, 19, 40, 1, 25, 0, 0, 10, 
    0, 10, 0, 0, 44, 0, 0, 0, 17, 29, 19, 23, 0, 0, 20, 
    0, 1, 0, 0, 15, 0, 0, 0, 11, 23, 15, 37, 0, 0, 7, 
    0, 1, 0, 13, 3, 21, 0, 12, 0, 16, 15, 29, 0, 0, 0, 
    0, 1, 0, 48, 0, 0, 0, 0, 16, 0, 0, 15, 17, 0, 2, 
    0, 15, 0, 9, 0, 0, 0, 0, 29, 0, 0, 0, 51, 6, 34, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 15, 0, 8, 5, 0, 17, 
    0, 0, 22, 0, 0, 0, 23, 0, 0, 0, 10, 9, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 25, 0, 6, 0, 0, 
    0, 0, 26, 0, 0, 2, 10, 0, 0, 0, 20, 0, 0, 4, 0, 
    0, 0, 34, 8, 0, 0, 0, 0, 0, 1, 17, 4, 0, 23, 6, 
    0, 5, 22, 22, 0, 0, 0, 2, 0, 22, 10, 7, 0, 9, 8, 
    
    -- channel=515
    0, 10, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 11, 4, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 15, 35, 40, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 
    0, 0, 0, 0, 0, 1, 0, 4, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 3, 0, 0, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 12, 2, 0, 0, 0, 0, 0, 6, 2, 13, 63, 31, 11, 2, 
    0, 3, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 32, 49, 24, 
    0, 0, 0, 0, 0, 22, 10, 0, 0, 0, 10, 1, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 4, 10, 3, 6, 9, 0, 0, 2, 7, 
    3, 0, 0, 0, 3, 12, 0, 0, 1, 6, 0, 4, 0, 0, 0, 
    2, 7, 3, 0, 8, 22, 3, 12, 16, 11, 2, 7, 19, 14, 0, 
    6, 8, 9, 0, 0, 0, 5, 15, 17, 12, 0, 1, 5, 0, 0, 
    23, 4, 13, 8, 0, 4, 27, 16, 12, 1, 3, 0, 0, 0, 8, 
    
    -- channel=516
    0, 21, 41, 26, 23, 35, 33, 40, 31, 0, 42, 48, 45, 44, 39, 
    0, 0, 37, 29, 37, 18, 34, 43, 27, 0, 75, 48, 44, 43, 41, 
    0, 0, 47, 29, 50, 0, 0, 5, 1, 29, 53, 40, 45, 54, 53, 
    0, 27, 72, 11, 49, 26, 20, 2, 8, 41, 35, 65, 56, 32, 45, 
    33, 60, 36, 0, 44, 30, 19, 0, 10, 29, 44, 69, 48, 13, 36, 
    35, 37, 29, 15, 47, 27, 2, 0, 20, 31, 34, 67, 50, 22, 27, 
    32, 32, 0, 38, 14, 19, 6, 33, 21, 31, 33, 67, 51, 49, 35, 
    24, 33, 0, 69, 31, 28, 19, 11, 29, 21, 17, 25, 60, 36, 45, 
    15, 23, 38, 53, 44, 53, 29, 0, 26, 11, 27, 0, 13, 5, 51, 
    31, 37, 45, 39, 29, 24, 37, 33, 15, 34, 6, 21, 30, 21, 16, 
    39, 17, 47, 40, 44, 9, 33, 28, 25, 4, 14, 33, 30, 8, 12, 
    36, 16, 51, 45, 34, 21, 45, 35, 22, 0, 34, 18, 31, 14, 7, 
    30, 18, 46, 37, 1, 0, 38, 23, 7, 0, 23, 12, 7, 11, 11, 
    24, 11, 37, 45, 24, 46, 19, 10, 0, 0, 16, 9, 0, 18, 22, 
    11, 17, 20, 45, 28, 17, 0, 11, 0, 10, 9, 13, 8, 17, 13, 
    
    -- channel=517
    0, 0, 0, 0, 0, 0, 5, 8, 27, 5, 0, 21, 13, 9, 6, 
    0, 0, 0, 0, 23, 4, 0, 7, 0, 4, 36, 10, 4, 2, 1, 
    1, 0, 0, 0, 1, 2, 0, 0, 0, 4, 21, 0, 0, 11, 16, 
    63, 58, 71, 0, 0, 12, 38, 13, 0, 0, 0, 4, 14, 0, 0, 
    34, 50, 5, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 15, 5, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 12, 3, 0, 0, 0, 11, 18, 
    0, 0, 0, 6, 8, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 8, 5, 33, 16, 2, 0, 0, 3, 0, 0, 0, 0, 
    2, 10, 0, 2, 0, 0, 0, 18, 25, 4, 0, 0, 13, 5, 0, 
    0, 0, 0, 1, 8, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    
    -- channel=518
    0, 3, 12, 18, 14, 12, 22, 20, 16, 25, 0, 39, 32, 33, 29, 
    0, 0, 2, 5, 16, 27, 11, 26, 27, 0, 44, 34, 30, 29, 27, 
    0, 0, 0, 27, 14, 18, 3, 0, 0, 0, 55, 17, 25, 28, 33, 
    46, 12, 81, 27, 9, 5, 30, 22, 4, 20, 22, 26, 41, 42, 18, 
    23, 67, 34, 14, 22, 10, 14, 9, 2, 12, 16, 46, 34, 28, 33, 
    28, 33, 27, 12, 32, 19, 5, 0, 17, 19, 24, 30, 35, 32, 38, 
    32, 25, 21, 9, 21, 0, 13, 7, 26, 23, 17, 39, 36, 32, 44, 
    30, 20, 9, 19, 29, 27, 0, 35, 0, 25, 22, 13, 9, 36, 23, 
    31, 16, 1, 47, 12, 39, 35, 8, 20, 9, 17, 25, 12, 0, 18, 
    27, 37, 27, 28, 25, 12, 3, 14, 44, 16, 16, 3, 20, 28, 24, 
    29, 32, 13, 29, 30, 26, 14, 15, 5, 30, 0, 23, 23, 6, 14, 
    31, 24, 28, 22, 27, 8, 32, 24, 22, 0, 23, 16, 14, 16, 6, 
    32, 23, 30, 22, 16, 0, 16, 16, 7, 3, 13, 8, 9, 0, 14, 
    29, 24, 24, 20, 10, 38, 27, 7, 0, 0, 14, 7, 2, 8, 10, 
    12, 18, 26, 12, 18, 21, 3, 3, 0, 1, 7, 8, 5, 22, 6, 
    
    -- channel=519
    0, 0, 42, 30, 32, 33, 35, 30, 24, 13, 0, 38, 35, 36, 36, 
    0, 0, 47, 10, 22, 29, 41, 38, 40, 22, 0, 38, 35, 36, 39, 
    0, 0, 16, 5, 23, 35, 19, 35, 43, 4, 31, 33, 38, 38, 38, 
    0, 0, 31, 41, 28, 28, 11, 18, 10, 5, 48, 26, 44, 63, 39, 
    38, 28, 42, 27, 13, 28, 39, 32, 15, 6, 35, 40, 44, 49, 38, 
    42, 37, 52, 19, 32, 38, 35, 3, 17, 4, 27, 42, 51, 52, 42, 
    44, 33, 46, 31, 14, 0, 33, 11, 36, 21, 17, 42, 49, 52, 38, 
    50, 38, 35, 32, 41, 35, 23, 29, 30, 21, 47, 64, 56, 66, 36, 
    52, 21, 21, 27, 30, 29, 16, 34, 14, 17, 46, 12, 24, 52, 43, 
    49, 29, 37, 36, 29, 44, 36, 20, 13, 21, 46, 27, 8, 40, 33, 
    47, 42, 29, 29, 34, 39, 26, 28, 42, 53, 13, 26, 31, 26, 33, 
    46, 50, 26, 40, 50, 36, 33, 30, 41, 29, 19, 30, 35, 31, 21, 
    48, 52, 30, 35, 51, 0, 42, 37, 41, 28, 27, 24, 39, 25, 23, 
    49, 51, 26, 38, 37, 13, 48, 32, 32, 13, 25, 19, 23, 14, 26, 
    45, 48, 24, 39, 34, 45, 42, 33, 31, 9, 21, 24, 15, 25, 26, 
    
    -- channel=520
    0, 0, 8, 15, 16, 6, 18, 10, 35, 21, 0, 26, 29, 26, 30, 
    0, 0, 0, 0, 26, 17, 7, 14, 26, 48, 0, 33, 33, 30, 32, 
    0, 0, 0, 0, 8, 56, 1, 0, 7, 2, 0, 15, 31, 30, 34, 
    33, 0, 0, 18, 0, 49, 41, 22, 0, 0, 23, 7, 40, 38, 13, 
    39, 2, 26, 35, 0, 23, 37, 31, 0, 0, 6, 11, 38, 46, 0, 
    24, 13, 26, 30, 0, 20, 39, 16, 10, 0, 4, 1, 38, 51, 8, 
    23, 17, 30, 17, 20, 9, 35, 0, 28, 2, 5, 6, 31, 50, 34, 
    24, 14, 58, 0, 32, 22, 25, 23, 7, 2, 21, 0, 9, 37, 19, 
    38, 5, 40, 0, 33, 39, 36, 53, 0, 19, 23, 26, 0, 9, 0, 
    37, 13, 24, 23, 14, 17, 28, 47, 41, 5, 28, 12, 10, 19, 0, 
    27, 29, 11, 31, 28, 44, 2, 15, 43, 30, 7, 7, 15, 23, 6, 
    20, 37, 0, 31, 38, 34, 21, 24, 33, 39, 0, 12, 14, 24, 21, 
    23, 24, 0, 29, 53, 4, 12, 20, 28, 18, 0, 8, 5, 9, 13, 
    24, 21, 0, 21, 53, 24, 24, 15, 15, 2, 0, 5, 13, 0, 8, 
    12, 15, 0, 9, 35, 34, 20, 4, 14, 0, 0, 4, 12, 0, 3, 
    
    -- channel=521
    0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 1, 18, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 9, 0, 11, 0, 0, 12, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 3, 7, 5, 0, 0, 5, 
    0, 0, 0, 0, 5, 5, 0, 0, 0, 1, 5, 3, 0, 0, 0, 
    0, 0, 0, 0, 2, 5, 0, 0, 0, 0, 1, 13, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 8, 0, 2, 0, 0, 11, 0, 7, 26, 29, 3, 1, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 18, 17, 
    0, 0, 0, 0, 0, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 2, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=522
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=523
    0, 0, 43, 38, 32, 33, 41, 48, 63, 10, 50, 65, 64, 60, 56, 
    0, 0, 12, 41, 74, 37, 37, 56, 48, 34, 85, 73, 65, 62, 58, 
    0, 0, 19, 49, 77, 47, 0, 0, 0, 56, 65, 57, 71, 79, 78, 
    67, 87, 79, 25, 54, 80, 81, 34, 27, 50, 55, 91, 93, 54, 60, 
    78, 85, 62, 28, 55, 60, 54, 21, 27, 40, 57, 86, 83, 47, 41, 
    60, 56, 47, 58, 60, 50, 35, 36, 54, 59, 49, 74, 79, 63, 39, 
    52, 53, 15, 65, 45, 57, 43, 55, 53, 51, 61, 78, 80, 91, 69, 
    43, 48, 43, 65, 65, 55, 55, 49, 46, 42, 38, 0, 62, 55, 75, 
    44, 38, 78, 64, 86, 100, 82, 46, 22, 44, 48, 38, 0, 3, 45, 
    62, 64, 68, 65, 50, 41, 70, 87, 72, 59, 16, 37, 63, 37, 11, 
    63, 47, 67, 76, 80, 46, 46, 55, 60, 18, 36, 49, 48, 31, 23, 
    55, 47, 63, 74, 63, 49, 72, 65, 51, 25, 44, 34, 48, 42, 34, 
    50, 35, 53, 69, 32, 25, 50, 40, 26, 20, 29, 28, 9, 24, 32, 
    44, 27, 38, 69, 67, 91, 28, 24, 13, 12, 23, 28, 17, 27, 42, 
    19, 30, 20, 60, 64, 42, 7, 15, 2, 25, 19, 30, 34, 28, 21, 
    
    -- channel=524
    0, 104, 14, 0, 0, 0, 0, 0, 0, 0, 72, 5, 0, 0, 0, 
    2, 65, 41, 4, 0, 0, 0, 0, 0, 0, 101, 0, 0, 0, 0, 
    1, 23, 75, 19, 20, 0, 0, 14, 0, 0, 42, 0, 0, 0, 0, 
    0, 55, 75, 0, 30, 0, 0, 0, 4, 58, 0, 25, 0, 0, 0, 
    0, 26, 0, 0, 50, 0, 0, 0, 5, 35, 14, 22, 0, 0, 13, 
    0, 0, 0, 0, 20, 0, 0, 0, 1, 28, 16, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 11, 0, 6, 18, 30, 0, 0, 0, 
    0, 0, 0, 51, 0, 0, 0, 0, 0, 8, 0, 26, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 0, 0, 43, 0, 0, 0, 57, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 6, 0, 16, 
    0, 0, 6, 0, 0, 0, 17, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 29, 0, 0, 0, 4, 0, 0, 0, 29, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 6, 9, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 5, 0, 0, 0, 0, 8, 0, 0, 18, 0, 
    0, 0, 14, 9, 0, 0, 0, 0, 0, 17, 0, 0, 0, 11, 0, 
    
    -- channel=525
    0, 27, 42, 21, 16, 29, 26, 25, 20, 0, 35, 28, 32, 29, 30, 
    0, 11, 50, 24, 10, 0, 17, 19, 14, 0, 36, 14, 19, 23, 26, 
    1, 3, 54, 22, 18, 0, 5, 15, 12, 19, 12, 8, 8, 11, 10, 
    0, 20, 24, 0, 24, 1, 0, 4, 14, 19, 6, 15, 0, 0, 6, 
    0, 9, 0, 0, 23, 5, 0, 0, 12, 14, 10, 15, 0, 0, 0, 
    0, 0, 0, 0, 14, 0, 0, 1, 10, 10, 6, 16, 0, 0, 0, 
    0, 3, 0, 27, 4, 7, 0, 12, 0, 9, 2, 15, 0, 0, 0, 
    0, 5, 8, 45, 0, 1, 1, 0, 19, 0, 0, 3, 14, 0, 0, 
    0, 5, 26, 16, 5, 6, 0, 0, 13, 4, 16, 7, 16, 2, 11, 
    0, 0, 9, 9, 1, 0, 5, 0, 0, 20, 4, 24, 17, 11, 11, 
    0, 0, 13, 3, 5, 0, 14, 5, 3, 0, 16, 18, 16, 8, 10, 
    0, 0, 12, 4, 1, 6, 12, 8, 3, 0, 22, 9, 19, 6, 9, 
    0, 0, 6, 3, 0, 17, 23, 9, 5, 5, 20, 10, 8, 15, 13, 
    0, 0, 3, 6, 0, 19, 7, 13, 8, 8, 18, 12, 6, 19, 16, 
    0, 0, 0, 10, 0, 0, 1, 18, 7, 17, 12, 14, 11, 14, 14, 
    
    -- channel=526
    0, 25, 43, 33, 31, 43, 38, 37, 21, 1, 28, 25, 36, 39, 40, 
    0, 15, 47, 31, 5, 12, 29, 28, 21, 5, 19, 24, 30, 35, 37, 
    0, 5, 43, 24, 8, 0, 17, 33, 34, 21, 11, 27, 24, 24, 23, 
    0, 0, 5, 20, 18, 0, 0, 1, 11, 15, 13, 20, 6, 11, 27, 
    11, 9, 16, 15, 14, 8, 5, 5, 11, 14, 17, 23, 16, 17, 31, 
    21, 20, 23, 17, 11, 6, 8, 7, 1, 6, 14, 29, 19, 19, 29, 
    26, 24, 23, 30, 9, 10, 1, 7, 0, 7, 10, 24, 20, 15, 16, 
    25, 28, 18, 31, 4, 6, 3, 0, 20, 9, 14, 39, 41, 22, 26, 
    21, 26, 16, 12, 9, 0, 0, 0, 20, 19, 17, 17, 38, 40, 40, 
    21, 16, 16, 14, 14, 15, 11, 0, 0, 19, 18, 29, 18, 17, 32, 
    22, 15, 20, 11, 12, 6, 20, 14, 12, 14, 28, 19, 19, 19, 21, 
    23, 18, 20, 12, 11, 15, 15, 13, 13, 17, 23, 19, 20, 16, 17, 
    23, 26, 26, 11, 10, 24, 26, 23, 22, 20, 26, 21, 21, 26, 18, 
    23, 29, 33, 14, 10, 8, 18, 28, 25, 24, 22, 20, 17, 24, 20, 
    30, 30, 29, 17, 11, 15, 24, 29, 21, 25, 21, 20, 17, 18, 23, 
    
    -- channel=527
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 12, 0, 0, 3, 4, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 19, 20, 0, 0, 0, 0, 11, 5, 10, 8, 5, 
    0, 0, 0, 0, 2, 17, 12, 8, 2, 0, 6, 1, 4, 0, 0, 
    0, 0, 0, 0, 6, 16, 12, 5, 3, 0, 2, 6, 8, 0, 0, 
    0, 0, 0, 0, 1, 6, 11, 12, 11, 10, 1, 1, 7, 9, 0, 
    0, 0, 0, 0, 11, 13, 22, 0, 12, 0, 3, 2, 13, 7, 1, 
    0, 0, 0, 0, 19, 15, 9, 13, 0, 0, 0, 0, 0, 6, 0, 
    1, 0, 4, 5, 7, 17, 26, 16, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 10, 3, 5, 6, 5, 8, 14, 0, 0, 0, 0, 0, 0, 
    0, 3, 3, 15, 11, 9, 0, 1, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=528
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 15, 10, 14, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 3, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 14, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 11, 17, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 14, 22, 0, 0, 4, 2, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 3, 0, 0, 
    4, 0, 0, 0, 0, 0, 1, 0, 9, 0, 0, 0, 0, 0, 0, 
    
    -- channel=529
    0, 30, 14, 0, 0, 5, 1, 0, 0, 0, 5, 0, 0, 0, 1, 
    0, 18, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 29, 0, 0, 0, 5, 13, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 22, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 3, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 1, 7, 3, 0, 1, 0, 0, 0, 3, 
    
    -- channel=530
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=531
    0, 0, 17, 17, 22, 12, 22, 15, 49, 30, 0, 36, 30, 26, 29, 
    0, 0, 1, 0, 43, 25, 16, 22, 33, 53, 0, 43, 39, 31, 31, 
    0, 0, 0, 0, 22, 66, 9, 0, 11, 14, 24, 28, 42, 43, 45, 
    60, 2, 22, 24, 6, 62, 53, 40, 15, 0, 41, 20, 49, 52, 24, 
    59, 24, 42, 43, 1, 33, 49, 42, 12, 0, 23, 29, 52, 57, 10, 
    39, 26, 42, 33, 18, 30, 46, 23, 32, 6, 19, 20, 53, 70, 29, 
    37, 28, 31, 30, 31, 19, 51, 9, 44, 24, 18, 23, 44, 68, 49, 
    37, 23, 54, 2, 44, 34, 40, 30, 22, 8, 30, 0, 15, 52, 32, 
    57, 17, 51, 4, 46, 59, 48, 72, 0, 17, 43, 30, 0, 15, 0, 
    56, 27, 37, 37, 25, 26, 38, 58, 52, 19, 35, 19, 15, 31, 0, 
    44, 42, 27, 40, 40, 53, 15, 20, 54, 40, 10, 19, 25, 29, 16, 
    36, 56, 12, 41, 46, 37, 29, 31, 41, 42, 3, 19, 27, 29, 27, 
    40, 42, 8, 42, 64, 0, 22, 24, 32, 24, 7, 15, 13, 14, 24, 
    40, 39, 0, 39, 63, 27, 28, 19, 19, 4, 11, 13, 21, 0, 20, 
    24, 39, 0, 27, 46, 43, 23, 11, 22, 0, 8, 16, 21, 10, 11, 
    
    -- channel=532
    5, 89, 20, 12, 15, 22, 18, 21, 0, 0, 60, 22, 20, 22, 19, 
    7, 62, 28, 27, 0, 19, 16, 19, 10, 0, 75, 14, 15, 19, 17, 
    8, 26, 48, 39, 15, 0, 16, 24, 0, 8, 37, 21, 10, 11, 10, 
    0, 47, 54, 10, 24, 0, 0, 0, 13, 54, 1, 34, 9, 0, 20, 
    0, 38, 12, 0, 40, 6, 0, 0, 12, 40, 19, 32, 7, 0, 38, 
    9, 23, 6, 6, 24, 8, 0, 0, 6, 33, 25, 34, 7, 0, 24, 
    14, 22, 10, 3, 11, 19, 0, 22, 0, 16, 28, 35, 15, 0, 13, 
    11, 23, 0, 30, 1, 5, 0, 13, 3, 33, 6, 44, 19, 1, 18, 
    0, 27, 0, 40, 0, 0, 6, 0, 53, 13, 0, 9, 60, 5, 43, 
    0, 25, 13, 4, 21, 11, 0, 0, 8, 21, 0, 10, 26, 10, 38, 
    9, 6, 19, 13, 10, 0, 25, 17, 0, 0, 12, 21, 14, 2, 14, 
    16, 0, 37, 7, 1, 0, 18, 13, 3, 0, 35, 13, 9, 5, 2, 
    12, 3, 38, 6, 0, 37, 12, 13, 0, 0, 24, 13, 13, 7, 9, 
    9, 5, 45, 9, 0, 23, 6, 10, 3, 14, 20, 15, 3, 29, 12, 
    11, 3, 48, 15, 0, 0, 0, 10, 0, 28, 18, 13, 7, 24, 15, 
    
    -- channel=533
    23, 36, 16, 15, 7, 10, 11, 9, 9, 8, 18, 15, 12, 10, 10, 
    23, 28, 24, 18, 6, 4, 8, 8, 8, 0, 25, 0, 1, 4, 7, 
    25, 25, 30, 17, 12, 0, 10, 9, 6, 4, 8, 0, 0, 0, 0, 
    12, 16, 24, 2, 18, 0, 4, 13, 14, 19, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 19, 0, 0, 5, 12, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 4, 0, 1, 12, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 2, 0, 0, 12, 8, 9, 0, 0, 0, 0, 0, 
    0, 0, 3, 25, 0, 4, 0, 9, 4, 3, 0, 1, 0, 0, 0, 
    0, 0, 10, 24, 0, 2, 0, 0, 16, 0, 5, 1, 7, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 5, 9, 10, 10, 9, 7, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 9, 3, 14, 12, 4, 9, 
    0, 0, 2, 0, 0, 1, 7, 3, 0, 0, 15, 9, 10, 4, 8, 
    0, 0, 0, 0, 0, 11, 7, 2, 1, 2, 13, 7, 12, 7, 9, 
    0, 0, 0, 0, 0, 17, 13, 4, 3, 8, 14, 8, 8, 16, 8, 
    0, 0, 0, 0, 0, 0, 2, 13, 9, 10, 13, 10, 9, 15, 12, 
    
    -- channel=534
    1, 0, 0, 0, 0, 0, 0, 0, 13, 13, 13, 3, 1, 1, 1, 
    1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 18, 4, 6, 3, 0, 
    0, 0, 9, 14, 0, 0, 0, 0, 0, 4, 11, 1, 0, 0, 1, 
    69, 68, 12, 0, 0, 2, 16, 9, 10, 0, 0, 2, 0, 0, 0, 
    0, 0, 1, 0, 10, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 9, 13, 9, 0, 0, 0, 3, 1, 
    0, 0, 0, 6, 21, 25, 2, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 5, 9, 0, 0, 7, 14, 6, 0, 0, 0, 18, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 6, 25, 7, 0, 0, 10, 0, 0, 
    0, 0, 0, 5, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 0, 0, 
    
    -- channel=535
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=536
    21, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=537
    8, 0, 0, 11, 7, 0, 5, 0, 3, 68, 0, 0, 1, 1, 5, 
    7, 0, 0, 0, 0, 25, 0, 0, 11, 43, 0, 0, 3, 1, 5, 
    9, 0, 0, 0, 0, 46, 22, 2, 10, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 37, 0, 0, 13, 29, 0, 0, 0, 0, 0, 27, 0, 
    0, 0, 0, 39, 0, 0, 16, 42, 0, 0, 0, 0, 0, 32, 0, 
    0, 0, 2, 4, 0, 6, 24, 5, 0, 0, 0, 0, 0, 18, 0, 
    2, 0, 40, 0, 7, 0, 29, 0, 16, 0, 0, 0, 0, 0, 8, 
    13, 0, 38, 0, 18, 1, 0, 25, 0, 7, 7, 5, 0, 14, 0, 
    21, 0, 0, 0, 0, 0, 12, 34, 0, 1, 0, 14, 0, 0, 0, 
    1, 0, 0, 0, 0, 4, 0, 0, 25, 0, 34, 0, 0, 16, 1, 
    0, 21, 0, 0, 0, 33, 0, 0, 3, 49, 0, 0, 0, 16, 14, 
    0, 15, 0, 0, 11, 12, 0, 0, 14, 32, 0, 7, 0, 15, 8, 
    1, 10, 0, 0, 42, 0, 0, 6, 22, 20, 0, 4, 18, 0, 7, 
    7, 13, 0, 0, 14, 0, 30, 7, 20, 5, 0, 0, 18, 0, 0, 
    6, 0, 0, 0, 2, 25, 32, 2, 30, 0, 0, 0, 1, 3, 0, 
    
    -- channel=538
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=539
    1, 72, 30, 0, 0, 5, 0, 3, 0, 0, 66, 21, 1, 0, 0, 
    1, 30, 62, 1, 5, 0, 3, 5, 0, 0, 90, 0, 0, 0, 0, 
    1, 7, 99, 1, 29, 0, 0, 2, 0, 5, 39, 1, 0, 0, 0, 
    0, 66, 83, 0, 37, 0, 0, 0, 10, 41, 2, 29, 0, 0, 0, 
    0, 21, 0, 0, 47, 0, 0, 0, 5, 20, 25, 26, 0, 0, 1, 
    0, 0, 0, 0, 24, 0, 0, 0, 10, 17, 10, 37, 0, 0, 0, 
    0, 0, 0, 6, 0, 1, 0, 11, 0, 9, 10, 35, 0, 0, 0, 
    0, 0, 0, 71, 0, 0, 0, 0, 11, 0, 0, 8, 7, 0, 0, 
    0, 0, 0, 25, 0, 3, 0, 0, 27, 0, 7, 0, 30, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 3, 2, 0, 0, 
    0, 0, 18, 0, 0, 0, 16, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 29, 0, 0, 0, 7, 0, 0, 0, 26, 0, 7, 0, 0, 
    0, 0, 14, 0, 0, 0, 15, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 9, 4, 0, 0, 0, 0, 0, 0, 10, 0, 0, 13, 4, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 6, 0, 0, 0, 7, 0, 
    
    -- channel=540
    0, 0, 34, 8, 0, 13, 11, 8, 33, 0, 0, 9, 12, 11, 13, 
    0, 0, 32, 0, 18, 0, 15, 16, 9, 37, 0, 13, 9, 7, 11, 
    0, 0, 19, 0, 13, 12, 0, 0, 18, 31, 0, 6, 11, 13, 13, 
    0, 0, 0, 0, 15, 37, 2, 0, 0, 0, 25, 6, 8, 11, 18, 
    39, 0, 10, 9, 0, 7, 17, 12, 1, 0, 14, 6, 16, 16, 0, 
    17, 0, 19, 8, 0, 0, 17, 3, 4, 0, 0, 8, 17, 28, 0, 
    9, 4, 0, 39, 0, 0, 5, 4, 9, 2, 0, 7, 11, 35, 0, 
    4, 6, 19, 21, 2, 5, 22, 0, 42, 0, 8, 0, 45, 17, 21, 
    21, 0, 37, 0, 32, 19, 0, 30, 0, 1, 31, 0, 0, 23, 8, 
    28, 0, 8, 17, 0, 0, 32, 25, 0, 4, 7, 21, 0, 2, 0, 
    18, 0, 18, 0, 10, 6, 0, 0, 37, 0, 20, 0, 5, 8, 0, 
    7, 29, 0, 11, 9, 21, 4, 5, 7, 21, 0, 1, 19, 5, 13, 
    9, 20, 0, 11, 17, 0, 16, 5, 15, 10, 2, 2, 0, 21, 5, 
    11, 16, 0, 18, 29, 0, 2, 7, 6, 2, 0, 0, 5, 0, 12, 
    11, 31, 0, 20, 13, 4, 10, 15, 10, 0, 0, 6, 10, 0, 6, 
    
    -- channel=541
    5, 0, 0, 19, 14, 4, 19, 6, 44, 63, 0, 11, 21, 17, 23, 
    3, 0, 0, 0, 10, 22, 0, 0, 20, 75, 0, 15, 22, 18, 21, 
    5, 0, 0, 0, 0, 67, 11, 0, 7, 0, 0, 0, 11, 10, 19, 
    71, 0, 0, 33, 0, 37, 45, 40, 3, 0, 0, 0, 13, 26, 0, 
    38, 0, 9, 58, 0, 1, 30, 51, 0, 0, 0, 0, 11, 44, 0, 
    11, 0, 12, 31, 0, 6, 37, 23, 7, 0, 0, 0, 7, 46, 4, 
    12, 4, 34, 0, 15, 0, 38, 0, 23, 0, 0, 0, 0, 23, 28, 
    17, 0, 67, 0, 25, 9, 18, 22, 0, 0, 7, 0, 0, 16, 0, 
    39, 0, 30, 0, 7, 18, 28, 61, 0, 15, 12, 36, 0, 0, 0, 
    26, 6, 4, 10, 0, 0, 0, 31, 48, 0, 32, 5, 2, 18, 0, 
    7, 28, 0, 10, 7, 44, 0, 0, 29, 40, 0, 1, 7, 27, 10, 
    2, 36, 0, 6, 19, 29, 0, 8, 21, 52, 0, 9, 0, 25, 25, 
    9, 20, 0, 5, 53, 0, 0, 10, 26, 29, 0, 9, 5, 4, 17, 
    14, 21, 0, 0, 46, 17, 21, 12, 21, 10, 0, 7, 23, 0, 4, 
    7, 12, 0, 0, 20, 29, 30, 5, 32, 0, 2, 4, 18, 0, 0, 
    
    -- channel=542
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=543
    15, 0, 0, 9, 11, 0, 4, 2, 27, 31, 0, 6, 5, 2, 3, 
    14, 0, 0, 6, 30, 19, 6, 6, 15, 50, 0, 17, 15, 10, 9, 
    13, 0, 0, 3, 21, 53, 20, 3, 17, 20, 1, 13, 21, 20, 21, 
    36, 4, 0, 18, 10, 50, 37, 32, 18, 0, 23, 6, 31, 30, 12, 
    27, 0, 15, 35, 3, 33, 38, 41, 17, 6, 14, 4, 28, 33, 0, 
    16, 10, 16, 23, 11, 29, 42, 36, 23, 12, 14, 1, 25, 30, 1, 
    13, 10, 18, 10, 29, 29, 42, 18, 35, 20, 16, 2, 20, 29, 20, 
    14, 7, 35, 0, 33, 27, 41, 23, 20, 12, 18, 0, 1, 24, 12, 
    25, 8, 33, 11, 34, 36, 40, 54, 0, 20, 19, 17, 0, 12, 0, 
    23, 10, 19, 28, 21, 26, 34, 46, 30, 9, 25, 11, 9, 14, 0, 
    17, 23, 14, 26, 24, 38, 13, 23, 38, 25, 14, 10, 15, 27, 11, 
    14, 28, 2, 29, 31, 32, 15, 23, 26, 37, 0, 16, 15, 21, 23, 
    15, 16, 0, 29, 45, 18, 13, 18, 27, 22, 2, 15, 14, 17, 17, 
    15, 10, 0, 22, 45, 17, 23, 14, 19, 15, 6, 13, 21, 2, 12, 
    12, 8, 0, 15, 33, 27, 22, 9, 22, 0, 9, 11, 18, 4, 11, 
    
    -- channel=544
    0, 132, 33, 0, 0, 13, 0, 5, 0, 0, 108, 9, 0, 0, 0, 
    1, 75, 74, 24, 0, 0, 15, 11, 0, 0, 116, 0, 0, 0, 0, 
    1, 25, 120, 16, 37, 0, 0, 27, 0, 20, 36, 17, 0, 0, 0, 
    0, 50, 63, 0, 64, 0, 0, 0, 7, 72, 0, 50, 0, 0, 23, 
    0, 24, 0, 0, 65, 2, 0, 0, 13, 51, 31, 42, 0, 0, 26, 
    0, 3, 0, 0, 32, 0, 0, 0, 0, 35, 24, 57, 0, 0, 0, 
    0, 0, 0, 12, 0, 14, 0, 31, 0, 21, 22, 51, 0, 0, 0, 
    0, 9, 0, 78, 0, 0, 0, 0, 25, 10, 0, 55, 49, 0, 5, 
    0, 13, 0, 28, 0, 0, 0, 0, 52, 0, 0, 0, 68, 3, 64, 
    0, 0, 6, 0, 8, 2, 2, 0, 0, 18, 0, 6, 7, 0, 25, 
    0, 0, 33, 0, 0, 0, 35, 8, 0, 0, 10, 11, 2, 0, 0, 
    0, 0, 52, 0, 0, 0, 9, 0, 0, 0, 37, 0, 10, 0, 0, 
    0, 0, 43, 0, 0, 19, 19, 0, 0, 0, 26, 0, 0, 4, 0, 
    0, 0, 46, 11, 0, 0, 0, 0, 0, 0, 15, 0, 0, 30, 5, 
    0, 0, 27, 36, 0, 0, 0, 4, 0, 24, 6, 3, 0, 10, 9, 
    
    -- channel=545
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=546
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=547
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 0, 0, 4, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 5, 0, 4, 0, 0, 4, 5, 0, 0, 
    15, 0, 0, 10, 0, 23, 11, 10, 0, 0, 16, 0, 14, 29, 7, 
    13, 0, 12, 22, 0, 14, 20, 24, 0, 0, 1, 0, 21, 35, 3, 
    13, 8, 17, 10, 0, 14, 28, 10, 3, 0, 3, 0, 23, 35, 13, 
    14, 7, 20, 0, 15, 5, 23, 0, 19, 4, 2, 0, 20, 25, 19, 
    19, 3, 17, 0, 17, 17, 16, 15, 4, 4, 18, 0, 5, 31, 15, 
    31, 2, 0, 0, 14, 14, 19, 32, 0, 7, 7, 10, 0, 19, 0, 
    24, 5, 4, 10, 13, 20, 18, 19, 14, 0, 14, 0, 0, 2, 0, 
    19, 26, 2, 11, 10, 31, 3, 11, 20, 19, 0, 0, 0, 7, 0, 
    18, 32, 0, 13, 20, 13, 2, 7, 16, 19, 0, 2, 0, 6, 5, 
    21, 25, 0, 18, 36, 0, 0, 8, 15, 8, 0, 1, 4, 0, 1, 
    22, 23, 0, 13, 23, 0, 9, 4, 7, 0, 0, 0, 5, 0, 0, 
    19, 16, 0, 8, 20, 17, 12, 0, 8, 0, 0, 0, 0, 0, 0, 
    
    -- channel=548
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 1, 9, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 21, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 
    0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=549
    0, 2, 36, 35, 29, 35, 33, 33, 23, 2, 16, 34, 42, 40, 40, 
    0, 0, 32, 37, 28, 25, 37, 36, 38, 12, 25, 39, 42, 43, 45, 
    0, 0, 15, 34, 47, 24, 20, 35, 38, 23, 29, 38, 43, 45, 42, 
    0, 0, 14, 30, 50, 34, 15, 11, 13, 30, 38, 45, 52, 46, 42, 
    19, 23, 28, 16, 37, 43, 38, 21, 19, 28, 36, 47, 48, 27, 31, 
    32, 33, 32, 23, 40, 43, 32, 16, 18, 25, 32, 49, 45, 24, 18, 
    30, 31, 28, 38, 26, 27, 28, 30, 25, 27, 30, 46, 47, 38, 18, 
    28, 36, 33, 50, 39, 37, 31, 31, 32, 27, 34, 49, 57, 48, 36, 
    22, 25, 40, 47, 42, 37, 31, 22, 26, 28, 32, 11, 32, 39, 41, 
    24, 26, 44, 43, 39, 51, 50, 29, 17, 33, 28, 29, 24, 27, 31, 
    32, 27, 39, 39, 42, 30, 39, 46, 38, 32, 24, 29, 35, 27, 27, 
    34, 25, 39, 50, 49, 40, 39, 41, 38, 20, 26, 31, 36, 29, 19, 
    29, 22, 34, 45, 40, 35, 47, 41, 35, 23, 27, 27, 32, 28, 22, 
    27, 16, 26, 44, 35, 41, 38, 33, 28, 16, 22, 22, 17, 21, 27, 
    24, 14, 19, 44, 38, 37, 30, 29, 18, 15, 18, 22, 15, 21, 25, 
    
    -- channel=550
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 10, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 7, 0, 6, 16, 0, 
    0, 0, 0, 0, 0, 6, 8, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 13, 8, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 7, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 9, 9, 7, 5, 0, 0, 9, 21, 8, 12, 0, 
    0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 1, 17, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 4, 0, 4, 6, 4, 0, 0, 0, 0, 0, 
    0, 1, 0, 8, 11, 5, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 9, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 9, 3, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=551
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=552
    14, 0, 0, 9, 0, 6, 8, 9, 20, 11, 0, 3, 6, 7, 8, 
    14, 0, 0, 8, 2, 3, 2, 4, 4, 31, 0, 6, 5, 3, 4, 
    15, 3, 0, 1, 0, 10, 0, 0, 0, 13, 0, 0, 2, 4, 9, 
    35, 26, 0, 13, 0, 11, 15, 10, 2, 0, 0, 0, 2, 2, 4, 
    32, 10, 8, 28, 0, 0, 2, 12, 0, 0, 0, 0, 1, 21, 4, 
    13, 7, 9, 20, 0, 0, 2, 12, 0, 0, 0, 0, 4, 23, 18, 
    14, 10, 8, 0, 0, 0, 1, 5, 6, 0, 0, 0, 4, 16, 27, 
    15, 7, 9, 0, 6, 0, 9, 0, 2, 6, 0, 0, 0, 1, 13, 
    20, 8, 8, 0, 6, 6, 3, 11, 0, 9, 0, 9, 0, 0, 0, 
    23, 17, 0, 0, 0, 0, 0, 15, 5, 0, 6, 4, 6, 3, 0, 
    14, 13, 0, 1, 3, 8, 0, 0, 9, 1, 10, 2, 0, 8, 1, 
    9, 20, 0, 0, 0, 10, 0, 1, 0, 19, 0, 3, 0, 6, 12, 
    12, 22, 6, 0, 0, 0, 0, 0, 4, 10, 0, 5, 0, 6, 5, 
    14, 21, 11, 0, 17, 0, 0, 0, 4, 13, 0, 4, 9, 0, 4, 
    15, 19, 14, 0, 4, 0, 8, 3, 8, 2, 6, 3, 13, 1, 3, 
    
    -- channel=553
    0, 0, 0, 0, 0, 0, 4, 6, 28, 9, 0, 23, 14, 10, 7, 
    0, 0, 0, 0, 19, 4, 0, 4, 0, 6, 29, 10, 6, 3, 1, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 21, 0, 0, 11, 15, 
    77, 61, 71, 0, 0, 13, 41, 15, 0, 0, 0, 2, 12, 0, 0, 
    38, 45, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 1, 4, 0, 0, 0, 18, 1, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 13, 0, 0, 0, 0, 12, 15, 
    0, 0, 0, 0, 10, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 4, 4, 32, 18, 8, 0, 0, 7, 0, 0, 0, 0, 
    6, 9, 1, 0, 0, 0, 0, 15, 30, 6, 0, 0, 11, 5, 0, 
    0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    
    -- channel=554
    5, 48, 75, 65, 60, 68, 74, 72, 54, 39, 47, 83, 85, 86, 84, 
    6, 32, 67, 53, 48, 56, 58, 69, 66, 28, 84, 76, 77, 80, 80, 
    8, 18, 59, 64, 52, 35, 37, 46, 36, 33, 78, 60, 64, 69, 72, 
    45, 41, 100, 57, 51, 37, 49, 42, 37, 56, 58, 68, 70, 69, 63, 
    58, 85, 68, 41, 58, 44, 45, 33, 35, 46, 58, 81, 71, 62, 73, 
    66, 68, 65, 49, 62, 48, 36, 24, 43, 47, 57, 73, 71, 64, 72, 
    69, 65, 57, 58, 47, 35, 39, 39, 48, 48, 54, 78, 73, 68, 68, 
    66, 63, 48, 70, 54, 50, 30, 54, 42, 55, 55, 64, 66, 71, 65, 
    61, 55, 49, 78, 48, 59, 51, 33, 59, 47, 57, 54, 61, 43, 71, 
    62, 66, 63, 60, 56, 49, 42, 43, 60, 58, 52, 53, 59, 63, 64, 
    65, 59, 56, 61, 62, 50, 54, 53, 44, 59, 41, 61, 60, 45, 53, 
    67, 55, 66, 57, 59, 46, 67, 59, 57, 37, 63, 53, 56, 53, 44, 
    66, 60, 67, 56, 45, 36, 63, 58, 49, 43, 56, 47, 50, 41, 50, 
    65, 62, 63, 56, 44, 73, 62, 52, 45, 38, 53, 47, 40, 51, 52, 
    54, 60, 58, 53, 51, 56, 44, 49, 39, 46, 46, 49, 43, 57, 48, 
    
    -- channel=555
    8, 0, 0, 8, 7, 0, 6, 0, 33, 82, 0, 0, 6, 5, 10, 
    6, 0, 0, 0, 3, 26, 0, 0, 12, 73, 0, 8, 13, 7, 7, 
    7, 0, 0, 0, 0, 73, 8, 0, 0, 0, 0, 0, 4, 2, 13, 
    101, 0, 0, 36, 0, 29, 52, 42, 0, 0, 0, 0, 9, 26, 0, 
    35, 0, 9, 61, 0, 0, 25, 50, 0, 0, 0, 0, 9, 53, 0, 
    10, 0, 9, 34, 0, 1, 33, 22, 5, 0, 0, 0, 7, 54, 12, 
    13, 2, 35, 0, 20, 0, 40, 0, 23, 0, 0, 0, 0, 21, 38, 
    23, 0, 61, 0, 26, 7, 10, 30, 0, 0, 5, 0, 0, 16, 0, 
    47, 0, 9, 0, 0, 13, 36, 58, 0, 13, 0, 41, 0, 0, 0, 
    29, 11, 0, 4, 0, 0, 0, 27, 61, 0, 26, 0, 0, 13, 0, 
    7, 37, 0, 9, 2, 48, 0, 0, 17, 39, 0, 0, 0, 21, 4, 
    4, 40, 0, 0, 14, 14, 0, 2, 17, 48, 0, 3, 0, 21, 21, 
    12, 24, 0, 1, 50, 0, 0, 1, 18, 23, 0, 2, 0, 0, 12, 
    17, 27, 0, 0, 39, 12, 16, 3, 15, 4, 0, 2, 20, 0, 0, 
    8, 11, 0, 0, 17, 28, 23, 0, 27, 0, 0, 0, 13, 0, 0, 
    
    -- channel=556
    17, 60, 3, 0, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 
    18, 48, 25, 0, 4, 2, 6, 6, 0, 0, 55, 0, 0, 0, 0, 
    16, 30, 40, 0, 25, 0, 8, 21, 3, 1, 40, 17, 3, 1, 0, 
    0, 11, 42, 0, 36, 0, 0, 0, 7, 39, 20, 27, 9, 11, 21, 
    0, 27, 11, 0, 38, 15, 0, 0, 16, 31, 26, 32, 12, 0, 29, 
    6, 16, 9, 0, 25, 16, 0, 0, 14, 28, 30, 39, 16, 0, 16, 
    7, 8, 0, 6, 7, 14, 0, 17, 7, 25, 27, 40, 18, 2, 1, 
    7, 10, 0, 25, 3, 18, 0, 19, 17, 17, 19, 41, 33, 14, 20, 
    0, 11, 0, 21, 7, 7, 4, 0, 26, 0, 4, 0, 41, 16, 41, 
    0, 11, 11, 8, 21, 23, 14, 0, 0, 12, 0, 0, 0, 0, 25, 
    12, 7, 21, 8, 10, 0, 27, 18, 0, 0, 0, 4, 6, 0, 3, 
    19, 0, 33, 12, 8, 0, 14, 6, 3, 0, 18, 3, 8, 0, 0, 
    16, 5, 30, 15, 0, 0, 15, 4, 0, 0, 15, 2, 9, 0, 0, 
    11, 6, 31, 21, 0, 0, 0, 0, 0, 0, 10, 4, 0, 14, 3, 
    12, 9, 27, 34, 5, 0, 0, 0, 0, 14, 5, 5, 0, 11, 6, 
    
    -- channel=557
    2, 0, 0, 6, 4, 0, 1, 0, 14, 73, 0, 0, 0, 0, 4, 
    2, 0, 0, 0, 0, 22, 0, 0, 5, 70, 0, 0, 5, 3, 4, 
    3, 0, 0, 0, 0, 65, 13, 0, 1, 0, 0, 0, 0, 0, 3, 
    57, 0, 0, 37, 0, 19, 38, 25, 0, 0, 0, 0, 3, 21, 0, 
    20, 0, 0, 59, 0, 0, 20, 48, 0, 0, 0, 0, 5, 48, 0, 
    4, 0, 3, 39, 0, 2, 31, 25, 0, 0, 0, 0, 3, 45, 6, 
    9, 3, 38, 0, 10, 0, 28, 0, 5, 0, 0, 0, 0, 11, 31, 
    22, 0, 62, 0, 19, 5, 6, 30, 0, 4, 8, 0, 0, 11, 0, 
    37, 0, 0, 0, 0, 0, 26, 37, 0, 28, 0, 44, 0, 0, 0, 
    17, 10, 0, 1, 0, 0, 0, 17, 52, 0, 18, 0, 0, 3, 0, 
    3, 36, 0, 4, 0, 40, 0, 0, 13, 29, 0, 0, 0, 20, 5, 
    2, 32, 0, 0, 10, 22, 0, 1, 14, 47, 0, 3, 0, 22, 17, 
    10, 18, 0, 0, 39, 18, 0, 7, 20, 29, 0, 7, 0, 0, 7, 
    17, 24, 0, 0, 27, 15, 8, 8, 20, 14, 0, 4, 19, 0, 0, 
    17, 6, 0, 0, 16, 22, 33, 0, 27, 0, 0, 0, 10, 0, 0, 
    
    -- channel=558
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=559
    6, 0, 7, 27, 29, 20, 28, 17, 42, 42, 0, 9, 22, 23, 29, 
    2, 0, 0, 0, 20, 24, 22, 16, 27, 88, 0, 30, 31, 27, 32, 
    2, 0, 0, 0, 0, 77, 21, 6, 44, 16, 0, 18, 32, 29, 34, 
    15, 0, 0, 43, 0, 53, 35, 29, 0, 0, 27, 0, 28, 53, 23, 
    55, 0, 29, 71, 0, 20, 46, 64, 3, 0, 5, 0, 37, 78, 7, 
    36, 19, 44, 48, 0, 25, 58, 33, 1, 0, 2, 0, 44, 82, 31, 
    39, 27, 54, 17, 15, 0, 44, 0, 30, 0, 0, 0, 32, 58, 52, 
    50, 28, 76, 0, 36, 25, 36, 16, 19, 3, 35, 6, 26, 53, 37, 
    71, 16, 33, 0, 32, 18, 21, 69, 0, 36, 26, 39, 0, 48, 0, 
    60, 21, 19, 26, 9, 23, 35, 46, 32, 0, 49, 20, 3, 23, 1, 
    42, 51, 6, 21, 22, 57, 0, 13, 59, 48, 26, 2, 13, 40, 20, 
    36, 69, 0, 27, 38, 52, 7, 19, 37, 74, 0, 22, 15, 36, 38, 
    44, 59, 0, 26, 67, 6, 5, 30, 50, 47, 0, 24, 21, 31, 23, 
    51, 61, 0, 18, 66, 4, 35, 32, 40, 31, 3, 18, 35, 0, 14, 
    54, 53, 0, 5, 43, 44, 59, 26, 47, 0, 14, 14, 27, 0, 17, 
    
    -- channel=560
    0, 0, 0, 0, 0, 0, 0, 0, 19, 12, 2, 6, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 1, 
    97, 91, 52, 0, 0, 0, 36, 8, 0, 0, 0, 0, 0, 0, 0, 
    15, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 16, 15, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 37, 2, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=561
    4, 40, 0, 0, 0, 0, 0, 2, 5, 0, 49, 10, 1, 0, 0, 
    5, 23, 0, 8, 20, 0, 0, 0, 0, 0, 76, 1, 0, 0, 0, 
    5, 9, 28, 19, 29, 0, 0, 0, 0, 16, 32, 0, 0, 4, 2, 
    43, 95, 67, 0, 18, 1, 18, 0, 11, 35, 0, 27, 5, 0, 0, 
    1, 37, 0, 0, 36, 0, 0, 0, 7, 21, 8, 19, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 0, 0, 20, 29, 7, 15, 0, 0, 0, 
    0, 0, 0, 6, 1, 18, 0, 23, 0, 15, 16, 14, 0, 0, 0, 
    0, 0, 0, 35, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 11, 24, 8, 25, 17, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 5, 3, 1, 0, 0, 0, 8, 10, 19, 0, 0, 20, 0, 0, 
    0, 0, 11, 5, 8, 0, 6, 0, 0, 0, 0, 10, 2, 0, 0, 
    0, 0, 21, 0, 0, 0, 10, 2, 0, 0, 20, 0, 1, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 2, 4, 0, 31, 0, 0, 0, 0, 0, 0, 0, 6, 3, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 8, 0, 0, 0, 5, 0, 
    
    -- channel=562
    0, 0, 15, 28, 25, 21, 23, 22, 29, 15, 0, 26, 29, 26, 28, 
    0, 0, 7, 24, 36, 27, 28, 24, 32, 36, 0, 33, 34, 31, 33, 
    0, 0, 0, 14, 38, 44, 22, 22, 32, 25, 14, 32, 40, 39, 38, 
    0, 0, 0, 26, 34, 50, 29, 23, 17, 12, 35, 29, 47, 43, 32, 
    30, 8, 27, 29, 20, 43, 44, 36, 19, 17, 30, 27, 43, 36, 14, 
    28, 25, 29, 27, 28, 41, 43, 29, 21, 18, 26, 28, 41, 33, 10, 
    25, 25, 31, 26, 27, 30, 40, 27, 34, 24, 27, 26, 40, 43, 25, 
    26, 28, 41, 26, 42, 35, 43, 27, 29, 24, 31, 27, 35, 42, 28, 
    26, 20, 46, 28, 44, 41, 39, 45, 13, 26, 30, 12, 9, 32, 19, 
    30, 21, 38, 37, 33, 43, 48, 47, 23, 22, 34, 24, 18, 24, 14, 
    30, 28, 32, 38, 37, 40, 29, 38, 48, 33, 24, 23, 28, 31, 22, 
    28, 30, 24, 47, 46, 46, 31, 36, 38, 36, 11, 27, 30, 29, 24, 
    26, 23, 18, 43, 49, 31, 33, 35, 37, 27, 16, 24, 27, 27, 21, 
    26, 17, 9, 40, 50, 29, 35, 27, 27, 19, 15, 19, 22, 12, 22, 
    22, 14, 4, 35, 42, 38, 32, 23, 22, 5, 16, 18, 19, 13, 21, 
    
    -- channel=563
    0, 0, 19, 27, 24, 17, 26, 31, 37, 31, 2, 42, 34, 36, 32, 
    0, 0, 4, 16, 44, 39, 26, 39, 38, 18, 50, 51, 42, 37, 33, 
    0, 0, 0, 30, 41, 44, 7, 4, 4, 14, 66, 42, 50, 54, 56, 
    56, 27, 80, 42, 31, 41, 53, 33, 16, 28, 47, 56, 67, 64, 46, 
    57, 78, 57, 31, 37, 36, 39, 27, 18, 23, 38, 71, 62, 55, 51, 
    54, 53, 51, 39, 49, 41, 29, 13, 39, 36, 39, 57, 68, 66, 58, 
    55, 45, 29, 37, 38, 22, 38, 24, 49, 41, 39, 62, 68, 73, 70, 
    56, 42, 25, 30, 55, 49, 28, 50, 20, 38, 44, 17, 46, 65, 58, 
    60, 34, 26, 50, 49, 67, 58, 33, 17, 26, 37, 32, 7, 12, 40, 
    63, 60, 52, 47, 44, 38, 40, 48, 57, 33, 25, 16, 32, 37, 25, 
    61, 59, 42, 52, 56, 46, 31, 37, 36, 37, 9, 35, 35, 19, 24, 
    59, 56, 50, 51, 51, 25, 52, 43, 42, 16, 31, 28, 31, 32, 22, 
    58, 52, 52, 51, 36, 0, 32, 31, 23, 16, 23, 20, 19, 10, 24, 
    54, 50, 46, 51, 42, 48, 32, 18, 13, 5, 22, 20, 15, 16, 26, 
    36, 45, 43, 44, 46, 42, 14, 13, 10, 14, 16, 22, 20, 28, 17, 
    
    -- channel=564
    9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=565
    0, 48, 15, 0, 0, 6, 0, 0, 0, 0, 40, 0, 0, 0, 0, 
    0, 27, 51, 18, 0, 0, 10, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 7, 56, 0, 12, 0, 16, 51, 44, 11, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 0, 0, 20, 6, 9, 0, 0, 25, 
    0, 0, 0, 0, 23, 9, 0, 0, 7, 20, 18, 4, 0, 0, 21, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 11, 32, 0, 0, 0, 
    0, 0, 0, 12, 0, 12, 0, 2, 0, 0, 5, 20, 3, 0, 0, 
    0, 9, 0, 34, 0, 0, 0, 0, 29, 0, 5, 76, 59, 5, 10, 
    0, 11, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 73, 66, 54, 
    0, 0, 0, 0, 12, 29, 16, 0, 0, 0, 0, 8, 0, 0, 32, 
    0, 0, 19, 0, 0, 0, 28, 17, 0, 0, 19, 0, 0, 0, 0, 
    4, 0, 20, 0, 0, 0, 0, 0, 0, 0, 2, 1, 4, 0, 0, 
    0, 0, 21, 2, 0, 35, 21, 11, 8, 0, 15, 6, 18, 22, 0, 
    0, 0, 30, 10, 0, 0, 0, 15, 11, 13, 7, 3, 0, 14, 0, 
    21, 4, 20, 31, 0, 0, 8, 18, 0, 12, 7, 1, 0, 0, 14, 
    
    -- channel=566
    0, 0, 27, 34, 35, 30, 39, 35, 40, 33, 0, 53, 50, 50, 48, 
    0, 0, 12, 19, 42, 49, 37, 47, 52, 34, 19, 61, 56, 53, 52, 
    0, 0, 0, 27, 38, 59, 22, 17, 23, 13, 55, 51, 61, 63, 64, 
    29, 0, 53, 54, 30, 53, 50, 36, 16, 20, 55, 52, 78, 80, 53, 
    60, 61, 62, 48, 26, 47, 55, 41, 16, 20, 45, 67, 75, 73, 52, 
    60, 57, 62, 45, 46, 54, 47, 20, 31, 27, 44, 57, 80, 79, 60, 
    63, 55, 58, 34, 41, 25, 49, 27, 53, 38, 40, 63, 78, 82, 76, 
    66, 52, 50, 27, 65, 54, 39, 53, 28, 46, 53, 45, 54, 82, 62, 
    69, 39, 39, 50, 54, 67, 61, 51, 26, 36, 45, 35, 19, 37, 46, 
    71, 59, 58, 55, 53, 54, 51, 56, 57, 32, 48, 26, 30, 47, 36, 
    68, 67, 45, 62, 62, 64, 39, 47, 55, 57, 16, 37, 42, 35, 33, 
    67, 66, 45, 63, 69, 52, 54, 53, 57, 39, 26, 38, 38, 42, 30, 
    67, 63, 48, 60, 63, 10, 42, 48, 44, 30, 25, 30, 34, 22, 31, 
    66, 59, 40, 57, 62, 46, 52, 34, 29, 15, 24, 25, 24, 16, 30, 
    49, 48, 40, 47, 59, 58, 39, 24, 24, 8, 22, 25, 24, 28, 26, 
    
    -- channel=567
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=568
    5, 0, 7, 37, 30, 24, 38, 27, 46, 71, 0, 20, 37, 38, 41, 
    4, 0, 0, 10, 10, 32, 12, 17, 30, 69, 0, 28, 36, 36, 39, 
    6, 0, 0, 20, 0, 61, 20, 0, 19, 1, 0, 8, 25, 23, 31, 
    65, 0, 0, 48, 0, 26, 44, 39, 6, 0, 8, 0, 19, 38, 4, 
    42, 16, 23, 65, 0, 3, 28, 50, 2, 0, 0, 0, 24, 59, 11, 
    29, 18, 29, 45, 0, 10, 35, 23, 8, 0, 0, 0, 25, 64, 35, 
    35, 25, 48, 12, 24, 0, 34, 0, 20, 0, 0, 0, 18, 36, 50, 
    42, 20, 69, 0, 29, 18, 11, 30, 0, 9, 22, 0, 0, 34, 19, 
    59, 17, 20, 0, 10, 16, 29, 45, 0, 33, 17, 57, 0, 12, 0, 
    42, 28, 11, 22, 7, 5, 3, 24, 58, 6, 35, 16, 19, 29, 12, 
    27, 48, 0, 19, 18, 46, 0, 7, 25, 46, 11, 12, 17, 32, 23, 
    25, 51, 0, 12, 25, 29, 9, 17, 28, 52, 0, 21, 8, 34, 32, 
    32, 40, 0, 12, 50, 8, 0, 22, 33, 39, 3, 21, 15, 13, 27, 
    37, 47, 2, 2, 36, 29, 29, 26, 33, 23, 9, 20, 30, 1, 14, 
    32, 36, 15, 0, 26, 35, 40, 19, 41, 7, 15, 15, 26, 14, 12, 
    
    -- channel=569
    0, 17, 34, 24, 28, 23, 22, 26, 20, 7, 32, 44, 31, 31, 27, 
    0, 7, 43, 31, 53, 41, 44, 48, 51, 14, 50, 56, 45, 42, 38, 
    0, 1, 36, 30, 77, 48, 37, 49, 43, 33, 72, 72, 67, 63, 56, 
    0, 3, 53, 39, 78, 63, 33, 29, 33, 54, 79, 80, 85, 83, 78, 
    45, 51, 66, 30, 69, 75, 63, 36, 39, 51, 77, 88, 88, 65, 69, 
    64, 67, 68, 36, 68, 73, 57, 34, 45, 52, 71, 96, 93, 67, 60, 
    64, 61, 54, 53, 57, 60, 56, 48, 60, 60, 68, 95, 96, 85, 62, 
    64, 59, 28, 69, 67, 68, 61, 53, 61, 59, 66, 83, 92, 94, 78, 
    60, 52, 41, 67, 74, 74, 64, 50, 50, 39, 57, 21, 67, 74, 83, 
    68, 56, 67, 66, 78, 88, 81, 62, 35, 49, 47, 35, 31, 45, 55, 
    78, 63, 75, 72, 74, 62, 74, 75, 65, 50, 32, 41, 48, 38, 38, 
    79, 63, 77, 81, 80, 57, 65, 65, 64, 30, 40, 45, 54, 39, 29, 
    74, 64, 71, 81, 66, 34, 69, 59, 51, 30, 42, 39, 49, 39, 34, 
    70, 56, 62, 84, 58, 31, 54, 43, 36, 23, 37, 34, 28, 33, 40, 
    60, 53, 52, 88, 70, 60, 37, 33, 23, 22, 31, 35, 25, 34, 39, 
    
    -- channel=570
    0, 0, 14, 16, 13, 11, 10, 3, 0, 2, 0, 0, 5, 6, 10, 
    0, 0, 25, 7, 0, 5, 14, 5, 19, 21, 0, 8, 11, 12, 16, 
    0, 0, 0, 0, 1, 26, 28, 38, 54, 0, 0, 17, 15, 7, 5, 
    0, 0, 0, 20, 17, 12, 0, 4, 0, 0, 24, 0, 7, 31, 18, 
    0, 0, 7, 23, 0, 21, 23, 29, 4, 0, 9, 1, 17, 31, 11, 
    11, 7, 24, 4, 0, 22, 41, 10, 0, 0, 7, 10, 21, 21, 7, 
    16, 10, 41, 14, 18, 4, 23, 0, 12, 0, 0, 7, 19, 14, 0, 
    20, 16, 34, 2, 10, 18, 15, 3, 19, 0, 29, 47, 38, 40, 6, 
    25, 12, 9, 0, 8, 0, 0, 29, 0, 13, 16, 6, 31, 63, 15, 
    15, 0, 12, 12, 21, 39, 25, 4, 0, 0, 39, 16, 0, 12, 28, 
    16, 17, 11, 8, 4, 32, 17, 22, 28, 37, 14, 0, 10, 24, 14, 
    18, 26, 0, 18, 28, 27, 3, 11, 24, 34, 0, 17, 14, 13, 14, 
    18, 26, 4, 21, 53, 23, 22, 29, 40, 23, 9, 16, 33, 26, 11, 
    22, 24, 3, 17, 25, 0, 33, 31, 32, 17, 9, 10, 18, 3, 5, 
    32, 19, 1, 22, 20, 29, 38, 27, 31, 0, 12, 8, 5, 0, 20, 
    
    -- channel=571
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 5, 9, 0, 
    0, 0, 0, 0, 0, 8, 1, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 2, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 4, 0, 0, 
    0, 0, 0, 0, 1, 4, 1, 4, 0, 0, 2, 13, 1, 7, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 6, 17, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=572
    3, 9, 6, 15, 14, 7, 6, 7, 0, 16, 5, 6, 8, 9, 9, 
    3, 11, 9, 23, 17, 22, 20, 15, 24, 14, 0, 14, 15, 15, 15, 
    3, 7, 0, 18, 35, 30, 31, 39, 39, 10, 15, 27, 23, 19, 15, 
    0, 0, 0, 26, 40, 26, 7, 12, 15, 25, 31, 24, 34, 39, 31, 
    0, 0, 18, 16, 30, 40, 34, 27, 20, 27, 27, 23, 33, 27, 25, 
    20, 25, 23, 17, 27, 41, 39, 25, 14, 22, 30, 29, 31, 15, 10, 
    19, 21, 34, 17, 29, 32, 32, 20, 26, 22, 30, 28, 35, 20, 8, 
    23, 25, 25, 21, 32, 34, 31, 35, 25, 32, 37, 54, 40, 41, 24, 
    16, 21, 15, 34, 28, 18, 28, 24, 27, 26, 19, 9, 45, 47, 30, 
    14, 14, 29, 28, 40, 55, 43, 23, 10, 18, 30, 16, 10, 17, 33, 
    22, 26, 27, 29, 27, 33, 36, 45, 30, 32, 20, 15, 22, 25, 23, 
    27, 20, 28, 38, 41, 33, 25, 31, 34, 24, 12, 26, 23, 23, 16, 
    24, 19, 24, 39, 42, 45, 34, 35, 35, 23, 19, 24, 35, 25, 16, 
    23, 15, 19, 33, 25, 13, 34, 29, 29, 20, 16, 20, 21, 17, 17, 
    27, 8, 21, 37, 32, 34, 32, 23, 22, 12, 18, 17, 12, 15, 23, 
    
    -- channel=573
    7, 16, 69, 61, 48, 65, 68, 64, 59, 30, 32, 66, 77, 76, 78, 
    8, 5, 62, 52, 34, 37, 50, 55, 56, 47, 33, 56, 64, 68, 72, 
    11, 6, 49, 47, 31, 29, 31, 37, 41, 38, 36, 44, 49, 50, 54, 
    29, 27, 46, 45, 32, 36, 33, 36, 33, 27, 40, 41, 44, 45, 45, 
    55, 43, 47, 47, 30, 30, 37, 34, 27, 24, 42, 45, 47, 51, 45, 
    51, 45, 50, 44, 37, 31, 33, 28, 27, 21, 33, 45, 46, 52, 51, 
    52, 50, 54, 50, 32, 25, 31, 30, 33, 27, 30, 46, 48, 52, 49, 
    49, 47, 53, 56, 37, 28, 32, 21, 41, 35, 35, 48, 48, 50, 44, 
    49, 41, 55, 43, 37, 38, 27, 38, 39, 38, 51, 42, 42, 47, 49, 
    51, 41, 41, 44, 34, 31, 32, 36, 32, 43, 50, 54, 45, 52, 42, 
    48, 39, 40, 41, 43, 40, 36, 34, 45, 48, 44, 47, 44, 46, 45, 
    45, 46, 37, 38, 42, 51, 43, 44, 43, 48, 44, 44, 46, 44, 44, 
    46, 51, 40, 36, 42, 39, 49, 48, 48, 44, 44, 42, 42, 44, 44, 
    48, 51, 39, 37, 44, 43, 52, 48, 46, 41, 44, 40, 41, 40, 46, 
    45, 52, 35, 33, 38, 43, 47, 48, 44, 35, 41, 43, 42, 42, 43, 
    
    -- channel=574
    0, 55, 0, 0, 0, 0, 0, 0, 0, 3, 45, 0, 0, 0, 0, 
    1, 48, 0, 19, 0, 4, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    1, 15, 0, 19, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 46, 0, 0, 0, 0, 10, 0, 0, 23, 0, 5, 0, 0, 0, 
    0, 6, 0, 3, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 16, 0, 18, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 13, 0, 25, 0, 0, 10, 0, 0, 0, 10, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 18, 
    0, 6, 0, 0, 0, 0, 2, 0, 15, 29, 0, 16, 0, 0, 5, 
    0, 14, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 59, 0, 0, 0, 1, 0, 2, 0, 0, 0, 
    0, 0, 16, 0, 0, 31, 0, 0, 0, 19, 0, 2, 0, 3, 0, 
    0, 0, 25, 0, 0, 0, 0, 0, 0, 18, 0, 0, 4, 0, 0, 
    
    -- channel=575
    0, 0, 0, 0, 1, 0, 0, 0, 11, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 7, 1, 0, 0, 0, 0, 4, 0, 0, 1, 0, 0, 
    0, 0, 16, 0, 0, 0, 7, 0, 3, 18, 0, 6, 0, 0, 0, 
    17, 28, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 5, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 19, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 7, 0, 0, 0, 0, 5, 0, 2, 0, 10, 5, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 10, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 
    
    -- channel=576
    1, 5, 0, 0, 3, 14, 14, 21, 16, 1, 0, 8, 0, 5, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 12, 0, 16, 2, 0, 18, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 44, 13, 0, 0, 25, 
    0, 0, 0, 0, 30, 7, 0, 0, 0, 0, 0, 29, 4, 0, 1, 
    2, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 37, 19, 0, 16, 
    16, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 19, 41, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 6, 18, 
    0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 9, 60, 
    0, 0, 36, 0, 19, 0, 5, 0, 26, 32, 0, 17, 25, 0, 61, 
    0, 0, 14, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 73, 
    0, 0, 4, 0, 0, 9, 26, 0, 36, 0, 0, 29, 0, 19, 51, 
    0, 0, 23, 6, 0, 0, 3, 0, 36, 1, 2, 0, 0, 0, 70, 
    0, 0, 0, 0, 0, 0, 0, 6, 18, 77, 0, 0, 0, 20, 61, 
    0, 0, 0, 0, 0, 0, 4, 10, 15, 14, 1, 0, 0, 24, 51, 
    0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 4, 0, 0, 20, 64, 
    
    -- channel=577
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 9, 0, 0, 0, 0, 0, 31, 23, 23, 34, 34, 2, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 4, 0, 0, 29, 0, 7, 0, 0, 10, 0, 0, 
    0, 0, 0, 12, 13, 5, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 32, 1, 0, 16, 1, 0, 0, 0, 2, 19, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 5, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 4, 1, 0, 0, 0, 7, 0, 0, 
    
    -- channel=578
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 5, 2, 9, 11, 5, 7, 0, 0, 17, 
    0, 0, 0, 0, 36, 11, 6, 0, 11, 23, 54, 2, 0, 0, 34, 
    0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 
    0, 0, 0, 0, 33, 2, 0, 0, 0, 0, 0, 31, 0, 0, 0, 
    5, 0, 0, 0, 39, 15, 0, 0, 4, 14, 6, 26, 43, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 26, 31, 14, 0, 
    0, 0, 39, 0, 0, 9, 22, 0, 8, 19, 4, 12, 47, 31, 63, 
    0, 0, 25, 0, 26, 0, 0, 0, 11, 4, 0, 3, 19, 0, 50, 
    0, 0, 31, 0, 30, 4, 33, 37, 0, 23, 3, 17, 16, 0, 80, 
    0, 0, 6, 0, 9, 37, 34, 0, 65, 2, 20, 49, 0, 20, 46, 
    0, 0, 49, 2, 0, 22, 39, 0, 55, 0, 2, 0, 0, 35, 84, 
    0, 0, 1, 0, 0, 0, 22, 29, 37, 68, 0, 0, 0, 39, 73, 
    0, 0, 0, 0, 2, 0, 23, 26, 25, 45, 30, 0, 0, 48, 63, 
    0, 0, 0, 0, 10, 0, 17, 21, 24, 25, 25, 0, 0, 46, 80, 
    
    -- channel=579
    0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 41, 47, 59, 75, 72, 47, 22, 0, 2, 5, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 6, 5, 0, 1, 19, 16, 
    0, 0, 3, 10, 0, 0, 0, 5, 0, 0, 0, 22, 0, 0, 8, 
    0, 0, 40, 32, 0, 20, 23, 2, 7, 8, 0, 0, 0, 0, 0, 
    11, 14, 0, 0, 16, 0, 0, 17, 18, 7, 25, 16, 0, 0, 0, 
    4, 26, 21, 0, 0, 0, 10, 0, 5, 20, 20, 30, 52, 58, 7, 
    10, 40, 3, 0, 16, 0, 0, 9, 38, 33, 26, 49, 42, 23, 5, 
    0, 1, 0, 49, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 15, 28, 8, 17, 11, 18, 36, 26, 27, 37, 31, 30, 26, 8, 
    0, 1, 0, 0, 0, 8, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    8, 28, 11, 0, 0, 5, 50, 41, 28, 31, 0, 27, 44, 29, 18, 
    2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 7, 0, 2, 2, 0, 0, 0, 0, 28, 38, 16, 7, 0, 0, 
    7, 0, 0, 9, 3, 0, 0, 0, 0, 0, 13, 14, 0, 0, 0, 
    
    -- channel=580
    49, 51, 42, 10, 34, 44, 56, 71, 67, 51, 43, 50, 44, 47, 32, 
    57, 58, 41, 0, 1, 6, 0, 0, 14, 29, 30, 51, 44, 21, 53, 
    52, 52, 34, 0, 11, 14, 16, 7, 0, 0, 53, 57, 31, 8, 42, 
    52, 44, 30, 0, 44, 49, 6, 5, 14, 27, 16, 45, 40, 31, 22, 
    53, 42, 0, 0, 23, 1, 0, 4, 9, 12, 13, 61, 67, 46, 63, 
    52, 28, 14, 0, 0, 0, 0, 0, 0, 0, 0, 14, 63, 52, 53, 
    39, 0, 0, 0, 22, 1, 0, 0, 8, 9, 0, 8, 20, 32, 59, 
    25, 0, 39, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 71, 
    35, 0, 31, 0, 5, 8, 19, 7, 40, 57, 37, 38, 51, 17, 67, 
    28, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 54, 
    33, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 12, 0, 15, 47, 
    25, 0, 4, 13, 0, 0, 0, 0, 13, 3, 16, 7, 0, 0, 39, 
    20, 0, 17, 0, 0, 0, 0, 0, 0, 84, 53, 0, 0, 0, 53, 
    27, 6, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 41, 
    9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 
    
    -- channel=581
    12, 12, 3, 0, 0, 22, 44, 61, 30, 3, 0, 0, 21, 19, 10, 
    4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 28, 28, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 14, 23, 4, 0, 5, 25, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 10, 21, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 49, 0, 0, 0, 8, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 10, 0, 0, 0, 4, 21, 52, 99, 106, 113, 109, 78, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 2, 0, 0, 0, 29, 0, 0, 0, 0, 2, 0, 13, 3, 
    0, 0, 0, 37, 17, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 50, 52, 0, 9, 9, 0, 0, 0, 64, 67, 39, 0, 0, 10, 
    0, 0, 0, 0, 0, 5, 10, 11, 18, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 10, 8, 0, 0, 0, 0, 4, 0, 7, 
    
    -- channel=582
    31, 41, 29, 20, 8, 20, 35, 59, 59, 35, 38, 24, 28, 51, 25, 
    34, 35, 30, 4, 0, 0, 0, 0, 0, 0, 8, 26, 26, 29, 27, 
    29, 28, 18, 0, 0, 0, 0, 2, 0, 0, 0, 34, 33, 13, 19, 
    28, 30, 10, 0, 0, 10, 22, 0, 0, 0, 34, 0, 9, 35, 37, 
    26, 25, 14, 0, 0, 0, 0, 0, 0, 0, 0, 19, 34, 24, 41, 
    12, 20, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 29, 
    17, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    21, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 1, 26, 0, 0, 3, 0, 1, 31, 46, 46, 43, 56, 25, 17, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 4, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 25, 
    3, 0, 0, 4, 1, 0, 0, 0, 5, 0, 4, 18, 0, 0, 0, 
    0, 0, 45, 0, 0, 0, 0, 0, 0, 18, 53, 26, 0, 0, 21, 
    7, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    
    -- channel=583
    33, 29, 36, 32, 33, 31, 36, 40, 50, 49, 47, 40, 32, 41, 28, 
    41, 41, 56, 42, 42, 36, 29, 46, 61, 55, 41, 40, 43, 52, 37, 
    40, 40, 45, 11, 0, 0, 0, 0, 0, 1, 20, 41, 49, 51, 36, 
    38, 46, 20, 30, 10, 28, 21, 3, 0, 0, 28, 34, 30, 49, 40, 
    39, 47, 43, 6, 9, 2, 5, 0, 8, 0, 16, 28, 40, 33, 8, 
    34, 59, 5, 8, 0, 0, 0, 1, 0, 0, 9, 2, 20, 39, 39, 
    28, 39, 16, 0, 0, 1, 12, 0, 7, 38, 16, 17, 41, 40, 43, 
    47, 18, 0, 46, 0, 0, 0, 0, 5, 0, 1, 16, 0, 0, 27, 
    30, 11, 27, 6, 0, 22, 8, 0, 0, 0, 8, 0, 0, 18, 20, 
    27, 16, 34, 0, 3, 0, 0, 0, 20, 0, 7, 0, 26, 0, 0, 
    27, 13, 4, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    29, 19, 2, 0, 2, 0, 4, 2, 13, 25, 19, 51, 0, 13, 0, 
    10, 0, 0, 29, 0, 0, 0, 0, 0, 13, 43, 58, 1, 0, 0, 
    14, 23, 9, 34, 4, 4, 0, 0, 4, 20, 1, 44, 0, 0, 0, 
    12, 6, 15, 8, 4, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    
    -- channel=584
    39, 34, 44, 34, 20, 23, 26, 27, 29, 35, 32, 29, 49, 26, 35, 
    43, 42, 53, 39, 3, 0, 0, 0, 0, 3, 16, 24, 32, 36, 9, 
    42, 41, 53, 72, 0, 19, 16, 28, 15, 1, 0, 30, 40, 35, 0, 
    42, 46, 39, 70, 0, 17, 38, 18, 23, 18, 21, 0, 44, 47, 10, 
    39, 51, 29, 43, 0, 0, 20, 8, 11, 9, 36, 0, 28, 64, 44, 
    22, 52, 46, 50, 0, 1, 10, 0, 1, 0, 0, 0, 0, 43, 41, 
    22, 45, 15, 39, 0, 4, 19, 6, 0, 4, 6, 0, 0, 0, 35, 
    34, 29, 0, 34, 2, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 42, 0, 13, 0, 0, 11, 34, 21, 13, 53, 28, 1, 9, 0, 
    49, 49, 0, 6, 0, 0, 0, 0, 22, 0, 6, 0, 0, 15, 0, 
    35, 65, 2, 0, 0, 0, 0, 10, 0, 12, 4, 0, 3, 2, 0, 
    35, 58, 0, 16, 17, 0, 0, 7, 0, 5, 8, 0, 24, 0, 0, 
    26, 76, 0, 17, 21, 0, 0, 0, 0, 0, 36, 63, 0, 0, 0, 
    20, 34, 37, 12, 0, 17, 0, 0, 0, 0, 0, 60, 0, 0, 0, 
    24, 25, 38, 9, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 
    
    -- channel=585
    0, 0, 0, 0, 8, 0, 0, 0, 3, 4, 2, 6, 0, 0, 0, 
    5, 4, 6, 0, 33, 44, 37, 45, 58, 41, 8, 12, 6, 0, 6, 
    9, 10, 1, 0, 15, 3, 3, 0, 0, 13, 33, 2, 0, 0, 8, 
    9, 10, 1, 0, 50, 35, 12, 37, 30, 19, 10, 36, 0, 0, 0, 
    11, 8, 6, 13, 39, 36, 36, 34, 37, 34, 26, 26, 12, 0, 0, 
    22, 14, 1, 0, 24, 26, 23, 35, 33, 36, 38, 28, 33, 9, 9, 
    12, 2, 7, 0, 4, 25, 35, 20, 35, 41, 21, 34, 45, 44, 28, 
    10, 0, 21, 0, 20, 0, 0, 18, 31, 24, 25, 40, 38, 32, 49, 
    0, 0, 18, 0, 29, 22, 18, 0, 0, 0, 0, 0, 0, 13, 35, 
    0, 0, 27, 0, 12, 10, 13, 44, 17, 26, 26, 24, 38, 6, 38, 
    6, 0, 0, 0, 0, 7, 0, 0, 19, 0, 2, 0, 0, 26, 12, 
    17, 0, 18, 0, 0, 2, 33, 13, 34, 28, 10, 34, 7, 15, 38, 
    18, 0, 0, 15, 0, 0, 0, 0, 0, 39, 0, 0, 0, 2, 21, 
    21, 15, 6, 15, 10, 0, 0, 0, 10, 20, 34, 7, 0, 8, 26, 
    20, 16, 5, 0, 10, 0, 0, 0, 0, 6, 21, 8, 0, 3, 29, 
    
    -- channel=586
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=587
    96, 94, 89, 46, 64, 81, 96, 119, 101, 85, 75, 83, 101, 80, 79, 
    100, 101, 83, 15, 2, 7, 0, 0, 0, 23, 48, 79, 75, 49, 75, 
    94, 94, 77, 45, 63, 83, 89, 82, 52, 25, 57, 87, 63, 34, 37, 
    94, 85, 78, 31, 74, 89, 70, 61, 80, 91, 45, 52, 85, 75, 34, 
    93, 86, 17, 24, 48, 39, 40, 54, 57, 64, 72, 72, 98, 105, 131, 
    80, 64, 90, 28, 4, 46, 38, 25, 20, 38, 21, 38, 87, 95, 94, 
    66, 29, 25, 69, 73, 46, 44, 37, 47, 31, 19, 14, 5, 30, 93, 
    47, 0, 64, 36, 22, 27, 17, 0, 0, 0, 0, 0, 0, 23, 75, 
    81, 40, 41, 0, 47, 32, 67, 75, 127, 136, 120, 122, 115, 60, 60, 
    79, 10, 0, 15, 0, 2, 0, 17, 11, 8, 0, 2, 6, 4, 63, 
    74, 35, 23, 12, 0, 0, 69, 0, 25, 28, 30, 74, 0, 73, 59, 
    63, 0, 8, 72, 9, 0, 0, 0, 0, 26, 48, 6, 0, 0, 57, 
    67, 111, 61, 29, 30, 0, 0, 0, 6, 108, 102, 52, 0, 16, 65, 
    72, 49, 45, 13, 21, 3, 0, 5, 15, 0, 15, 2, 0, 13, 61, 
    54, 60, 49, 0, 9, 4, 7, 9, 8, 10, 6, 7, 0, 9, 88, 
    
    -- channel=588
    0, 0, 0, 0, 0, 0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 4, 
    0, 0, 0, 0, 14, 4, 0, 0, 0, 18, 48, 0, 0, 0, 26, 
    0, 0, 0, 0, 61, 0, 0, 0, 0, 0, 5, 29, 0, 0, 0, 
    0, 0, 0, 0, 31, 13, 0, 0, 0, 0, 0, 47, 0, 0, 0, 
    6, 0, 0, 0, 28, 0, 0, 0, 0, 9, 3, 18, 48, 0, 0, 
    8, 0, 0, 0, 11, 3, 0, 0, 10, 0, 0, 29, 27, 9, 0, 
    0, 0, 34, 0, 0, 0, 3, 0, 0, 0, 0, 6, 23, 31, 64, 
    0, 0, 41, 0, 22, 11, 0, 0, 17, 30, 0, 2, 49, 3, 75, 
    0, 0, 8, 0, 22, 0, 17, 52, 0, 10, 0, 0, 0, 0, 111, 
    0, 0, 1, 0, 0, 16, 22, 0, 33, 0, 0, 26, 0, 10, 88, 
    0, 0, 18, 0, 0, 15, 41, 0, 89, 0, 0, 18, 0, 12, 106, 
    0, 0, 26, 0, 0, 0, 1, 9, 28, 88, 0, 0, 0, 17, 112, 
    2, 0, 0, 0, 0, 0, 3, 16, 26, 40, 8, 0, 0, 48, 85, 
    0, 0, 0, 0, 0, 0, 0, 4, 11, 16, 23, 0, 0, 34, 103, 
    
    -- channel=589
    0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 4, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 19, 5, 0, 0, 3, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 10, 5, 0, 5, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 
    10, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 5, 
    13, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 30, 
    2, 0, 22, 0, 9, 0, 0, 0, 9, 2, 0, 5, 8, 0, 18, 
    1, 0, 19, 0, 2, 0, 0, 5, 0, 0, 0, 0, 5, 0, 25, 
    3, 0, 0, 0, 0, 6, 14, 0, 25, 0, 3, 23, 0, 11, 7, 
    0, 0, 23, 3, 0, 0, 0, 0, 9, 0, 3, 0, 0, 3, 23, 
    0, 0, 0, 3, 0, 0, 0, 2, 3, 36, 0, 0, 0, 10, 21, 
    0, 0, 0, 3, 0, 0, 0, 2, 6, 7, 5, 0, 0, 12, 17, 
    0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 6, 0, 0, 12, 25, 
    
    -- channel=590
    2, 4, 1, 3, 9, 0, 0, 0, 0, 7, 9, 12, 1, 5, 6, 
    0, 1, 0, 0, 1, 1, 5, 11, 17, 26, 22, 14, 13, 16, 22, 
    2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 21, 7, 8, 20, 34, 
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 9, 3, 16, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 2, 
    7, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 20, 10, 
    7, 4, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 4, 0, 1, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=591
    18, 14, 19, 11, 22, 20, 23, 14, 17, 21, 14, 20, 16, 2, 10, 
    28, 27, 30, 37, 52, 56, 51, 56, 55, 33, 20, 15, 18, 5, 7, 
    30, 30, 37, 36, 61, 59, 60, 59, 59, 41, 26, 19, 11, 7, 1, 
    30, 31, 29, 61, 57, 69, 70, 84, 78, 73, 32, 25, 21, 5, 0, 
    29, 32, 44, 71, 67, 63, 84, 79, 75, 74, 73, 33, 27, 26, 5, 
    27, 35, 36, 48, 52, 67, 65, 70, 70, 62, 65, 42, 27, 30, 30, 
    19, 31, 20, 43, 54, 66, 79, 64, 66, 71, 49, 39, 42, 46, 36, 
    18, 17, 15, 28, 58, 42, 37, 36, 40, 42, 33, 36, 50, 46, 38, 
    17, 21, 4, 38, 38, 35, 50, 40, 9, 12, 28, 9, 15, 40, 35, 
    27, 20, 28, 17, 35, 36, 31, 35, 56, 48, 55, 51, 56, 45, 23, 
    29, 34, 10, 25, 12, 29, 32, 15, 36, 26, 31, 27, 23, 38, 20, 
    46, 31, 32, 26, 16, 8, 19, 38, 13, 44, 38, 30, 35, 32, 21, 
    53, 41, 13, 42, 32, 9, 10, 12, 11, 24, 36, 40, 15, 22, 23, 
    46, 55, 42, 43, 35, 21, 6, 9, 16, 33, 48, 49, 13, 17, 35, 
    60, 56, 48, 36, 31, 23, 12, 15, 18, 24, 31, 47, 9, 18, 31, 
    
    -- channel=592
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 10, 13, 18, 22, 8, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 24, 4, 0, 0, 0, 16, 26, 0, 0, 0, 10, 0, 
    0, 0, 3, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 24, 0, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 11, 9, 2, 0, 11, 8, 0, 12, 0, 0, 0, 
    0, 17, 13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 12, 2, 0, 
    0, 32, 0, 0, 12, 39, 32, 12, 6, 16, 8, 0, 20, 19, 0, 
    0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 2, 10, 0, 21, 27, 0, 30, 33, 37, 37, 12, 32, 0, 
    0, 5, 0, 5, 7, 1, 0, 4, 21, 24, 26, 12, 17, 0, 0, 
    0, 33, 0, 0, 0, 2, 14, 29, 0, 0, 0, 0, 26, 23, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 5, 0, 0, 5, 0, 0, 0, 13, 29, 30, 9, 0, 0, 
    2, 1, 3, 8, 0, 2, 0, 0, 0, 1, 3, 12, 1, 0, 0, 
    
    -- channel=593
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 0, 10, 10, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 0, 4, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=594
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=595
    55, 49, 61, 39, 36, 36, 45, 49, 47, 51, 45, 42, 64, 43, 50, 
    55, 54, 66, 40, 18, 12, 0, 0, 8, 15, 28, 38, 44, 49, 29, 
    52, 51, 65, 73, 24, 46, 41, 54, 40, 18, 4, 49, 50, 45, 1, 
    52, 59, 42, 83, 4, 34, 50, 37, 47, 41, 36, 13, 52, 64, 19, 
    48, 62, 35, 50, 16, 11, 33, 28, 29, 21, 59, 17, 42, 82, 61, 
    26, 62, 48, 62, 0, 21, 27, 17, 18, 16, 13, 8, 19, 52, 52, 
    25, 46, 14, 43, 25, 19, 43, 23, 14, 31, 17, 0, 0, 0, 43, 
    41, 17, 0, 53, 17, 27, 13, 15, 0, 0, 0, 0, 0, 0, 10, 
    50, 42, 5, 4, 11, 2, 24, 57, 54, 36, 91, 64, 31, 28, 0, 
    56, 48, 5, 10, 0, 13, 0, 0, 29, 1, 16, 11, 22, 14, 0, 
    42, 68, 17, 20, 0, 0, 14, 27, 0, 29, 23, 27, 13, 25, 0, 
    43, 56, 0, 40, 33, 0, 0, 18, 0, 12, 33, 9, 16, 0, 0, 
    37, 93, 24, 43, 40, 20, 0, 0, 0, 6, 61, 95, 9, 0, 0, 
    35, 44, 49, 41, 19, 36, 1, 0, 0, 0, 0, 81, 7, 0, 0, 
    35, 41, 58, 21, 14, 21, 6, 6, 1, 0, 0, 48, 11, 0, 0, 
    
    -- channel=596
    4, 13, 0, 0, 0, 5, 6, 16, 18, 5, 10, 10, 0, 20, 2, 
    4, 5, 0, 0, 0, 0, 9, 0, 0, 6, 11, 16, 7, 0, 23, 
    4, 5, 0, 0, 0, 0, 0, 0, 0, 11, 34, 10, 2, 0, 41, 
    4, 0, 3, 0, 17, 0, 0, 0, 0, 0, 12, 25, 0, 0, 25, 
    5, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 30, 12, 0, 10, 
    14, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 18, 31, 4, 4, 
    17, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 22, 23, 18, 3, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 20, 30, 
    0, 0, 28, 0, 1, 9, 0, 0, 3, 22, 0, 0, 28, 2, 54, 
    0, 0, 0, 0, 14, 0, 15, 36, 0, 6, 0, 0, 0, 0, 75, 
    0, 0, 4, 0, 7, 12, 8, 0, 15, 0, 0, 6, 5, 0, 73, 
    0, 0, 3, 0, 0, 17, 34, 0, 60, 0, 0, 10, 0, 6, 78, 
    0, 0, 22, 0, 0, 0, 4, 8, 25, 33, 0, 0, 0, 12, 77, 
    0, 0, 0, 0, 0, 0, 6, 13, 18, 30, 6, 0, 0, 31, 58, 
    0, 0, 0, 0, 0, 0, 4, 4, 10, 11, 14, 0, 0, 21, 62, 
    
    -- channel=597
    0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 13, 7, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 27, 24, 20, 23, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 35, 25, 22, 15, 17, 20, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 37, 20, 11, 24, 21, 17, 8, 12, 0, 0, 0, 
    0, 0, 0, 15, 34, 24, 21, 25, 24, 19, 17, 13, 0, 0, 0, 
    10, 0, 11, 4, 40, 34, 28, 30, 32, 33, 18, 17, 9, 0, 0, 
    16, 3, 16, 23, 23, 18, 18, 17, 28, 28, 21, 30, 34, 19, 7, 
    9, 5, 33, 8, 26, 27, 28, 26, 24, 30, 26, 25, 39, 30, 28, 
    0, 0, 28, 5, 38, 18, 26, 16, 23, 12, 10, 12, 15, 8, 23, 
    3, 0, 28, 19, 23, 28, 31, 22, 28, 16, 17, 21, 16, 21, 33, 
    9, 0, 27, 26, 18, 27, 27, 3, 40, 17, 26, 26, 0, 32, 20, 
    15, 0, 32, 26, 11, 18, 27, 29, 28, 30, 24, 14, 20, 30, 41, 
    15, 14, 9, 24, 22, 13, 25, 28, 32, 40, 8, 0, 11, 37, 36, 
    15, 13, 11, 19, 23, 18, 24, 26, 28, 29, 30, 15, 19, 34, 35, 
    
    -- channel=598
    4, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 22, 28, 22, 27, 22, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 8, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 39, 40, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 8, 47, 25, 14, 43, 32, 0, 0, 
    0, 0, 0, 1, 0, 1, 5, 0, 0, 5, 0, 0, 0, 0, 2, 
    0, 0, 9, 3, 5, 0, 23, 4, 25, 38, 37, 56, 13, 13, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 29, 10, 0, 5, 3, 0, 0, 8, 0, 0, 0, 0, 4, 5, 
    0, 0, 0, 0, 0, 0, 7, 2, 0, 0, 0, 0, 0, 1, 1, 
    0, 0, 0, 0, 0, 0, 6, 7, 6, 4, 0, 0, 0, 7, 22, 
    
    -- channel=599
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=600
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 26, 12, 37, 6, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 66, 2, 11, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 14, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=601
    0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 74, 14, 0, 10, 16, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 15, 84, 0, 0, 0, 3, 8, 1, 0, 0, 20, 18, 0, 
    0, 3, 0, 93, 0, 0, 43, 0, 0, 0, 18, 0, 0, 23, 12, 
    0, 6, 63, 43, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 1, 87, 0, 0, 18, 8, 4, 0, 2, 0, 0, 0, 0, 
    0, 40, 16, 3, 2, 14, 11, 10, 0, 14, 16, 0, 0, 0, 0, 
    22, 68, 0, 64, 11, 2, 13, 33, 20, 3, 22, 13, 0, 0, 0, 
    19, 58, 0, 72, 0, 12, 0, 2, 0, 0, 7, 0, 0, 22, 0, 
    9, 98, 0, 23, 7, 9, 6, 0, 17, 1, 15, 3, 6, 27, 0, 
    1, 81, 12, 12, 24, 0, 0, 79, 0, 27, 0, 0, 67, 0, 0, 
    10, 110, 0, 0, 53, 16, 5, 13, 0, 0, 0, 31, 34, 18, 0, 
    0, 6, 21, 15, 15, 42, 7, 0, 0, 0, 10, 65, 49, 0, 0, 
    0, 21, 29, 24, 7, 36, 4, 0, 0, 0, 0, 65, 20, 0, 0, 
    7, 2, 27, 44, 6, 16, 6, 1, 0, 0, 0, 22, 36, 0, 0, 
    
    -- channel=602
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=603
    0, 0, 0, 0, 0, 5, 13, 18, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 9, 
    0, 0, 0, 0, 27, 13, 1, 0, 0, 0, 43, 10, 0, 0, 16, 
    0, 0, 0, 0, 66, 17, 0, 0, 0, 9, 0, 28, 0, 0, 0, 
    0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 47, 5, 0, 5, 
    4, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 2, 45, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 7, 0, 0, 10, 12, 0, 0, 
    0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 73, 
    0, 0, 32, 0, 26, 4, 0, 0, 39, 40, 1, 31, 50, 0, 66, 
    0, 0, 23, 0, 19, 0, 0, 18, 0, 0, 0, 0, 0, 0, 78, 
    0, 0, 0, 0, 0, 17, 31, 0, 40, 0, 0, 37, 0, 20, 51, 
    0, 0, 40, 11, 0, 0, 5, 0, 60, 0, 7, 5, 0, 10, 62, 
    0, 0, 11, 2, 0, 0, 0, 6, 17, 115, 0, 0, 0, 22, 76, 
    0, 0, 0, 0, 0, 0, 5, 14, 20, 28, 0, 0, 0, 37, 59, 
    0, 0, 0, 0, 0, 0, 0, 5, 7, 8, 9, 0, 0, 30, 81, 
    
    -- channel=604
    11, 0, 12, 0, 20, 12, 21, 8, 1, 16, 4, 17, 23, 0, 17, 
    9, 7, 13, 0, 0, 0, 0, 0, 11, 25, 14, 7, 13, 11, 19, 
    6, 5, 20, 0, 3, 0, 0, 0, 0, 0, 5, 14, 0, 18, 0, 
    6, 10, 0, 20, 0, 23, 0, 0, 4, 0, 0, 10, 28, 13, 0, 
    8, 13, 0, 22, 0, 0, 8, 0, 0, 0, 16, 0, 13, 36, 1, 
    8, 16, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 6, 
    0, 9, 0, 28, 0, 0, 17, 0, 0, 9, 0, 0, 0, 2, 28, 
    12, 0, 18, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    3, 0, 0, 0, 10, 0, 26, 26, 0, 0, 36, 0, 0, 0, 0, 
    16, 0, 17, 0, 0, 0, 0, 0, 5, 0, 0, 0, 1, 0, 0, 
    5, 16, 0, 6, 0, 0, 2, 0, 12, 0, 0, 4, 0, 23, 0, 
    0, 0, 27, 7, 0, 0, 0, 44, 0, 37, 17, 0, 14, 0, 0, 
    3, 47, 0, 17, 17, 0, 0, 0, 0, 29, 20, 46, 0, 0, 0, 
    0, 6, 6, 21, 0, 10, 0, 0, 0, 0, 0, 41, 0, 0, 0, 
    0, 0, 8, 0, 0, 7, 0, 0, 0, 0, 0, 46, 0, 0, 0, 
    
    -- channel=605
    11, 9, 20, 32, 4, 2, 3, 0, 0, 5, 8, 0, 26, 6, 21, 
    7, 6, 27, 60, 0, 0, 0, 0, 0, 0, 0, 0, 1, 24, 0, 
    4, 3, 32, 108, 0, 8, 8, 26, 12, 0, 0, 0, 21, 26, 0, 
    5, 15, 14, 109, 0, 0, 35, 0, 6, 0, 0, 0, 13, 40, 3, 
    0, 20, 38, 63, 0, 0, 13, 0, 0, 0, 13, 0, 0, 43, 21, 
    0, 31, 38, 84, 0, 0, 9, 0, 0, 0, 0, 0, 0, 5, 3, 
    0, 41, 10, 39, 4, 1, 17, 9, 0, 0, 9, 0, 0, 0, 0, 
    21, 49, 0, 59, 7, 18, 6, 16, 0, 0, 0, 0, 0, 0, 0, 
    34, 70, 0, 52, 0, 0, 2, 45, 21, 6, 66, 37, 0, 8, 0, 
    32, 92, 0, 37, 0, 14, 0, 0, 16, 0, 3, 0, 0, 25, 0, 
    13, 107, 10, 23, 12, 0, 0, 50, 0, 27, 7, 0, 36, 0, 0, 
    15, 110, 0, 16, 57, 0, 0, 33, 0, 0, 5, 0, 52, 0, 0, 
    4, 82, 15, 16, 42, 39, 2, 0, 0, 0, 27, 89, 37, 0, 0, 
    0, 24, 42, 24, 8, 51, 6, 0, 0, 0, 0, 81, 27, 0, 0, 
    9, 13, 43, 33, 4, 24, 9, 4, 0, 0, 0, 36, 34, 0, 0, 
    
    -- channel=606
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=607
    36, 31, 41, 41, 29, 33, 28, 19, 19, 31, 27, 27, 41, 19, 30, 
    41, 39, 47, 60, 42, 42, 39, 40, 31, 22, 22, 21, 30, 30, 8, 
    43, 42, 56, 89, 60, 73, 75, 81, 74, 48, 11, 29, 35, 29, 0, 
    43, 46, 49, 101, 34, 57, 79, 80, 80, 73, 44, 14, 42, 36, 10, 
    40, 49, 56, 91, 50, 57, 83, 74, 69, 68, 77, 26, 30, 57, 37, 
    30, 51, 61, 88, 44, 67, 74, 66, 68, 61, 59, 40, 22, 43, 42, 
    32, 58, 39, 72, 53, 66, 79, 68, 55, 58, 52, 24, 21, 27, 35, 
    38, 55, 17, 56, 65, 72, 62, 56, 41, 44, 42, 28, 31, 40, 19, 
    48, 63, 8, 69, 37, 33, 50, 70, 43, 34, 65, 45, 30, 50, 10, 
    54, 71, 24, 46, 29, 51, 36, 20, 63, 50, 61, 55, 51, 65, 0, 
    48, 86, 31, 44, 34, 30, 40, 54, 33, 62, 55, 46, 62, 41, 9, 
    58, 87, 25, 44, 54, 18, 9, 57, 0, 41, 42, 24, 61, 31, 0, 
    63, 92, 34, 52, 60, 39, 20, 20, 19, 0, 45, 73, 43, 23, 0, 
    55, 69, 70, 54, 46, 54, 22, 18, 14, 17, 42, 83, 38, 10, 14, 
    67, 68, 73, 58, 41, 45, 28, 28, 28, 31, 32, 68, 39, 17, 7, 
    
    -- channel=608
    0, 0, 0, 0, 0, 0, 2, 5, 8, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 19, 14, 30, 30, 7, 16, 0, 0, 27, 
    0, 0, 0, 0, 32, 0, 0, 0, 0, 9, 81, 11, 0, 0, 49, 
    0, 0, 0, 0, 79, 29, 0, 0, 0, 8, 0, 62, 0, 0, 0, 
    0, 0, 0, 0, 52, 21, 0, 9, 11, 13, 0, 65, 19, 0, 0, 
    29, 0, 0, 0, 54, 16, 0, 5, 7, 19, 21, 50, 73, 0, 0, 
    17, 0, 0, 0, 4, 0, 0, 0, 19, 1, 0, 49, 59, 50, 19, 
    0, 0, 70, 0, 0, 0, 0, 0, 13, 22, 0, 26, 75, 48, 107, 
    0, 0, 47, 0, 38, 15, 5, 0, 0, 7, 0, 0, 21, 0, 120, 
    0, 0, 39, 0, 40, 0, 27, 74, 0, 19, 0, 7, 14, 0, 149, 
    0, 0, 0, 0, 0, 41, 38, 0, 78, 0, 0, 39, 0, 24, 108, 
    0, 0, 59, 0, 0, 10, 56, 0, 102, 2, 3, 14, 0, 28, 153, 
    1, 0, 0, 0, 0, 0, 3, 15, 37, 118, 0, 0, 0, 40, 134, 
    4, 0, 0, 0, 0, 0, 0, 15, 34, 63, 38, 0, 0, 60, 119, 
    0, 0, 0, 0, 0, 0, 0, 3, 13, 21, 35, 0, 0, 47, 132, 
    
    -- channel=609
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=610
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=611
    21, 18, 25, 27, 10, 8, 9, 7, 16, 25, 25, 18, 25, 17, 23, 
    25, 24, 34, 42, 22, 15, 17, 25, 20, 20, 21, 14, 22, 34, 8, 
    27, 27, 36, 64, 11, 24, 20, 29, 25, 17, 0, 14, 28, 31, 1, 
    27, 33, 28, 66, 0, 20, 50, 41, 38, 24, 27, 5, 22, 25, 13, 
    25, 35, 40, 54, 13, 27, 43, 35, 33, 32, 38, 0, 12, 30, 4, 
    13, 40, 33, 59, 13, 25, 36, 35, 36, 32, 34, 18, 1, 28, 26, 
    11, 38, 18, 33, 5, 27, 37, 27, 14, 26, 27, 6, 10, 12, 23, 
    19, 34, 0, 32, 34, 36, 26, 35, 27, 24, 26, 20, 4, 8, 0, 
    12, 29, 0, 40, 5, 8, 16, 19, 0, 0, 18, 0, 0, 18, 0, 
    26, 50, 1, 19, 6, 21, 12, 0, 35, 20, 33, 25, 22, 36, 0, 
    19, 53, 7, 16, 12, 0, 0, 35, 1, 32, 24, 8, 30, 6, 0, 
    26, 66, 0, 8, 27, 4, 4, 32, 0, 16, 13, 13, 41, 16, 0, 
    25, 38, 0, 26, 25, 17, 1, 0, 0, 0, 18, 51, 23, 0, 0, 
    20, 37, 38, 26, 17, 27, 0, 0, 0, 3, 13, 61, 13, 0, 0, 
    32, 28, 37, 29, 16, 16, 2, 2, 2, 5, 9, 35, 15, 0, 0, 
    
    -- channel=612
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 34, 37, 47, 61, 53, 36, 4, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 
    0, 0, 0, 16, 0, 2, 1, 23, 7, 0, 0, 8, 0, 0, 0, 
    0, 0, 22, 50, 3, 23, 44, 18, 17, 22, 7, 0, 0, 0, 0, 
    0, 0, 4, 6, 29, 21, 13, 33, 38, 25, 34, 26, 0, 0, 0, 
    0, 19, 17, 9, 0, 9, 27, 15, 11, 20, 27, 21, 34, 40, 0, 
    0, 33, 2, 0, 35, 20, 4, 20, 49, 51, 34, 54, 52, 28, 0, 
    0, 1, 0, 57, 6, 1, 10, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 12, 22, 21, 16, 27, 26, 30, 39, 31, 46, 39, 29, 42, 2, 
    0, 11, 0, 9, 9, 18, 0, 0, 27, 0, 3, 0, 0, 0, 0, 
    4, 40, 15, 0, 0, 10, 44, 61, 1, 39, 0, 1, 67, 30, 18, 
    9, 0, 0, 0, 5, 0, 7, 6, 2, 0, 0, 0, 15, 5, 0, 
    0, 13, 9, 5, 9, 7, 0, 0, 0, 20, 42, 23, 18, 0, 0, 
    14, 7, 0, 16, 10, 9, 0, 0, 0, 4, 17, 23, 0, 0, 0, 
    
    -- channel=613
    43, 42, 47, 34, 40, 38, 33, 35, 44, 47, 46, 48, 35, 30, 23, 
    56, 56, 56, 38, 44, 50, 49, 55, 63, 50, 41, 51, 51, 34, 40, 
    60, 61, 54, 23, 23, 22, 24, 19, 20, 24, 39, 50, 49, 31, 34, 
    59, 59, 51, 33, 46, 55, 46, 41, 38, 35, 29, 54, 44, 33, 27, 
    60, 58, 53, 34, 38, 41, 44, 38, 42, 44, 38, 47, 57, 41, 33, 
    65, 60, 40, 19, 21, 29, 29, 31, 29, 32, 36, 33, 57, 60, 60, 
    58, 49, 43, 20, 25, 34, 33, 23, 32, 37, 23, 34, 55, 66, 64, 
    56, 33, 39, 39, 27, 7, 8, 11, 13, 8, 9, 16, 27, 37, 61, 
    50, 21, 38, 19, 22, 31, 27, 0, 0, 5, 0, 0, 14, 34, 55, 
    49, 17, 28, 2, 13, 9, 11, 35, 36, 36, 34, 32, 42, 19, 42, 
    54, 14, 5, 3, 0, 2, 7, 2, 15, 8, 8, 10, 6, 23, 33, 
    56, 12, 14, 12, 0, 0, 16, 0, 23, 31, 24, 42, 10, 13, 34, 
    48, 11, 9, 27, 0, 0, 0, 0, 0, 33, 36, 22, 0, 0, 31, 
    49, 46, 25, 24, 13, 0, 0, 0, 4, 27, 40, 21, 0, 4, 32, 
    45, 38, 27, 9, 8, 0, 0, 0, 0, 9, 23, 14, 0, 0, 34, 
    
    -- channel=614
    4, 1, 6, 10, 9, 9, 10, 7, 12, 15, 11, 8, 2, 1, 0, 
    17, 15, 25, 42, 48, 47, 46, 57, 56, 33, 10, 7, 11, 8, 0, 
    18, 19, 25, 25, 22, 24, 25, 25, 27, 26, 9, 6, 12, 9, 0, 
    17, 21, 14, 50, 37, 49, 55, 58, 49, 44, 32, 12, 4, 5, 3, 
    17, 22, 46, 52, 43, 50, 60, 55, 54, 52, 46, 20, 15, 4, 0, 
    16, 33, 17, 43, 29, 35, 46, 53, 49, 41, 52, 25, 8, 18, 18, 
    11, 25, 14, 14, 36, 52, 61, 45, 51, 66, 40, 31, 37, 38, 21, 
    16, 19, 0, 29, 39, 9, 7, 28, 36, 27, 31, 41, 28, 29, 16, 
    9, 18, 2, 32, 18, 34, 32, 7, 0, 0, 0, 0, 0, 34, 22, 
    13, 26, 21, 9, 24, 21, 17, 25, 40, 30, 39, 31, 42, 29, 2, 
    15, 26, 3, 11, 6, 7, 0, 21, 0, 4, 4, 0, 13, 13, 7, 
    33, 36, 8, 6, 12, 7, 23, 23, 19, 34, 24, 42, 30, 25, 0, 
    32, 6, 5, 28, 13, 6, 4, 2, 0, 2, 28, 39, 16, 0, 2, 
    29, 40, 29, 32, 22, 13, 0, 0, 10, 27, 27, 43, 4, 3, 9, 
    40, 34, 31, 26, 19, 11, 0, 1, 4, 10, 20, 29, 4, 1, 0, 
    
    -- channel=615
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=616
    2, 1, 0, 5, 2, 2, 14, 8, 0, 3, 2, 1, 14, 8, 22, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 5, 0, 0, 9, 8, 
    0, 0, 1, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 4, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 
    0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 17, 0, 0, 7, 23, 12, 16, 29, 22, 0, 0, 0, 
    0, 12, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 31, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 16, 0, 0, 14, 0, 4, 0, 0, 15, 0, 0, 
    0, 19, 0, 0, 9, 12, 9, 6, 4, 0, 11, 12, 13, 4, 0, 
    0, 0, 0, 0, 0, 15, 12, 7, 0, 0, 0, 0, 15, 0, 0, 
    0, 0, 0, 4, 0, 10, 9, 4, 0, 0, 0, 2, 15, 0, 0, 
    
    -- channel=617
    11, 10, 6, 0, 0, 19, 39, 57, 27, 0, 0, 0, 20, 19, 9, 
    1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 22, 24, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 9, 14, 0, 0, 2, 17, 0, 0, 0, 25, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 20, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 2, 0, 0, 0, 0, 10, 43, 104, 106, 111, 114, 83, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 23, 0, 0, 0, 0, 4, 0, 13, 0, 
    0, 0, 0, 41, 16, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 51, 51, 0, 6, 12, 0, 0, 0, 60, 62, 46, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 9, 9, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 8, 7, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=618
    58, 61, 55, 44, 41, 47, 55, 73, 75, 62, 64, 58, 54, 72, 52, 
    58, 59, 54, 17, 5, 2, 1, 1, 14, 36, 46, 61, 60, 60, 66, 
    55, 56, 42, 0, 0, 0, 0, 0, 0, 3, 34, 65, 61, 49, 63, 
    55, 53, 38, 0, 16, 17, 7, 0, 0, 0, 34, 42, 47, 60, 61, 
    55, 51, 24, 0, 0, 0, 0, 0, 0, 0, 0, 43, 60, 48, 61, 
    52, 46, 17, 0, 0, 0, 0, 0, 0, 0, 0, 14, 50, 55, 56, 
    51, 25, 25, 0, 5, 0, 0, 0, 0, 0, 0, 13, 24, 25, 49, 
    51, 12, 27, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 
    47, 14, 53, 0, 3, 19, 6, 2, 32, 41, 32, 36, 44, 26, 48, 
    38, 6, 16, 0, 4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 34, 
    39, 0, 20, 0, 0, 0, 3, 10, 0, 0, 0, 6, 0, 4, 42, 
    23, 0, 1, 16, 1, 6, 4, 0, 32, 0, 17, 35, 0, 0, 18, 
    10, 0, 33, 11, 0, 2, 1, 1, 3, 50, 51, 22, 0, 0, 34, 
    21, 6, 0, 6, 0, 0, 5, 8, 17, 19, 0, 0, 0, 11, 18, 
    1, 0, 0, 0, 0, 0, 5, 4, 4, 4, 6, 0, 0, 7, 25, 
    
    -- channel=619
    12, 11, 18, 38, 0, 0, 0, 0, 0, 3, 11, 0, 28, 14, 27, 
    4, 3, 25, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 
    1, 0, 26, 129, 0, 11, 11, 34, 18, 0, 0, 0, 23, 29, 0, 
    1, 13, 13, 117, 0, 0, 46, 0, 2, 0, 12, 0, 6, 43, 9, 
    0, 18, 42, 60, 0, 0, 6, 0, 0, 0, 7, 0, 0, 38, 23, 
    0, 26, 37, 101, 0, 0, 14, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 34, 5, 39, 6, 2, 9, 7, 0, 0, 6, 0, 0, 0, 0, 
    6, 56, 0, 59, 5, 22, 13, 24, 0, 0, 4, 0, 0, 0, 0, 
    30, 78, 0, 57, 0, 0, 0, 40, 27, 15, 67, 45, 6, 9, 0, 
    26, 113, 0, 48, 0, 14, 0, 0, 10, 0, 0, 0, 0, 30, 0, 
    5, 117, 16, 21, 19, 0, 0, 72, 0, 40, 11, 0, 55, 0, 0, 
    7, 127, 0, 16, 70, 2, 0, 24, 0, 0, 0, 0, 57, 0, 0, 
    0, 84, 27, 9, 42, 50, 3, 0, 0, 0, 24, 89, 48, 0, 0, 
    0, 19, 46, 13, 7, 56, 9, 0, 0, 0, 0, 77, 32, 0, 0, 
    5, 9, 41, 37, 2, 24, 13, 6, 0, 0, 0, 24, 45, 0, 0, 
    
    -- channel=620
    13, 18, 10, 2, 12, 15, 16, 29, 34, 21, 21, 19, 2, 22, 4, 
    19, 19, 10, 0, 33, 42, 45, 44, 48, 48, 21, 30, 19, 11, 26, 
    21, 22, 2, 0, 34, 32, 29, 24, 29, 49, 59, 19, 13, 5, 41, 
    21, 18, 11, 0, 71, 41, 22, 45, 40, 36, 52, 47, 3, 0, 21, 
    22, 12, 8, 0, 59, 57, 29, 48, 49, 50, 30, 56, 29, 0, 0, 
    29, 9, 0, 0, 51, 38, 38, 46, 44, 53, 50, 55, 55, 20, 21, 
    24, 0, 11, 0, 32, 44, 30, 34, 45, 45, 33, 57, 60, 44, 33, 
    6, 0, 26, 0, 31, 20, 24, 30, 40, 35, 35, 50, 51, 53, 69, 
    0, 0, 43, 0, 42, 33, 24, 0, 6, 16, 0, 0, 34, 31, 72, 
    0, 0, 32, 0, 40, 21, 42, 58, 21, 40, 30, 32, 38, 13, 84, 
    9, 0, 20, 10, 24, 29, 28, 18, 42, 13, 23, 31, 5, 32, 71, 
    18, 0, 27, 14, 0, 35, 59, 0, 73, 21, 23, 49, 0, 40, 77, 
    23, 0, 28, 21, 0, 7, 22, 26, 31, 65, 15, 0, 7, 27, 81, 
    32, 15, 6, 17, 22, 0, 17, 25, 37, 58, 38, 0, 4, 45, 71, 
    25, 23, 8, 8, 26, 8, 17, 21, 27, 32, 43, 0, 6, 38, 77, 
    
    -- channel=621
    4, 3, 7, 43, 0, 0, 0, 0, 0, 0, 10, 0, 21, 2, 24, 
    0, 0, 15, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 
    1, 0, 22, 132, 0, 0, 0, 17, 2, 0, 0, 0, 20, 34, 0, 
    0, 7, 22, 110, 0, 0, 43, 0, 0, 0, 10, 0, 5, 29, 14, 
    0, 12, 60, 76, 0, 0, 17, 0, 0, 0, 2, 0, 0, 21, 4, 
    0, 23, 50, 95, 0, 0, 12, 1, 0, 0, 0, 0, 0, 2, 0, 
    0, 39, 17, 44, 0, 1, 9, 9, 0, 0, 22, 0, 0, 0, 0, 
    6, 77, 0, 48, 12, 24, 11, 24, 3, 0, 13, 0, 0, 0, 0, 
    22, 90, 0, 77, 0, 0, 0, 23, 0, 0, 22, 0, 0, 6, 0, 
    23, 125, 0, 70, 0, 21, 0, 0, 12, 0, 12, 0, 0, 47, 0, 
    6, 123, 3, 20, 23, 0, 0, 65, 0, 30, 4, 0, 54, 0, 0, 
    10, 144, 0, 0, 63, 7, 0, 44, 0, 0, 0, 0, 94, 0, 0, 
    0, 72, 6, 0, 41, 40, 1, 0, 0, 0, 3, 57, 54, 0, 0, 
    0, 15, 46, 0, 5, 51, 1, 0, 0, 0, 0, 58, 42, 0, 0, 
    6, 9, 31, 34, 0, 22, 6, 0, 0, 0, 0, 12, 46, 0, 0, 
    
    -- channel=622
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=623
    29, 19, 31, 52, 25, 14, 15, 2, 8, 35, 34, 26, 48, 19, 47, 
    28, 27, 48, 89, 29, 15, 17, 34, 29, 39, 37, 11, 31, 62, 11, 
    28, 26, 58, 103, 0, 0, 0, 0, 0, 0, 0, 13, 41, 69, 0, 
    28, 36, 36, 114, 0, 4, 30, 7, 4, 0, 10, 0, 46, 52, 25, 
    25, 43, 61, 88, 0, 0, 32, 0, 0, 0, 29, 0, 12, 60, 8, 
    5, 57, 52, 71, 0, 0, 0, 0, 3, 0, 0, 0, 0, 29, 26, 
    0, 67, 20, 49, 0, 0, 25, 4, 0, 15, 29, 0, 0, 15, 23, 
    31, 72, 0, 45, 9, 8, 0, 7, 4, 4, 4, 0, 0, 0, 0, 
    34, 78, 0, 77, 0, 0, 18, 33, 0, 0, 29, 0, 0, 0, 0, 
    44, 96, 0, 45, 0, 20, 0, 0, 39, 0, 25, 10, 6, 42, 0, 
    25, 117, 0, 23, 0, 0, 0, 18, 0, 0, 0, 0, 7, 0, 0, 
    29, 128, 0, 0, 45, 0, 0, 77, 0, 41, 7, 0, 97, 0, 0, 
    12, 77, 0, 13, 46, 24, 1, 0, 0, 0, 21, 84, 38, 0, 0, 
    0, 35, 47, 25, 11, 55, 0, 0, 0, 0, 0, 99, 35, 0, 0, 
    17, 19, 41, 35, 6, 30, 0, 0, 0, 0, 0, 56, 27, 0, 0, 
    
    -- channel=624
    0, 5, 0, 0, 0, 0, 6, 27, 0, 0, 0, 0, 9, 2, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 26, 29, 34, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 28, 106, 93, 82, 108, 75, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 29, 0, 0, 3, 1, 33, 0, 16, 0, 
    0, 0, 0, 34, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 57, 41, 0, 6, 7, 0, 0, 0, 33, 11, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 9, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 0, 0, 0, 0, 16, 
    
    -- channel=625
    12, 15, 8, 0, 3, 15, 25, 39, 17, 0, 0, 1, 7, 8, 0, 
    7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 10, 
    2, 2, 0, 0, 53, 57, 61, 50, 37, 13, 22, 12, 0, 0, 0, 
    3, 0, 0, 0, 59, 25, 6, 19, 32, 47, 1, 3, 0, 0, 0, 
    2, 0, 0, 0, 39, 16, 0, 25, 20, 24, 16, 29, 15, 6, 50, 
    5, 0, 6, 0, 17, 30, 18, 9, 5, 22, 4, 9, 36, 2, 3, 
    4, 0, 0, 11, 60, 23, 12, 17, 29, 3, 0, 3, 0, 0, 0, 
    0, 0, 35, 0, 13, 14, 26, 0, 0, 0, 0, 0, 4, 17, 34, 
    6, 0, 19, 0, 40, 13, 20, 35, 96, 96, 60, 89, 95, 28, 31, 
    0, 0, 0, 0, 11, 0, 3, 25, 0, 1, 0, 0, 0, 0, 69, 
    3, 0, 11, 5, 3, 19, 63, 0, 35, 19, 24, 65, 2, 46, 59, 
    0, 0, 21, 41, 0, 5, 0, 0, 28, 0, 19, 0, 0, 0, 71, 
    13, 27, 53, 2, 4, 0, 5, 12, 27, 94, 28, 0, 0, 29, 85, 
    24, 0, 0, 0, 9, 0, 17, 24, 28, 0, 0, 0, 0, 40, 68, 
    5, 14, 1, 0, 6, 0, 17, 20, 21, 19, 11, 0, 0, 34, 92, 
    
    -- channel=626
    47, 39, 50, 43, 41, 41, 37, 32, 38, 47, 41, 44, 45, 28, 32, 
    56, 55, 61, 60, 47, 51, 51, 56, 55, 41, 39, 41, 47, 36, 27, 
    58, 58, 66, 58, 43, 47, 49, 50, 49, 38, 23, 47, 46, 36, 17, 
    58, 59, 57, 77, 42, 65, 69, 65, 61, 63, 41, 38, 52, 42, 22, 
    58, 62, 64, 71, 43, 53, 67, 59, 60, 60, 67, 40, 50, 58, 39, 
    54, 65, 56, 60, 31, 49, 52, 50, 50, 45, 49, 38, 40, 59, 58, 
    50, 62, 43, 55, 41, 51, 62, 47, 47, 55, 41, 32, 44, 56, 56, 
    54, 51, 30, 47, 50, 37, 34, 31, 25, 25, 23, 20, 29, 39, 41, 
    56, 49, 20, 48, 31, 36, 42, 41, 18, 19, 36, 17, 16, 46, 38, 
    58, 50, 27, 22, 23, 27, 20, 28, 54, 43, 50, 46, 49, 45, 20, 
    58, 59, 17, 23, 8, 15, 21, 23, 21, 31, 29, 23, 35, 32, 22, 
    64, 53, 21, 29, 21, 0, 9, 32, 3, 40, 37, 36, 38, 21, 13, 
    61, 58, 19, 42, 32, 9, 0, 0, 2, 15, 48, 53, 17, 9, 10, 
    55, 64, 52, 40, 31, 22, 0, 0, 6, 22, 44, 60, 11, 2, 20, 
    62, 58, 54, 36, 24, 20, 6, 8, 10, 17, 26, 49, 10, 3, 16, 
    
    -- channel=627
    67, 71, 62, 42, 43, 49, 67, 93, 89, 68, 69, 59, 68, 76, 63, 
    70, 71, 69, 35, 18, 10, 2, 0, 11, 23, 43, 58, 56, 55, 60, 
    64, 65, 54, 42, 12, 37, 36, 40, 25, 17, 22, 64, 58, 43, 41, 
    63, 65, 44, 31, 35, 42, 59, 27, 34, 41, 53, 25, 47, 65, 51, 
    61, 63, 36, 1, 27, 24, 10, 24, 28, 30, 36, 41, 66, 64, 74, 
    44, 55, 39, 31, 0, 8, 15, 11, 5, 12, 10, 19, 42, 65, 64, 
    38, 18, 10, 13, 49, 27, 19, 16, 23, 30, 16, 13, 11, 11, 56, 
    32, 0, 2, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 26, 
    48, 24, 36, 0, 10, 25, 32, 28, 62, 75, 76, 69, 75, 46, 29, 
    42, 23, 0, 3, 0, 0, 0, 0, 11, 0, 0, 0, 2, 0, 11, 
    39, 19, 24, 4, 0, 0, 18, 23, 0, 9, 1, 12, 1, 25, 26, 
    36, 4, 0, 40, 18, 1, 0, 0, 10, 10, 32, 35, 0, 0, 0, 
    27, 39, 51, 25, 8, 9, 0, 0, 0, 53, 83, 61, 2, 0, 29, 
    38, 26, 23, 17, 10, 4, 4, 7, 17, 8, 0, 10, 0, 9, 17, 
    25, 26, 27, 1, 7, 0, 8, 7, 5, 4, 2, 0, 5, 4, 31, 
    
    -- channel=628
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 6, 17, 15, 14, 22, 24, 17, 18, 13, 0, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 6, 6, 11, 15, 0, 3, 5, 10, 8, 0, 15, 0, 
    0, 0, 0, 4, 13, 10, 0, 4, 10, 4, 6, 0, 9, 0, 0, 
    0, 15, 1, 0, 2, 9, 19, 26, 0, 0, 0, 0, 19, 18, 0, 
    0, 0, 0, 0, 0, 5, 9, 9, 6, 0, 0, 0, 12, 2, 0, 
    0, 0, 0, 0, 0, 7, 3, 0, 0, 1, 2, 5, 14, 0, 0, 
    0, 0, 0, 8, 1, 6, 1, 0, 2, 3, 4, 8, 8, 0, 0, 
    
    -- channel=629
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 41, 57, 68, 86, 86, 69, 31, 11, 8, 0, 13, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 19, 54, 0, 0, 6, 46, 
    0, 0, 3, 0, 21, 0, 0, 12, 0, 0, 0, 65, 0, 0, 0, 
    5, 0, 8, 6, 23, 25, 28, 10, 11, 14, 0, 16, 0, 0, 0, 
    33, 0, 0, 0, 54, 20, 0, 24, 32, 30, 44, 47, 45, 0, 0, 
    18, 15, 26, 0, 0, 0, 0, 0, 0, 3, 6, 44, 82, 83, 26, 
    3, 15, 39, 0, 25, 9, 12, 9, 49, 55, 30, 59, 84, 52, 73, 
    0, 0, 10, 33, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    0, 0, 53, 0, 36, 14, 42, 64, 31, 54, 52, 55, 50, 24, 70, 
    0, 0, 0, 0, 0, 32, 0, 0, 66, 0, 6, 0, 0, 0, 26, 
    3, 0, 45, 0, 0, 8, 78, 36, 49, 29, 0, 17, 12, 58, 82, 
    11, 0, 0, 0, 0, 0, 1, 5, 11, 0, 0, 0, 0, 15, 29, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 61, 75, 0, 0, 16, 42, 
    9, 0, 0, 0, 6, 0, 0, 0, 0, 11, 35, 12, 0, 15, 33, 
    
    -- channel=630
    73, 74, 70, 60, 46, 53, 66, 80, 87, 79, 78, 68, 74, 77, 64, 
    81, 82, 86, 59, 32, 22, 23, 30, 37, 48, 56, 66, 70, 73, 57, 
    79, 79, 77, 55, 0, 23, 22, 26, 18, 19, 31, 70, 77, 61, 47, 
    78, 80, 61, 57, 19, 55, 61, 29, 34, 35, 60, 38, 61, 77, 59, 
    75, 80, 64, 22, 16, 24, 22, 25, 31, 30, 38, 50, 72, 76, 67, 
    58, 81, 47, 42, 0, 3, 19, 12, 9, 9, 17, 20, 43, 79, 78, 
    53, 53, 31, 11, 29, 27, 20, 14, 15, 33, 24, 18, 33, 41, 67, 
    58, 30, 2, 58, 2, 0, 0, 1, 0, 0, 0, 0, 0, 3, 33, 
    60, 42, 28, 10, 0, 24, 24, 24, 26, 39, 56, 36, 39, 44, 35, 
    59, 44, 4, 0, 0, 0, 0, 0, 25, 3, 10, 3, 16, 7, 0, 
    54, 45, 13, 0, 0, 0, 0, 28, 0, 8, 0, 0, 16, 2, 19, 
    53, 39, 0, 20, 18, 0, 0, 0, 0, 15, 27, 39, 5, 0, 0, 
    36, 35, 37, 25, 7, 4, 0, 0, 0, 15, 76, 68, 5, 0, 0, 
    44, 45, 29, 24, 6, 6, 0, 0, 0, 8, 0, 36, 0, 0, 0, 
    36, 32, 36, 15, 2, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    
    -- channel=631
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=632
    17, 19, 20, 38, 7, 0, 2, 6, 7, 14, 23, 6, 31, 22, 33, 
    10, 10, 23, 60, 0, 0, 0, 0, 0, 0, 10, 0, 12, 41, 2, 
    8, 6, 24, 90, 0, 0, 0, 0, 0, 0, 0, 0, 30, 44, 0, 
    8, 16, 13, 74, 0, 0, 11, 0, 0, 0, 0, 0, 14, 42, 29, 
    4, 18, 39, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 21, 
    0, 26, 29, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 
    0, 31, 8, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 49, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 59, 0, 35, 0, 0, 0, 9, 0, 0, 33, 12, 0, 0, 0, 
    23, 83, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    7, 83, 0, 11, 5, 0, 0, 36, 0, 6, 0, 0, 14, 0, 0, 
    2, 92, 0, 0, 40, 0, 0, 16, 0, 0, 0, 0, 48, 0, 0, 
    0, 46, 5, 0, 21, 27, 0, 0, 0, 0, 12, 57, 27, 0, 0, 
    0, 0, 19, 0, 0, 32, 1, 0, 0, 0, 0, 43, 21, 0, 0, 
    0, 0, 12, 11, 0, 9, 2, 0, 0, 0, 0, 1, 26, 0, 0, 
    
    -- channel=633
    88, 84, 88, 67, 67, 71, 76, 83, 97, 97, 91, 93, 78, 82, 67, 
    104, 104, 101, 59, 76, 82, 83, 94, 102, 98, 85, 95, 95, 81, 82, 
    108, 109, 97, 40, 68, 76, 69, 67, 72, 79, 90, 94, 89, 70, 82, 
    107, 106, 90, 55, 95, 100, 91, 101, 94, 91, 89, 101, 83, 70, 62, 
    107, 104, 82, 56, 91, 93, 87, 95, 99, 96, 94, 99, 98, 81, 65, 
    105, 101, 62, 49, 70, 74, 79, 81, 81, 87, 95, 89, 111, 108, 108, 
    90, 77, 65, 46, 56, 78, 75, 64, 71, 81, 59, 74, 101, 106, 111, 
    76, 42, 53, 53, 63, 51, 52, 51, 49, 45, 45, 50, 62, 77, 120, 
    64, 25, 62, 34, 55, 59, 54, 33, 27, 34, 33, 23, 51, 70, 107, 
    76, 29, 55, 8, 50, 36, 48, 64, 72, 76, 75, 72, 83, 51, 86, 
    83, 26, 34, 23, 18, 31, 38, 35, 54, 49, 50, 56, 45, 53, 76, 
    88, 27, 39, 41, 13, 16, 49, 18, 53, 51, 57, 79, 16, 55, 63, 
    88, 35, 41, 67, 25, 9, 6, 11, 18, 71, 71, 54, 14, 21, 67, 
    88, 85, 57, 60, 43, 13, 5, 12, 25, 73, 78, 59, 3, 29, 70, 
    87, 78, 64, 42, 40, 20, 12, 18, 24, 38, 57, 49, 5, 27, 75, 
    
    -- channel=634
    4, 0, 14, 25, 12, 0, 0, 0, 0, 16, 17, 17, 0, 0, 0, 
    14, 13, 31, 50, 55, 52, 57, 80, 75, 52, 34, 18, 25, 31, 3, 
    23, 24, 37, 37, 0, 0, 0, 0, 4, 19, 0, 14, 29, 42, 16, 
    23, 32, 26, 54, 0, 4, 22, 22, 5, 0, 15, 31, 23, 7, 17, 
    25, 33, 56, 53, 7, 20, 40, 15, 17, 13, 22, 0, 9, 13, 0, 
    28, 49, 7, 29, 22, 13, 15, 25, 33, 19, 32, 25, 4, 24, 23, 
    27, 63, 39, 9, 0, 6, 21, 7, 0, 19, 24, 21, 60, 55, 33, 
    41, 62, 0, 26, 26, 21, 11, 23, 37, 36, 26, 37, 36, 23, 16, 
    11, 8, 6, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    25, 34, 41, 0, 18, 21, 25, 0, 64, 39, 58, 50, 45, 43, 0, 
    25, 26, 0, 6, 0, 1, 0, 7, 12, 8, 9, 0, 11, 0, 0, 
    34, 59, 6, 0, 0, 0, 33, 46, 0, 30, 2, 28, 44, 48, 0, 
    24, 0, 0, 30, 2, 0, 0, 0, 0, 0, 0, 22, 10, 0, 0, 
    9, 40, 23, 33, 8, 8, 0, 0, 0, 42, 43, 73, 0, 0, 0, 
    31, 18, 21, 29, 10, 5, 0, 0, 0, 1, 17, 45, 0, 0, 0, 
    
    -- channel=635
    6, 5, 8, 12, 0, 2, 0, 0, 6, 12, 11, 8, 0, 0, 0, 
    19, 18, 19, 32, 28, 35, 44, 46, 39, 24, 8, 8, 12, 6, 0, 
    24, 25, 21, 21, 23, 29, 32, 32, 35, 36, 8, 6, 13, 3, 0, 
    24, 24, 25, 29, 32, 35, 51, 57, 47, 43, 37, 15, 7, 0, 0, 
    24, 22, 42, 38, 35, 59, 53, 54, 54, 56, 43, 21, 14, 1, 0, 
    23, 25, 19, 34, 35, 39, 48, 52, 50, 49, 54, 41, 22, 24, 24, 
    19, 23, 20, 15, 23, 46, 46, 38, 38, 41, 29, 28, 35, 37, 23, 
    12, 23, 0, 12, 40, 25, 24, 27, 29, 26, 26, 30, 31, 42, 24, 
    7, 8, 2, 26, 13, 23, 17, 0, 0, 0, 0, 0, 0, 29, 31, 
    14, 22, 4, 4, 18, 16, 23, 33, 33, 40, 42, 37, 34, 33, 28, 
    19, 13, 0, 0, 3, 4, 0, 21, 10, 20, 16, 3, 27, 9, 29, 
    32, 29, 0, 0, 0, 0, 25, 7, 12, 13, 8, 28, 20, 17, 25, 
    36, 2, 1, 13, 2, 0, 0, 0, 0, 0, 5, 4, 5, 0, 19, 
    32, 35, 26, 11, 12, 0, 0, 0, 0, 23, 33, 18, 0, 0, 25, 
    41, 35, 22, 18, 8, 0, 0, 0, 0, 7, 21, 11, 0, 0, 18, 
    
    -- channel=636
    31, 28, 36, 41, 30, 28, 16, 12, 27, 37, 38, 38, 23, 21, 19, 
    45, 43, 49, 61, 61, 65, 75, 83, 76, 53, 40, 40, 42, 34, 24, 
    52, 53, 51, 49, 44, 43, 41, 40, 50, 57, 27, 36, 45, 35, 30, 
    51, 53, 55, 60, 52, 53, 71, 73, 60, 55, 54, 47, 37, 23, 29, 
    52, 53, 72, 70, 56, 78, 77, 71, 72, 74, 58, 39, 38, 24, 7, 
    57, 60, 44, 62, 62, 59, 67, 73, 72, 71, 77, 62, 48, 52, 52, 
    57, 62, 58, 44, 37, 65, 64, 56, 56, 59, 51, 53, 70, 72, 53, 
    50, 65, 30, 38, 67, 50, 52, 56, 61, 56, 57, 63, 64, 66, 50, 
    39, 35, 34, 67, 41, 47, 37, 9, 0, 0, 0, 0, 6, 48, 56, 
    45, 51, 38, 30, 46, 42, 50, 59, 67, 71, 73, 68, 62, 64, 49, 
    51, 37, 27, 25, 28, 31, 15, 42, 40, 45, 42, 23, 53, 32, 45, 
    61, 56, 22, 18, 18, 24, 61, 39, 42, 44, 31, 59, 50, 53, 47, 
    63, 15, 15, 43, 22, 13, 12, 13, 19, 3, 21, 26, 30, 17, 36, 
    56, 64, 52, 38, 37, 18, 4, 9, 14, 58, 67, 53, 17, 21, 44, 
    67, 56, 46, 44, 35, 21, 10, 13, 20, 34, 51, 43, 16, 19, 38, 
    
    -- channel=637
    35, 31, 34, 31, 29, 30, 35, 32, 32, 37, 35, 37, 37, 39, 36, 
    31, 31, 33, 13, 0, 0, 0, 0, 6, 22, 34, 34, 39, 43, 43, 
    29, 28, 33, 0, 0, 0, 0, 0, 0, 0, 19, 39, 37, 41, 40, 
    29, 29, 22, 6, 0, 0, 0, 0, 0, 0, 0, 28, 38, 45, 36, 
    30, 30, 11, 0, 0, 0, 0, 0, 0, 0, 0, 11, 30, 39, 35, 
    30, 31, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 29, 29, 
    26, 31, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 25, 
    40, 18, 24, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    32, 16, 18, 8, 0, 1, 0, 6, 9, 5, 18, 14, 0, 0, 9, 
    29, 6, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 14, 1, 0, 0, 0, 0, 0, 3, 6, 3, 0, 0, 0, 
    0, 2, 0, 6, 0, 2, 2, 0, 0, 15, 20, 17, 0, 0, 0, 
    0, 1, 0, 8, 0, 2, 5, 1, 1, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 10, 0, 0, 0, 
    
    -- channel=638
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 11, 
    0, 0, 0, 16, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 11, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 4, 
    0, 0, 0, 9, 0, 12, 0, 0, 0, 18, 0, 0, 0, 0, 12, 
    0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 2, 24, 10, 0, 0, 2, 1, 0, 11, 6, 0, 6, 0, 
    0, 16, 27, 0, 2, 4, 0, 0, 0, 0, 0, 0, 7, 16, 0, 
    0, 40, 0, 19, 1, 3, 20, 8, 8, 36, 0, 0, 0, 0, 9, 
    0, 23, 0, 58, 0, 5, 0, 43, 0, 0, 0, 0, 0, 25, 54, 
    0, 24, 0, 0, 12, 11, 19, 0, 1, 0, 0, 0, 9, 1, 61, 
    0, 19, 0, 0, 8, 8, 1, 12, 6, 9, 0, 0, 62, 0, 97, 
    0, 20, 2, 0, 9, 0, 0, 2, 28, 0, 0, 0, 18, 17, 49, 
    0, 0, 0, 0, 0, 0, 3, 7, 8, 0, 5, 0, 30, 8, 49, 
    0, 0, 0, 0, 0, 1, 6, 0, 2, 0, 0, 0, 21, 2, 41, 
    
    -- channel=639
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 8, 25, 13, 11, 15, 25, 20, 1, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 15, 0, 0, 6, 0, 0, 0, 0, 0, 0, 11, 1, 
    0, 0, 0, 0, 15, 15, 0, 0, 5, 5, 0, 18, 1, 0, 0, 
    0, 4, 4, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 7, 0, 10, 45, 31, 0, 0, 9, 0, 0, 22, 14, 4, 
    0, 0, 0, 26, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 16, 19, 0, 26, 21, 24, 29, 0, 27, 5, 
    0, 0, 0, 5, 1, 10, 15, 0, 45, 22, 29, 39, 5, 0, 0, 
    0, 3, 5, 0, 0, 0, 0, 22, 0, 0, 0, 0, 15, 11, 16, 
    5, 17, 0, 0, 8, 0, 0, 1, 10, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 7, 25, 5, 7, 0, 4, 
    2, 4, 0, 3, 0, 2, 2, 2, 2, 2, 0, 9, 0, 5, 5, 
    
    
    others => 0);
end gold_package;
