library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    324, 249, 301, 
    153, 153, 66, 
    79, 244, 268, 
    
    -- channel=1
    0, 0, 0, 
    20, 0, 0, 
    100, 179, 158, 
    
    -- channel=2
    120, 27, 81, 
    352, 153, 283, 
    323, 324, 138, 
    
    -- channel=3
    372, 449, 297, 
    278, 294, 269, 
    126, 0, 0, 
    
    -- channel=4
    405, 324, 240, 
    235, 159, 72, 
    73, 0, 6, 
    
    -- channel=5
    250, 399, 531, 
    402, 533, 410, 
    378, 62, 85, 
    
    -- channel=6
    84, 13, 0, 
    0, 0, 0, 
    0, 0, 12, 
    
    -- channel=7
    348, 180, 151, 
    250, 220, 86, 
    541, 338, 265, 
    
    -- channel=8
    302, 547, 351, 
    585, 525, 346, 
    521, 435, 391, 
    
    -- channel=9
    0, 0, 0, 
    0, 76, 0, 
    23, 119, 105, 
    
    -- channel=10
    272, 394, 518, 
    364, 281, 388, 
    253, 58, 20, 
    
    -- channel=11
    57, 0, 0, 
    0, 0, 0, 
    0, 196, 121, 
    
    -- channel=12
    102, 0, 0, 
    50, 101, 86, 
    268, 382, 347, 
    
    -- channel=13
    215, 335, 292, 
    257, 278, 249, 
    313, 240, 221, 
    
    -- channel=14
    0, 113, 190, 
    232, 243, 55, 
    447, 111, 50, 
    
    -- channel=15
    0, 0, 4, 
    0, 0, 102, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
