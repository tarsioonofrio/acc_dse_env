LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE ifmap_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_map: padroes := ( 

			179, 140, 78, 255, 244, 190, 27, 167, 247, 56, 133, 248, 112, 23, 144, 
			36, 206, 222, 69, 85, 166, 176, 159, 229, 151, 0, 119, 217, 170, 27, 
			212, 229, 76, 143, 43, 142, 175, 124, 0, 0, 0, 0, 0, 0, 23, 
			49, 0, 255, 12, 103, 27, 0, 0, 0, 0, 142, 0, 211, 0, 129, 
			165, 0, 43, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 
			0, 0, 170, 0, 65, 0, 0, 141, 16, 0, 0, 182, 0, 0, 0, 
			0, 0, 240, 205, 0, 0, 0, 0, 244, 0, 8, 67, 0, 0, 0, 
			0, 0, 0, 88, 0, 0, 0, 0, 98, 0, 99, 176, 0, 0, 156, 
			0, 0, 0, 0, 0, 80, 107, 0, 0, 254, 0, 96, 0, 225, 4, 
			0, 0, 245, 0, 0, 0, 179, 0, 0, 0, 66, 48, 0, 0, 62, 
			0, 0, 48, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 162, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 224, 0, 0, 0, 0, 0, 0, 125, 0, 0, 
			0, 0, 0, 116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 166, 58, 131, 
			186, 101, 0, 0, 0, 151, 4, 220, 95, 247, 144, 210, 1, 102, 62, 
			79, 1, 0, 0, 106, 57, 142, 129, 155, 203, 164, 139, 134, 52, 16, 
			123, 96, 115, 57, 226, 59, 234, 4, 71, 236, 105, 113, 156, 104, 39, 
			224, 195, 193, 131, 201, 131, 66, 113, 102, 223, 243, 98, 59, 121, 70, 
			

			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 184, 157, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 138, 63, 60, 11, 0, 0, 0, 
			0, 250, 0, 0, 0, 0, 79, 121, 235, 219, 0, 6, 0, 0, 0, 
			0, 6, 0, 89, 31, 245, 241, 31, 105, 43, 57, 232, 23, 0, 211, 
			223, 207, 0, 0, 149, 160, 30, 80, 0, 58, 209, 0, 34, 90, 203, 
			17, 80, 0, 0, 34, 120, 6, 178, 0, 223, 89, 28, 189, 130, 22, 
			130, 225, 35, 0, 229, 21, 0, 117, 0, 82, 39, 212, 35, 193, 0, 
			24, 156, 110, 133, 253, 243, 200, 91, 2, 0, 248, 0, 234, 179, 0, 
			60, 17, 28, 208, 152, 215, 96, 30, 223, 160, 0, 108, 6, 101, 0, 
			181, 75, 226, 170, 231, 214, 82, 42, 64, 212, 1, 192, 246, 208, 115, 
			49, 130, 103, 46, 194, 201, 94, 31, 64, 120, 140, 93, 230, 47, 155, 
			199, 32, 36, 6, 13, 240, 103, 126, 174, 255, 152, 130, 212, 60, 69, 
			227, 96, 192, 130, 210, 65, 206, 92, 246, 117, 103, 135, 250, 9, 242, 
			54, 88, 185, 243, 21, 127, 142, 2, 185, 225, 205, 83, 100, 249, 175, 
			

			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 67, 53, 171, 0, 170, 127, 0, 0, 0, 
			234, 0, 0, 0, 0, 0, 115, 112, 0, 0, 46, 173, 250, 0, 0, 
			235, 0, 0, 0, 17, 0, 244, 166, 127, 0, 119, 218, 126, 15, 0, 
			243, 0, 159, 0, 39, 149, 247, 209, 236, 0, 8, 143, 123, 97, 0, 
			30, 245, 109, 0, 0, 246, 156, 155, 140, 0, 196, 198, 245, 57, 245, 
			236, 130, 241, 26, 0, 0, 107, 107, 242, 0, 212, 242, 167, 143, 32, 
			9, 228, 173, 174, 0, 0, 215, 169, 184, 0, 76, 114, 0, 85, 238, 
			174, 219, 40, 225, 248, 79, 228, 107, 0, 155, 101, 65, 0, 0, 0, 
			82, 82, 164, 0, 127, 97, 0, 202, 169, 52, 249, 27, 0, 0, 78, 
			5, 111, 86, 0, 243, 27, 237, 182, 163, 34, 195, 177, 209, 34, 227, 
			69, 186, 83, 0, 114, 151, 75, 56, 231, 87, 21, 200, 99, 1, 212, 
			115, 103, 0, 204, 107, 40, 5, 86, 175, 178, 18, 152, 90, 19, 249, 
			254, 145, 0, 172, 151, 73, 10, 106, 244, 128, 200, 32, 16, 179, 238, 
			20, 54, 77, 130, 43, 139, 61, 190, 77, 142, 228, 220, 96, 236, 18, 
			

			0, 0, 74, 185, 79, 52, 192, 0, 132, 0, 0, 0, 0, 159, 145, 
			55, 184, 46, 38, 28, 157, 52, 0, 0, 0, 144, 25, 0, 0, 214, 
			0, 0, 168, 5, 49, 0, 0, 0, 134, 17, 213, 43, 43, 0, 0, 
			19, 85, 157, 41, 142, 0, 80, 196, 98, 0, 0, 0, 0, 184, 0, 
			189, 214, 51, 145, 201, 124, 172, 28, 0, 0, 29, 184, 77, 34, 0, 
			0, 0, 48, 0, 0, 0, 79, 13, 202, 188, 0, 0, 0, 166, 62, 
			207, 157, 0, 82, 0, 57, 0, 187, 181, 157, 0, 20, 0, 246, 220, 
			112, 147, 39, 131, 86, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			204, 229, 109, 62, 164, 0, 0, 252, 159, 0, 0, 0, 0, 90, 181, 
			0, 0, 76, 130, 60, 0, 0, 108, 212, 0, 0, 0, 173, 55, 0, 
			0, 0, 0, 54, 242, 107, 150, 0, 0, 0, 194, 248, 234, 0, 0, 
			0, 0, 189, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			213, 0, 0, 0, 0, 0, 0, 0, 0, 159, 150, 183, 0, 0, 30, 
			0, 0, 0, 0, 0, 0, 245, 125, 0, 0, 0, 0, 0, 30, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 59, 4, 149, 0, 28, 24, 0, 
			

			8, 102, 200, 3, 147, 122, 88, 190, 194, 112, 38, 143, 129, 84, 191, 
			76, 247, 57, 223, 6, 240, 164, 58, 46, 6, 100, 241, 33, 252, 172, 
			5, 69, 104, 157, 212, 105, 28, 193, 235, 0, 204, 169, 110, 68, 187, 
			126, 115, 210, 138, 24, 12, 170, 203, 24, 124, 40, 60, 54, 42, 247, 
			166, 198, 235, 175, 193, 128, 76, 241, 57, 0, 154, 223, 141, 227, 206, 
			107, 116, 15, 99, 202, 49, 137, 216, 45, 0, 42, 41, 209, 131, 126, 
			210, 17, 138, 48, 200, 92, 103, 85, 244, 0, 45, 180, 194, 211, 88, 
			227, 44, 223, 88, 3, 194, 66, 61, 245, 92, 160, 203, 253, 65, 171, 
			143, 0, 179, 141, 206, 243, 17, 226, 114, 248, 99, 12, 42, 244, 127, 
			67, 0, 75, 0, 117, 157, 0, 239, 9, 91, 109, 0, 253, 210, 139, 
			0, 188, 179, 0, 252, 160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 252, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			

			17, 219, 160, 106, 6, 98, 140, 139, 123, 229, 89, 245, 78, 223, 100, 
			244, 149, 150, 124, 230, 66, 0, 114, 0, 44, 0, 0, 122, 172, 31, 
			0, 254, 180, 132, 224, 38, 0, 0, 66, 154, 0, 0, 0, 144, 3, 
			0, 9, 196, 66, 0, 213, 0, 0, 0, 41, 0, 0, 0, 0, 35, 
			0, 247, 0, 41, 0, 0, 0, 0, 0, 249, 0, 0, 0, 0, 244, 
			0, 0, 0, 213, 78, 190, 0, 0, 0, 212, 0, 0, 104, 0, 0, 
			0, 0, 211, 0, 248, 152, 0, 0, 0, 151, 0, 0, 0, 2, 0, 
			0, 0, 0, 0, 246, 160, 0, 0, 0, 254, 0, 0, 83, 0, 0, 
			0, 0, 0, 173, 0, 80, 0, 0, 204, 0, 207, 0, 97, 181, 202, 
			0, 0, 0, 229, 0, 0, 112, 0, 0, 0, 0, 0, 130, 54, 180, 
			224, 0, 0, 63, 0, 0, 121, 0, 0, 0, 0, 0, 0, 0, 0, 
			46, 130, 0, 112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 149, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			

			90, 172, 38, 221, 206, 118, 17, 118, 141, 51, 183, 38, 63, 99, 161, 
			114, 194, 56, 115, 103, 0, 106, 116, 51, 0, 0, 0, 0, 229, 7, 
			101, 195, 117, 177, 71, 166, 41, 236, 0, 0, 0, 0, 0, 0, 112, 
			0, 0, 125, 65, 99, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 246, 0, 0, 0, 0, 0, 148, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			

			237, 105, 126, 203, 131, 140, 22, 170, 32, 68, 36, 210, 7, 57, 140, 
			182, 35, 178, 238, 141, 0, 90, 45, 153, 223, 0, 0, 86, 176, 50, 
			48, 106, 225, 56, 171, 217, 177, 165, 0, 0, 253, 0, 0, 233, 244, 
			0, 0, 21, 66, 181, 103, 0, 138, 0, 196, 154, 148, 172, 0, 127, 
			132, 0, 251, 220, 0, 0, 237, 0, 187, 0, 0, 0, 0, 0, 0, 
			117, 42, 164, 105, 54, 201, 0, 0, 0, 0, 193, 144, 206, 245, 0, 
			0, 0, 163, 230, 73, 0, 87, 0, 140, 0, 129, 0, 0, 0, 0, 
			0, 0, 0, 46, 146, 104, 233, 14, 212, 0, 90, 0, 178, 228, 0, 
			0, 81, 0, 91, 0, 73, 103, 0, 0, 0, 121, 20, 223, 0, 0, 
			249, 148, 24, 0, 165, 243, 0, 0, 0, 166, 30, 120, 0, 0, 166, 
			48, 69, 202, 0, 0, 0, 72, 151, 180, 0, 0, 0, 0, 94, 209, 
			64, 47, 161, 0, 74, 249, 123, 78, 91, 104, 0, 0, 0, 0, 0, 
			0, 169, 0, 187, 161, 0, 0, 0, 0, 0, 0, 0, 0, 101, 0, 
			0, 0, 213, 115, 137, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 
			0, 0, 0, 247, 202, 130, 248, 0, 0, 0, 0, 0, 0, 0, 0, 
			

			146, 78, 90, 41, 170, 210, 158, 129, 5, 70, 5, 169, 202, 201, 168, 
			158, 75, 105, 169, 126, 221, 11, 227, 90, 111, 47, 50, 42, 133, 87, 
			173, 197, 124, 134, 142, 5, 49, 59, 157, 134, 109, 203, 13, 238, 102, 
			5, 169, 75, 50, 85, 149, 2, 192, 6, 88, 182, 202, 166, 136, 199, 
			181, 40, 213, 78, 236, 133, 252, 211, 229, 13, 61, 189, 84, 43, 210, 
			6, 44, 119, 72, 80, 54, 92, 215, 15, 240, 129, 25, 58, 10, 16, 
			102, 230, 253, 33, 124, 112, 25, 22, 238, 113, 121, 140, 24, 30, 83, 
			123, 29, 242, 34, 102, 234, 190, 233, 75, 250, 135, 181, 31, 132, 227, 
			213, 196, 129, 223, 170, 207, 159, 141, 255, 217, 28, 147, 250, 63, 228, 
			183, 175, 233, 205, 201, 49, 93, 42, 156, 175, 100, 79, 111, 65, 150, 
			111, 185, 193, 128, 253, 21, 21, 221, 162, 68, 67, 58, 67, 105, 106, 
			168, 35, 163, 240, 52, 32, 132, 184, 195, 82, 174, 255, 139, 112, 242, 
			56, 175, 167, 29, 75, 73, 134, 86, 233, 36, 4, 202, 97, 189, 130, 
			66, 131, 183, 209, 193, 30, 245, 136, 230, 26, 203, 189, 87, 201, 128, 
			85, 226, 48, 83, 141, 7, 98, 109, 198, 109, 251, 96, 174, 3, 138, 
			

			0, 0, 0, 0, 0, 0, 0, 0, 0, 129, 115, 159, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 46, 203, 185, 0, 0, 220, 59, 0, 0, 
			69, 0, 0, 0, 0, 244, 39, 209, 0, 0, 0, 0, 61, 161, 0, 
			173, 0, 0, 0, 166, 0, 0, 120, 0, 0, 224, 237, 173, 34, 0, 
			0, 0, 183, 0, 0, 0, 213, 153, 96, 0, 0, 237, 0, 0, 53, 
			118, 0, 197, 75, 121, 42, 0, 0, 101, 0, 26, 133, 0, 0, 0, 
			60, 145, 45, 157, 0, 0, 9, 0, 78, 0, 196, 227, 0, 0, 0, 
			79, 0, 112, 0, 0, 0, 34, 24, 0, 0, 0, 69, 0, 94, 0, 
			0, 0, 2, 0, 25, 118, 15, 0, 0, 200, 32, 60, 30, 0, 0, 
			0, 0, 20, 0, 116, 172, 0, 0, 87, 226, 159, 158, 0, 0, 95, 
			0, 0, 73, 0, 0, 0, 0, 213, 241, 166, 0, 0, 0, 186, 205, 
			210, 0, 0, 0, 208, 150, 52, 246, 141, 167, 0, 151, 0, 0, 99, 
			143, 182, 0, 34, 128, 0, 183, 152, 0, 0, 0, 0, 235, 0, 0, 
			253, 209, 236, 90, 140, 0, 0, 22, 0, 0, 51, 33, 0, 0, 232, 
			91, 0, 75, 126, 85, 182, 158, 0, 0, 0, 42, 0, 0, 0, 20, 
			

			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 92, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 134, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 114, 0, 0, 0, 0, 131, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 215, 0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 21, 0, 0, 0, 4, 0, 0, 168, 0, 0, 
			0, 175, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 105, 0, 0, 
			0, 30, 0, 237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			232, 0, 0, 96, 0, 0, 174, 0, 0, 0, 189, 207, 18, 77, 211, 
			99, 206, 0, 44, 0, 91, 32, 101, 27, 194, 207, 32, 209, 109, 98, 
			71, 35, 37, 0, 0, 129, 193, 123, 92, 90, 224, 93, 185, 33, 1, 
			4, 135, 174, 0, 41, 194, 61, 113, 67, 75, 71, 200, 119, 0, 221, 
			62, 188, 2, 156, 140, 232, 167, 54, 105, 141, 33, 169, 185, 103, 183, 
			

			136, 34, 192, 135, 233, 157, 67, 75, 109, 204, 107, 53, 96, 106, 145, 
			206, 33, 74, 2, 123, 123, 0, 118, 0, 78, 0, 0, 13, 169, 44, 
			150, 147, 252, 150, 198, 87, 0, 0, 91, 83, 0, 0, 0, 166, 98, 
			0, 166, 47, 176, 178, 114, 58, 0, 0, 206, 0, 0, 0, 0, 115, 
			0, 161, 0, 194, 79, 70, 0, 0, 0, 10, 0, 0, 253, 0, 162, 
			0, 82, 0, 212, 205, 0, 0, 0, 0, 211, 0, 0, 129, 0, 0, 
			0, 0, 0, 0, 42, 66, 0, 0, 0, 65, 0, 0, 239, 140, 0, 
			0, 0, 0, 0, 73, 44, 0, 0, 0, 142, 0, 0, 212, 197, 0, 
			0, 0, 0, 119, 0, 0, 0, 217, 166, 0, 208, 0, 18, 131, 221, 
			0, 117, 0, 122, 0, 180, 21, 0, 0, 0, 0, 0, 213, 50, 105, 
			202, 0, 0, 57, 0, 0, 225, 0, 0, 0, 0, 47, 114, 206, 0, 
			69, 168, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 146, 186, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 129, 0, 
			0, 0, 35, 0, 0, 0, 0, 0, 115, 0, 0, 0, 140, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 133, 0, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 246, 0, 0, 0, 0, 217, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 192, 0, 0, 0, 0, 204, 0, 0, 
			0, 0, 0, 236, 105, 244, 0, 0, 0, 0, 88, 38, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 191, 0, 0, 
			

			66, 85, 17, 99, 110, 252, 233, 140, 204, 43, 237, 232, 232, 213, 138, 
			240, 157, 38, 39, 73, 250, 150, 203, 49, 167, 178, 99, 213, 19, 202, 
			252, 221, 46, 59, 173, 103, 124, 49, 25, 155, 22, 137, 99, 145, 5, 
			111, 124, 209, 143, 92, 227, 101, 79, 178, 85, 78, 166, 76, 54, 114, 
			122, 180, 32, 200, 43, 65, 240, 61, 144, 9, 252, 27, 131, 104, 78, 
			204, 136, 226, 191, 126, 70, 114, 210, 225, 196, 109, 37, 184, 122, 166, 
			243, 169, 209, 183, 61, 232, 11, 103, 243, 127, 32, 169, 237, 34, 16, 
			229, 80, 66, 144, 144, 94, 178, 73, 132, 118, 162, 4, 5, 31, 237, 
			217, 41, 158, 236, 194, 139, 227, 69, 21, 85, 59, 202, 128, 127, 255, 
			125, 250, 83, 82, 13, 255, 72, 32, 99, 190, 114, 10, 252, 217, 38, 
			46, 184, 72, 192, 55, 209, 238, 102, 243, 22, 91, 179, 233, 205, 1, 
			121, 237, 112, 227, 212, 20, 182, 185, 0, 0, 0, 0, 0, 0, 0, 
			0, 208, 128, 27, 138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 240, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 95, 
			0, 0, 0, 139, 0, 0, 0, 0, 0, 0, 0, 0, 0, 226, 0, 
			

			63, 130, 150, 251, 163, 94, 32, 202, 229, 245, 233, 0, 168, 24, 167, 
			150, 3, 60, 94, 202, 0, 10, 121, 133, 0, 209, 18, 0, 0, 207, 
			77, 0, 96, 233, 25, 89, 88, 75, 0, 0, 0, 0, 89, 0, 0, 
			114, 0, 24, 219, 166, 0, 184, 4, 0, 0, 16, 0, 0, 218, 0, 
			86, 0, 1, 0, 0, 12, 220, 89, 42, 0, 0, 90, 0, 171, 0, 
			54, 0, 30, 18, 0, 0, 0, 0, 148, 0, 3, 147, 0, 0, 151, 
			0, 214, 0, 196, 0, 0, 0, 0, 255, 0, 215, 179, 0, 0, 41, 
			0, 0, 107, 192, 0, 0, 116, 0, 0, 0, 0, 109, 0, 0, 0, 
			0, 0, 72, 0, 82, 0, 0, 0, 0, 9, 0, 46, 0, 0, 0, 
			0, 0, 180, 0, 219, 0, 0, 0, 146, 0, 136, 0, 0, 0, 4, 
			0, 0, 251, 0, 52, 98, 0, 0, 201, 114, 0, 0, 0, 0, 133, 
			0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 224, 212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
			
		others=>0 );
END ifmap_package;
