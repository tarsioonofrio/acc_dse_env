library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    18, 18, 15, 20, 23, 13, 15, 29, 29, 10, 0, 1, 6, 12, 21, 
    22, 18, 15, 19, 19, 4, 8, 3, 0, 4, 0, 0, 0, 5, 11, 
    0, 11, 19, 27, 18, 27, 32, 30, 0, 0, 0, 0, 0, 0, 1, 
    1, 0, 12, 25, 11, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 4, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 4, 7, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 26, 15, 
    63, 10, 0, 0, 0, 50, 58, 56, 37, 32, 34, 41, 37, 39, 32, 
    44, 58, 0, 0, 30, 29, 29, 32, 32, 31, 36, 30, 34, 40, 33, 
    48, 47, 47, 14, 15, 33, 25, 29, 34, 35, 47, 51, 52, 40, 58, 
    41, 51, 49, 65, 42, 48, 42, 31, 23, 28, 33, 45, 26, 28, 41, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 14, 6, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 2, 1, 0, 27, 0, 6, 0, 0, 0, 
    0, 30, 0, 0, 17, 20, 5, 3, 0, 29, 16, 0, 8, 0, 3, 
    15, 23, 0, 0, 26, 10, 6, 4, 0, 68, 3, 0, 11, 0, 2, 
    23, 11, 0, 0, 12, 30, 11, 0, 0, 55, 0, 4, 10, 17, 2, 
    32, 20, 6, 0, 6, 45, 0, 0, 0, 32, 0, 0, 17, 8, 0, 
    29, 40, 4, 17, 8, 0, 0, 11, 11, 0, 16, 0, 6, 0, 0, 
    24, 36, 0, 39, 14, 9, 18, 18, 21, 0, 0, 0, 12, 0, 0, 
    43, 35, 0, 88, 13, 40, 45, 17, 0, 0, 27, 34, 31, 11, 0, 
    54, 35, 18, 69, 0, 7, 31, 33, 26, 30, 34, 40, 46, 47, 47, 
    42, 56, 51, 37, 0, 39, 37, 36, 36, 42, 47, 54, 47, 46, 58, 
    44, 46, 82, 0, 19, 43, 38, 42, 42, 47, 46, 47, 42, 69, 40, 
    43, 51, 44, 25, 25, 40, 35, 36, 46, 49, 45, 46, 67, 58, 31, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 8, 23, 0, 31, 28, 3, 0, 0, 
    42, 0, 0, 0, 0, 0, 43, 17, 0, 0, 66, 45, 63, 0, 0, 
    113, 0, 0, 0, 14, 0, 40, 44, 37, 0, 90, 38, 59, 42, 0, 
    108, 5, 35, 0, 52, 36, 93, 72, 60, 0, 47, 82, 30, 62, 0, 
    89, 49, 55, 0, 0, 44, 97, 62, 96, 0, 115, 92, 18, 49, 37, 
    72, 115, 21, 56, 0, 0, 90, 74, 106, 0, 117, 71, 18, 12, 55, 
    77, 101, 40, 49, 0, 6, 139, 56, 70, 0, 79, 80, 6, 37, 19, 
    104, 66, 132, 11, 42, 19, 46, 44, 0, 41, 22, 91, 4, 0, 0, 
    74, 58, 159, 0, 100, 24, 0, 77, 48, 59, 90, 23, 0, 0, 12, 
    15, 60, 148, 0, 147, 76, 32, 113, 131, 65, 26, 29, 35, 32, 49, 
    29, 43, 78, 0, 216, 115, 58, 60, 71, 56, 61, 60, 62, 64, 79, 
    95, 18, 0, 130, 175, 66, 73, 63, 62, 57, 56, 64, 80, 72, 61, 
    106, 69, 0, 203, 90, 57, 77, 66, 60, 65, 72, 77, 78, 56, 123, 
    118, 75, 62, 84, 72, 53, 67, 68, 56, 68, 85, 58, 26, 111, 128, 
    
    -- channel=4
    0, 0, 8, 8, 6, 3, 5, 0, 4, 0, 0, 0, 0, 6, 5, 
    7, 10, 12, 7, 10, 73, 26, 0, 0, 0, 36, 6, 0, 0, 4, 
    0, 0, 4, 4, 7, 0, 0, 0, 13, 26, 21, 7, 23, 0, 0, 
    40, 37, 9, 5, 13, 0, 55, 27, 5, 0, 0, 0, 0, 1, 0, 
    38, 90, 19, 11, 128, 86, 6, 14, 0, 0, 37, 37, 15, 24, 0, 
    0, 0, 8, 0, 0, 0, 42, 26, 31, 58, 0, 0, 0, 9, 39, 
    6, 7, 0, 4, 0, 33, 0, 10, 9, 17, 0, 11, 0, 23, 29, 
    21, 7, 28, 16, 25, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 4, 11, 4, 28, 0, 0, 26, 4, 0, 0, 0, 0, 3, 47, 
    0, 0, 9, 4, 17, 0, 0, 74, 12, 0, 0, 0, 27, 31, 0, 
    0, 0, 0, 70, 156, 133, 40, 0, 0, 0, 32, 65, 27, 0, 0, 
    0, 0, 15, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 18, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 19, 4, 0, 40, 34, 0, 
    
    -- channel=5
    157, 163, 162, 165, 164, 157, 172, 183, 173, 148, 124, 124, 132, 146, 146, 
    162, 173, 168, 172, 160, 140, 169, 160, 122, 58, 46, 62, 78, 110, 139, 
    137, 106, 172, 176, 175, 142, 115, 72, 45, 7, 30, 10, 39, 58, 103, 
    77, 43, 164, 170, 162, 89, 77, 39, 21, 12, 51, 45, 27, 37, 58, 
    23, 31, 148, 96, 78, 71, 67, 47, 31, 0, 49, 57, 23, 28, 47, 
    22, 18, 142, 153, 37, 59, 69, 49, 45, 0, 62, 42, 16, 18, 23, 
    14, 42, 98, 159, 47, 50, 62, 45, 47, 0, 50, 40, 16, 14, 38, 
    28, 10, 44, 98, 55, 38, 46, 39, 41, 30, 47, 45, 9, 34, 65, 
    20, 0, 43, 14, 85, 34, 54, 48, 13, 84, 66, 38, 15, 45, 121, 
    16, 5, 36, 0, 53, 32, 8, 40, 45, 52, 29, 6, 9, 98, 138, 
    0, 21, 35, 0, 23, 26, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    34, 35, 37, 32, 30, 39, 38, 36, 29, 23, 26, 38, 36, 30, 24, 
    35, 44, 42, 31, 40, 32, 15, 29, 14, 29, 0, 9, 32, 43, 28, 
    6, 57, 40, 33, 39, 26, 0, 6, 33, 46, 0, 0, 0, 37, 44, 
    0, 76, 33, 41, 15, 36, 4, 0, 0, 72, 0, 9, 0, 0, 74, 
    0, 38, 2, 86, 9, 11, 0, 0, 0, 89, 0, 0, 6, 0, 43, 
    0, 10, 0, 26, 62, 19, 0, 0, 0, 142, 0, 0, 20, 0, 0, 
    0, 0, 32, 0, 63, 54, 0, 0, 0, 102, 0, 0, 10, 21, 0, 
    0, 0, 0, 0, 56, 66, 0, 0, 0, 66, 0, 0, 29, 15, 8, 
    0, 2, 0, 33, 4, 17, 0, 0, 36, 0, 37, 0, 30, 33, 35, 
    0, 0, 0, 44, 0, 15, 39, 0, 2, 5, 0, 12, 48, 52, 20, 
    42, 4, 0, 120, 0, 0, 34, 0, 0, 0, 8, 9, 1, 0, 0, 
    32, 20, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=7
    43, 48, 45, 44, 47, 41, 48, 58, 55, 42, 37, 38, 39, 42, 49, 
    44, 53, 48, 46, 45, 0, 31, 41, 59, 12, 0, 0, 14, 31, 37, 
    28, 41, 46, 53, 50, 59, 45, 35, 0, 0, 0, 0, 0, 4, 26, 
    0, 0, 35, 50, 37, 25, 0, 0, 0, 0, 0, 0, 6, 0, 17, 
    0, 0, 18, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 11, 56, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 58, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 26, 5, 0, 0, 15, 3, 24, 4, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 17, 10, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    10, 17, 8, 8, 4, 12, 12, 11, 11, 33, 45, 35, 17, 8, 6, 
    0, 10, 10, 12, 8, 0, 5, 35, 66, 0, 0, 0, 10, 23, 10, 
    53, 51, 5, 8, 5, 55, 22, 9, 0, 0, 0, 0, 0, 14, 12, 
    0, 0, 5, 8, 8, 0, 0, 2, 0, 26, 4, 16, 6, 0, 14, 
    1, 0, 2, 14, 0, 0, 9, 0, 7, 0, 0, 0, 0, 0, 0, 
    15, 0, 6, 3, 62, 40, 0, 0, 0, 0, 20, 21, 7, 0, 0, 
    0, 0, 28, 24, 18, 0, 49, 0, 17, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 53, 53, 33, 14, 0, 9, 0, 5, 14, 0, 
    0, 1, 0, 0, 0, 38, 0, 0, 0, 0, 38, 48, 0, 0, 0, 
    12, 0, 4, 0, 35, 9, 0, 0, 0, 78, 54, 17, 0, 0, 24, 
    3, 0, 7, 0, 0, 0, 30, 81, 55, 0, 0, 0, 0, 5, 10, 
    53, 33, 12, 0, 86, 40, 4, 5, 3, 0, 0, 0, 0, 0, 0, 
    0, 22, 0, 24, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 79, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 34, 0, 3, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    13, 19, 10, 14, 9, 21, 8, 6, 12, 28, 34, 27, 19, 6, 2, 
    8, 11, 9, 13, 15, 54, 15, 26, 31, 52, 53, 36, 33, 26, 10, 
    38, 36, 11, 10, 8, 81, 51, 40, 32, 83, 94, 75, 43, 25, 26, 
    51, 20, 14, 18, 25, 46, 69, 47, 54, 91, 93, 66, 59, 21, 27, 
    113, 94, 21, 53, 126, 68, 100, 59, 51, 59, 103, 56, 57, 37, 1, 
    127, 158, 40, 19, 189, 126, 125, 75, 46, 91, 127, 80, 71, 60, 21, 
    122, 148, 67, 23, 90, 117, 168, 101, 78, 120, 129, 70, 59, 76, 51, 
    142, 165, 64, 57, 57, 165, 133, 106, 80, 95, 120, 76, 72, 75, 38, 
    176, 184, 102, 115, 56, 102, 89, 78, 81, 51, 101, 65, 44, 43, 14, 
    192, 179, 134, 117, 111, 51, 95, 121, 66, 90, 64, 37, 47, 39, 39, 
    199, 171, 139, 162, 158, 101, 145, 185, 121, 60, 64, 71, 90, 113, 104, 
    193, 203, 157, 201, 231, 165, 138, 133, 124, 111, 120, 128, 136, 138, 142, 
    140, 161, 177, 229, 175, 122, 117, 112, 113, 118, 132, 140, 149, 154, 163, 
    157, 133, 166, 239, 136, 128, 121, 115, 119, 130, 140, 155, 147, 163, 171, 
    151, 143, 127, 167, 116, 127, 137, 126, 124, 136, 134, 133, 154, 175, 141, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 28, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 20, 51, 0, 0, 20, 30, 0, 0, 
    63, 0, 0, 0, 0, 62, 28, 40, 0, 0, 0, 0, 7, 30, 0, 
    25, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 26, 6, 14, 0, 
    0, 0, 9, 0, 0, 0, 15, 4, 29, 0, 0, 8, 0, 0, 37, 
    47, 0, 2, 79, 3, 0, 0, 0, 6, 0, 38, 28, 0, 0, 0, 
    0, 24, 13, 13, 0, 0, 5, 0, 9, 0, 24, 8, 0, 0, 0, 
    2, 0, 7, 0, 0, 0, 61, 30, 0, 0, 0, 28, 0, 16, 0, 
    0, 0, 46, 0, 34, 50, 3, 0, 0, 54, 38, 58, 13, 0, 0, 
    0, 0, 10, 0, 18, 21, 0, 0, 46, 31, 49, 1, 0, 0, 8, 
    0, 0, 34, 0, 0, 0, 0, 25, 15, 13, 0, 0, 0, 22, 33, 
    65, 0, 0, 0, 162, 82, 63, 55, 12, 6, 0, 2, 0, 0, 0, 
    13, 54, 0, 65, 86, 0, 2, 0, 0, 0, 0, 0, 3, 0, 0, 
    2, 0, 37, 62, 6, 0, 0, 1, 0, 0, 7, 10, 0, 0, 66, 
    12, 0, 24, 54, 36, 19, 9, 0, 0, 0, 5, 0, 0, 0, 4, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 31, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 5, 45, 0, 7, 0, 2, 1, 
    0, 2, 0, 0, 0, 0, 0, 0, 2, 59, 0, 0, 3, 0, 16, 
    1, 6, 0, 0, 44, 0, 0, 0, 0, 93, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 28, 15, 0, 0, 0, 82, 0, 0, 18, 19, 0, 
    4, 0, 0, 0, 12, 23, 0, 5, 0, 45, 0, 0, 29, 3, 0, 
    0, 22, 0, 17, 0, 18, 0, 0, 8, 0, 17, 0, 27, 0, 0, 
    9, 25, 0, 59, 0, 3, 16, 0, 5, 0, 0, 18, 18, 0, 0, 
    51, 13, 0, 88, 0, 0, 45, 4, 0, 2, 40, 51, 62, 44, 29, 
    112, 54, 0, 59, 0, 46, 78, 78, 68, 73, 79, 86, 88, 90, 83, 
    90, 111, 72, 8, 0, 73, 72, 74, 76, 84, 91, 91, 87, 93, 94, 
    90, 96, 138, 0, 49, 80, 69, 77, 83, 87, 97, 100, 97, 116, 94, 
    80, 103, 103, 65, 73, 95, 85, 73, 82, 82, 82, 94, 107, 83, 69, 
    
    -- channel=12
    47, 46, 51, 46, 47, 47, 49, 47, 43, 35, 28, 39, 38, 39, 36, 
    50, 50, 53, 45, 52, 85, 19, 37, 4, 33, 19, 21, 36, 45, 40, 
    26, 59, 52, 46, 56, 44, 0, 0, 26, 79, 10, 11, 4, 39, 57, 
    0, 121, 44, 54, 37, 35, 26, 8, 24, 83, 0, 18, 0, 14, 83, 
    0, 99, 10, 73, 44, 26, 0, 0, 8, 95, 11, 0, 30, 0, 57, 
    0, 56, 0, 46, 73, 0, 0, 0, 0, 191, 0, 0, 35, 4, 13, 
    0, 21, 12, 0, 97, 80, 10, 0, 0, 164, 0, 0, 30, 39, 13, 
    0, 0, 1, 0, 69, 104, 0, 8, 0, 124, 0, 0, 42, 34, 18, 
    0, 23, 0, 60, 17, 3, 0, 28, 49, 6, 34, 0, 38, 58, 68, 
    10, 24, 0, 74, 0, 25, 42, 14, 23, 10, 0, 5, 72, 86, 28, 
    81, 17, 0, 163, 0, 11, 86, 0, 0, 0, 20, 40, 45, 30, 0, 
    64, 40, 0, 152, 0, 0, 0, 0, 0, 9, 16, 16, 14, 17, 0, 
    3, 65, 72, 31, 0, 9, 5, 10, 8, 16, 20, 23, 16, 8, 23, 
    0, 16, 116, 0, 0, 17, 0, 9, 13, 16, 13, 9, 0, 38, 0, 
    0, 13, 25, 0, 0, 22, 12, 9, 24, 16, 0, 11, 49, 3, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 18, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 39, 0, 0, 56, 8, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 17, 0, 0, 
    0, 0, 0, 30, 48, 62, 0, 0, 0, 0, 28, 36, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 
    
    -- channel=14
    47, 54, 51, 53, 53, 48, 57, 59, 54, 43, 32, 32, 37, 40, 39, 
    48, 56, 54, 57, 51, 66, 59, 57, 35, 2, 2, 6, 6, 17, 39, 
    48, 19, 54, 57, 55, 61, 30, 0, 0, 0, 4, 0, 1, 0, 23, 
    21, 0, 50, 55, 64, 18, 30, 0, 0, 0, 23, 0, 0, 0, 0, 
    0, 18, 52, 16, 68, 51, 37, 6, 0, 0, 16, 9, 0, 0, 0, 
    0, 15, 49, 56, 11, 13, 43, 8, 11, 0, 42, 0, 0, 0, 0, 
    0, 44, 7, 61, 14, 17, 46, 23, 8, 3, 19, 0, 0, 0, 0, 
    4, 25, 0, 37, 0, 34, 46, 10, 0, 19, 15, 0, 0, 2, 0, 
    21, 17, 9, 0, 28, 0, 0, 12, 0, 44, 0, 0, 0, 0, 33, 
    22, 14, 20, 0, 3, 0, 0, 31, 6, 5, 0, 0, 0, 30, 40, 
    5, 20, 21, 0, 44, 6, 17, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    39, 34, 35, 41, 44, 32, 40, 43, 47, 50, 41, 29, 30, 41, 46, 
    40, 36, 36, 44, 33, 14, 67, 48, 46, 5, 33, 41, 25, 21, 44, 
    63, 2, 40, 41, 42, 32, 40, 36, 16, 0, 28, 12, 50, 26, 11, 
    92, 0, 46, 36, 56, 12, 39, 37, 25, 0, 35, 24, 26, 38, 0, 
    44, 5, 65, 0, 19, 39, 42, 36, 37, 0, 20, 56, 18, 43, 26, 
    36, 0, 55, 47, 0, 0, 22, 37, 67, 0, 52, 42, 7, 29, 32, 
    17, 36, 14, 70, 0, 0, 21, 28, 57, 0, 43, 40, 13, 0, 37, 
    11, 6, 41, 52, 2, 0, 53, 11, 24, 0, 17, 44, 0, 17, 13, 
    13, 0, 63, 0, 52, 0, 14, 27, 0, 63, 5, 43, 0, 0, 26, 
    0, 0, 57, 0, 42, 20, 0, 29, 44, 15, 47, 15, 0, 16, 47, 
    0, 0, 56, 0, 41, 50, 0, 5, 39, 43, 15, 8, 8, 17, 33, 
    0, 0, 0, 0, 82, 5, 0, 0, 0, 7, 3, 0, 0, 0, 3, 
    20, 0, 0, 34, 46, 0, 6, 2, 5, 1, 0, 0, 2, 0, 0, 
    9, 0, 0, 34, 13, 0, 9, 6, 0, 0, 1, 0, 0, 0, 21, 
    19, 0, 0, 4, 20, 0, 0, 0, 0, 0, 12, 0, 0, 18, 26, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 31, 18, 0, 
    0, 0, 0, 0, 0, 0, 19, 9, 0, 0, 0, 0, 0, 0, 0, 
    66, 69, 13, 0, 0, 4, 31, 10, 0, 0, 0, 3, 0, 14, 16, 
    37, 0, 9, 9, 0, 0, 0, 0, 25, 23, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 39, 32, 
    27, 55, 64, 62, 58, 49, 42, 33, 28, 20, 38, 33, 18, 10, 11, 
    55, 65, 63, 75, 80, 85, 86, 76, 66, 62, 50, 41, 30, 0, 0, 
    2, 10, 0, 0, 3, 11, 1, 0, 8, 2, 0, 0, 0, 0, 0, 
    0, 16, 24, 10, 6, 6, 34, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 3, 6, 4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    43, 43, 43, 43, 44, 43, 43, 43, 43, 44, 45, 42, 43, 43, 44, 
    43, 43, 43, 43, 43, 43, 44, 41, 43, 28, 40, 49, 44, 43, 44, 
    41, 43, 43, 43, 45, 44, 43, 35, 28, 26, 44, 43, 43, 43, 44, 
    50, 45, 44, 43, 44, 31, 47, 32, 44, 45, 51, 70, 43, 43, 43, 
    25, 34, 46, 41, 44, 32, 50, 41, 51, 49, 32, 20, 23, 41, 43, 
    50, 56, 47, 33, 37, 18, 19, 23, 29, 30, 43, 50, 38, 75, 46, 
    22, 31, 41, 39, 27, 5, 33, 59, 85, 45, 32, 21, 25, 20, 38, 
    30, 59, 21, 52, 39, 46, 67, 33, 25, 28, 32, 42, 47, 53, 59, 
    107, 42, 48, 55, 50, 35, 40, 23, 39, 35, 37, 30, 24, 20, 25, 
    46, 29, 37, 39, 41, 43, 39, 44, 48, 40, 40, 31, 41, 36, 36, 
    12, 23, 26, 23, 20, 25, 33, 34, 29, 28, 31, 35, 41, 44, 37, 
    0, 18, 1, 0, 0, 13, 43, 47, 45, 49, 54, 60, 33, 24, 36, 
    0, 0, 2, 0, 0, 0, 63, 33, 38, 32, 14, 14, 31, 25, 38, 
    0, 0, 0, 0, 0, 0, 27, 39, 18, 7, 21, 23, 13, 26, 35, 
    0, 0, 0, 0, 0, 0, 3, 6, 10, 21, 13, 8, 17, 26, 36, 
    
    -- channel=19
    82, 79, 79, 79, 78, 79, 79, 81, 77, 82, 81, 79, 79, 79, 78, 
    82, 79, 79, 80, 78, 79, 77, 79, 84, 128, 49, 58, 80, 78, 78, 
    81, 78, 78, 79, 76, 86, 74, 111, 100, 113, 49, 39, 81, 78, 79, 
    69, 81, 76, 78, 80, 121, 42, 111, 67, 80, 55, 17, 82, 79, 78, 
    63, 34, 33, 75, 79, 100, 53, 87, 72, 106, 122, 104, 91, 9, 72, 
    73, 52, 75, 84, 84, 127, 94, 88, 62, 100, 75, 67, 96, 0, 68, 
    81, 28, 58, 41, 124, 128, 3, 0, 0, 98, 116, 116, 95, 102, 37, 
    0, 20, 55, 0, 57, 76, 40, 118, 80, 72, 64, 39, 22, 35, 42, 
    0, 93, 69, 64, 77, 109, 97, 133, 89, 105, 100, 124, 98, 85, 73, 
    32, 94, 85, 90, 85, 84, 97, 77, 76, 91, 77, 83, 60, 55, 40, 
    43, 15, 56, 52, 48, 46, 74, 78, 84, 84, 69, 51, 24, 43, 28, 
    46, 0, 58, 55, 29, 2, 0, 44, 23, 15, 0, 29, 58, 44, 6, 
    55, 0, 10, 35, 18, 8, 0, 70, 68, 82, 73, 27, 13, 12, 6, 
    117, 9, 6, 15, 9, 7, 0, 34, 61, 6, 0, 1, 28, 11, 16, 
    98, 10, 4, 5, 2, 0, 0, 0, 0, 0, 24, 29, 19, 19, 21, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 40, 58, 74, 45, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 5, 23, 8, 0, 0, 0, 0, 0, 
    118, 124, 23, 0, 0, 0, 0, 0, 0, 0, 50, 95, 98, 86, 0, 
    0, 0, 0, 0, 22, 0, 0, 35, 78, 0, 0, 0, 0, 0, 0, 
    0, 114, 0, 0, 0, 121, 163, 23, 0, 0, 0, 19, 40, 68, 61, 
    111, 36, 102, 78, 11, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 9, 
    0, 0, 25, 32, 4, 0, 77, 142, 83, 85, 99, 112, 29, 0, 28, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 28, 30, 
    25, 3, 0, 0, 0, 0, 0, 0, 0, 0, 66, 68, 5, 10, 3, 
    0, 34, 29, 20, 22, 25, 12, 0, 73, 80, 29, 0, 11, 16, 14, 
    
    -- channel=21
    23, 21, 21, 21, 21, 21, 21, 24, 23, 22, 16, 21, 22, 21, 21, 
    23, 22, 22, 22, 21, 22, 21, 23, 26, 33, 0, 14, 22, 22, 22, 
    21, 22, 21, 23, 22, 25, 15, 31, 7, 0, 0, 0, 22, 22, 21, 
    7, 12, 18, 24, 24, 39, 7, 19, 0, 0, 0, 0, 12, 15, 17, 
    0, 0, 0, 23, 22, 18, 17, 17, 8, 10, 1, 0, 2, 0, 9, 
    0, 0, 11, 31, 17, 25, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 13, 1, 0, 0, 0, 16, 12, 8, 0, 0, 0, 
    0, 0, 1, 2, 0, 0, 0, 20, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 7, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    34, 10, 21, 22, 10, 9, 0, 82, 89, 87, 68, 32, 29, 8, 0, 
    48, 11, 13, 12, 10, 9, 50, 188, 167, 76, 45, 34, 19, 7, 0, 
    33, 20, 13, 10, 11, 7, 27, 65, 50, 40, 39, 20, 12, 3, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 29, 0, 0, 0, 
    0, 20, 25, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 37, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 49, 0, 
    0, 27, 18, 9, 0, 0, 8, 32, 62, 0, 0, 0, 0, 0, 22, 
    54, 21, 0, 52, 0, 0, 11, 0, 0, 0, 0, 0, 8, 6, 13, 
    162, 0, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 
    0, 19, 5, 11, 16, 18, 6, 7, 0, 0, 0, 8, 19, 10, 18, 
    0, 53, 0, 0, 6, 31, 56, 0, 0, 13, 29, 28, 13, 5, 30, 
    0, 27, 32, 9, 12, 19, 157, 57, 50, 33, 19, 27, 35, 22, 26, 
    0, 16, 22, 17, 18, 18, 108, 129, 87, 67, 55, 38, 5, 20, 17, 
    0, 3, 9, 9, 15, 15, 40, 63, 59, 53, 12, 0, 12, 11, 12, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 26, 27, 35, 38, 37, 15, 4, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 1, 18, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 23, 48, 46, 29, 26, 14, 67, 57, 56, 64, 50, 0, 0, 0, 
    0, 23, 28, 30, 26, 25, 31, 153, 165, 89, 0, 0, 0, 0, 0, 
    1, 7, 9, 10, 14, 12, 11, 69, 10, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    2, 1, 1, 1, 2, 3, 2, 2, 1, 3, 4, 2, 2, 1, 1, 
    2, 1, 1, 1, 1, 0, 1, 0, 2, 28, 14, 0, 0, 0, 0, 
    10, 7, 1, 0, 0, 4, 6, 17, 42, 36, 37, 22, 1, 1, 1, 
    0, 0, 0, 2, 2, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 49, 12, 9, 4, 1, 0, 2, 0, 12, 57, 64, 67, 42, 0, 
    0, 0, 0, 45, 40, 130, 137, 120, 71, 0, 0, 0, 0, 0, 1, 
    77, 68, 52, 2, 0, 0, 0, 0, 0, 37, 85, 102, 105, 82, 57, 
    8, 0, 0, 0, 0, 0, 0, 4, 28, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 26, 36, 56, 75, 32, 71, 65, 79, 86, 63, 28, 
    60, 91, 74, 72, 53, 39, 18, 0, 8, 5, 17, 18, 5, 13, 0, 
    10, 0, 24, 50, 71, 86, 95, 94, 76, 64, 43, 17, 0, 0, 0, 
    18, 19, 8, 0, 0, 1, 0, 0, 0, 0, 0, 0, 23, 1, 0, 
    0, 0, 28, 23, 3, 0, 36, 93, 77, 89, 87, 26, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 5, 96, 120, 26, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    239, 239, 239, 239, 239, 240, 240, 239, 237, 241, 243, 239, 240, 239, 240, 
    241, 240, 240, 240, 240, 240, 240, 239, 239, 233, 238, 241, 239, 240, 241, 
    241, 240, 240, 241, 240, 240, 242, 237, 236, 222, 207, 243, 242, 242, 243, 
    247, 245, 246, 242, 242, 235, 235, 229, 205, 196, 181, 215, 250, 248, 248, 
    210, 222, 253, 240, 241, 242, 224, 241, 234, 243, 240, 233, 224, 243, 252, 
    170, 172, 211, 220, 238, 230, 243, 247, 252, 245, 210, 185, 162, 183, 247, 
    189, 201, 223, 208, 211, 117, 107, 131, 182, 236, 238, 228, 231, 219, 233, 
    86, 117, 130, 173, 222, 177, 169, 190, 207, 194, 160, 143, 142, 163, 174, 
    80, 209, 177, 192, 228, 244, 255, 233, 193, 198, 212, 201, 198, 199, 194, 
    146, 203, 209, 213, 212, 212, 201, 174, 180, 155, 154, 143, 128, 127, 138, 
    49, 72, 76, 81, 92, 112, 139, 139, 138, 122, 111, 104, 107, 104, 117, 
    0, 23, 26, 0, 0, 0, 48, 26, 39, 41, 46, 66, 86, 107, 121, 
    0, 0, 5, 0, 0, 0, 58, 69, 37, 41, 59, 81, 83, 106, 151, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 14, 31, 63, 103, 127, 173, 
    30, 0, 0, 0, 0, 0, 0, 1, 0, 33, 79, 106, 118, 140, 179, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 30, 53, 23, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    115, 73, 0, 0, 0, 0, 0, 0, 0, 0, 50, 79, 97, 0, 0, 
    0, 0, 1, 47, 23, 117, 84, 59, 9, 0, 0, 0, 0, 0, 0, 
    123, 87, 31, 0, 3, 52, 0, 0, 0, 18, 58, 81, 39, 76, 24, 
    0, 0, 31, 7, 0, 0, 0, 43, 70, 41, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 37, 0, 0, 12, 0, 36, 51, 76, 42, 
    47, 84, 89, 83, 71, 49, 47, 30, 32, 25, 46, 23, 1, 2, 0, 
    94, 48, 95, 102, 110, 107, 100, 93, 80, 73, 47, 22, 0, 0, 0, 
    6, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 24, 37, 26, 3, 3, 20, 0, 0, 7, 62, 17, 0, 0, 0, 
    24, 0, 3, 4, 0, 0, 0, 21, 70, 2, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    8, 10, 10, 10, 11, 10, 10, 8, 10, 11, 13, 9, 10, 10, 11, 
    9, 11, 11, 10, 11, 11, 12, 10, 11, 6, 43, 26, 10, 11, 12, 
    10, 11, 11, 10, 11, 9, 16, 9, 26, 16, 50, 42, 10, 12, 12, 
    26, 16, 14, 10, 10, 0, 34, 0, 21, 16, 27, 54, 16, 15, 14, 
    73, 75, 49, 12, 12, 0, 22, 4, 20, 15, 26, 39, 45, 67, 21, 
    4, 16, 18, 18, 24, 21, 44, 40, 42, 12, 12, 9, 0, 64, 24, 
    73, 92, 54, 29, 0, 0, 69, 70, 68, 16, 19, 24, 29, 32, 62, 
    81, 50, 26, 71, 25, 0, 21, 13, 43, 41, 36, 39, 43, 33, 45, 
    127, 2, 2, 12, 25, 17, 32, 0, 19, 30, 35, 29, 48, 55, 50, 
    89, 67, 80, 78, 78, 71, 57, 61, 66, 51, 65, 52, 58, 53, 52, 
    60, 84, 75, 84, 87, 97, 98, 91, 78, 72, 73, 71, 69, 43, 43, 
    11, 52, 0, 3, 19, 42, 74, 31, 52, 52, 46, 30, 26, 22, 35, 
    0, 39, 30, 11, 17, 24, 95, 0, 0, 0, 0, 18, 19, 26, 39, 
    0, 18, 22, 17, 18, 19, 36, 0, 0, 0, 3, 15, 12, 32, 41, 
    0, 5, 15, 16, 16, 20, 34, 3, 0, 9, 4, 10, 20, 27, 37, 
    
    -- channel=28
    16, 19, 19, 19, 20, 19, 19, 18, 20, 19, 20, 20, 20, 19, 21, 
    15, 19, 19, 18, 19, 18, 19, 18, 16, 0, 33, 31, 18, 19, 20, 
    16, 18, 20, 18, 20, 17, 20, 1, 0, 0, 49, 51, 18, 19, 20, 
    26, 19, 23, 20, 19, 0, 43, 0, 17, 9, 28, 76, 19, 21, 22, 
    0, 13, 63, 18, 19, 0, 47, 10, 31, 12, 2, 0, 0, 44, 29, 
    40, 63, 49, 3, 25, 0, 14, 18, 26, 0, 7, 25, 3, 107, 31, 
    0, 10, 17, 38, 1, 0, 21, 53, 92, 20, 2, 0, 7, 5, 33, 
    44, 98, 1, 73, 10, 14, 80, 14, 0, 0, 0, 8, 30, 36, 59, 
    197, 27, 43, 57, 42, 8, 21, 0, 30, 18, 28, 8, 14, 2, 0, 
    96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 21, 33, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 28, 45, 
    0, 65, 11, 4, 11, 29, 88, 5, 15, 22, 40, 53, 37, 17, 55, 
    0, 39, 16, 0, 12, 25, 136, 0, 0, 0, 0, 0, 33, 53, 71, 
    0, 24, 28, 15, 23, 25, 85, 7, 0, 0, 44, 68, 36, 53, 62, 
    0, 26, 31, 28, 29, 30, 62, 24, 38, 83, 46, 31, 46, 53, 61, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 0, 0, 0, 
    0, 27, 0, 0, 0, 45, 63, 0, 0, 0, 0, 0, 0, 16, 0, 
    77, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 18, 7, 0, 69, 98, 63, 62, 74, 61, 0, 0, 0, 
    19, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 11, 3, 1, 9, 9, 0, 0, 0, 0, 32, 12, 0, 0, 0, 
    0, 32, 28, 25, 27, 28, 12, 0, 44, 36, 0, 0, 0, 0, 0, 
    
    -- channel=30
    44, 44, 44, 44, 44, 44, 44, 45, 44, 45, 42, 44, 44, 44, 44, 
    44, 44, 44, 44, 43, 44, 43, 43, 46, 48, 17, 32, 44, 43, 44, 
    43, 44, 44, 44, 44, 47, 39, 49, 23, 9, 13, 23, 43, 44, 44, 
    31, 38, 41, 45, 46, 57, 25, 41, 14, 15, 10, 21, 39, 40, 42, 
    0, 0, 16, 43, 43, 42, 42, 40, 38, 39, 31, 17, 9, 0, 38, 
    17, 27, 54, 32, 36, 25, 14, 16, 15, 31, 11, 18, 26, 17, 36, 
    0, 0, 0, 7, 49, 0, 0, 0, 0, 43, 34, 25, 12, 30, 0, 
    0, 3, 0, 4, 6, 5, 23, 49, 12, 0, 0, 0, 0, 0, 12, 
    0, 38, 20, 41, 41, 40, 29, 12, 17, 12, 7, 14, 1, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 44, 56, 48, 28, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 74, 52, 1, 0, 6, 4, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 0, 0, 3, 9, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 5, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 16, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 30, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 42, 0, 0, 1, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 19, 43, 34, 12, 0, 36, 7, 0, 0, 0, 0, 0, 0, 
    73, 22, 5, 22, 26, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    93, 30, 25, 28, 29, 28, 0, 0, 0, 0, 0, 11, 11, 0, 0, 
    75, 44, 39, 36, 31, 31, 11, 0, 0, 2, 18, 13, 3, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 24, 46, 46, 61, 22, 0, 0, 
    32, 23, 30, 26, 20, 15, 16, 11, 5, 4, 15, 0, 0, 0, 9, 
    10, 0, 0, 8, 0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 
    12, 7, 19, 18, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 16, 0, 0, 0, 0, 
    13, 37, 33, 10, 8, 21, 25, 7, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 19, 16, 0, 0, 0, 12, 0, 0, 0, 2, 17, 22, 
    27, 13, 8, 11, 27, 28, 9, 30, 17, 4, 18, 24, 9, 13, 7, 
    30, 21, 21, 30, 15, 7, 7, 3, 15, 15, 10, 27, 10, 15, 13, 
    26, 27, 31, 25, 36, 40, 16, 5, 19, 29, 9, 14, 14, 14, 10, 
    38, 37, 25, 18, 15, 21, 27, 20, 5, 0, 18, 11, 13, 10, 5, 
    8, 9, 11, 11, 7, 3, 10, 12, 20, 10, 11, 11, 11, 11, 8, 
    
    -- channel=34
    47, 60, 63, 58, 58, 53, 50, 42, 51, 51, 40, 47, 45, 47, 51, 
    41, 52, 56, 47, 47, 43, 45, 41, 47, 25, 47, 50, 43, 44, 50, 
    33, 43, 46, 36, 37, 35, 32, 34, 42, 0, 60, 39, 31, 35, 45, 
    23, 42, 39, 33, 26, 33, 23, 25, 7, 11, 26, 28, 37, 21, 25, 
    15, 15, 16, 21, 14, 18, 21, 14, 22, 25, 25, 39, 30, 13, 21, 
    32, 35, 17, 29, 36, 38, 39, 28, 27, 27, 48, 45, 13, 22, 5, 
    36, 27, 24, 42, 50, 42, 52, 47, 49, 45, 54, 34, 11, 25, 0, 
    46, 46, 56, 63, 59, 55, 53, 46, 41, 17, 25, 32, 27, 0, 35, 
    49, 28, 57, 58, 53, 40, 33, 33, 46, 25, 43, 33, 28, 27, 18, 
    45, 66, 49, 44, 46, 50, 45, 31, 22, 33, 38, 28, 12, 4, 9, 
    46, 49, 49, 33, 36, 35, 21, 15, 45, 30, 13, 8, 5, 3, 3, 
    53, 42, 26, 30, 38, 55, 17, 13, 20, 19, 9, 1, 12, 5, 2, 
    39, 24, 16, 18, 13, 17, 21, 19, 10, 6, 10, 13, 1, 8, 7, 
    13, 12, 10, 15, 11, 5, 9, 9, 21, 8, 7, 9, 6, 10, 9, 
    4, 8, 8, 10, 12, 12, 10, 3, 21, 0, 10, 9, 9, 10, 0, 
    
    -- channel=35
    120, 43, 68, 85, 87, 81, 81, 103, 66, 85, 86, 72, 86, 87, 67, 
    114, 39, 56, 87, 80, 81, 84, 83, 67, 143, 17, 60, 90, 90, 62, 
    111, 34, 44, 78, 74, 75, 103, 65, 51, 186, 0, 52, 97, 78, 55, 
    108, 35, 68, 60, 80, 61, 92, 100, 102, 90, 25, 26, 0, 78, 43, 
    66, 46, 57, 37, 58, 53, 57, 107, 80, 78, 48, 26, 14, 86, 32, 
    18, 24, 80, 14, 39, 47, 62, 92, 62, 61, 0, 29, 115, 27, 91, 
    46, 56, 64, 9, 38, 67, 65, 62, 51, 52, 10, 51, 107, 68, 113, 
    58, 59, 49, 56, 71, 79, 88, 99, 83, 124, 24, 33, 64, 104, 21, 
    86, 80, 32, 66, 100, 96, 81, 70, 49, 93, 26, 56, 64, 76, 68, 
    73, 38, 69, 84, 63, 66, 79, 97, 56, 62, 63, 95, 91, 89, 43, 
    51, 76, 84, 101, 74, 49, 115, 77, 0, 63, 86, 86, 71, 54, 59, 
    14, 67, 111, 57, 39, 28, 115, 76, 41, 56, 68, 51, 52, 42, 45, 
    34, 81, 96, 68, 56, 47, 49, 51, 56, 49, 48, 31, 62, 32, 31, 
    37, 34, 36, 29, 41, 38, 33, 42, 4, 71, 37, 37, 35, 26, 33, 
    30, 17, 20, 18, 23, 29, 35, 48, 0, 81, 30, 33, 28, 22, 62, 
    
    -- channel=36
    8, 5, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 13, 0, 0, 
    10, 29, 12, 0, 50, 33, 15, 0, 0, 8, 45, 105, 69, 0, 6, 
    3, 0, 0, 0, 0, 16, 32, 50, 79, 64, 52, 0, 0, 0, 0, 
    35, 58, 94, 89, 47, 31, 22, 7, 0, 0, 0, 0, 0, 16, 114, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 32, 64, 12, 0, 2, 0, 
    0, 67, 23, 0, 0, 25, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 5, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 1, 10, 2, 11, 13, 13, 15, 14, 11, 
    0, 0, 0, 0, 1, 13, 18, 9, 10, 37, 0, 15, 25, 22, 17, 
    0, 0, 0, 19, 26, 23, 33, 17, 9, 36, 0, 0, 29, 30, 22, 
    16, 7, 33, 31, 49, 36, 35, 36, 19, 0, 0, 16, 0, 35, 36, 
    1, 4, 13, 20, 31, 28, 9, 1, 0, 0, 0, 0, 2, 46, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 20, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 35, 52, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 24, 26, 24, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 8, 20, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 9, 12, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    
    -- channel=38
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 12, 4, 0, 0, 0, 0, 0, 0, 0, 35, 9, 0, 0, 5, 
    0, 15, 11, 0, 0, 0, 0, 1, 13, 0, 70, 14, 0, 0, 9, 
    0, 25, 14, 15, 0, 4, 0, 0, 0, 0, 5, 21, 65, 0, 23, 
    1, 9, 3, 25, 13, 16, 6, 0, 0, 0, 0, 21, 25, 0, 18, 
    14, 17, 0, 12, 0, 0, 0, 0, 0, 0, 37, 18, 0, 24, 0, 
    1, 0, 0, 23, 10, 0, 0, 0, 0, 0, 33, 7, 0, 4, 0, 
    0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 20, 23, 0, 0, 8, 
    0, 0, 18, 0, 0, 0, 0, 0, 2, 0, 20, 0, 0, 0, 0, 
    0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 
    0, 2, 0, 6, 0, 0, 0, 0, 17, 0, 0, 1, 0, 5, 3, 
    2, 8, 3, 4, 2, 0, 0, 0, 34, 0, 6, 4, 4, 8, 0, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    1, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 9, 10, 1, 21, 14, 3, 5, 8, 0, 
    4, 0, 0, 0, 1, 4, 10, 35, 30, 30, 18, 45, 17, 15, 9, 
    38, 15, 45, 44, 37, 21, 29, 15, 36, 26, 0, 18, 78, 63, 59, 
    63, 39, 38, 53, 66, 71, 58, 57, 22, 9, 3, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 13, 1, 0, 0, 0, 0, 13, 12, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 5, 27, 47, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 28, 16, 12, 10, 0, 0, 
    22, 35, 0, 1, 19, 26, 1, 0, 0, 0, 0, 0, 1, 14, 47, 
    0, 0, 0, 0, 0, 0, 0, 40, 43, 4, 0, 28, 51, 46, 24, 
    0, 0, 0, 35, 48, 19, 0, 0, 0, 38, 50, 34, 28, 18, 23, 
    0, 0, 0, 0, 0, 0, 66, 30, 0, 4, 28, 5, 0, 3, 4, 
    27, 55, 67, 40, 18, 6, 4, 7, 27, 9, 2, 5, 14, 0, 0, 
    4, 10, 4, 5, 15, 16, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 2, 7, 0, 0, 0, 0, 13, 
    
    -- channel=41
    223, 195, 243, 245, 251, 241, 248, 249, 244, 256, 246, 251, 245, 253, 244, 
    221, 191, 236, 233, 244, 229, 239, 249, 240, 238, 222, 248, 243, 254, 241, 
    212, 176, 218, 218, 228, 219, 224, 218, 230, 208, 189, 243, 237, 238, 236, 
    195, 156, 193, 203, 204, 203, 206, 185, 168, 165, 122, 140, 211, 210, 200, 
    151, 126, 147, 151, 164, 169, 178, 184, 141, 121, 116, 100, 104, 141, 125, 
    96, 94, 108, 99, 121, 121, 145, 144, 125, 124, 115, 142, 107, 157, 88, 
    116, 105, 111, 116, 160, 160, 162, 146, 134, 139, 143, 176, 173, 115, 83, 
    134, 128, 138, 153, 184, 198, 207, 194, 196, 165, 152, 162, 162, 101, 71, 
    160, 159, 176, 207, 210, 208, 200, 186, 168, 156, 129, 150, 161, 145, 150, 
    139, 144, 169, 181, 187, 181, 181, 175, 170, 180, 170, 167, 150, 127, 100, 
    175, 176, 176, 169, 169, 187, 171, 121, 111, 164, 158, 139, 104, 80, 61, 
    148, 169, 158, 121, 117, 144, 157, 110, 102, 115, 102, 89, 65, 48, 34, 
    124, 142, 141, 109, 106, 111, 100, 87, 88, 85, 68, 56, 53, 34, 27, 
    57, 61, 60, 60, 63, 65, 69, 64, 64, 55, 49, 36, 33, 28, 27, 
    24, 22, 31, 35, 43, 44, 50, 44, 55, 57, 31, 26, 27, 30, 12, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 31, 7, 69, 0, 3, 11, 0, 0, 
    18, 1, 18, 0, 10, 0, 1, 11, 110, 70, 70, 139, 16, 29, 31, 
    70, 64, 74, 81, 80, 79, 61, 61, 4, 3, 0, 0, 0, 27, 71, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 11, 0, 39, 
    0, 10, 17, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 80, 56, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 54, 17, 0, 0, 0, 0, 
    20, 39, 5, 0, 17, 28, 21, 0, 0, 0, 0, 0, 2, 0, 31, 
    0, 0, 0, 26, 0, 0, 0, 34, 15, 0, 0, 23, 54, 66, 44, 
    0, 0, 5, 23, 46, 0, 37, 44, 2, 28, 58, 54, 35, 19, 35, 
    0, 2, 28, 14, 0, 3, 32, 5, 15, 22, 36, 22, 16, 19, 11, 
    14, 45, 40, 27, 44, 41, 6, 7, 35, 26, 7, 11, 20, 3, 0, 
    44, 31, 16, 5, 12, 21, 21, 16, 0, 22, 7, 11, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 18, 0, 24, 5, 2, 0, 0, 35, 
    
    -- channel=43
    36, 69, 59, 46, 39, 32, 25, 9, 29, 20, 14, 19, 12, 14, 20, 
    26, 57, 48, 26, 25, 20, 20, 17, 23, 2, 50, 22, 7, 10, 21, 
    13, 45, 36, 9, 11, 10, 3, 27, 33, 0, 83, 37, 2, 8, 23, 
    3, 33, 17, 9, 0, 6, 0, 4, 31, 30, 73, 75, 71, 7, 16, 
    42, 51, 40, 50, 31, 36, 38, 18, 32, 40, 53, 28, 32, 0, 40, 
    54, 44, 20, 45, 37, 38, 52, 37, 44, 36, 51, 17, 0, 11, 0, 
    59, 46, 38, 77, 65, 49, 54, 45, 43, 38, 51, 20, 0, 2, 0, 
    50, 38, 43, 53, 52, 51, 49, 46, 48, 17, 48, 26, 7, 0, 4, 
    64, 62, 85, 73, 62, 62, 59, 45, 44, 0, 28, 18, 19, 9, 8, 
    53, 71, 61, 60, 62, 53, 42, 34, 47, 35, 31, 16, 23, 19, 35, 
    80, 65, 61, 48, 66, 68, 31, 37, 75, 47, 36, 28, 28, 26, 27, 
    95, 66, 44, 58, 61, 75, 22, 32, 49, 40, 35, 37, 32, 35, 23, 
    75, 56, 43, 53, 58, 57, 46, 42, 44, 42, 33, 42, 25, 36, 32, 
    56, 55, 49, 51, 44, 44, 48, 40, 48, 22, 35, 36, 33, 36, 31, 
    29, 37, 38, 40, 38, 37, 39, 28, 65, 13, 37, 33, 37, 37, 13, 
    
    -- channel=44
    0, 31, 40, 18, 25, 17, 25, 9, 35, 25, 7, 26, 9, 22, 22, 
    0, 30, 42, 12, 30, 14, 23, 23, 27, 0, 31, 35, 5, 20, 27, 
    0, 22, 45, 12, 33, 14, 12, 19, 30, 0, 89, 40, 3, 23, 34, 
    0, 24, 34, 24, 13, 23, 0, 14, 0, 0, 18, 2, 55, 26, 25, 
    0, 7, 0, 24, 3, 10, 0, 0, 0, 8, 18, 34, 59, 14, 19, 
    42, 33, 10, 28, 35, 21, 28, 0, 16, 15, 62, 70, 0, 49, 0, 
    35, 9, 0, 49, 27, 3, 13, 6, 27, 31, 76, 33, 0, 12, 0, 
    20, 24, 39, 50, 34, 25, 19, 12, 15, 0, 34, 32, 9, 0, 37, 
    11, 0, 33, 26, 7, 2, 4, 3, 28, 0, 61, 27, 11, 7, 12, 
    0, 51, 37, 7, 10, 26, 27, 12, 13, 23, 22, 3, 0, 0, 4, 
    35, 15, 15, 0, 21, 28, 0, 0, 47, 31, 0, 0, 0, 0, 11, 
    65, 12, 0, 0, 17, 62, 0, 4, 24, 8, 3, 0, 3, 11, 0, 
    47, 8, 0, 11, 10, 4, 4, 23, 13, 7, 5, 27, 0, 15, 15, 
    10, 8, 13, 26, 25, 20, 16, 10, 37, 5, 12, 14, 11, 23, 23, 
    18, 26, 26, 26, 26, 29, 26, 11, 57, 0, 20, 13, 21, 26, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 2, 0, 0, 7, 0, 0, 0, 0, 0, 24, 34, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 30, 19, 0, 0, 0, 0, 0, 
    3, 18, 44, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    5, 0, 8, 15, 25, 25, 36, 44, 36, 42, 38, 41, 40, 47, 36, 
    13, 0, 16, 25, 36, 33, 42, 41, 36, 55, 0, 42, 43, 50, 39, 
    22, 0, 22, 33, 46, 35, 49, 28, 21, 48, 0, 27, 45, 46, 39, 
    28, 0, 38, 36, 51, 38, 41, 39, 16, 0, 0, 0, 0, 42, 28, 
    0, 0, 0, 0, 6, 7, 0, 4, 0, 0, 0, 0, 8, 39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 44, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 23, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 9, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 20, 10, 6, 20, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 1, 8, 13, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 2, 0, 0, 56, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 16, 29, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 12, 0, 0, 1, 19, 0, 
    0, 1, 25, 0, 0, 11, 0, 10, 4, 8, 0, 0, 64, 0, 56, 
    0, 7, 7, 0, 0, 0, 0, 0, 6, 6, 0, 0, 7, 38, 38, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 27, 0, 0, 0, 38, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 4, 0, 5, 7, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 8, 14, 19, 2, 
    0, 0, 0, 1, 0, 0, 25, 15, 0, 0, 7, 12, 19, 18, 28, 
    0, 0, 19, 0, 0, 0, 12, 8, 5, 9, 24, 17, 22, 22, 23, 
    0, 0, 2, 2, 5, 0, 0, 14, 20, 11, 18, 15, 27, 17, 21, 
    10, 2, 10, 7, 16, 16, 13, 18, 0, 48, 15, 20, 19, 18, 22, 
    21, 18, 20, 18, 18, 21, 24, 27, 0, 41, 18, 16, 20, 14, 45, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 36, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 41, 20, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 5, 45, 66, 38, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 17, 22, 27, 32, 13, 1, 19, 31, 4, 17, 1, 20, 31, 22, 
    0, 0, 0, 0, 0, 0, 0, 6, 9, 15, 20, 24, 27, 26, 33, 
    10, 17, 15, 11, 4, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    
    -- channel=50
    50, 53, 41, 42, 48, 46, 43, 46, 45, 46, 46, 44, 51, 50, 46, 
    52, 57, 49, 35, 66, 50, 40, 48, 42, 45, 39, 46, 57, 52, 52, 
    52, 54, 54, 38, 29, 42, 27, 43, 32, 33, 40, 44, 40, 51, 54, 
    53, 56, 39, 69, 61, 59, 52, 60, 67, 58, 61, 56, 76, 55, 55, 
    50, 56, 53, 38, 40, 40, 42, 48, 43, 38, 41, 54, 52, 51, 53, 
    46, 49, 38, 46, 52, 53, 57, 56, 53, 51, 52, 55, 51, 51, 55, 
    47, 35, 31, 45, 42, 47, 58, 58, 56, 53, 54, 52, 51, 51, 53, 
    51, 52, 42, 13, 30, 48, 41, 48, 53, 50, 52, 52, 53, 52, 56, 
    50, 50, 48, 41, 0, 16, 24, 34, 30, 35, 50, 55, 53, 51, 55, 
    48, 49, 50, 43, 0, 8, 12, 12, 11, 12, 32, 25, 26, 36, 52, 
    51, 51, 50, 25, 45, 20, 38, 69, 37, 33, 38, 35, 71, 57, 59, 
    27, 26, 19, 18, 17, 10, 20, 32, 34, 35, 38, 39, 42, 48, 46, 
    23, 32, 29, 21, 19, 17, 23, 29, 21, 22, 19, 22, 23, 19, 19, 
    3, 11, 9, 6, 0, 4, 7, 6, 3, 0, 2, 1, 0, 0, 21, 
    0, 4, 3, 3, 0, 9, 7, 6, 3, 5, 2, 0, 4, 24, 0, 
    
    -- channel=51
    29, 74, 100, 65, 50, 68, 71, 57, 63, 60, 65, 64, 49, 66, 72, 
    38, 69, 98, 112, 57, 65, 79, 56, 75, 73, 72, 45, 68, 80, 75, 
    39, 71, 103, 84, 84, 55, 67, 42, 64, 75, 66, 59, 53, 84, 76, 
    49, 68, 118, 66, 59, 60, 73, 56, 62, 85, 55, 66, 21, 78, 76, 
    70, 69, 85, 112, 71, 69, 64, 67, 78, 82, 63, 41, 81, 80, 80, 
    68, 96, 92, 71, 83, 78, 75, 84, 89, 82, 76, 73, 82, 80, 74, 
    58, 101, 99, 47, 35, 67, 78, 86, 87, 93, 83, 89, 85, 85, 80, 
    51, 83, 100, 132, 68, 7, 35, 77, 89, 90, 81, 84, 83, 85, 79, 
    51, 77, 86, 98, 205, 21, 4, 27, 57, 78, 62, 85, 86, 84, 80, 
    49, 77, 83, 126, 210, 22, 15, 24, 22, 40, 8, 56, 58, 65, 76, 
    43, 81, 80, 120, 67, 100, 0, 0, 57, 52, 19, 24, 0, 40, 61, 
    62, 105, 104, 101, 94, 122, 89, 60, 97, 96, 86, 92, 85, 88, 86, 
    41, 59, 66, 62, 57, 58, 56, 52, 78, 67, 70, 64, 68, 78, 63, 
    37, 34, 40, 25, 32, 26, 26, 24, 31, 28, 20, 23, 20, 10, 0, 
    34, 25, 24, 19, 22, 8, 22, 8, 19, 17, 23, 22, 0, 5, 59, 
    
    -- channel=52
    1, 7, 9, 1, 0, 4, 6, 5, 12, 6, 8, 2, 13, 24, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 49, 18, 36, 46, 52, 47, 40, 0, 0, 0, 
    6, 0, 0, 32, 6, 5, 18, 9, 1, 0, 0, 6, 15, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    8, 0, 0, 0, 48, 46, 44, 39, 43, 39, 34, 24, 0, 0, 3, 
    2, 8, 26, 0, 0, 0, 0, 2, 5, 5, 0, 0, 0, 0, 0, 
    1, 3, 33, 126, 20, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    1, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 126, 183, 103, 125, 163, 116, 163, 117, 109, 47, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 7, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    0, 0, 0, 0, 0, 12, 24, 20, 19, 24, 16, 4, 19, 78, 0, 
    
    -- channel=53
    0, 0, 0, 7, 0, 0, 7, 2, 5, 5, 7, 5, 0, 5, 0, 
    0, 0, 0, 72, 70, 51, 59, 55, 60, 54, 48, 32, 0, 0, 0, 
    0, 0, 0, 57, 57, 60, 74, 61, 50, 57, 49, 49, 0, 0, 0, 
    0, 0, 13, 90, 55, 45, 61, 63, 58, 73, 65, 55, 34, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 29, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 63, 18, 21, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 2, 27, 47, 19, 15, 21, 26, 30, 6, 4, 0, 0, 0, 
    0, 1, 0, 7, 12, 35, 12, 0, 15, 15, 6, 18, 0, 4, 0, 
    0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 21, 18, 18, 27, 22, 19, 19, 21, 21, 19, 18, 17, 8, 0, 
    32, 17, 17, 20, 21, 13, 21, 19, 22, 22, 24, 24, 0, 0, 2, 
    
    -- channel=54
    17, 0, 0, 2, 6, 0, 0, 3, 0, 0, 0, 0, 11, 5, 0, 
    15, 0, 0, 0, 63, 38, 21, 46, 30, 27, 27, 37, 6, 0, 0, 
    15, 0, 0, 20, 12, 45, 38, 51, 29, 28, 28, 34, 16, 0, 0, 
    8, 0, 0, 57, 43, 41, 24, 51, 43, 30, 49, 33, 64, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 21, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 41, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 61, 34, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 22, 35, 46, 28, 2, 7, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 20, 29, 21, 11, 5, 52, 33, 22, 5, 0, 
    14, 0, 0, 0, 0, 0, 15, 79, 0, 0, 6, 0, 72, 14, 12, 
    15, 0, 0, 0, 0, 0, 0, 18, 0, 0, 1, 0, 0, 3, 7, 
    6, 7, 2, 1, 2, 0, 7, 14, 0, 4, 1, 7, 5, 0, 4, 
    0, 12, 8, 11, 3, 8, 13, 12, 5, 3, 10, 9, 8, 8, 23, 
    0, 8, 10, 13, 7, 16, 8, 15, 4, 7, 6, 3, 15, 14, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 11, 18, 18, 16, 15, 10, 10, 7, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 15, 3, 0, 3, 29, 31, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 
    20, 24, 20, 15, 15, 16, 12, 11, 5, 5, 4, 0, 1, 0, 0, 
    6, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 36, 66, 61, 56, 63, 64, 63, 51, 10, 6, 3, 
    0, 0, 5, 58, 26, 18, 26, 29, 19, 16, 17, 19, 26, 4, 4, 
    0, 0, 1, 0, 6, 1, 1, 0, 0, 4, 1, 0, 0, 4, 5, 
    0, 0, 0, 5, 0, 3, 0, 0, 11, 6, 0, 1, 0, 0, 0, 
    0, 19, 48, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 97, 23, 0, 0, 0, 0, 4, 8, 7, 8, 8, 
    0, 0, 0, 0, 0, 69, 73, 10, 2, 6, 0, 1, 0, 0, 0, 
    0, 1, 0, 4, 3, 0, 9, 90, 117, 69, 19, 0, 0, 1, 1, 
    0, 5, 3, 26, 52, 19, 14, 5, 0, 12, 71, 130, 116, 55, 9, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    110, 122, 128, 131, 132, 139, 112, 82, 87, 81, 72, 74, 52, 58, 64, 
    12, 12, 16, 24, 25, 31, 34, 39, 52, 58, 60, 62, 67, 67, 63, 
    10, 11, 12, 4, 4, 3, 2, 0, 2, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    
    -- channel=57
    192, 213, 188, 167, 179, 192, 187, 184, 181, 185, 188, 186, 191, 203, 212, 
    197, 225, 224, 133, 138, 146, 142, 141, 145, 152, 150, 158, 210, 223, 219, 
    195, 222, 224, 116, 129, 115, 101, 108, 126, 131, 129, 132, 192, 226, 228, 
    190, 219, 205, 114, 144, 148, 142, 141, 151, 153, 149, 162, 158, 226, 227, 
    199, 216, 216, 192, 177, 178, 180, 181, 186, 184, 176, 204, 203, 220, 223, 
    214, 214, 207, 214, 195, 195, 197, 202, 198, 197, 198, 204, 223, 221, 222, 
    219, 197, 139, 152, 210, 221, 221, 225, 222, 218, 218, 221, 222, 224, 227, 
    225, 231, 215, 125, 73, 159, 218, 226, 223, 220, 217, 218, 219, 219, 222, 
    225, 233, 230, 222, 100, 60, 93, 169, 206, 212, 216, 216, 218, 220, 223, 
    225, 227, 231, 221, 117, 41, 53, 55, 62, 95, 139, 191, 211, 216, 218, 
    225, 222, 228, 209, 127, 44, 42, 83, 101, 67, 64, 53, 115, 163, 202, 
    206, 208, 207, 205, 204, 198, 163, 174, 203, 186, 185, 188, 184, 201, 200, 
    107, 107, 100, 93, 87, 88, 88, 101, 113, 112, 112, 116, 123, 123, 112, 
    70, 73, 72, 61, 55, 53, 51, 51, 51, 40, 39, 37, 34, 38, 64, 
    36, 35, 36, 33, 33, 35, 30, 32, 34, 30, 28, 29, 45, 80, 83, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 23, 24, 32, 19, 26, 20, 22, 3, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 6, 0, 0, 3, 1, 0, 0, 0, 0, 0, 
    0, 11, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 116, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 76, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 45, 7, 77, 97, 42, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 79, 30, 0, 0, 36, 112, 124, 95, 33, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    63, 82, 92, 95, 99, 60, 31, 43, 72, 26, 42, 13, 48, 59, 49, 
    0, 0, 0, 0, 0, 0, 0, 16, 30, 32, 40, 45, 47, 52, 57, 
    58, 50, 41, 28, 32, 30, 23, 18, 10, 12, 5, 3, 3, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 
    
    -- channel=59
    54, 43, 19, 23, 39, 29, 24, 28, 25, 28, 27, 25, 29, 22, 23, 
    59, 59, 26, 0, 7, 5, 0, 8, 0, 0, 2, 19, 31, 28, 29, 
    60, 57, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 30, 32, 
    54, 55, 11, 0, 6, 9, 0, 8, 13, 0, 9, 6, 38, 36, 38, 
    42, 55, 39, 18, 37, 39, 38, 35, 35, 26, 34, 44, 28, 34, 39, 
    36, 36, 42, 36, 25, 27, 28, 23, 22, 23, 24, 38, 36, 33, 38, 
    37, 16, 11, 62, 74, 46, 38, 34, 30, 27, 33, 31, 34, 35, 39, 
    43, 34, 0, 0, 18, 82, 63, 34, 28, 26, 30, 31, 33, 32, 41, 
    39, 29, 23, 2, 0, 29, 61, 70, 53, 38, 42, 30, 32, 34, 40, 
    35, 24, 24, 7, 0, 27, 23, 15, 30, 50, 91, 65, 53, 41, 37, 
    43, 25, 27, 0, 0, 0, 21, 38, 0, 0, 3, 3, 54, 32, 40, 
    50, 37, 37, 40, 46, 17, 29, 57, 45, 39, 44, 36, 49, 56, 53, 
    26, 26, 20, 18, 20, 18, 26, 42, 35, 43, 44, 51, 52, 47, 57, 
    22, 34, 30, 28, 17, 23, 24, 24, 17, 14, 18, 17, 17, 22, 37, 
    3, 17, 15, 15, 11, 16, 9, 12, 6, 7, 6, 7, 30, 32, 16, 
    
    -- channel=60
    52, 21, 0, 11, 24, 13, 8, 13, 12, 13, 13, 9, 23, 27, 21, 
    49, 28, 1, 0, 14, 0, 0, 6, 0, 0, 0, 4, 29, 12, 14, 
    47, 26, 5, 0, 0, 27, 0, 25, 15, 16, 23, 28, 33, 18, 17, 
    41, 24, 0, 0, 3, 2, 0, 6, 0, 0, 5, 5, 31, 15, 15, 
    30, 26, 11, 0, 11, 8, 8, 14, 7, 1, 16, 35, 14, 16, 13, 
    31, 14, 1, 21, 19, 21, 25, 17, 13, 19, 23, 29, 13, 13, 17, 
    37, 0, 0, 13, 31, 26, 15, 11, 10, 8, 15, 11, 13, 12, 12, 
    47, 16, 0, 0, 0, 60, 45, 18, 5, 3, 13, 11, 14, 10, 14, 
    52, 22, 13, 0, 0, 38, 46, 31, 25, 18, 20, 9, 9, 11, 12, 
    50, 19, 13, 2, 0, 12, 31, 28, 27, 1, 27, 21, 29, 25, 16, 
    49, 13, 15, 0, 0, 0, 30, 83, 33, 0, 45, 17, 98, 43, 24, 
    32, 0, 0, 0, 0, 0, 17, 38, 0, 0, 8, 0, 8, 0, 0, 
    20, 11, 11, 16, 24, 18, 23, 29, 5, 12, 8, 13, 10, 1, 4, 
    0, 6, 4, 12, 8, 11, 16, 20, 18, 17, 24, 24, 24, 28, 69, 
    2, 20, 21, 27, 20, 32, 24, 33, 22, 26, 24, 29, 45, 77, 17, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 81, 94, 72, 100, 84, 81, 101, 73, 59, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 0, 0, 0, 3, 3, 2, 7, 0, 0, 5, 36, 0, 
    
    -- channel=62
    7, 14, 16, 17, 14, 17, 20, 13, 19, 18, 20, 19, 17, 30, 28, 
    1, 5, 12, 48, 39, 40, 42, 38, 47, 45, 39, 26, 30, 26, 27, 
    0, 3, 22, 37, 53, 48, 56, 52, 51, 58, 55, 56, 31, 25, 25, 
    1, 2, 24, 42, 30, 25, 33, 38, 30, 36, 32, 34, 22, 18, 20, 
    10, 4, 7, 28, 10, 7, 4, 14, 13, 13, 15, 7, 29, 21, 18, 
    15, 16, 6, 7, 19, 16, 20, 24, 21, 19, 21, 22, 18, 20, 18, 
    20, 13, 13, 0, 0, 12, 19, 22, 22, 24, 21, 21, 21, 21, 20, 
    21, 20, 19, 37, 11, 0, 0, 25, 27, 22, 22, 21, 20, 19, 16, 
    24, 27, 30, 29, 29, 0, 0, 0, 0, 18, 15, 24, 22, 18, 17, 
    27, 31, 31, 46, 16, 0, 0, 0, 0, 0, 0, 0, 0, 13, 22, 
    26, 29, 28, 31, 0, 27, 0, 0, 25, 0, 0, 0, 0, 26, 16, 
    12, 16, 14, 11, 8, 0, 5, 12, 7, 0, 8, 1, 15, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 47, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 99, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 79, 12, 0, 1, 14, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 76, 16, 0, 23, 42, 15, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 3, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 3, 5, 5, 19, 15, 12, 12, 19, 26, 20, 22, 20, 15, 6, 
    29, 20, 18, 20, 22, 11, 23, 17, 27, 25, 30, 29, 9, 28, 62, 
    
    -- channel=64
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 7, 0, 21, 0, 0, 
    0, 0, 0, 0, 13, 0, 7, 0, 0, 0, 14, 0, 44, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    19, 0, 0, 0, 7, 0, 0, 50, 0, 21, 0, 0, 7, 0, 0, 
    0, 0, 4, 0, 0, 0, 36, 0, 0, 0, 0, 1, 0, 0, 31, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 8, 0, 4, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 2, 3, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 7, 7, 8, 17, 33, 0, 0, 0, 0, 18, 0, 43, 
    9, 9, 0, 0, 3, 0, 4, 16, 0, 0, 0, 23, 13, 13, 0, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 27, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 17, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 18, 0, 0, 1, 0, 0, 0, 
    0, 14, 0, 0, 1, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 4, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 8, 2, 0, 0, 0, 0, 6, 5, 6, 6, 10, 0, 0, 0, 
    0, 2, 7, 0, 0, 2, 5, 13, 0, 11, 19, 15, 2, 0, 0, 
    0, 1, 0, 0, 18, 0, 20, 8, 11, 11, 5, 13, 5, 0, 0, 
    2, 0, 0, 0, 0, 21, 10, 20, 20, 8, 9, 4, 0, 0, 5, 
    0, 1, 0, 0, 7, 0, 34, 15, 12, 12, 8, 4, 0, 0, 0, 
    8, 8, 0, 0, 0, 11, 13, 14, 16, 7, 15, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 1, 0, 6, 12, 15, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 12, 9, 1, 0, 3, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 20, 
    
    -- channel=67
    27, 21, 0, 8, 82, 0, 24, 0, 15, 0, 62, 0, 145, 0, 0, 
    16, 16, 27, 13, 78, 0, 8, 0, 29, 0, 63, 0, 124, 0, 43, 
    51, 12, 14, 30, 57, 0, 0, 34, 0, 61, 0, 0, 96, 12, 49, 
    51, 0, 47, 41, 0, 0, 44, 37, 0, 37, 0, 0, 70, 27, 132, 
    48, 0, 93, 45, 0, 6, 86, 0, 8, 0, 29, 0, 41, 37, 171, 
    71, 0, 32, 76, 0, 3, 43, 0, 26, 9, 31, 0, 65, 21, 169, 
    56, 0, 0, 51, 48, 16, 17, 14, 25, 20, 16, 4, 42, 6, 132, 
    43, 0, 0, 42, 32, 34, 0, 26, 31, 14, 24, 3, 80, 22, 115, 
    1, 4, 29, 23, 6, 72, 8, 32, 29, 23, 39, 23, 82, 50, 74, 
    33, 39, 45, 4, 22, 0, 34, 28, 37, 59, 31, 50, 82, 25, 0, 
    92, 0, 50, 0, 7, 30, 0, 52, 56, 64, 36, 41, 54, 3, 24, 
    0, 5, 65, 0, 47, 0, 7, 39, 44, 70, 28, 49, 55, 0, 23, 
    23, 0, 46, 40, 38, 0, 34, 89, 0, 42, 41, 60, 73, 0, 30, 
    69, 0, 0, 8, 53, 16, 11, 32, 0, 31, 33, 73, 103, 0, 0, 
    90, 25, 0, 0, 21, 35, 30, 8, 37, 34, 50, 37, 37, 0, 0, 
    
    -- channel=68
    28, 24, 57, 10, 0, 27, 13, 0, 0, 0, 0, 5, 5, 0, 18, 
    10, 49, 3, 10, 0, 0, 0, 20, 12, 21, 0, 17, 25, 88, 33, 
    0, 0, 0, 0, 0, 52, 82, 19, 0, 0, 0, 23, 31, 23, 21, 
    0, 57, 30, 1, 23, 76, 0, 0, 30, 7, 70, 40, 0, 14, 0, 
    7, 18, 37, 0, 43, 13, 0, 78, 42, 64, 17, 0, 0, 0, 0, 
    0, 0, 0, 66, 72, 0, 25, 59, 30, 0, 0, 55, 0, 0, 0, 
    37, 20, 0, 1, 0, 0, 35, 12, 0, 0, 16, 27, 0, 16, 0, 
    0, 2, 19, 0, 42, 0, 0, 16, 25, 58, 31, 0, 46, 0, 0, 
    29, 35, 0, 0, 0, 50, 17, 0, 23, 0, 0, 9, 0, 0, 10, 
    18, 0, 0, 0, 0, 0, 5, 37, 1, 10, 1, 0, 0, 22, 10, 
    0, 19, 13, 5, 21, 11, 2, 3, 14, 0, 0, 0, 17, 11, 61, 
    55, 149, 87, 38, 0, 0, 1, 0, 0, 1, 20, 6, 0, 17, 0, 
    0, 0, 19, 59, 20, 13, 0, 0, 0, 2, 0, 0, 9, 0, 0, 
    0, 0, 0, 1, 54, 33, 0, 25, 45, 0, 1, 0, 0, 24, 0, 
    0, 25, 0, 0, 0, 59, 51, 4, 0, 0, 0, 0, 62, 46, 79, 
    
    -- channel=69
    15, 12, 7, 0, 17, 0, 16, 0, 24, 8, 30, 0, 76, 2, 13, 
    2, 20, 7, 0, 21, 2, 3, 3, 13, 9, 25, 0, 56, 5, 17, 
    31, 7, 3, 3, 16, 0, 6, 25, 0, 37, 0, 0, 50, 10, 22, 
    11, 0, 34, 15, 1, 9, 39, 12, 10, 6, 12, 21, 31, 13, 48, 
    14, 0, 23, 38, 0, 17, 46, 2, 11, 21, 36, 7, 37, 10, 49, 
    27, 0, 0, 17, 24, 46, 51, 9, 35, 39, 43, 21, 47, 0, 60, 
    24, 0, 0, 21, 62, 70, 70, 70, 68, 63, 53, 60, 45, 6, 38, 
    17, 0, 9, 21, 49, 83, 62, 82, 67, 76, 83, 45, 76, 20, 42, 
    1, 11, 9, 2, 40, 56, 65, 64, 82, 81, 80, 71, 68, 27, 20, 
    18, 10, 27, 11, 15, 37, 50, 63, 71, 76, 69, 79, 67, 29, 0, 
    30, 9, 25, 0, 19, 23, 34, 64, 69, 78, 67, 76, 66, 5, 6, 
    0, 37, 58, 14, 12, 12, 48, 78, 61, 69, 67, 87, 81, 25, 0, 
    32, 9, 45, 60, 37, 11, 44, 92, 32, 59, 71, 80, 89, 9, 12, 
    38, 36, 5, 36, 61, 42, 44, 30, 38, 68, 66, 91, 70, 13, 0, 
    39, 21, 21, 15, 34, 47, 48, 44, 69, 55, 61, 38, 40, 2, 30, 
    
    -- channel=70
    0, 0, 0, 0, 0, 45, 0, 10, 0, 0, 0, 56, 0, 25, 0, 
    0, 0, 0, 0, 0, 28, 0, 27, 0, 0, 0, 72, 0, 29, 0, 
    0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 4, 62, 0, 0, 0, 
    0, 32, 0, 0, 8, 8, 0, 0, 43, 0, 15, 21, 0, 0, 0, 
    0, 43, 0, 0, 37, 0, 0, 42, 0, 0, 0, 5, 0, 0, 0, 
    0, 50, 0, 0, 9, 2, 1, 11, 0, 0, 0, 32, 0, 0, 0, 
    0, 24, 11, 0, 0, 14, 15, 13, 14, 22, 22, 21, 0, 0, 0, 
    0, 12, 0, 0, 5, 3, 39, 27, 9, 18, 18, 39, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 38, 20, 15, 22, 14, 21, 0, 0, 0, 
    0, 0, 0, 5, 0, 55, 13, 23, 23, 0, 20, 0, 0, 0, 17, 
    0, 23, 0, 1, 0, 0, 71, 2, 3, 5, 14, 10, 0, 0, 0, 
    6, 0, 0, 0, 0, 10, 28, 19, 9, 0, 20, 13, 0, 9, 0, 
    0, 28, 0, 0, 0, 15, 1, 0, 52, 12, 20, 0, 0, 15, 0, 
    0, 29, 36, 0, 0, 0, 0, 0, 37, 26, 19, 0, 0, 33, 0, 
    0, 0, 63, 28, 0, 0, 0, 0, 0, 19, 14, 0, 0, 0, 54, 
    
    -- channel=71
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 13, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 10, 0, 16, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 20, 
    12, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 16, 11, 0, 0, 1, 21, 1, 0, 10, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 22, 0, 0, 15, 
    0, 0, 11, 4, 24, 0, 6, 14, 0, 0, 18, 0, 56, 45, 0, 
    0, 14, 0, 0, 0, 59, 0, 0, 9, 3, 0, 9, 5, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 2, 24, 5, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 13, 9, 0, 16, 17, 5, 0, 
    32, 57, 0, 0, 0, 8, 21, 74, 54, 3, 21, 0, 20, 4, 0, 
    0, 32, 38, 0, 0, 0, 0, 0, 0, 18, 7, 25, 48, 0, 0, 
    15, 0, 3, 30, 3, 0, 0, 0, 12, 51, 79, 20, 0, 0, 0, 
    
    -- channel=73
    58, 18, 35, 60, 36, 10, 48, 42, 71, 79, 80, 65, 78, 36, 48, 
    75, 42, 69, 67, 26, 9, 47, 36, 78, 62, 75, 69, 98, 45, 77, 
    82, 70, 73, 58, 17, 9, 46, 62, 76, 50, 75, 82, 133, 95, 112, 
    55, 60, 69, 44, 8, 58, 91, 40, 47, 52, 59, 101, 165, 121, 114, 
    55, 108, 111, 48, 49, 94, 55, 24, 78, 84, 107, 109, 141, 136, 95, 
    49, 105, 152, 71, 65, 87, 62, 79, 87, 90, 83, 78, 134, 143, 79, 
    52, 82, 126, 143, 85, 71, 62, 70, 81, 81, 78, 77, 112, 124, 93, 
    74, 96, 108, 147, 106, 45, 83, 95, 82, 71, 76, 120, 92, 117, 71, 
    86, 95, 114, 125, 131, 101, 82, 103, 92, 110, 107, 96, 125, 93, 66, 
    110, 103, 85, 99, 109, 132, 106, 113, 121, 117, 99, 103, 81, 62, 84, 
    98, 81, 74, 93, 87, 90, 128, 136, 130, 122, 102, 98, 77, 85, 112, 
    104, 100, 87, 92, 118, 107, 120, 134, 134, 110, 103, 95, 81, 89, 133, 
    125, 182, 156, 114, 105, 126, 130, 109, 125, 118, 119, 92, 71, 60, 124, 
    72, 55, 155, 167, 118, 107, 119, 102, 75, 117, 117, 94, 59, 59, 103, 
    79, 20, 43, 159, 179, 131, 118, 121, 104, 112, 111, 96, 52, 58, 104, 
    
    -- channel=74
    0, 0, 0, 0, 29, 0, 0, 0, 20, 6, 18, 0, 41, 0, 0, 
    0, 0, 2, 0, 28, 6, 3, 0, 0, 0, 6, 0, 0, 0, 0, 
    56, 0, 0, 23, 18, 0, 0, 24, 0, 69, 0, 0, 0, 0, 0, 
    3, 0, 16, 0, 0, 0, 36, 40, 0, 0, 0, 0, 0, 0, 60, 
    10, 0, 0, 36, 0, 0, 30, 0, 0, 0, 6, 2, 0, 0, 66, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 21, 0, 39, 
    0, 0, 0, 0, 7, 0, 0, 3, 3, 0, 0, 0, 1, 0, 12, 
    8, 0, 0, 0, 0, 53, 0, 0, 0, 0, 4, 0, 0, 0, 79, 
    0, 0, 32, 6, 34, 0, 0, 0, 0, 1, 0, 9, 35, 44, 0, 
    9, 35, 33, 0, 0, 40, 0, 0, 0, 0, 0, 2, 7, 0, 0, 
    51, 0, 0, 0, 12, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 0, 0, 
    77, 1, 0, 0, 0, 0, 7, 87, 8, 0, 0, 0, 17, 23, 24, 
    24, 109, 0, 0, 0, 0, 0, 0, 0, 5, 0, 35, 69, 0, 0, 
    26, 0, 56, 0, 0, 0, 0, 0, 36, 19, 53, 0, 0, 0, 0, 
    
    -- channel=75
    3, 0, 25, 27, 0, 46, 6, 24, 10, 17, 0, 52, 0, 37, 14, 
    7, 1, 6, 24, 0, 41, 18, 37, 0, 19, 0, 66, 0, 30, 1, 
    15, 18, 17, 17, 0, 32, 20, 9, 29, 0, 18, 60, 0, 12, 0, 
    0, 43, 0, 2, 14, 28, 0, 0, 53, 0, 25, 44, 0, 6, 0, 
    0, 61, 0, 0, 33, 0, 0, 32, 0, 14, 0, 16, 0, 13, 0, 
    0, 68, 9, 0, 24, 0, 0, 4, 0, 0, 0, 29, 0, 23, 0, 
    0, 45, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 40, 30, 6, 0, 0, 0, 0, 0, 0, 0, 5, 0, 13, 0, 
    12, 17, 18, 14, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 8, 10, 32, 15, 28, 0, 0, 0, 0, 0, 0, 0, 11, 24, 
    0, 31, 0, 26, 15, 3, 31, 0, 0, 0, 0, 0, 0, 10, 24, 
    0, 0, 0, 34, 1, 18, 8, 0, 0, 0, 0, 0, 0, 21, 15, 
    31, 35, 0, 0, 0, 33, 0, 0, 22, 0, 0, 0, 0, 26, 16, 
    0, 49, 46, 0, 0, 0, 5, 0, 23, 0, 0, 0, 0, 43, 13, 
    0, 0, 57, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 49, 
    
    -- channel=76
    38, 10, 74, 49, 0, 98, 43, 57, 58, 48, 11, 106, 0, 69, 39, 
    32, 28, 30, 48, 0, 77, 29, 76, 39, 65, 10, 132, 0, 96, 39, 
    29, 34, 34, 21, 0, 88, 82, 47, 50, 0, 71, 123, 5, 53, 44, 
    0, 112, 24, 15, 25, 117, 45, 0, 112, 0, 107, 118, 20, 46, 0, 
    8, 136, 0, 10, 100, 56, 0, 96, 66, 94, 68, 63, 37, 41, 0, 
    0, 131, 45, 0, 103, 44, 3, 90, 45, 41, 12, 115, 20, 50, 0, 
    0, 99, 66, 32, 14, 38, 24, 41, 21, 36, 30, 51, 5, 71, 0, 
    8, 79, 65, 45, 38, 0, 53, 34, 25, 35, 34, 46, 5, 47, 0, 
    47, 68, 27, 36, 59, 11, 45, 20, 37, 26, 9, 44, 0, 10, 0, 
    52, 14, 12, 74, 40, 47, 34, 45, 19, 23, 17, 16, 0, 29, 67, 
    0, 79, 13, 70, 63, 38, 93, 28, 18, 2, 24, 13, 7, 32, 81, 
    48, 98, 14, 81, 17, 66, 73, 31, 15, 0, 47, 18, 3, 63, 40, 
    63, 78, 31, 41, 38, 79, 49, 0, 42, 19, 27, 0, 1, 39, 56, 
    12, 72, 111, 54, 32, 59, 62, 18, 84, 41, 30, 0, 0, 99, 58, 
    0, 41, 120, 122, 51, 43, 50, 58, 25, 42, 27, 0, 2, 54, 158, 
    
    -- channel=77
    8, 21, 23, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    2, 15, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 52, 0, 
    0, 0, 0, 0, 0, 42, 49, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 41, 0, 0, 24, 27, 0, 0, 1, 2, 31, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 53, 19, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 24, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 66, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 42, 15, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 26, 
    0, 0, 1, 0, 0, 0, 4, 0, 0, 0, 5, 0, 13, 0, 14, 
    0, 0, 0, 0, 0, 2, 0, 9, 7, 7, 3, 0, 23, 0, 13, 
    0, 0, 0, 2, 19, 23, 12, 26, 11, 16, 13, 23, 5, 0, 0, 
    0, 0, 0, 0, 23, 15, 18, 26, 32, 30, 30, 12, 42, 0, 0, 
    0, 0, 0, 0, 12, 24, 25, 28, 42, 31, 22, 35, 26, 3, 0, 
    0, 0, 0, 0, 0, 0, 31, 33, 33, 50, 22, 35, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 48, 37, 35, 29, 28, 19, 0, 0, 
    0, 28, 14, 0, 0, 0, 29, 42, 34, 29, 40, 36, 27, 0, 0, 
    0, 0, 20, 15, 0, 0, 26, 43, 0, 28, 39, 35, 28, 0, 0, 
    0, 0, 0, 8, 26, 0, 0, 0, 0, 35, 26, 37, 12, 0, 0, 
    0, 0, 0, 0, 13, 28, 9, 7, 0, 19, 22, 0, 0, 0, 0, 
    
    -- channel=79
    43, 52, 44, 44, 84, 3, 55, 24, 58, 31, 70, 0, 122, 14, 29, 
    38, 54, 64, 41, 81, 26, 31, 19, 49, 44, 70, 0, 93, 25, 64, 
    52, 18, 36, 46, 64, 10, 49, 77, 17, 81, 7, 0, 70, 47, 52, 
    65, 3, 70, 44, 24, 46, 94, 64, 9, 37, 32, 27, 44, 38, 94, 
    69, 0, 72, 69, 0, 54, 99, 2, 64, 42, 71, 29, 52, 35, 115, 
    72, 0, 23, 79, 49, 23, 24, 18, 55, 46, 48, 7, 75, 21, 120, 
    63, 16, 11, 41, 42, 13, 14, 30, 15, 3, 0, 21, 43, 35, 95, 
    51, 13, 26, 30, 0, 55, 0, 6, 10, 17, 26, 0, 48, 29, 98, 
    24, 45, 42, 29, 10, 1, 6, 0, 14, 1, 9, 15, 21, 40, 59, 
    45, 40, 57, 17, 21, 0, 0, 0, 3, 15, 6, 22, 41, 37, 10, 
    76, 0, 68, 18, 54, 30, 0, 9, 2, 19, 0, 10, 35, 20, 49, 
    3, 41, 101, 51, 48, 20, 0, 0, 0, 19, 0, 17, 42, 18, 53, 
    32, 0, 47, 92, 77, 12, 20, 43, 0, 0, 7, 22, 46, 22, 67, 
    69, 37, 0, 26, 97, 80, 54, 42, 22, 0, 0, 37, 67, 15, 13, 
    85, 55, 24, 0, 26, 81, 92, 70, 53, 1, 10, 7, 59, 49, 15, 
    
    -- channel=80
    23, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 31, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 9, 0, 0, 0, 0, 5, 
    0, 0, 0, 53, 0, 7, 13, 0, 24, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 8, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 8, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 9, 3, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 8, 
    0, 4, 0, 0, 0, 0, 0, 7, 0, 5, 0, 0, 2, 0, 3, 
    21, 0, 11, 0, 0, 10, 0, 3, 0, 8, 0, 0, 4, 0, 7, 
    39, 6, 0, 0, 6, 9, 0, 0, 27, 19, 0, 0, 5, 3, 4, 
    2, 32, 0, 1, 14, 3, 6, 16, 11, 4, 0, 0, 2, 10, 0, 
    11, 28, 12, 0, 3, 8, 0, 0, 0, 0, 0, 0, 17, 22, 0, 
    1, 37, 12, 0, 15, 9, 0, 15, 0, 0, 2, 3, 12, 32, 0, 
    8, 25, 3, 0, 12, 1, 0, 17, 0, 0, 0, 0, 12, 33, 0, 
    3, 20, 3, 5, 0, 15, 18, 0, 0, 0, 0, 0, 7, 17, 0, 
    15, 14, 15, 2, 0, 0, 15, 4, 1, 1, 0, 3, 11, 0, 21, 
    10, 19, 2, 7, 0, 12, 22, 1, 11, 8, 7, 15, 6, 15, 0, 
    13, 26, 10, 19, 10, 15, 9, 3, 3, 11, 12, 12, 8, 0, 15, 
    
    -- channel=83
    44, 0, 16, 10, 18, 9, 17, 0, 51, 9, 11, 16, 1, 0, 43, 
    20, 38, 3, 9, 7, 10, 20, 2, 38, 18, 0, 13, 11, 31, 12, 
    58, 5, 6, 6, 7, 12, 21, 0, 12, 38, 0, 28, 18, 15, 15, 
    40, 10, 13, 0, 17, 11, 26, 17, 2, 14, 10, 47, 17, 0, 12, 
    15, 5, 14, 3, 11, 19, 24, 16, 40, 0, 11, 92, 1, 17, 14, 
    0, 19, 0, 19, 22, 0, 75, 54, 63, 0, 42, 69, 0, 11, 4, 
    0, 0, 43, 40, 0, 25, 47, 47, 0, 17, 79, 50, 0, 3, 14, 
    36, 0, 52, 19, 0, 49, 32, 21, 45, 47, 108, 65, 0, 0, 56, 
    39, 0, 41, 57, 24, 0, 92, 37, 39, 62, 107, 34, 0, 0, 121, 
    44, 0, 45, 167, 0, 17, 98, 0, 85, 30, 17, 32, 0, 0, 165, 
    55, 0, 55, 143, 0, 1, 22, 0, 81, 33, 20, 7, 0, 0, 144, 
    35, 16, 14, 52, 41, 5, 7, 57, 24, 9, 20, 0, 0, 0, 24, 
    13, 22, 22, 3, 66, 46, 4, 50, 36, 16, 17, 0, 0, 0, 0, 
    45, 0, 62, 3, 54, 7, 0, 55, 16, 30, 17, 1, 18, 3, 36, 
    15, 9, 35, 14, 24, 27, 28, 32, 27, 21, 10, 8, 27, 39, 0, 
    
    -- channel=84
    24, 95, 5, 25, 11, 12, 9, 11, 3, 0, 0, 14, 11, 20, 6, 
    17, 0, 8, 16, 20, 28, 25, 24, 28, 9, 0, 0, 8, 11, 3, 
    5, 0, 17, 6, 16, 10, 19, 8, 24, 73, 72, 34, 0, 0, 16, 
    0, 0, 0, 14, 3, 1, 0, 7, 0, 0, 17, 20, 0, 11, 1, 
    0, 12, 11, 4, 10, 15, 3, 46, 13, 0, 2, 0, 0, 0, 0, 
    0, 9, 32, 13, 0, 31, 42, 0, 0, 6, 0, 0, 0, 0, 0, 
    46, 0, 0, 4, 25, 16, 0, 64, 102, 58, 1, 0, 3, 6, 0, 
    9, 5, 0, 0, 27, 18, 37, 15, 1, 8, 39, 0, 0, 47, 22, 
    25, 30, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 22, 
    3, 18, 3, 0, 0, 0, 0, 60, 24, 0, 15, 42, 3, 21, 40, 
    16, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 
    0, 26, 0, 72, 45, 79, 69, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 11, 0, 39, 0, 15, 55, 58, 54, 47, 39, 21, 0, 0, 
    1, 0, 0, 0, 0, 15, 11, 12, 33, 50, 52, 79, 68, 59, 0, 
    3, 51, 7, 35, 37, 26, 5, 0, 0, 0, 22, 17, 23, 17, 32, 
    
    -- channel=85
    116, 120, 137, 139, 143, 147, 140, 116, 105, 74, 75, 81, 75, 82, 79, 
    128, 137, 138, 141, 150, 154, 161, 149, 138, 89, 69, 84, 86, 98, 83, 
    133, 117, 143, 149, 150, 160, 166, 157, 145, 110, 97, 108, 102, 94, 93, 
    100, 116, 141, 144, 154, 166, 165, 153, 144, 142, 135, 135, 96, 96, 96, 
    94, 119, 139, 146, 157, 157, 128, 125, 142, 136, 131, 127, 81, 91, 92, 
    41, 123, 137, 145, 147, 97, 102, 102, 94, 98, 120, 90, 67, 85, 89, 
    74, 90, 122, 123, 104, 118, 99, 84, 78, 86, 100, 70, 54, 81, 89, 
    102, 75, 119, 103, 91, 115, 134, 95, 84, 82, 110, 69, 36, 71, 100, 
    125, 77, 109, 118, 92, 91, 153, 113, 102, 106, 86, 51, 38, 66, 103, 
    130, 86, 86, 138, 34, 92, 119, 92, 137, 69, 54, 65, 47, 51, 99, 
    137, 94, 92, 100, 60, 69, 81, 110, 104, 65, 50, 47, 67, 57, 87, 
    120, 119, 80, 103, 101, 79, 92, 93, 57, 35, 26, 33, 44, 87, 63, 
    132, 118, 117, 88, 127, 109, 103, 110, 69, 45, 38, 26, 55, 60, 85, 
    131, 103, 126, 105, 104, 102, 113, 130, 96, 90, 80, 82, 86, 93, 79, 
    112, 126, 125, 118, 109, 127, 135, 121, 121, 115, 118, 118, 122, 119, 98, 
    
    -- channel=86
    4, 51, 42, 57, 41, 50, 44, 51, 3, 35, 43, 32, 44, 57, 19, 
    38, 20, 49, 46, 52, 51, 45, 59, 14, 23, 56, 52, 53, 32, 44, 
    3, 45, 46, 52, 51, 48, 40, 65, 49, 5, 57, 33, 53, 51, 45, 
    8, 39, 43, 57, 47, 53, 50, 47, 64, 51, 39, 16, 42, 61, 51, 
    35, 51, 43, 45, 51, 41, 41, 47, 29, 78, 55, 0, 54, 44, 47, 
    127, 24, 58, 42, 34, 61, 0, 28, 4, 61, 32, 0, 54, 43, 54, 
    107, 72, 21, 18, 52, 33, 8, 0, 44, 30, 0, 3, 44, 45, 44, 
    21, 113, 18, 35, 52, 17, 34, 38, 16, 8, 0, 0, 51, 52, 8, 
    45, 92, 28, 10, 35, 52, 7, 36, 34, 21, 0, 9, 80, 71, 0, 
    32, 107, 21, 0, 104, 49, 0, 73, 0, 14, 29, 25, 74, 96, 0, 
    37, 86, 11, 0, 45, 45, 44, 81, 8, 19, 29, 45, 61, 115, 0, 
    47, 61, 37, 12, 14, 51, 49, 0, 9, 24, 13, 38, 73, 76, 32, 
    68, 56, 43, 56, 13, 25, 68, 23, 11, 13, 11, 28, 51, 41, 62, 
    43, 87, 29, 52, 17, 53, 74, 32, 46, 35, 35, 48, 29, 50, 22, 
    60, 68, 50, 64, 42, 53, 52, 54, 47, 55, 65, 63, 47, 32, 64, 
    
    -- channel=87
    35, 1, 54, 47, 56, 60, 67, 54, 48, 42, 44, 41, 38, 33, 40, 
    20, 34, 50, 47, 54, 51, 63, 65, 72, 44, 44, 48, 44, 47, 45, 
    26, 25, 39, 50, 46, 58, 62, 61, 62, 29, 24, 45, 54, 57, 43, 
    26, 22, 43, 44, 43, 67, 66, 64, 58, 61, 57, 54, 60, 49, 48, 
    35, 24, 33, 46, 44, 56, 38, 26, 42, 64, 50, 47, 42, 49, 48, 
    35, 34, 21, 34, 49, 13, 0, 20, 44, 35, 44, 59, 36, 47, 46, 
    0, 33, 15, 22, 14, 0, 30, 6, 0, 0, 30, 40, 25, 40, 46, 
    48, 18, 18, 25, 0, 0, 17, 4, 0, 0, 5, 30, 25, 17, 32, 
    56, 15, 3, 23, 6, 32, 27, 55, 48, 55, 81, 56, 20, 15, 23, 
    69, 26, 0, 37, 36, 12, 56, 19, 47, 62, 27, 29, 27, 9, 0, 
    54, 42, 13, 65, 28, 63, 72, 75, 88, 50, 43, 48, 29, 24, 11, 
    71, 42, 31, 0, 40, 26, 28, 63, 47, 37, 32, 30, 44, 43, 42, 
    54, 63, 33, 39, 14, 52, 53, 46, 27, 21, 19, 15, 23, 49, 31, 
    59, 57, 54, 48, 53, 41, 48, 65, 42, 31, 32, 19, 24, 24, 50, 
    62, 39, 59, 45, 35, 45, 62, 67, 61, 62, 54, 52, 50, 52, 40, 
    
    -- channel=88
    0, 0, 24, 17, 15, 13, 23, 4, 18, 19, 10, 0, 0, 4, 18, 
    17, 25, 11, 6, 13, 10, 16, 10, 2, 1, 11, 31, 20, 13, 12, 
    23, 8, 7, 19, 13, 16, 11, 21, 21, 0, 0, 8, 23, 30, 11, 
    18, 15, 18, 17, 23, 29, 38, 30, 36, 25, 0, 9, 15, 1, 15, 
    34, 7, 13, 5, 17, 30, 16, 0, 11, 37, 31, 43, 21, 30, 19, 
    4, 0, 0, 18, 28, 0, 1, 79, 55, 13, 26, 38, 21, 19, 16, 
    0, 35, 23, 13, 0, 7, 33, 0, 0, 0, 16, 12, 0, 2, 20, 
    3, 7, 27, 32, 0, 16, 9, 16, 18, 7, 9, 31, 7, 0, 10, 
    25, 0, 12, 34, 24, 12, 48, 71, 73, 99, 103, 21, 0, 0, 11, 
    13, 0, 17, 37, 102, 45, 66, 12, 13, 27, 0, 0, 6, 0, 0, 
    28, 24, 35, 48, 0, 42, 54, 48, 98, 26, 32, 31, 0, 26, 33, 
    47, 7, 23, 0, 1, 0, 0, 17, 0, 4, 11, 6, 10, 33, 44, 
    20, 24, 0, 62, 35, 35, 3, 0, 0, 0, 0, 0, 0, 0, 3, 
    31, 35, 48, 9, 45, 0, 16, 23, 0, 0, 0, 0, 0, 0, 33, 
    10, 0, 24, 13, 0, 10, 33, 49, 25, 21, 14, 16, 14, 15, 3, 
    
    -- channel=89
    26, 3, 21, 18, 17, 6, 2, 0, 11, 3, 5, 0, 0, 7, 10, 
    56, 53, 20, 25, 23, 16, 0, 0, 0, 0, 6, 10, 11, 8, 8, 
    60, 59, 30, 34, 36, 25, 15, 8, 13, 0, 0, 0, 4, 13, 8, 
    62, 54, 43, 39, 44, 26, 29, 13, 26, 27, 8, 8, 4, 2, 14, 
    51, 54, 45, 38, 44, 39, 51, 41, 21, 30, 31, 31, 12, 14, 17, 
    40, 45, 58, 56, 44, 79, 81, 86, 55, 38, 35, 22, 9, 5, 14, 
    7, 77, 87, 73, 57, 90, 88, 56, 49, 59, 42, 7, 0, 2, 10, 
    7, 53, 88, 76, 95, 105, 56, 101, 110, 105, 60, 13, 7, 24, 3, 
    18, 48, 95, 55, 115, 96, 79, 78, 90, 85, 65, 0, 0, 52, 29, 
    19, 54, 120, 47, 95, 83, 72, 47, 8, 3, 0, 0, 0, 65, 63, 
    32, 47, 107, 46, 0, 36, 38, 38, 43, 0, 7, 9, 0, 62, 100, 
    37, 29, 74, 38, 0, 0, 0, 0, 0, 0, 0, 0, 7, 17, 85, 
    21, 41, 34, 82, 39, 23, 20, 0, 0, 0, 0, 0, 0, 0, 28, 
    31, 40, 43, 17, 48, 17, 29, 17, 9, 0, 0, 0, 0, 0, 21, 
    30, 21, 30, 19, 22, 26, 22, 31, 15, 12, 9, 21, 18, 12, 7, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 32, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 4, 53, 2, 0, 28, 44, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 24, 13, 0, 0, 4, 
    4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 23, 0, 0, 27, 
    0, 0, 0, 47, 3, 0, 48, 57, 33, 90, 94, 18, 0, 0, 29, 
    0, 0, 0, 87, 0, 15, 28, 0, 47, 24, 0, 0, 0, 0, 13, 
    1, 0, 23, 38, 20, 89, 33, 63, 53, 33, 33, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 28, 33, 12, 10, 31, 0, 48, 0, 
    0, 0, 18, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    16, 0, 10, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 3, 0, 
    0, 12, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 13, 16, 0, 
    0, 0, 0, 0, 27, 25, 0, 4, 0, 0, 8, 0, 0, 33, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 25, 15, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    0, 72, 21, 34, 20, 26, 11, 30, 0, 21, 22, 16, 22, 42, 0, 
    31, 17, 20, 29, 29, 27, 16, 28, 0, 5, 37, 19, 32, 13, 13, 
    0, 44, 32, 28, 30, 21, 13, 32, 14, 0, 52, 10, 25, 15, 23, 
    0, 41, 26, 38, 28, 21, 10, 17, 30, 16, 10, 0, 11, 32, 22, 
    14, 43, 32, 31, 31, 24, 12, 29, 4, 38, 23, 0, 38, 22, 23, 
    89, 12, 47, 27, 12, 56, 7, 16, 0, 46, 5, 0, 42, 24, 32, 
    134, 50, 19, 16, 35, 49, 0, 0, 60, 46, 0, 0, 36, 33, 25, 
    6, 104, 9, 17, 65, 9, 20, 44, 22, 16, 0, 0, 39, 54, 0, 
    3, 92, 17, 0, 71, 23, 0, 20, 20, 0, 0, 0, 73, 78, 0, 
    0, 90, 24, 0, 82, 52, 0, 66, 0, 0, 5, 21, 67, 105, 0, 
    0, 56, 16, 0, 62, 14, 0, 49, 0, 0, 18, 20, 53, 103, 0, 
    0, 37, 19, 0, 0, 27, 42, 0, 0, 11, 14, 43, 49, 51, 17, 
    25, 9, 24, 27, 0, 12, 23, 0, 1, 15, 14, 39, 60, 14, 60, 
    8, 33, 0, 28, 0, 29, 43, 0, 12, 12, 17, 46, 22, 46, 3, 
    7, 46, 0, 25, 13, 24, 19, 3, 11, 5, 29, 28, 10, 2, 31, 
    
    -- channel=93
    0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 47, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 10, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 14, 44, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 25, 32, 31, 38, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 24, 37, 30, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    36, 40, 49, 52, 54, 53, 43, 34, 24, 1, 7, 10, 1, 13, 10, 
    46, 57, 46, 54, 58, 57, 61, 53, 42, 1, 1, 11, 23, 28, 9, 
    54, 43, 54, 56, 60, 63, 65, 51, 55, 34, 24, 30, 30, 20, 23, 
    31, 50, 54, 54, 65, 69, 67, 57, 53, 55, 46, 37, 18, 17, 23, 
    24, 41, 57, 60, 60, 67, 49, 52, 50, 46, 45, 46, 11, 20, 22, 
    0, 52, 49, 63, 56, 37, 57, 37, 36, 32, 42, 12, 0, 12, 19, 
    13, 29, 64, 57, 31, 66, 32, 33, 29, 40, 34, 0, 0, 10, 17, 
    37, 19, 58, 39, 45, 56, 65, 54, 48, 46, 46, 3, 0, 16, 22, 
    46, 33, 52, 43, 56, 27, 69, 51, 40, 36, 15, 0, 0, 21, 30, 
    53, 26, 46, 64, 0, 48, 46, 45, 68, 0, 0, 3, 0, 18, 51, 
    60, 35, 46, 27, 0, 0, 0, 33, 8, 0, 0, 0, 0, 14, 46, 
    43, 54, 24, 32, 33, 11, 30, 33, 0, 0, 0, 0, 0, 13, 18, 
    46, 50, 46, 20, 44, 50, 32, 33, 3, 0, 0, 0, 0, 0, 24, 
    54, 31, 52, 34, 24, 33, 43, 50, 23, 24, 15, 22, 20, 23, 20, 
    36, 54, 47, 46, 41, 56, 52, 42, 43, 30, 40, 43, 44, 41, 21, 
    
    -- channel=95
    37, 23, 13, 4, 13, 16, 12, 8, 35, 12, 2, 15, 4, 0, 17, 
    9, 24, 9, 10, 7, 11, 22, 5, 33, 37, 0, 0, 0, 12, 3, 
    43, 0, 12, 6, 7, 13, 18, 8, 10, 35, 2, 20, 2, 0, 2, 
    19, 13, 10, 0, 12, 4, 11, 13, 1, 0, 16, 40, 6, 0, 0, 
    5, 0, 8, 10, 5, 16, 7, 5, 34, 0, 0, 59, 0, 5, 0, 
    0, 19, 0, 17, 22, 0, 46, 17, 12, 0, 22, 44, 0, 7, 0, 
    0, 0, 17, 15, 0, 24, 2, 15, 6, 17, 45, 33, 7, 7, 7, 
    22, 0, 12, 4, 0, 12, 19, 0, 6, 5, 56, 41, 0, 0, 50, 
    3, 0, 5, 40, 0, 0, 37, 0, 0, 14, 37, 19, 0, 0, 72, 
    9, 0, 0, 98, 0, 0, 24, 0, 64, 18, 11, 28, 0, 0, 91, 
    10, 0, 6, 70, 16, 1, 0, 0, 18, 30, 16, 0, 0, 0, 53, 
    0, 0, 0, 22, 42, 0, 7, 40, 36, 23, 27, 19, 0, 0, 0, 
    0, 0, 11, 0, 37, 15, 0, 26, 30, 30, 36, 15, 13, 0, 3, 
    5, 0, 10, 0, 9, 0, 0, 7, 0, 14, 7, 5, 18, 12, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 4, 15, 0, 
    
    -- channel=96
    0, 11, 12, 19, 22, 16, 11, 17, 0, 27, 6, 3, 0, 0, 0, 
    19, 9, 8, 7, 4, 1, 0, 3, 0, 0, 4, 0, 4, 0, 0, 
    0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 30, 18, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 4, 0, 0, 0, 0, 64, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 28, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 2, 0, 0, 13, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 8, 37, 52, 31, 22, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 9, 7, 27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 4, 10, 11, 0, 0, 0, 20, 0, 0, 0, 0, 
    0, 32, 0, 2, 7, 1, 0, 0, 0, 59, 53, 58, 1, 7, 43, 
    0, 0, 2, 0, 0, 3, 5, 0, 0, 1, 0, 40, 14, 5, 0, 
    0, 3, 13, 0, 0, 0, 0, 0, 0, 3, 0, 0, 39, 14, 3, 
    0, 0, 26, 29, 63, 87, 88, 89, 46, 24, 17, 0, 44, 13, 7, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 25, 6, 7, 1, 0, 0, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 14, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 1, 9, 0, 
    0, 5, 4, 2, 4, 5, 11, 5, 2, 4, 0, 10, 5, 0, 0, 
    7, 8, 7, 6, 9, 10, 0, 7, 24, 33, 10, 10, 6, 0, 0, 
    9, 8, 5, 4, 9, 31, 44, 18, 5, 0, 21, 0, 5, 0, 2, 
    8, 8, 5, 5, 32, 0, 0, 0, 0, 57, 76, 0, 8, 1, 0, 
    8, 6, 18, 25, 3, 18, 0, 25, 72, 90, 53, 0, 0, 6, 33, 
    9, 12, 14, 13, 0, 1, 43, 72, 43, 44, 25, 0, 44, 68, 44, 
    12, 75, 0, 23, 0, 19, 57, 52, 50, 29, 19, 20, 51, 36, 23, 
    49, 12, 0, 6, 0, 23, 82, 47, 17, 0, 24, 55, 23, 19, 0, 
    20, 21, 21, 0, 11, 41, 71, 48, 0, 11, 7, 45, 33, 0, 0, 
    16, 19, 26, 1, 49, 52, 74, 48, 0, 25, 12, 17, 29, 0, 2, 
    15, 23, 10, 0, 11, 6, 2, 0, 0, 22, 0, 0, 0, 0, 0, 
    12, 6, 14, 15, 9, 10, 9, 6, 2, 24, 0, 0, 0, 0, 1, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 3, 3, 50, 0, 10, 
    0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 34, 38, 0, 9, 
    6, 14, 3, 6, 0, 0, 0, 0, 0, 0, 15, 60, 13, 0, 21, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 82, 0, 2, 7, 9, 
    0, 0, 0, 4, 0, 3, 3, 0, 0, 39, 63, 4, 25, 10, 3, 
    0, 1, 4, 4, 0, 0, 10, 69, 83, 97, 56, 164, 0, 47, 10, 
    0, 4, 15, 0, 0, 27, 73, 68, 32, 0, 0, 251, 36, 19, 21, 
    1, 7, 0, 26, 58, 6, 47, 0, 0, 0, 78, 253, 108, 0, 0, 
    7, 0, 29, 19, 92, 0, 0, 0, 87, 87, 150, 173, 0, 0, 30, 
    0, 0, 183, 9, 80, 0, 0, 52, 76, 152, 65, 122, 47, 76, 116, 
    0, 54, 164, 64, 36, 0, 0, 65, 194, 113, 0, 0, 127, 128, 146, 
    0, 16, 62, 100, 0, 0, 0, 81, 268, 13, 44, 0, 45, 180, 19, 
    0, 14, 34, 74, 0, 11, 0, 72, 245, 0, 78, 17, 0, 143, 0, 
    1, 15, 59, 65, 21, 56, 66, 78, 144, 0, 69, 65, 5, 34, 1, 
    14, 27, 13, 39, 15, 15, 20, 22, 22, 0, 65, 52, 7, 5, 0, 
    
    -- channel=100
    58, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 7, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 8, 12, 30, 0, 13, 14, 
    0, 0, 0, 0, 0, 2, 7, 11, 17, 17, 50, 0, 26, 39, 14, 
    0, 4, 7, 12, 13, 15, 29, 40, 38, 36, 0, 0, 1, 0, 0, 
    9, 10, 6, 9, 9, 32, 6, 14, 66, 128, 75, 41, 9, 3, 0, 
    10, 12, 10, 7, 12, 60, 130, 70, 0, 0, 100, 68, 0, 4, 0, 
    12, 9, 10, 4, 56, 0, 0, 0, 0, 0, 37, 79, 46, 0, 0, 
    5, 10, 34, 69, 0, 13, 3, 115, 243, 250, 17, 0, 0, 12, 97, 
    6, 24, 18, 0, 0, 0, 0, 107, 0, 0, 0, 0, 47, 168, 59, 
    21, 171, 48, 0, 0, 0, 6, 0, 0, 0, 0, 96, 134, 24, 0, 
    32, 0, 0, 0, 0, 46, 76, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 27, 36, 15, 12, 0, 9, 4, 0, 0, 0, 0, 
    1, 0, 0, 22, 95, 120, 77, 0, 0, 15, 51, 8, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 11, 18, 74, 35, 38, 31, 17, 10, 0, 0, 0, 7, 8, 12, 
    
    -- channel=101
    303, 316, 325, 331, 321, 295, 281, 268, 240, 187, 186, 156, 92, 62, 138, 
    308, 294, 288, 279, 258, 236, 228, 219, 202, 185, 157, 132, 45, 71, 156, 
    227, 223, 222, 216, 204, 196, 197, 193, 188, 178, 109, 41, 70, 121, 163, 
    179, 185, 187, 189, 192, 195, 191, 194, 188, 168, 71, 23, 126, 165, 169, 
    175, 189, 191, 191, 189, 185, 163, 161, 141, 140, 41, 49, 138, 162, 161, 
    186, 190, 191, 189, 167, 110, 79, 60, 46, 0, 0, 85, 25, 111, 147, 
    192, 192, 190, 162, 124, 56, 34, 28, 23, 0, 0, 51, 39, 31, 95, 
    190, 190, 133, 112, 49, 30, 11, 0, 0, 3, 0, 53, 23, 0, 17, 
    189, 144, 92, 6, 17, 0, 0, 0, 0, 0, 32, 69, 19, 7, 0, 
    152, 66, 52, 0, 19, 0, 0, 0, 0, 27, 0, 0, 0, 0, 34, 
    117, 8, 0, 9, 7, 0, 0, 0, 42, 0, 14, 0, 0, 10, 25, 
    107, 1, 0, 14, 0, 0, 0, 0, 42, 0, 9, 0, 0, 31, 17, 
    78, 0, 0, 0, 0, 0, 0, 0, 43, 0, 13, 15, 0, 17, 25, 
    76, 16, 0, 0, 0, 0, 0, 0, 0, 0, 2, 23, 1, 6, 10, 
    69, 24, 0, 2, 0, 0, 0, 0, 6, 0, 6, 7, 7, 6, 2, 
    
    -- channel=102
    130, 120, 136, 131, 119, 117, 121, 102, 110, 74, 81, 70, 21, 65, 68, 
    135, 120, 115, 122, 119, 109, 112, 98, 97, 90, 85, 47, 8, 75, 78, 
    101, 98, 110, 107, 106, 102, 101, 96, 93, 95, 59, 1, 40, 79, 66, 
    99, 105, 101, 99, 106, 103, 107, 96, 93, 80, 0, 58, 73, 73, 81, 
    101, 107, 106, 102, 111, 102, 83, 89, 87, 36, 0, 41, 66, 87, 83, 
    105, 106, 101, 100, 106, 99, 74, 33, 18, 0, 0, 0, 63, 40, 80, 
    107, 105, 95, 100, 95, 35, 0, 0, 14, 114, 54, 0, 2, 34, 61, 
    108, 99, 99, 62, 5, 47, 0, 18, 59, 68, 0, 0, 0, 31, 54, 
    104, 101, 34, 32, 0, 23, 91, 62, 0, 0, 0, 0, 60, 76, 24, 
    115, 124, 0, 31, 0, 49, 115, 6, 0, 0, 12, 0, 13, 0, 0, 
    149, 24, 0, 0, 0, 48, 114, 0, 0, 0, 33, 105, 0, 0, 0, 
    93, 21, 0, 0, 30, 51, 86, 0, 0, 18, 0, 93, 6, 0, 21, 
    80, 24, 6, 0, 59, 11, 47, 0, 0, 43, 0, 23, 47, 0, 38, 
    62, 41, 0, 0, 23, 8, 3, 0, 0, 44, 0, 0, 20, 2, 27, 
    53, 11, 6, 0, 8, 8, 7, 6, 7, 52, 0, 0, 16, 17, 26, 
    
    -- channel=103
    172, 191, 196, 205, 204, 191, 182, 177, 167, 139, 136, 122, 65, 50, 104, 
    196, 177, 186, 193, 184, 168, 161, 155, 143, 134, 114, 83, 50, 38, 114, 
    156, 170, 164, 162, 154, 144, 145, 136, 131, 130, 54, 24, 39, 64, 113, 
    137, 141, 139, 139, 140, 141, 129, 122, 116, 111, 57, 24, 85, 122, 130, 
    130, 143, 143, 143, 141, 121, 96, 104, 70, 24, 0, 0, 78, 115, 120, 
    142, 144, 141, 141, 134, 66, 0, 0, 0, 0, 0, 0, 31, 52, 109, 
    144, 143, 143, 134, 62, 49, 38, 49, 52, 0, 0, 0, 0, 37, 66, 
    143, 145, 104, 43, 18, 3, 5, 0, 0, 0, 0, 0, 10, 25, 0, 
    144, 130, 46, 15, 5, 17, 0, 0, 0, 0, 0, 31, 21, 0, 0, 
    149, 0, 0, 0, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    104, 17, 0, 0, 28, 0, 0, 0, 0, 45, 18, 0, 0, 0, 47, 
    118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 25, 
    89, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 33, 
    68, 22, 0, 10, 8, 32, 34, 39, 46, 0, 12, 17, 33, 34, 23, 
    53, 30, 0, 0, 0, 0, 0, 2, 11, 11, 12, 28, 18, 16, 10, 
    
    -- channel=104
    38, 63, 76, 85, 89, 81, 76, 74, 64, 66, 43, 48, 47, 27, 26, 
    76, 69, 79, 83, 79, 70, 63, 59, 50, 41, 20, 26, 10, 0, 28, 
    87, 83, 71, 65, 52, 44, 43, 36, 35, 31, 44, 37, 0, 1, 37, 
    43, 42, 41, 40, 38, 40, 28, 18, 21, 30, 41, 0, 16, 39, 43, 
    37, 43, 45, 46, 44, 48, 40, 19, 0, 0, 0, 0, 26, 38, 39, 
    42, 44, 43, 44, 32, 0, 10, 84, 138, 151, 0, 0, 46, 15, 35, 
    43, 45, 50, 37, 39, 58, 41, 36, 19, 0, 0, 0, 0, 50, 34, 
    46, 46, 30, 10, 6, 7, 0, 0, 0, 0, 0, 107, 14, 0, 0, 
    49, 22, 1, 33, 37, 3, 0, 0, 31, 19, 0, 6, 0, 0, 0, 
    29, 0, 0, 0, 20, 15, 0, 0, 3, 109, 140, 0, 0, 0, 34, 
    47, 134, 35, 0, 6, 0, 0, 0, 48, 49, 1, 83, 46, 55, 86, 
    41, 0, 0, 4, 0, 0, 0, 0, 48, 0, 0, 6, 15, 39, 1, 
    29, 3, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 44, 53, 7, 
    9, 31, 62, 71, 79, 126, 139, 144, 122, 0, 14, 5, 18, 16, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 16, 51, 14, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 73, 99, 134, 171, 157, 2, 28, 0, 0, 
    0, 0, 0, 0, 0, 54, 100, 65, 45, 64, 217, 120, 0, 34, 0, 
    0, 0, 0, 0, 44, 36, 48, 31, 47, 118, 232, 186, 22, 0, 31, 
    0, 0, 5, 73, 54, 32, 69, 191, 238, 258, 225, 81, 22, 34, 126, 
    0, 60, 62, 39, 12, 9, 83, 223, 230, 214, 241, 152, 121, 159, 145, 
    0, 152, 135, 28, 0, 10, 86, 214, 197, 95, 55, 206, 199, 165, 82, 
    0, 41, 119, 22, 0, 64, 152, 216, 147, 23, 18, 44, 168, 91, 0, 
    0, 46, 117, 34, 52, 103, 158, 215, 126, 46, 35, 0, 117, 50, 0, 
    0, 28, 84, 59, 86, 141, 157, 162, 114, 49, 67, 0, 14, 0, 0, 
    0, 3, 25, 8, 0, 4, 0, 0, 0, 22, 41, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 17, 22, 21, 15, 17, 23, 38, 12, 0, 57, 1, 0, 
    8, 5, 24, 22, 18, 14, 10, 7, 3, 0, 0, 39, 0, 0, 0, 
    38, 40, 13, 13, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 59, 31, 0, 93, 0, 0, 3, 
    0, 0, 0, 0, 0, 79, 96, 116, 45, 0, 0, 0, 49, 14, 9, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 110, 0, 0, 0, 
    0, 0, 61, 12, 57, 24, 0, 0, 16, 0, 45, 62, 0, 0, 0, 
    0, 0, 57, 5, 42, 0, 0, 0, 0, 129, 0, 0, 0, 0, 66, 
    0, 119, 2, 30, 6, 0, 0, 0, 122, 89, 117, 0, 41, 76, 122, 
    20, 0, 0, 37, 0, 0, 0, 0, 93, 0, 1, 43, 0, 97, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 37, 24, 64, 5, 
    0, 2, 57, 56, 105, 147, 157, 165, 72, 0, 25, 33, 63, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 32, 11, 0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
    0, 0, 0, 0, 0, 13, 28, 29, 35, 105, 70, 0, 11, 19, 0, 
    0, 0, 0, 0, 0, 17, 2, 18, 17, 59, 31, 0, 0, 27, 13, 
    0, 0, 0, 29, 1, 46, 70, 60, 28, 26, 2, 0, 14, 29, 20, 
    0, 13, 0, 48, 0, 53, 118, 55, 40, 22, 39, 0, 20, 24, 10, 
    4, 44, 0, 20, 13, 54, 120, 46, 6, 5, 85, 129, 22, 17, 0, 
    0, 40, 31, 0, 37, 75, 105, 34, 0, 36, 11, 105, 53, 0, 8, 
    0, 38, 49, 0, 66, 38, 83, 43, 0, 49, 0, 38, 82, 0, 21, 
    0, 32, 45, 37, 84, 81, 79, 73, 0, 70, 16, 6, 49, 18, 25, 
    0, 11, 28, 16, 29, 28, 26, 24, 19, 57, 23, 2, 20, 21, 26, 
    
    -- channel=108
    43, 19, 25, 11, 0, 2, 12, 0, 8, 0, 0, 5, 0, 20, 8, 
    6, 2, 0, 0, 0, 0, 7, 0, 5, 7, 20, 0, 0, 61, 7, 
    4, 0, 0, 0, 3, 4, 7, 9, 12, 15, 48, 0, 9, 52, 5, 
    4, 6, 6, 3, 10, 10, 14, 17, 18, 21, 0, 32, 25, 10, 0, 
    11, 6, 4, 3, 12, 23, 28, 14, 26, 4, 0, 43, 13, 4, 8, 
    9, 4, 4, 4, 18, 42, 76, 51, 44, 0, 60, 0, 37, 8, 5, 
    5, 2, 0, 11, 52, 14, 0, 0, 0, 96, 108, 0, 0, 28, 7, 
    3, 0, 22, 25, 0, 37, 0, 46, 95, 156, 31, 0, 0, 27, 81, 
    1, 14, 3, 9, 0, 31, 65, 149, 34, 6, 0, 0, 34, 81, 67, 
    12, 128, 0, 35, 0, 54, 134, 55, 16, 0, 11, 0, 57, 21, 0, 
    69, 14, 0, 7, 0, 71, 147, 32, 0, 0, 43, 97, 0, 0, 0, 
    26, 14, 37, 0, 40, 96, 124, 23, 0, 30, 0, 103, 32, 0, 2, 
    18, 30, 50, 0, 90, 58, 106, 9, 0, 57, 0, 28, 83, 0, 34, 
    22, 34, 30, 0, 48, 8, 0, 0, 0, 77, 0, 0, 33, 0, 34, 
    19, 3, 9, 18, 25, 28, 24, 18, 16, 61, 4, 0, 26, 28, 39, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 43, 43, 39, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 59, 0, 0, 0, 42, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 109, 209, 110, 0, 0, 0, 12, 81, 
    0, 0, 0, 0, 0, 0, 13, 15, 0, 0, 0, 0, 49, 104, 16, 
    0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 42, 0, 0, 
    0, 0, 0, 0, 0, 48, 31, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 4, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 17, 80, 78, 0, 0, 0, 17, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 29, 56, 37, 36, 30, 18, 15, 0, 0, 0, 15, 15, 19, 
    
    -- channel=110
    128, 132, 137, 137, 133, 116, 109, 100, 90, 60, 56, 40, 14, 0, 31, 
    123, 118, 118, 108, 97, 85, 82, 75, 67, 54, 45, 33, 0, 0, 44, 
    86, 80, 73, 73, 67, 65, 66, 63, 60, 55, 36, 0, 0, 28, 54, 
    51, 57, 61, 60, 63, 66, 66, 68, 64, 58, 12, 0, 24, 50, 46, 
    54, 61, 63, 63, 62, 65, 63, 56, 46, 56, 0, 0, 39, 43, 44, 
    60, 63, 63, 62, 51, 32, 36, 53, 56, 13, 13, 25, 0, 38, 37, 
    64, 64, 64, 46, 40, 25, 0, 0, 0, 0, 21, 36, 0, 0, 8, 
    63, 63, 33, 40, 12, 0, 0, 0, 0, 26, 32, 42, 0, 0, 0, 
    63, 40, 18, 0, 0, 0, 0, 29, 46, 27, 53, 0, 0, 0, 20, 
    36, 37, 28, 0, 0, 0, 0, 21, 10, 33, 0, 21, 26, 15, 23, 
    28, 17, 0, 0, 0, 0, 0, 10, 48, 0, 0, 0, 12, 9, 0, 
    26, 0, 0, 0, 0, 0, 0, 16, 34, 0, 0, 0, 0, 5, 0, 
    4, 0, 0, 0, 0, 0, 2, 3, 16, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 0, 41, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 25, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 22, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 47, 20, 11, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 11, 0, 0, 138, 0, 15, 0, 
    0, 0, 0, 0, 0, 5, 10, 23, 0, 0, 0, 96, 68, 0, 3, 
    0, 0, 0, 14, 31, 0, 25, 0, 0, 0, 0, 93, 29, 2, 0, 
    0, 0, 37, 0, 51, 2, 0, 0, 0, 0, 26, 63, 0, 0, 0, 
    0, 0, 120, 0, 50, 0, 0, 0, 0, 34, 0, 1, 16, 8, 31, 
    0, 0, 30, 40, 25, 0, 0, 0, 64, 19, 9, 0, 8, 25, 57, 
    0, 0, 0, 66, 3, 0, 0, 0, 120, 4, 32, 0, 0, 89, 3, 
    0, 0, 0, 44, 0, 0, 0, 0, 109, 0, 48, 30, 0, 60, 10, 
    0, 0, 13, 12, 0, 0, 0, 0, 11, 0, 18, 49, 20, 16, 18, 
    0, 19, 17, 44, 30, 28, 32, 30, 32, 3, 18, 33, 29, 28, 19, 
    
    -- channel=112
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 16, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 23, 28, 37, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 31, 33, 29, 20, 21, 17, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 7, 5, 4, 20, 32, 30, 28, 23, 0, 0, 0, 
    0, 0, 7, 0, 12, 0, 19, 34, 27, 27, 31, 33, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 31, 20, 21, 31, 24, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 10, 10, 19, 33, 28, 29, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 20, 27, 28, 34, 25, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 24, 19, 22, 22, 34, 25, 22, 0, 
    0, 0, 17, 43, 7, 44, 20, 16, 11, 17, 22, 41, 24, 4, 0, 
    0, 19, 0, 0, 12, 28, 16, 0, 23, 32, 9, 20, 17, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 24, 3, 7, 0, 19, 22, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 1, 0, 18, 28, 23, 5, 0, 
    0, 0, 10, 0, 0, 0, 0, 6, 0, 0, 0, 0, 14, 0, 0, 
    
    -- channel=113
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=114
    2, 0, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 8, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    21, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    21, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 20, 14, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 28, 33, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 51, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    31, 34, 17, 38, 21, 12, 30, 27, 31, 29, 28, 30, 23, 10, 16, 
    31, 37, 24, 14, 22, 0, 14, 9, 17, 17, 9, 8, 8, 13, 24, 
    29, 31, 47, 5, 5, 0, 0, 0, 0, 13, 23, 26, 29, 39, 37, 
    22, 16, 43, 0, 0, 0, 0, 0, 0, 0, 8, 29, 21, 32, 21, 
    0, 8, 102, 36, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 17, 
    33, 46, 123, 35, 0, 0, 2, 1, 0, 0, 0, 0, 0, 19, 32, 
    47, 50, 58, 96, 0, 0, 16, 0, 0, 0, 0, 0, 0, 13, 47, 
    29, 29, 59, 49, 83, 0, 13, 0, 0, 13, 0, 0, 0, 0, 17, 
    21, 8, 30, 62, 60, 82, 13, 8, 0, 4, 0, 0, 0, 4, 41, 
    27, 56, 101, 163, 31, 105, 0, 23, 0, 0, 0, 0, 0, 22, 13, 
    81, 123, 151, 51, 20, 29, 0, 0, 0, 0, 0, 0, 0, 5, 24, 
    125, 97, 81, 56, 45, 0, 0, 25, 0, 0, 0, 5, 3, 0, 44, 
    52, 41, 33, 28, 51, 24, 0, 22, 0, 0, 10, 12, 18, 0, 4, 
    20, 21, 37, 39, 10, 14, 0, 4, 0, 0, 0, 1, 12, 3, 0, 
    39, 30, 11, 11, 0, 2, 17, 15, 0, 0, 0, 0, 11, 0, 7, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 3, 13, 
    0, 0, 0, 0, 2, 0, 0, 3, 0, 3, 21, 42, 53, 54, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 24, 50, 33, 24, 5, 0, 0, 
    0, 3, 27, 27, 0, 5, 15, 8, 0, 0, 0, 0, 0, 7, 11, 
    78, 100, 79, 7, 5, 7, 39, 20, 4, 0, 0, 0, 6, 27, 33, 
    27, 3, 0, 18, 26, 37, 0, 0, 7, 8, 5, 0, 0, 2, 5, 
    0, 0, 0, 59, 0, 0, 0, 0, 13, 16, 5, 0, 0, 0, 0, 
    0, 17, 15, 0, 84, 72, 31, 15, 13, 11, 5, 4, 0, 0, 11, 
    20, 37, 94, 107, 49, 63, 21, 27, 0, 0, 15, 11, 0, 0, 0, 
    123, 88, 0, 0, 0, 0, 0, 5, 5, 0, 11, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 
    0, 0, 0, 0, 0, 0, 3, 13, 0, 0, 18, 11, 0, 0, 16, 
    0, 0, 0, 1, 19, 35, 0, 0, 19, 10, 29, 0, 8, 1, 0, 
    0, 5, 0, 0, 0, 4, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    8, 12, 10, 16, 27, 37, 37, 17, 16, 18, 15, 14, 13, 11, 14, 
    8, 12, 17, 17, 45, 53, 51, 51, 31, 19, 27, 27, 26, 26, 29, 
    10, 10, 30, 21, 51, 65, 76, 81, 50, 33, 37, 43, 42, 39, 41, 
    13, 12, 27, 45, 51, 66, 79, 94, 95, 59, 45, 58, 41, 41, 48, 
    11, 14, 55, 46, 57, 40, 63, 90, 98, 95, 82, 71, 57, 67, 71, 
    23, 27, 39, 50, 42, 46, 66, 75, 82, 97, 103, 78, 79, 81, 78, 
    22, 24, 21, 61, 56, 40, 67, 71, 68, 80, 93, 81, 86, 68, 60, 
    19, 25, 44, 29, 55, 48, 76, 79, 64, 69, 85, 89, 71, 57, 54, 
    24, 21, 27, 73, 51, 85, 58, 88, 61, 61, 76, 85, 65, 73, 82, 
    25, 33, 45, 55, 46, 72, 56, 87, 62, 58, 70, 83, 73, 83, 80, 
    26, 45, 68, 52, 62, 63, 72, 66, 68, 69, 75, 81, 82, 76, 90, 
    30, 21, 34, 32, 60, 59, 46, 64, 55, 59, 61, 76, 96, 79, 93, 
    26, 20, 23, 37, 41, 52, 56, 57, 47, 42, 52, 69, 96, 98, 79, 
    28, 38, 53, 64, 63, 64, 60, 73, 67, 62, 43, 59, 91, 96, 90, 
    53, 62, 71, 83, 79, 73, 81, 90, 91, 81, 72, 78, 88, 99, 95, 
    
    -- channel=118
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 5, 
    0, 0, 5, 5, 0, 2, 0, 0, 0, 3, 6, 10, 13, 15, 9, 
    0, 0, 0, 9, 0, 0, 0, 0, 10, 3, 5, 6, 8, 7, 6, 
    0, 0, 0, 15, 0, 0, 0, 6, 0, 8, 0, 0, 13, 6, 12, 
    16, 14, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 17, 19, 21, 
    6, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 26, 25, 18, 
    0, 0, 0, 0, 24, 16, 0, 0, 0, 0, 0, 5, 0, 24, 3, 
    1, 7, 0, 0, 0, 36, 0, 2, 0, 0, 0, 0, 0, 9, 16, 
    7, 15, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 5, 6, 
    20, 8, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 14, 23, 
    0, 0, 0, 0, 0, 0, 10, 0, 7, 0, 0, 0, 0, 44, 0, 
    0, 0, 0, 9, 0, 0, 7, 0, 0, 9, 0, 0, 0, 35, 32, 
    8, 12, 1, 1, 20, 19, 15, 4, 1, 6, 0, 0, 0, 28, 42, 
    3, 9, 22, 26, 52, 34, 14, 18, 30, 23, 26, 18, 9, 38, 39, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 3, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 51, 
    0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 16, 38, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 36, 34, 
    0, 0, 0, 29, 43, 19, 6, 3, 8, 0, 0, 0, 1, 46, 46, 
    10, 39, 46, 43, 44, 29, 17, 41, 47, 33, 26, 30, 40, 54, 59, 
    
    -- channel=120
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 7, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 
    13, 9, 0, 0, 3, 30, 6, 0, 0, 0, 0, 0, 2, 24, 28, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 39, 
    0, 0, 61, 53, 26, 33, 0, 0, 0, 0, 0, 0, 0, 2, 14, 
    3, 30, 27, 19, 24, 37, 6, 26, 0, 0, 0, 0, 0, 0, 2, 
    106, 67, 33, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    29, 19, 0, 0, 18, 0, 11, 0, 0, 0, 0, 0, 0, 3, 18, 
    0, 0, 23, 37, 19, 1, 0, 2, 2, 8, 25, 0, 5, 19, 17, 
    32, 34, 15, 10, 10, 11, 3, 14, 7, 1, 3, 20, 18, 17, 21, 
    
    -- channel=121
    74, 68, 70, 73, 64, 66, 60, 59, 47, 42, 36, 25, 15, 8, 2, 
    72, 66, 64, 48, 49, 53, 56, 42, 42, 34, 25, 19, 17, 18, 20, 
    67, 66, 51, 31, 33, 22, 23, 28, 40, 51, 53, 52, 49, 49, 37, 
    57, 58, 34, 0, 18, 17, 12, 17, 25, 66, 67, 59, 50, 36, 22, 
    69, 85, 89, 6, 13, 44, 45, 22, 22, 23, 42, 58, 51, 32, 25, 
    129, 143, 136, 11, 19, 39, 60, 45, 34, 17, 17, 43, 53, 48, 44, 
    143, 139, 134, 34, 28, 56, 56, 40, 50, 36, 24, 28, 52, 60, 52, 
    126, 128, 129, 115, 39, 14, 32, 31, 65, 59, 29, 22, 49, 43, 35, 
    131, 145, 155, 101, 135, 80, 72, 29, 67, 68, 41, 29, 41, 42, 23, 
    179, 206, 224, 198, 147, 133, 73, 47, 60, 68, 54, 35, 35, 22, 0, 
    257, 251, 148, 137, 98, 91, 66, 52, 55, 64, 51, 36, 26, 20, 0, 
    232, 203, 130, 86, 34, 25, 51, 12, 35, 51, 55, 45, 17, 23, 6, 
    117, 101, 92, 77, 59, 16, 35, 46, 27, 56, 79, 63, 30, 4, 26, 
    69, 62, 61, 47, 28, 30, 7, 25, 12, 34, 75, 55, 38, 2, 1, 
    46, 30, 12, 0, 0, 19, 16, 2, 0, 0, 0, 13, 3, 0, 0, 
    
    -- channel=122
    0, 2, 0, 7, 3, 0, 5, 0, 0, 1, 4, 4, 0, 0, 0, 
    0, 0, 0, 9, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 34, 0, 4, 0, 9, 0, 0, 0, 0, 0, 0, 7, 12, 
    0, 0, 0, 13, 0, 0, 0, 0, 12, 1, 0, 6, 0, 0, 0, 
    0, 0, 0, 9, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 17, 0, 0, 0, 4, 0, 0, 0, 0, 
    10, 7, 0, 0, 25, 11, 2, 0, 0, 0, 1, 0, 5, 8, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 11, 37, 
    0, 0, 45, 4, 24, 3, 0, 2, 0, 0, 0, 0, 5, 19, 0, 
    0, 27, 123, 70, 46, 44, 26, 18, 0, 2, 9, 0, 0, 0, 2, 
    115, 94, 2, 0, 37, 15, 0, 26, 10, 0, 0, 0, 10, 0, 0, 
    31, 25, 5, 0, 0, 0, 11, 0, 0, 0, 0, 2, 0, 7, 0, 
    0, 0, 22, 42, 17, 0, 0, 8, 9, 35, 21, 3, 16, 7, 10, 
    30, 37, 9, 0, 0, 0, 1, 4, 1, 0, 13, 20, 7, 3, 7, 
    
    -- channel=123
    16, 13, 22, 14, 6, 0, 3, 13, 9, 9, 12, 11, 13, 17, 10, 
    16, 11, 18, 10, 0, 0, 0, 0, 9, 7, 3, 1, 0, 0, 0, 
    18, 14, 4, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 15, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 8, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 10, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 9, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 16, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    28, 24, 37, 23, 40, 39, 26, 25, 22, 26, 20, 16, 20, 27, 19, 
    27, 23, 38, 19, 45, 61, 43, 41, 23, 27, 28, 32, 36, 38, 28, 
    28, 26, 15, 43, 42, 61, 64, 63, 58, 51, 38, 35, 24, 18, 11, 
    30, 33, 3, 43, 58, 66, 68, 71, 64, 54, 50, 22, 21, 17, 22, 
    54, 62, 21, 0, 63, 88, 71, 50, 67, 68, 72, 50, 39, 25, 30, 
    46, 33, 0, 0, 51, 100, 51, 49, 68, 61, 66, 70, 53, 27, 17, 
    25, 18, 8, 0, 52, 71, 42, 63, 72, 53, 55, 81, 51, 35, 2, 
    36, 38, 30, 4, 0, 69, 43, 71, 77, 48, 52, 69, 59, 36, 21, 
    46, 48, 35, 22, 40, 19, 51, 42, 73, 51, 57, 58, 72, 42, 5, 
    67, 62, 14, 0, 38, 0, 60, 25, 73, 63, 61, 50, 63, 11, 13, 
    24, 1, 0, 3, 42, 24, 55, 36, 68, 62, 48, 46, 49, 34, 10, 
    0, 0, 0, 12, 10, 53, 71, 21, 63, 65, 65, 47, 26, 51, 1, 
    5, 18, 16, 29, 11, 39, 62, 29, 70, 88, 64, 48, 29, 40, 30, 
    24, 38, 29, 9, 12, 30, 36, 38, 45, 63, 50, 45, 35, 22, 38, 
    19, 8, 13, 17, 38, 41, 31, 14, 23, 33, 44, 34, 17, 28, 22, 
    
    -- channel=125
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 25, 35, 29, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 0, 0, 0, 0, 0, 
    0, 0, 10, 1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 52, 10, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 35, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 5, 0, 0, 0, 
    0, 0, 34, 0, 0, 0, 2, 2, 4, 1, 0, 1, 4, 8, 11, 
    16, 17, 24, 0, 0, 0, 0, 0, 1, 4, 7, 0, 6, 22, 18, 
    9, 9, 6, 9, 0, 0, 0, 0, 0, 0, 3, 0, 12, 10, 5, 
    2, 8, 23, 0, 24, 0, 11, 0, 1, 1, 0, 0, 0, 0, 0, 
    13, 16, 23, 34, 35, 41, 7, 11, 0, 0, 0, 0, 0, 3, 13, 
    38, 60, 54, 48, 20, 36, 2, 8, 0, 0, 0, 0, 0, 4, 0, 
    52, 59, 27, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 6, 10, 
    36, 9, 0, 6, 0, 0, 0, 0, 0, 0, 0, 7, 6, 7, 18, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 4, 0, 12, 13, 7, 
    0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 12, 
    2, 0, 0, 0, 0, 9, 8, 9, 6, 0, 0, 1, 6, 8, 11, 
    
    -- channel=127
    24, 28, 12, 20, 28, 33, 42, 24, 31, 31, 30, 32, 30, 22, 28, 
    25, 29, 21, 24, 47, 46, 49, 54, 34, 25, 29, 26, 26, 24, 28, 
    26, 25, 41, 19, 57, 65, 70, 62, 32, 28, 29, 28, 25, 24, 25, 
    26, 23, 38, 50, 65, 70, 68, 69, 66, 32, 30, 43, 14, 23, 23, 
    10, 13, 69, 64, 71, 37, 65, 88, 77, 74, 58, 49, 20, 18, 22, 
    7, 9, 54, 65, 52, 41, 77, 77, 70, 81, 84, 60, 24, 12, 21, 
    6, 6, 11, 74, 40, 29, 69, 68, 60, 77, 85, 65, 51, 14, 28, 
    6, 2, 23, 8, 74, 32, 68, 59, 60, 80, 87, 83, 57, 35, 19, 
    3, 0, 0, 65, 25, 64, 18, 81, 63, 73, 82, 92, 63, 50, 31, 
    0, 0, 14, 43, 29, 57, 31, 78, 67, 68, 75, 96, 75, 54, 13, 
    0, 9, 76, 35, 46, 55, 57, 46, 63, 67, 69, 83, 69, 25, 37, 
    15, 4, 11, 41, 83, 66, 35, 73, 46, 53, 56, 77, 63, 9, 38, 
    13, 15, 10, 15, 34, 56, 41, 54, 59, 44, 64, 75, 64, 29, 8, 
    15, 18, 32, 29, 10, 14, 40, 48, 52, 48, 38, 65, 69, 28, 16, 
    30, 22, 15, 23, 8, 13, 34, 31, 29, 32, 35, 34, 35, 21, 18, 
    
    -- channel=128
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=130
    0, 38, 9, 3, 7, 2, 0, 6, 0, 0, 35, 19, 10, 6, 3, 
    2, 23, 13, 16, 25, 18, 11, 11, 14, 0, 57, 15, 12, 12, 10, 
    2, 7, 23, 28, 47, 6, 10, 17, 0, 12, 37, 18, 17, 20, 15, 
    7, 39, 45, 1, 40, 23, 21, 10, 20, 46, 20, 41, 34, 12, 15, 
    1, 24, 13, 0, 48, 33, 21, 0, 21, 35, 27, 33, 23, 0, 11, 
    7, 14, 2, 4, 36, 29, 9, 14, 29, 40, 27, 35, 16, 0, 0, 
    2, 9, 0, 14, 20, 36, 20, 31, 22, 26, 35, 33, 21, 8, 0, 
    0, 10, 0, 42, 25, 22, 24, 32, 14, 28, 13, 16, 9, 9, 8, 
    0, 10, 24, 48, 27, 34, 36, 8, 33, 8, 15, 0, 27, 0, 15, 
    0, 13, 26, 20, 29, 31, 28, 22, 19, 29, 1, 10, 21, 12, 12, 
    5, 3, 26, 29, 28, 8, 33, 33, 13, 4, 7, 21, 18, 6, 12, 
    7, 0, 35, 31, 26, 12, 29, 26, 19, 0, 24, 14, 20, 11, 2, 
    1, 0, 19, 28, 9, 28, 27, 15, 5, 0, 15, 10, 13, 5, 9, 
    0, 0, 10, 28, 12, 39, 10, 6, 3, 0, 13, 10, 3, 17, 16, 
    0, 0, 8, 30, 18, 14, 0, 3, 0, 13, 8, 12, 5, 17, 8, 
    
    -- channel=131
    20, 0, 6, 37, 40, 14, 30, 16, 55, 88, 0, 25, 32, 29, 35, 
    17, 0, 0, 3, 47, 55, 32, 26, 58, 121, 0, 46, 46, 39, 44, 
    17, 0, 0, 1, 22, 134, 44, 23, 61, 11, 0, 28, 53, 49, 53, 
    53, 0, 0, 75, 2, 98, 75, 66, 23, 0, 60, 0, 73, 99, 29, 
    74, 1, 49, 93, 0, 60, 94, 106, 27, 0, 22, 9, 70, 104, 9, 
    53, 35, 62, 63, 20, 68, 101, 58, 39, 2, 22, 0, 68, 100, 31, 
    51, 34, 80, 30, 49, 24, 99, 16, 79, 27, 20, 2, 55, 79, 58, 
    65, 35, 113, 0, 84, 65, 72, 77, 31, 31, 69, 17, 20, 89, 37, 
    90, 20, 60, 10, 63, 62, 74, 120, 0, 51, 58, 52, 0, 56, 0, 
    73, 34, 50, 60, 43, 68, 70, 79, 75, 19, 80, 31, 14, 52, 10, 
    54, 79, 19, 54, 55, 101, 20, 50, 92, 95, 24, 22, 40, 64, 45, 
    50, 92, 0, 66, 86, 80, 38, 52, 77, 97, 0, 46, 40, 66, 54, 
    57, 69, 0, 63, 125, 16, 37, 57, 80, 68, 11, 41, 51, 39, 44, 
    63, 64, 0, 48, 103, 41, 70, 50, 64, 33, 18, 34, 57, 0, 33, 
    54, 48, 0, 28, 76, 87, 82, 39, 69, 0, 25, 31, 40, 22, 30, 
    
    -- channel=132
    0, 0, 0, 1, 4, 0, 13, 20, 44, 43, 0, 41, 31, 26, 20, 
    1, 0, 0, 0, 37, 19, 0, 9, 2, 7, 80, 26, 21, 16, 11, 
    3, 0, 0, 24, 10, 14, 0, 0, 0, 0, 58, 0, 5, 23, 31, 
    151, 125, 141, 0, 0, 18, 78, 33, 8, 10, 0, 14, 31, 1, 0, 
    52, 92, 18, 0, 6, 0, 1, 0, 0, 0, 0, 19, 11, 0, 0, 
    8, 5, 0, 10, 18, 0, 0, 0, 39, 23, 0, 0, 0, 14, 5, 
    0, 0, 0, 0, 0, 0, 7, 9, 24, 11, 7, 1, 0, 20, 34, 
    0, 0, 0, 8, 21, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 18, 36, 8, 58, 49, 8, 0, 0, 10, 18, 0, 0, 0, 
    8, 28, 6, 14, 0, 0, 0, 24, 76, 27, 0, 0, 34, 16, 0, 
    0, 2, 0, 14, 24, 0, 0, 0, 0, 0, 0, 22, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 6, 0, 0, 22, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 0, 
    
    -- channel=133
    6, 7, 85, 92, 83, 93, 103, 89, 78, 88, 7, 84, 110, 111, 116, 
    8, 13, 64, 63, 29, 69, 61, 65, 79, 71, 15, 73, 94, 102, 108, 
    12, 13, 24, 79, 14, 57, 56, 62, 62, 23, 38, 50, 63, 64, 70, 
    56, 1, 42, 85, 7, 32, 49, 56, 40, 21, 34, 29, 45, 60, 39, 
    58, 44, 55, 79, 20, 29, 49, 57, 32, 20, 24, 39, 54, 77, 58, 
    60, 53, 62, 69, 31, 34, 49, 38, 30, 20, 29, 33, 50, 76, 71, 
    70, 62, 91, 55, 49, 27, 52, 15, 33, 20, 26, 33, 49, 51, 62, 
    74, 62, 102, 32, 50, 32, 24, 54, 20, 44, 47, 53, 27, 65, 42, 
    76, 58, 63, 50, 26, 27, 40, 51, 45, 59, 57, 79, 61, 59, 38, 
    61, 55, 48, 48, 43, 41, 21, 26, 74, 56, 72, 67, 59, 73, 66, 
    52, 67, 27, 50, 47, 62, 36, 41, 46, 83, 49, 60, 60, 67, 70, 
    54, 65, 29, 41, 55, 56, 48, 51, 61, 73, 53, 60, 52, 69, 60, 
    58, 67, 37, 38, 77, 62, 57, 65, 70, 70, 54, 59, 62, 50, 64, 
    62, 73, 44, 31, 57, 70, 72, 73, 76, 56, 57, 59, 63, 49, 57, 
    59, 63, 56, 16, 46, 70, 76, 65, 75, 52, 54, 58, 56, 61, 53, 
    
    -- channel=134
    14, 126, 49, 12, 18, 36, 21, 27, 0, 0, 101, 29, 26, 23, 20, 
    17, 80, 73, 38, 6, 5, 27, 22, 3, 0, 108, 4, 9, 18, 18, 
    18, 36, 103, 43, 39, 0, 11, 38, 4, 26, 35, 11, 0, 5, 0, 
    0, 66, 67, 0, 50, 0, 0, 0, 24, 74, 0, 38, 0, 0, 8, 
    0, 25, 0, 0, 60, 7, 0, 0, 25, 52, 27, 22, 0, 0, 12, 
    0, 2, 0, 0, 31, 2, 0, 0, 13, 41, 25, 35, 0, 0, 0, 
    0, 1, 0, 12, 0, 22, 0, 40, 0, 16, 27, 32, 0, 0, 0, 
    0, 6, 0, 75, 0, 0, 0, 0, 19, 18, 0, 43, 15, 0, 0, 
    0, 9, 11, 48, 0, 0, 0, 0, 62, 0, 5, 0, 65, 0, 39, 
    0, 0, 7, 0, 5, 2, 0, 0, 0, 36, 0, 22, 30, 6, 27, 
    0, 0, 21, 0, 2, 0, 29, 13, 0, 0, 19, 27, 17, 0, 15, 
    0, 0, 37, 1, 0, 0, 15, 8, 0, 0, 47, 10, 19, 0, 0, 
    0, 0, 21, 0, 0, 47, 28, 5, 0, 0, 33, 11, 12, 13, 7, 
    0, 0, 22, 5, 0, 34, 0, 6, 0, 10, 27, 15, 0, 39, 21, 
    0, 0, 15, 19, 0, 0, 0, 17, 0, 39, 19, 19, 6, 29, 18, 
    
    -- channel=135
    13, 1, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 4, 9, 12, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    17, 11, 0, 0, 0, 0, 1, 5, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    0, 0, 11, 19, 3, 18, 6, 2, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 22, 22, 0, 0, 33, 7, 14, 16, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 15, 43, 59, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 19, 0, 0, 0, 0, 0, 7, 0, 2, 21, 12, 
    0, 0, 0, 8, 0, 8, 17, 22, 3, 0, 6, 0, 0, 0, 0, 
    0, 0, 7, 0, 3, 23, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 2, 15, 0, 0, 0, 0, 0, 0, 0, 
    5, 16, 16, 9, 11, 1, 16, 0, 20, 11, 17, 95, 41, 18, 0, 
    0, 0, 1, 0, 2, 0, 0, 0, 9, 9, 9, 0, 21, 57, 26, 
    0, 0, 0, 0, 0, 31, 27, 0, 0, 0, 28, 13, 0, 7, 11, 
    0, 0, 0, 0, 0, 0, 3, 15, 25, 24, 14, 0, 1, 12, 20, 
    0, 0, 0, 12, 16, 43, 0, 3, 11, 22, 0, 16, 11, 10, 1, 
    0, 9, 0, 0, 16, 23, 15, 24, 33, 24, 7, 17, 34, 27, 0, 
    5, 4, 0, 2, 8, 0, 22, 23, 30, 19, 3, 5, 13, 0, 6, 
    23, 0, 7, 10, 4, 13, 49, 33, 25, 0, 9, 5, 0, 1, 16, 
    
    -- channel=137
    0, 14, 98, 101, 97, 98, 94, 100, 98, 35, 76, 117, 110, 110, 107, 
    0, 0, 95, 107, 136, 108, 125, 127, 136, 85, 92, 157, 145, 135, 129, 
    0, 0, 73, 95, 174, 135, 93, 118, 128, 112, 139, 184, 182, 177, 166, 
    0, 10, 87, 118, 176, 171, 98, 79, 83, 110, 177, 192, 202, 195, 195, 
    142, 115, 161, 113, 144, 180, 162, 109, 96, 113, 170, 203, 218, 180, 167, 
    168, 162, 172, 125, 152, 170, 150, 105, 105, 114, 152, 216, 227, 187, 152, 
    169, 160, 136, 145, 138, 151, 144, 123, 135, 139, 153, 203, 229, 218, 163, 
    169, 163, 112, 149, 168, 159, 163, 114, 148, 132, 151, 174, 224, 225, 202, 
    167, 145, 147, 135, 194, 178, 156, 141, 102, 117, 141, 71, 128, 183, 187, 
    184, 150, 175, 167, 180, 203, 205, 166, 98, 125, 122, 107, 92, 110, 118, 
    196, 166, 186, 175, 179, 158, 168, 178, 177, 122, 107, 109, 124, 114, 101, 
    192, 174, 178, 202, 190, 157, 150, 160, 157, 110, 96, 120, 137, 113, 93, 
    183, 169, 173, 200, 174, 99, 158, 153, 141, 99, 103, 109, 118, 114, 96, 
    174, 149, 156, 204, 175, 105, 131, 122, 107, 80, 93, 95, 86, 85, 109, 
    159, 144, 131, 199, 181, 155, 115, 100, 79, 67, 86, 94, 82, 83, 103, 
    
    -- channel=138
    0, 0, 0, 0, 1, 0, 0, 0, 0, 45, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 16, 44, 44, 43, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 17, 0, 0, 0, 24, 0, 0, 0, 0, 0, 19, 4, 
    0, 0, 0, 0, 0, 6, 23, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 54, 0, 11, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 17, 0, 0, 0, 0, 19, 0, 7, 16, 67, 0, 21, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 1, 67, 45, 0, 
    0, 0, 0, 0, 12, 30, 0, 0, 0, 0, 32, 0, 0, 0, 43, 
    0, 17, 0, 0, 0, 24, 0, 6, 0, 45, 0, 0, 0, 7, 9, 
    0, 0, 0, 0, 7, 0, 0, 0, 4, 15, 0, 4, 0, 0, 0, 
    1, 7, 0, 0, 41, 33, 0, 14, 24, 13, 0, 3, 34, 0, 0, 
    7, 14, 0, 0, 0, 0, 27, 17, 26, 8, 0, 0, 10, 0, 0, 
    25, 0, 20, 0, 0, 20, 37, 6, 28, 0, 0, 0, 0, 0, 3, 
    
    -- channel=139
    19, 73, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 
    20, 56, 8, 0, 0, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 
    18, 34, 39, 0, 29, 0, 3, 14, 0, 0, 23, 0, 0, 0, 0, 
    0, 26, 25, 0, 43, 0, 0, 0, 5, 44, 0, 19, 0, 0, 4, 
    0, 1, 0, 0, 48, 9, 0, 0, 13, 36, 10, 15, 0, 0, 8, 
    0, 0, 0, 0, 19, 5, 0, 0, 7, 29, 18, 24, 0, 0, 0, 
    0, 0, 0, 0, 3, 21, 0, 16, 0, 22, 18, 20, 0, 0, 0, 
    0, 0, 0, 26, 0, 5, 0, 0, 7, 5, 0, 22, 9, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 24, 0, 0, 0, 43, 0, 19, 
    0, 0, 0, 0, 13, 14, 5, 0, 0, 1, 0, 0, 0, 0, 9, 
    0, 0, 13, 0, 0, 0, 23, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 20, 4, 0, 5, 1, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 12, 24, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    
    -- channel=140
    20, 123, 68, 15, 27, 36, 28, 38, 1, 0, 98, 54, 33, 35, 27, 
    22, 83, 98, 22, 29, 16, 36, 44, 21, 0, 156, 36, 25, 28, 23, 
    20, 46, 128, 40, 57, 0, 6, 38, 2, 19, 97, 39, 26, 33, 27, 
    5, 79, 145, 0, 71, 0, 2, 0, 28, 83, 39, 72, 26, 12, 41, 
    6, 86, 41, 0, 87, 18, 0, 0, 32, 57, 55, 83, 26, 0, 62, 
    27, 41, 26, 0, 62, 17, 0, 0, 40, 57, 51, 86, 29, 0, 42, 
    28, 29, 0, 45, 15, 21, 0, 30, 16, 45, 48, 88, 36, 17, 12, 
    18, 33, 0, 95, 7, 25, 0, 27, 33, 29, 28, 52, 61, 20, 36, 
    0, 31, 4, 66, 18, 30, 8, 0, 59, 1, 34, 4, 72, 10, 79, 
    12, 36, 40, 21, 32, 20, 13, 0, 9, 49, 0, 25, 37, 26, 50, 
    28, 7, 51, 24, 29, 0, 50, 24, 0, 0, 15, 44, 35, 0, 23, 
    34, 0, 76, 22, 13, 0, 49, 23, 12, 0, 67, 19, 38, 7, 2, 
    28, 13, 66, 25, 0, 0, 48, 15, 0, 0, 51, 14, 21, 11, 17, 
    19, 15, 65, 41, 0, 39, 11, 12, 0, 0, 42, 21, 0, 47, 32, 
    12, 29, 47, 59, 5, 6, 0, 20, 0, 46, 27, 31, 11, 44, 27, 
    
    -- channel=141
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    94, 115, 55, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=142
    0, 0, 42, 44, 37, 37, 48, 41, 43, 27, 0, 54, 60, 59, 61, 
    0, 0, 29, 22, 24, 35, 30, 41, 50, 22, 2, 51, 57, 58, 60, 
    0, 0, 0, 30, 21, 40, 13, 18, 27, 0, 37, 33, 46, 49, 52, 
    11, 0, 31, 46, 18, 28, 28, 25, 5, 2, 36, 30, 54, 57, 30, 
    32, 34, 40, 33, 15, 27, 36, 27, 3, 1, 19, 49, 48, 48, 32, 
    39, 35, 43, 29, 29, 32, 36, 2, 16, 6, 19, 38, 51, 50, 34, 
    43, 35, 48, 35, 32, 4, 33, 0, 33, 15, 12, 43, 50, 51, 41, 
    43, 35, 56, 30, 42, 35, 12, 37, 10, 18, 38, 24, 40, 60, 27, 
    47, 23, 36, 46, 28, 42, 34, 34, 9, 22, 36, 32, 15, 27, 22, 
    42, 31, 43, 38, 35, 36, 27, 28, 42, 22, 44, 27, 22, 40, 34, 
    40, 42, 24, 43, 39, 48, 23, 29, 35, 54, 8, 32, 36, 29, 27, 
    39, 42, 24, 42, 54, 33, 42, 38, 44, 30, 19, 30, 31, 33, 24, 
    38, 37, 25, 39, 58, 6, 39, 39, 38, 22, 21, 21, 29, 16, 25, 
    38, 35, 17, 34, 43, 35, 50, 33, 27, 6, 20, 18, 17, 11, 22, 
    25, 27, 16, 27, 35, 47, 30, 25, 23, 1, 15, 19, 15, 21, 21, 
    
    -- channel=143
    22, 0, 0, 13, 16, 0, 16, 6, 24, 75, 0, 3, 6, 10, 11, 
    20, 0, 0, 0, 0, 31, 0, 0, 12, 47, 0, 7, 12, 8, 8, 
    21, 9, 0, 1, 0, 46, 14, 0, 0, 0, 0, 0, 2, 2, 11, 
    81, 0, 0, 45, 0, 0, 28, 35, 0, 0, 0, 0, 0, 25, 0, 
    31, 9, 17, 53, 0, 0, 9, 37, 0, 0, 0, 0, 1, 52, 7, 
    15, 9, 19, 25, 0, 0, 18, 7, 1, 0, 0, 0, 8, 53, 39, 
    27, 10, 41, 0, 14, 0, 26, 0, 19, 0, 0, 0, 0, 16, 47, 
    38, 3, 36, 0, 19, 2, 0, 21, 0, 6, 9, 0, 0, 22, 0, 
    54, 7, 0, 0, 0, 0, 15, 33, 0, 7, 1, 33, 0, 0, 0, 
    36, 21, 0, 0, 0, 0, 0, 2, 42, 0, 29, 0, 0, 20, 3, 
    17, 42, 0, 2, 0, 36, 0, 0, 1, 42, 0, 0, 0, 15, 13, 
    17, 42, 0, 0, 5, 0, 0, 0, 10, 34, 0, 6, 0, 17, 17, 
    25, 41, 0, 0, 33, 0, 0, 1, 14, 20, 0, 5, 8, 0, 12, 
    30, 47, 0, 0, 20, 0, 22, 5, 17, 9, 1, 5, 20, 0, 0, 
    26, 32, 21, 0, 5, 24, 25, 0, 30, 0, 6, 3, 12, 8, 0, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 25, 30, 37, 21, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 9, 0, 1, 24, 30, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 28, 8, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 13, 26, 36, 29, 29, 24, 22, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 53, 31, 22, 40, 48, 40, 41, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 26, 21, 14, 13, 9, 13, 24, 3, 0, 
    0, 0, 0, 0, 34, 33, 24, 16, 42, 51, 31, 47, 69, 41, 0, 
    0, 0, 0, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 17, 0, 39, 23, 42, 18, 41, 39, 44, 45, 22, 30, 21, 
    0, 0, 0, 0, 5, 23, 0, 0, 47, 9, 20, 6, 3, 0, 6, 
    0, 0, 11, 0, 0, 9, 49, 26, 15, 5, 0, 0, 11, 50, 26, 
    4, 0, 0, 3, 0, 0, 6, 11, 13, 0, 0, 0, 1, 12, 10, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 53, 38, 4, 0, 10, 22, 
    10, 4, 0, 10, 10, 0, 0, 0, 5, 13, 24, 14, 0, 12, 12, 
    
    -- channel=146
    34, 34, 37, 18, 29, 40, 35, 43, 39, 28, 25, 30, 22, 25, 9, 
    43, 43, 35, 11, 31, 44, 43, 33, 34, 15, 15, 36, 28, 4, 21, 
    45, 46, 31, 12, 72, 80, 81, 74, 72, 62, 43, 39, 27, 0, 15, 
    45, 40, 40, 14, 96, 74, 66, 77, 77, 84, 52, 44, 25, 17, 8, 
    44, 39, 27, 24, 79, 77, 58, 80, 81, 78, 62, 68, 43, 24, 47, 
    50, 32, 34, 32, 63, 70, 76, 66, 61, 71, 64, 53, 67, 44, 46, 
    52, 21, 36, 34, 74, 77, 62, 62, 74, 55, 37, 53, 49, 44, 44, 
    33, 11, 49, 27, 52, 47, 64, 51, 34, 32, 40, 30, 47, 67, 71, 
    42, 10, 51, 3, 56, 56, 42, 31, 64, 71, 35, 51, 81, 67, 72, 
    35, 7, 26, 13, 41, 29, 43, 69, 31, 61, 43, 46, 50, 32, 87, 
    47, 0, 35, 19, 25, 37, 55, 36, 47, 50, 50, 62, 48, 60, 78, 
    52, 0, 32, 49, 13, 21, 38, 0, 62, 19, 39, 52, 0, 30, 83, 
    60, 32, 61, 41, 20, 13, 11, 17, 32, 78, 44, 14, 10, 32, 91, 
    69, 50, 39, 32, 37, 5, 15, 25, 34, 45, 51, 8, 6, 45, 83, 
    62, 58, 43, 27, 32, 16, 20, 25, 32, 42, 50, 20, 11, 37, 98, 
    
    -- channel=147
    70, 58, 85, 96, 61, 58, 51, 43, 52, 76, 74, 57, 82, 53, 64, 
    80, 77, 116, 153, 90, 73, 70, 86, 79, 56, 54, 47, 68, 93, 22, 
    83, 82, 117, 199, 37, 69, 70, 91, 75, 50, 0, 53, 93, 94, 0, 
    82, 99, 86, 218, 18, 86, 147, 108, 106, 85, 77, 16, 76, 101, 45, 
    77, 108, 134, 171, 45, 75, 124, 94, 94, 85, 115, 16, 53, 103, 48, 
    49, 131, 113, 181, 24, 69, 104, 93, 89, 72, 81, 31, 1, 84, 81, 
    54, 128, 74, 110, 58, 92, 125, 94, 75, 105, 94, 31, 37, 49, 67, 
    95, 128, 0, 141, 87, 78, 60, 99, 71, 54, 77, 58, 6, 30, 0, 
    98, 135, 14, 131, 30, 65, 73, 82, 25, 12, 97, 35, 8, 86, 0, 
    105, 175, 37, 85, 24, 73, 30, 4, 105, 58, 92, 70, 79, 103, 0, 
    85, 189, 49, 68, 49, 11, 6, 113, 0, 78, 57, 5, 90, 43, 0, 
    104, 209, 2, 60, 105, 25, 9, 105, 0, 78, 65, 74, 133, 39, 0, 
    87, 147, 41, 94, 96, 75, 28, 16, 0, 0, 96, 186, 86, 0, 0, 
    80, 122, 128, 102, 70, 104, 21, 13, 10, 6, 40, 191, 63, 0, 0, 
    102, 97, 128, 99, 61, 70, 32, 29, 25, 30, 34, 119, 66, 0, 0, 
    
    -- channel=148
    28, 33, 23, 0, 0, 29, 54, 97, 48, 7, 4, 0, 38, 46, 19, 
    13, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 1, 0, 50, 58, 61, 14, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 18, 0, 7, 0, 6, 29, 2, 0, 0, 42, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 33, 106, 
    0, 0, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 74, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 13, 9, 0, 0, 5, 6, 58, 184, 181, 171, 189, 160, 46, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 15, 0, 0, 0, 46, 28, 0, 4, 0, 30, 0, 31, 7, 
    0, 0, 0, 67, 31, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 83, 107, 0, 10, 26, 0, 0, 0, 98, 91, 58, 0, 0, 29, 
    6, 0, 0, 0, 0, 4, 19, 20, 26, 0, 0, 0, 0, 7, 0, 
    0, 0, 2, 0, 0, 0, 17, 15, 4, 0, 0, 0, 12, 0, 27, 
    
    -- channel=149
    29, 34, 39, 50, 27, 13, 6, 12, 20, 27, 41, 27, 32, 42, 34, 
    22, 23, 37, 40, 0, 0, 0, 0, 0, 4, 31, 31, 36, 58, 34, 
    23, 23, 29, 49, 0, 0, 0, 0, 0, 0, 0, 27, 57, 60, 36, 
    23, 30, 22, 28, 0, 0, 0, 0, 0, 0, 0, 12, 27, 61, 52, 
    21, 31, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 32, 36, 
    17, 41, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 23, 
    29, 45, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    51, 56, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 39, 20, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 58, 2, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 39, 7, 0, 4, 0, 0, 25, 0, 0, 0, 0, 15, 0, 0, 
    4, 51, 0, 0, 13, 4, 0, 0, 0, 0, 0, 11, 4, 0, 0, 
    0, 0, 5, 0, 0, 15, 0, 0, 0, 0, 0, 24, 9, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 21, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 2, 13, 5, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 20, 10, 15, 8, 0, 9, 0, 0, 8, 
    0, 0, 0, 0, 34, 12, 14, 0, 6, 25, 62, 2, 0, 0, 26, 
    0, 0, 0, 0, 74, 25, 0, 0, 0, 13, 0, 45, 0, 0, 0, 
    0, 0, 0, 0, 42, 22, 0, 10, 12, 12, 0, 60, 11, 0, 5, 
    23, 0, 0, 0, 43, 17, 7, 8, 4, 19, 15, 27, 57, 0, 0, 
    25, 0, 8, 0, 25, 15, 0, 5, 31, 6, 0, 45, 42, 36, 3, 
    1, 0, 74, 0, 6, 0, 18, 4, 14, 15, 12, 22, 46, 51, 80, 
    0, 0, 53, 0, 42, 31, 5, 0, 28, 39, 0, 9, 47, 15, 91, 
    0, 0, 35, 0, 37, 0, 31, 79, 0, 28, 0, 10, 19, 0, 129, 
    1, 0, 10, 0, 13, 41, 43, 0, 57, 0, 10, 41, 0, 32, 99, 
    0, 0, 52, 9, 0, 25, 53, 0, 101, 0, 8, 25, 0, 24, 133, 
    6, 0, 29, 0, 0, 0, 17, 26, 45, 106, 0, 0, 0, 41, 122, 
    17, 0, 0, 0, 7, 0, 18, 31, 45, 46, 35, 0, 0, 62, 101, 
    0, 0, 0, 0, 9, 0, 14, 20, 27, 32, 39, 0, 0, 50, 114, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 0, 0, 0, 20, 27, 3, 13, 13, 0, 0, 
    0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 14, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 1, 9, 0, 0, 7, 21, 34, 0, 0, 0, 0, 18, 18, 0, 
    0, 0, 0, 0, 0, 0, 12, 10, 1, 0, 0, 0, 6, 3, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=152
    0, 0, 0, 14, 18, 5, 0, 0, 0, 5, 0, 3, 0, 0, 0, 
    0, 0, 15, 70, 65, 65, 74, 99, 102, 62, 23, 0, 8, 6, 0, 
    2, 3, 23, 0, 0, 0, 0, 0, 0, 0, 11, 0, 7, 19, 12, 
    1, 4, 6, 49, 17, 46, 18, 20, 2, 2, 0, 27, 1, 0, 4, 
    5, 9, 65, 61, 9, 20, 49, 18, 22, 19, 9, 6, 1, 0, 0, 
    22, 36, 11, 12, 19, 4, 8, 31, 27, 2, 41, 1, 0, 2, 1, 
    9, 51, 33, 11, 0, 20, 40, 19, 36, 64, 38, 38, 62, 83, 14, 
    40, 55, 14, 26, 22, 0, 0, 11, 54, 41, 34, 65, 41, 14, 10, 
    8, 27, 0, 81, 0, 52, 26, 0, 0, 0, 0, 0, 0, 15, 24, 
    7, 29, 53, 8, 30, 10, 7, 48, 31, 20, 39, 27, 52, 28, 0, 
    14, 34, 0, 4, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 45, 35, 0, 0, 1, 47, 57, 42, 62, 10, 54, 54, 34, 0, 
    15, 0, 0, 14, 0, 0, 6, 0, 0, 0, 2, 14, 19, 0, 0, 
    6, 31, 9, 31, 14, 3, 0, 0, 10, 27, 41, 38, 11, 0, 0, 
    23, 9, 4, 29, 11, 9, 0, 0, 0, 0, 17, 41, 0, 0, 0, 
    
    -- channel=153
    213, 203, 214, 168, 176, 162, 169, 175, 207, 226, 215, 224, 199, 179, 176, 
    242, 240, 238, 165, 168, 181, 178, 202, 225, 215, 216, 218, 225, 195, 205, 
    251, 252, 239, 138, 140, 142, 141, 136, 140, 141, 187, 222, 206, 177, 183, 
    250, 248, 221, 174, 171, 210, 192, 201, 190, 185, 155, 222, 213, 174, 141, 
    248, 247, 203, 168, 161, 173, 196, 181, 190, 193, 201, 191, 225, 217, 171, 
    235, 239, 176, 120, 120, 152, 147, 150, 152, 158, 177, 172, 232, 252, 251, 
    198, 193, 151, 133, 106, 138, 153, 118, 132, 151, 120, 142, 204, 242, 255, 
    178, 123, 135, 129, 136, 105, 102, 91, 86, 85, 77, 82, 122, 146, 233, 
    170, 98, 111, 108, 112, 117, 123, 85, 56, 65, 80, 48, 84, 136, 193, 
    194, 100, 114, 48, 82, 79, 83, 126, 157, 155, 160, 154, 173, 119, 152, 
    201, 111, 57, 61, 29, 64, 79, 53, 110, 99, 100, 112, 87, 116, 123, 
    203, 96, 93, 86, 29, 20, 75, 75, 71, 129, 122, 140, 80, 93, 125, 
    194, 124, 62, 134, 71, 13, 8, 15, 28, 133, 156, 131, 29, 46, 105, 
    187, 189, 137, 125, 91, 37, 5, 17, 43, 115, 172, 144, 22, 44, 123, 
    190, 173, 146, 88, 80, 49, 24, 32, 43, 70, 103, 121, 12, 45, 131, 
    
    -- channel=154
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 82, 61, 49, 84, 105, 71, 28, 8, 0, 0, 17, 0, 
    0, 0, 1, 58, 0, 0, 0, 0, 0, 41, 0, 0, 22, 28, 2, 
    0, 0, 5, 61, 0, 0, 25, 0, 0, 0, 41, 0, 0, 0, 26, 
    0, 0, 93, 49, 0, 35, 22, 0, 3, 4, 0, 0, 0, 0, 0, 
    0, 27, 0, 62, 25, 0, 24, 26, 28, 12, 27, 3, 0, 0, 0, 
    10, 54, 44, 0, 0, 14, 0, 0, 0, 4, 30, 36, 71, 41, 0, 
    19, 101, 0, 29, 33, 14, 30, 50, 56, 36, 49, 58, 20, 28, 0, 
    0, 19, 0, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 84, 19, 14, 28, 23, 55, 9, 58, 57, 70, 54, 37, 61, 0, 
    0, 30, 3, 0, 32, 0, 0, 72, 0, 19, 0, 0, 67, 0, 0, 
    15, 111, 0, 0, 16, 31, 83, 20, 20, 0, 0, 56, 55, 72, 0, 
    0, 0, 0, 2, 0, 16, 0, 0, 0, 0, 0, 0, 43, 0, 0, 
    0, 22, 9, 9, 0, 4, 0, 0, 0, 67, 29, 59, 8, 0, 0, 
    14, 0, 4, 45, 2, 0, 0, 0, 0, 5, 26, 3, 15, 0, 0, 
    
    -- channel=155
    0, 1, 0, 0, 4, 0, 0, 0, 6, 0, 0, 4, 0, 0, 0, 
    4, 4, 0, 0, 36, 58, 55, 47, 46, 25, 7, 12, 1, 0, 10, 
    10, 11, 0, 0, 79, 66, 68, 57, 66, 67, 48, 11, 0, 0, 20, 
    10, 6, 8, 0, 97, 49, 42, 77, 67, 66, 47, 43, 0, 0, 0, 
    12, 0, 10, 3, 95, 92, 57, 84, 80, 81, 51, 53, 16, 0, 0, 
    27, 0, 0, 0, 97, 82, 69, 82, 81, 90, 84, 83, 63, 9, 11, 
    25, 0, 19, 2, 62, 69, 61, 59, 72, 56, 37, 70, 66, 46, 21, 
    0, 0, 41, 0, 67, 57, 66, 50, 67, 72, 56, 71, 101, 90, 77, 
    0, 0, 46, 0, 66, 44, 34, 4, 10, 17, 0, 0, 46, 45, 91, 
    0, 0, 41, 3, 72, 39, 74, 90, 39, 75, 56, 64, 60, 31, 124, 
    9, 0, 23, 20, 34, 61, 59, 22, 88, 44, 56, 69, 32, 56, 98, 
    21, 0, 53, 20, 0, 46, 86, 7, 93, 20, 32, 48, 0, 64, 130, 
    45, 0, 32, 30, 6, 3, 29, 38, 51, 75, 0, 0, 8, 51, 123, 
    45, 27, 15, 22, 37, 0, 24, 34, 47, 83, 67, 0, 10, 70, 116, 
    47, 43, 12, 17, 39, 15, 24, 31, 42, 53, 69, 8, 6, 62, 125, 
    
    -- channel=156
    23, 32, 16, 0, 21, 28, 37, 68, 66, 29, 27, 30, 5, 45, 8, 
    21, 23, 2, 0, 0, 9, 0, 0, 14, 29, 20, 49, 24, 1, 57, 
    17, 19, 0, 0, 19, 10, 0, 0, 0, 21, 71, 44, 9, 0, 67, 
    16, 10, 0, 0, 85, 20, 0, 0, 0, 3, 34, 61, 1, 4, 31, 
    20, 2, 0, 0, 49, 13, 0, 0, 3, 0, 0, 72, 45, 0, 31, 
    35, 0, 0, 0, 21, 0, 0, 0, 0, 7, 0, 33, 79, 16, 19, 
    31, 0, 0, 0, 18, 0, 0, 0, 15, 8, 0, 42, 46, 20, 38, 
    2, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 14, 30, 26, 96, 
    0, 0, 84, 0, 40, 23, 6, 0, 48, 60, 2, 38, 81, 17, 100, 
    0, 0, 33, 0, 32, 0, 12, 42, 0, 0, 0, 0, 0, 0, 119, 
    0, 0, 25, 0, 0, 17, 35, 0, 39, 0, 0, 38, 0, 38, 90, 
    0, 0, 32, 26, 0, 23, 42, 0, 105, 0, 20, 46, 0, 18, 102, 
    0, 0, 39, 10, 0, 0, 17, 23, 32, 148, 29, 0, 0, 31, 122, 
    13, 0, 0, 0, 0, 0, 20, 33, 49, 59, 2, 0, 0, 63, 91, 
    0, 0, 0, 0, 5, 0, 13, 19, 22, 24, 28, 0, 0, 49, 121, 
    
    -- channel=157
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 7, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 36, 131, 122, 106, 136, 84, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 32, 38, 0, 0, 6, 0, 0, 0, 53, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 2, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=158
    39, 44, 45, 32, 23, 24, 26, 37, 52, 43, 47, 39, 38, 42, 30, 
    48, 49, 58, 28, 15, 2, 0, 6, 16, 14, 27, 42, 43, 42, 28, 
    47, 48, 46, 34, 0, 0, 0, 0, 0, 0, 0, 46, 54, 40, 20, 
    47, 54, 30, 27, 0, 0, 19, 0, 0, 0, 21, 15, 34, 50, 38, 
    46, 54, 34, 0, 0, 0, 0, 0, 0, 0, 0, 11, 42, 47, 36, 
    35, 58, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 13, 48, 48, 
    41, 37, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 8, 42, 
    49, 18, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    44, 9, 25, 0, 0, 0, 0, 0, 0, 0, 13, 0, 6, 1, 0, 
    39, 15, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    34, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    7, 0, 4, 10, 0, 0, 0, 0, 0, 0, 35, 42, 0, 0, 0, 
    12, 15, 0, 6, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    4, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    0, 1, 0, 26, 0, 0, 0, 0, 0, 0, 9, 0, 9, 20, 21, 
    0, 0, 8, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 
    0, 0, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 15, 29, 0, 
    0, 0, 0, 61, 0, 0, 1, 0, 0, 0, 1, 0, 0, 35, 25, 
    0, 0, 23, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 6, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 32, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 42, 0, 38, 0, 0, 0, 0, 0, 0, 25, 15, 0, 0, 0, 
    0, 73, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 63, 10, 3, 14, 0, 0, 53, 0, 2, 0, 0, 28, 0, 0, 
    0, 81, 0, 0, 50, 11, 0, 0, 0, 0, 0, 0, 21, 0, 0, 
    0, 7, 16, 0, 8, 44, 12, 1, 0, 0, 5, 56, 38, 0, 0, 
    0, 0, 1, 0, 0, 34, 14, 2, 0, 0, 0, 40, 19, 0, 0, 
    0, 0, 3, 19, 0, 9, 12, 4, 0, 0, 0, 0, 36, 0, 0, 
    
    
    others => 0);
end gold_package;
