-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        INPUT_SIZE : integer := 8;
        ADDRESS_SIZE    : integer := 12;
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(ADDRESS_SIZE-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(4-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
          

    MEM_IWGHT_LAYER0_ENTITY0 : if BRAM_NAME = "iwght_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffff05b000004fefffffa57000008940000001d000008a40000112a00001869",
            INIT_01 => X"fffffcf0ffffdeecfffffeba000013d20000188d00000a4bffffcfa000001da3",
            INIT_02 => X"0000001f000000220000000afffffff7ffffffcaffffffe50000000000000004",
            INIT_03 => X"000000030000002c0000002effffffd300000038ffffffffffffffdd00000018",
            INIT_04 => X"00000035000000210000002000000018ffffffc9ffffffccffffffc3ffffffed",
            INIT_05 => X"ffffffc6ffffffda0000000bffffffe60000001b0000001fffffffd3ffffffc0",
            INIT_06 => X"ffffffc6ffffffe200000010fffffff50000001700000018000000250000000f",
            INIT_07 => X"ffffffd8ffffffd8fffffff6ffffffd3000000070000000700000032fffffff3",
            INIT_08 => X"000000260000001d00000033ffffffd8000000060000000cffffffcf00000013",
            INIT_09 => X"fffffff3000000200000000500000024fffffffffffffffb0000000bffffffeb",
            INIT_0A => X"ffffffdffffffffaffffffc1ffffffdcfffffff4ffffffec0000000effffffdb",
            INIT_0B => X"000000320000000900000027ffffffe100000006000000370000002d00000018",
            INIT_0C => X"000000240000001200000002ffffffe6000000210000002dffffffee00000016",
            INIT_0D => X"ffffffe7ffffffc6fffffff8fffffffbffffffc200000037fffffffcffffffd2",
            INIT_0E => X"ffffffe60000001effffffc2000000400000001f000000000000003400000010",
            INIT_0F => X"fffffff5000000520000001effffffccffffffe5ffffffc6ffffffe6fffffff6",
            INIT_10 => X"0000002bffffffeb0000004d0000002bfffffffaffffffbeffffffaffffffffc",
            INIT_11 => X"ffffffcdfffffffd0000002b000000220000004400000039ffffffe1ffffffc2",
            INIT_12 => X"ffffffe100000001000000390000000b00000033fffffffafffffff90000002c",
            INIT_13 => X"00000028000000260000001f0000002f0000003b000000450000002ffffffffa",
            INIT_14 => X"0000001bffffffeffffffff0ffffffe600000018ffffffe400000021fffffff8",
            INIT_15 => X"ffffffd5ffffffd6ffffffd200000004ffffffe5ffffffcaffffffc6fffffff4",
            INIT_16 => X"ffffffe9ffffffd600000019000000000000001c000000040000003000000033",
            INIT_17 => X"ffffffd60000000d00000044ffffffbefffffffc00000005ffffffb3ffffffc1",
            INIT_18 => X"00000022fffffff0ffffffd0fffffff500000009ffffffe40000001cffffffbc",
            INIT_19 => X"00000010000000250000000f000000000000000e000000260000004000000011",
            INIT_1A => X"000000330000002dffffffea0000001f0000003400000000fffffff0ffffffcd",
            INIT_1B => X"fffffff6fffffff500000009ffffffc9ffffffc4ffffffbbffffffd300000021",
            INIT_1C => X"0000001c0000000affffffc7ffffffba00000000fffffff2ffffffc600000028",
            INIT_1D => X"000000150000002dffffffff000000340000003c00000033fffffff7ffffffcb",
            INIT_1E => X"ffffffc70000002f00000003ffffffdefffffff8fffffff700000017ffffffd1",
            INIT_1F => X"ffffffc9ffffffc5fffffff80000000afffffffc0000000b000000390000001c",
            INIT_20 => X"fffffff7ffffffd5fffffff90000000300000002fffffffbfffffffafffffff8",
            INIT_21 => X"00000016ffffffc1ffffffc5fffffff00000002b0000001effffffdf0000001d",
            INIT_22 => X"0000001b00000017000000310000002dfffffff3000000200000003b00000028",
            INIT_23 => X"ffffffe90000002900000006fffffff70000002c00000027000000140000003d",
            INIT_24 => X"0000002500000025fffffff5ffffffd2fffffff1ffffffd8ffffffc80000001d",
            INIT_25 => X"00000010000000310000001effffffe40000001200000021ffffffbfffffffae",
            INIT_26 => X"ffffffe60000001d00000045fffffff3ffffffdcffffffda0000003500000010",
            INIT_27 => X"ffffffcbffffffedffffffdd0000001cffffffd0fffffff7ffffffe6ffffffd5",
            INIT_28 => X"ffffffecffffffe0ffffffd9fffffffd00000026ffffffe3ffffffe2fffffff9",
            INIT_29 => X"00000015000000010000001f0000002f0000001600000033ffffffea0000002c",
            INIT_2A => X"00000033ffffffe5fffffffb00000033ffffffc5ffffffdb0000003effffffe0",
            INIT_2B => X"fffffff90000001bffffffd700000028fffffff8ffffffd70000000500000026",
            INIT_2C => X"000000030000000a0000004bfffffff30000003a00000030ffffffd8fffffffe",
            INIT_2D => X"fffffff9ffffffc700000029ffffffffffffffd7ffffffebfffffffaffffffdd",
            INIT_2E => X"ffffffc9ffffffd9ffffffdfffffffe400000034fffffff90000004dfffffffe",
            INIT_2F => X"ffffffd6ffffffffffffffbfffffffec00000019000000130000003d00000003",
            INIT_30 => X"0000001bffffffdbfffffff2ffffffbcffffffe900000007ffffffff00000036",
            INIT_31 => X"ffffffe80000003efffffffb000000380000000f00000024000000120000000a",
            INIT_32 => X"000000230000002d0000000affffffe400000010fffffffa0000001500000029",
            INIT_33 => X"ffffffd1fffffff7fffffffdffffffd1ffffffdfffffffe00000000900000019",
            INIT_34 => X"ffffffda00000010fffffff70000001affffffebfffffff50000000dffffffdd",
            INIT_35 => X"00000018ffffffe1ffffffef00000013ffffffe4ffffffd20000000200000031",
            INIT_36 => X"000000140000004600000026fffffff0000000420000002bfffffff5ffffffdb",
            INIT_37 => X"ffffffcffffffff8fffffff7ffffffe4ffffffda00000023fffffff2ffffffcc",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY0 : if BRAM_NAME = "ifmap_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e0000009f000000a5000000a6000000a00000009c000000a20000009f",
            INIT_01 => X"0000009e0000009f000000a1000000a0000000a1000000a6000000a9000000aa",
            INIT_02 => X"000000a7000000a2000000a0000000a00000009c000000950000009600000094",
            INIT_03 => X"000000950000008f0000008c0000008d0000008f000000890000007e00000074",
            INIT_04 => X"00000098000000970000009f000000a6000000a2000000a0000000a4000000a2",
            INIT_05 => X"000000a30000009c0000009b0000009f000000a3000000aa000000ab000000ab",
            INIT_06 => X"000000a9000000a00000009a00000097000000910000008b0000008c0000008d",
            INIT_07 => X"0000009500000093000000910000008e0000008f000000880000007d00000077",
            INIT_08 => X"00000097000000970000009e000000a7000000a0000000a3000000a5000000a5",
            INIT_09 => X"000000a3000000a20000009e0000009d000000a1000000a6000000a7000000a9",
            INIT_0A => X"000000aa0000009f00000091000000790000006e000000620000006500000072",
            INIT_0B => X"00000078000000860000008f0000008c0000008e0000008b0000008200000078",
            INIT_0C => X"0000009b0000009b000000a0000000ae000000a7000000a7000000a9000000a9",
            INIT_0D => X"000000a5000000a5000000a7000000bf000000b10000009d000000a2000000a4",
            INIT_0E => X"0000009e000000950000006800000067000000620000005c000000500000004a",
            INIT_0F => X"000000560000005300000071000000840000008c0000008c000000880000007f",
            INIT_10 => X"0000009b0000009c000000a1000000aa000000a9000000a3000000a9000000a6",
            INIT_11 => X"000000a4000000a4000000ad000000f6000000c300000097000000920000008e",
            INIT_12 => X"0000006f0000004e0000005500000071000000700000006a000000610000005d",
            INIT_13 => X"0000004a000000540000005500000069000000800000008a0000008500000081",
            INIT_14 => X"00000094000000850000008200000093000000a1000000a5000000a7000000a7",
            INIT_15 => X"000000a3000000a5000000a3000000b40000009d000000800000006100000042",
            INIT_16 => X"000000450000004200000059000000760000007a00000077000000720000005e",
            INIT_17 => X"000000630000005b0000003a000000430000006c0000008c0000008a00000086",
            INIT_18 => X"0000007f0000006d0000002f0000005800000099000000aa000000a8000000aa",
            INIT_19 => X"000000a9000000a6000000a400000093000000810000007f0000006400000044",
            INIT_1A => X"0000004e000000480000005300000084000000920000007c000000690000006b",
            INIT_1B => X"00000073000000550000003f0000002e0000004f000000840000008d00000086",
            INIT_1C => X"00000083000000630000002a000000460000008f000000a7000000a5000000a8",
            INIT_1D => X"000000ab000000a10000008c0000007800000082000000900000007400000058",
            INIT_1E => X"0000005b000000550000004d0000007c000000a300000088000000660000006a",
            INIT_1F => X"00000064000000550000003600000031000000390000006b0000008a00000088",
            INIT_20 => X"000000aa00000067000000360000007c00000099000000a1000000a3000000a6",
            INIT_21 => X"000000a5000000ae000000710000007d0000009d0000009c0000007900000056",
            INIT_22 => X"000000520000005400000050000000510000008a000000920000007100000057",
            INIT_23 => X"00000053000000560000004700000038000000280000004a0000008500000089",
            INIT_24 => X"000000b4000000860000005e0000009a000000ae0000009e0000009c00000099",
            INIT_25 => X"000000cf000000ed000000cf0000009c000000ae000000940000007d0000005d",
            INIT_26 => X"000000560000004a0000003b0000004c000000890000008f000000850000006a",
            INIT_27 => X"0000005600000057000000540000004b00000032000000280000005f00000084",
            INIT_28 => X"000000b70000006c0000008e000000a5000000b10000009b0000009f0000007a",
            INIT_29 => X"000000d5000000ed000000dc000000a4000000b70000009c0000007d00000078",
            INIT_2A => X"0000004e000000500000002d0000005b000000af0000009d0000009b0000006b",
            INIT_2B => X"0000005700000067000000580000004e0000003b000000290000003b00000068",
            INIT_2C => X"000000bc0000006400000087000000aa000000bb000000a6000000ad00000086",
            INIT_2D => X"00000075000000c2000000c7000000aa000000b9000000bd0000008600000075",
            INIT_2E => X"0000006600000054000000260000007d000000d2000000a0000000920000005d",
            INIT_2F => X"000000530000005e000000680000005500000049000000370000003e0000004c",
            INIT_30 => X"000000bd0000005a0000007f000000af000000ae000000a6000000b20000009f",
            INIT_31 => X"00000061000000a8000000a800000089000000ba000000d8000000a00000007b",
            INIT_32 => X"00000078000000730000003200000096000000c20000009b0000007b0000005b",
            INIT_33 => X"00000054000000540000005f0000005600000054000000490000004f00000049",
            INIT_34 => X"000000bd0000005d00000098000000b90000007700000088000000ad000000a7",
            INIT_35 => X"000000670000009300000091000000a7000000bd000000e2000000b40000008d",
            INIT_36 => X"0000007e00000075000000470000009a000000ba000000950000007200000057",
            INIT_37 => X"00000050000000480000005000000063000000640000005a000000610000005e",
            INIT_38 => X"000000c20000006c000000a8000000ba00000069000000630000009c000000a7",
            INIT_39 => X"00000064000000730000008a000000c6000000be000000ac000000910000009a",
            INIT_3A => X"00000092000000670000004700000098000000b300000089000000820000006e",
            INIT_3B => X"000000550000005b0000005f0000006d00000073000000640000006100000075",
            INIT_3C => X"000000c500000084000000ac000000b8000000820000004e0000008c0000009b",
            INIT_3D => X"00000073000000820000008f000000e6000000f2000000910000008700000083",
            INIT_3E => X"000000790000006c0000005f00000090000000a8000000980000007000000057",
            INIT_3F => X"0000004700000057000000690000007000000078000000670000007900000088",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY1 : if BRAM_NAME = "ifmap_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cb00000092000000a8000000bf000000a80000004e0000007e0000008a",
            INIT_01 => X"0000008a000000600000009a000000ad000000a20000008c0000007100000071",
            INIT_02 => X"000000650000006900000070000000ab0000009c00000094000000870000006d",
            INIT_03 => X"0000004e0000004f0000005e000000650000006b0000007d0000009700000090",
            INIT_04 => X"000000d6000000a3000000a4000000b7000000b00000005e000000600000009c",
            INIT_05 => X"000000940000006a000000810000007600000072000000740000006600000073",
            INIT_06 => X"000000560000006500000090000000760000004400000080000000850000004b",
            INIT_07 => X"0000003c0000003a0000004700000066000000740000008f000000960000008c",
            INIT_08 => X"000000d4000000b2000000a7000000ad000000b00000007c000000560000008d",
            INIT_09 => X"0000009900000087000000680000004d000000860000007c0000008100000093",
            INIT_0A => X"000000550000005c0000009600000084000000750000006b0000004b00000040",
            INIT_0B => X"0000002c0000004100000056000000850000009b000000a00000009a00000097",
            INIT_0C => X"000000c7000000bb000000ab000000ae000000b1000000900000005600000077",
            INIT_0D => X"0000007a000000890000009000000046000000810000006c00000091000000b8",
            INIT_0E => X"0000007400000049000000830000008900000086000000590000003300000034",
            INIT_0F => X"0000002f0000005a00000079000000a3000000ab000000a40000009e00000095",
            INIT_10 => X"000000a5000000c3000000b3000000b1000000b5000000980000006300000083",
            INIT_11 => X"000000ab000000670000005d000000500000005d0000007a000000b2000000bf",
            INIT_12 => X"000000960000006400000059000000570000003c0000002e0000002600000018",
            INIT_13 => X"0000002e0000003c0000006c0000009000000090000000800000007f00000078",
            INIT_14 => X"00000075000000c3000000b1000000b2000000b50000008a0000005300000096",
            INIT_15 => X"000000f5000000db000000850000008600000095000000b0000000be000000c2",
            INIT_16 => X"000000a80000007d0000006e0000003d0000002300000022000000310000003a",
            INIT_17 => X"0000003d0000003a00000045000000480000004e000000450000003b00000037",
            INIT_18 => X"0000004f000000af000000ae000000b0000000b10000008c0000006d000000d3",
            INIT_19 => X"000000fd000000fc000000d00000007c000000720000007c000000740000007a",
            INIT_1A => X"0000006800000044000000440000003c00000034000000320000003300000038",
            INIT_1B => X"00000038000000330000002b000000330000003b000000300000002b0000002a",
            INIT_1C => X"000000290000006000000090000000a8000000b2000000a5000000a5000000f6",
            INIT_1D => X"000000fd000000e30000006e0000003c00000035000000310000003100000030",
            INIT_1E => X"0000002d0000002a0000002e0000002a000000260000002e0000002e0000002b",
            INIT_1F => X"0000002a0000002e0000002e000000320000003700000035000000330000002d",
            INIT_20 => X"0000001d0000001d0000003b00000083000000a600000084000000c2000000fe",
            INIT_21 => X"000000f10000008d0000003d0000003200000032000000330000003100000032",
            INIT_22 => X"0000002f0000002a00000027000000220000002300000027000000260000002a",
            INIT_23 => X"0000002d000000380000003e0000003b00000038000000320000002e00000033",
            INIT_24 => X"000000300000001e00000022000000490000008000000080000000d700000100",
            INIT_25 => X"000000bb00000042000000360000003200000034000000340000002e0000002d",
            INIT_26 => X"0000002b00000029000000240000002700000028000000280000002b0000002e",
            INIT_27 => X"0000003b0000003e000000400000003b00000036000000320000004600000053",
            INIT_28 => X"00000034000000230000001f000000290000004200000080000000e0000000f0",
            INIT_29 => X"0000007c0000003a0000003100000038000000360000002c0000002c0000002f",
            INIT_2A => X"0000002e0000002b0000002b0000002c0000002c0000002d000000360000003a",
            INIT_2B => X"000000360000002e0000002b000000240000003300000049000000550000004c",
            INIT_2C => X"00000032000000230000001d000000230000002c0000004e000000ca000000d3",
            INIT_2D => X"000000610000004100000036000000300000003a00000030000000280000002d",
            INIT_2E => X"0000002f000000300000002f0000002e00000033000000270000002700000030",
            INIT_2F => X"0000002f000000270000001c0000002800000043000000430000002e00000033",
            INIT_30 => X"00000032000000230000002000000021000000290000002e00000068000000aa",
            INIT_31 => X"000000400000003600000034000000350000003d0000003a000000360000002d",
            INIT_32 => X"0000002a000000290000002e000000310000002e0000002a0000002800000027",
            INIT_33 => X"00000025000000280000002c0000003f0000002f0000001f0000000f00000033",
            INIT_34 => X"000000440000002a0000001f00000026000000250000002b0000002a00000047",
            INIT_35 => X"000000310000001f0000001b0000002600000031000000380000003a00000035",
            INIT_36 => X"000000380000003c0000003900000035000000320000002d0000002700000021",
            INIT_37 => X"0000002a0000003e0000004f0000004900000038000000260000000d00000028",
            INIT_38 => X"0000003d00000031000000230000002b000000270000002a0000002c00000028",
            INIT_39 => X"0000002a0000001b000000170000001e0000001b0000001d000000240000002f",
            INIT_3A => X"000000380000003e000000420000004b00000045000000310000002b0000002b",
            INIT_3B => X"0000003c000000550000006d0000005d0000003c0000001a0000001d00000014",
            INIT_3C => X"00000036000000380000002d0000002b00000028000000280000002800000026",
            INIT_3D => X"000000240000001a000000160000001d000000190000001d0000001300000012",
            INIT_3E => X"000000200000002f0000003d0000004a0000004200000035000000340000002d",
            INIT_3F => X"0000004300000059000000690000005900000030000000180000002200000015",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY1;


    MEM_IFMAP_LAYER0_ENTITY2 : if BRAM_NAME = "ifmap_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000700000006f0000007400000076000000700000006d0000007300000071",
            INIT_01 => X"0000006f00000071000000740000006f0000006f000000750000007500000077",
            INIT_02 => X"00000075000000710000006f000000700000006d0000006b0000006b0000006a",
            INIT_03 => X"0000006b000000650000006200000061000000610000005f0000005b00000055",
            INIT_04 => X"000000700000006e000000720000007400000070000000710000007500000072",
            INIT_05 => X"000000740000006e0000006f0000006e00000071000000770000007500000073",
            INIT_06 => X"000000730000006f00000070000000730000006e000000680000006600000064",
            INIT_07 => X"00000069000000660000006600000061000000620000005f0000005b00000058",
            INIT_08 => X"0000006e0000006d0000006f0000006f0000006a000000730000007500000075",
            INIT_09 => X"0000007300000073000000720000006d0000006f000000730000007200000071",
            INIT_0A => X"00000074000000720000006f000000600000005a0000004e0000004d00000055",
            INIT_0B => X"0000005600000060000000670000006300000063000000620000005f00000059",
            INIT_0C => X"0000006b0000006e0000006d000000700000006e000000750000007800000077",
            INIT_0D => X"00000073000000750000007b00000092000000820000006f0000007300000072",
            INIT_0E => X"000000700000006f00000050000000570000005a0000005a0000004b0000003f",
            INIT_0F => X"000000460000003e00000055000000620000006600000065000000630000005e",
            INIT_10 => X"0000006b00000072000000730000007200000072000000710000007800000074",
            INIT_11 => X"000000710000007400000080000000d60000009c000000720000006f0000006c",
            INIT_12 => X"000000500000003500000045000000670000006e00000072000000660000005e",
            INIT_13 => X"000000480000004e000000490000005300000060000000650000005e0000005d",
            INIT_14 => X"0000006d00000068000000640000007000000073000000710000007400000073",
            INIT_15 => X"0000006f00000074000000760000008a0000007a000000660000004b00000032",
            INIT_16 => X"0000003a000000380000005300000071000000790000007a0000007400000060",
            INIT_17 => X"000000640000005b0000003a0000003a0000005400000069000000620000005f",
            INIT_18 => X"000000640000005f000000250000004a00000075000000760000007300000076",
            INIT_19 => X"0000007500000074000000780000006b000000620000006c0000005700000043",
            INIT_1A => X"000000530000004b00000054000000820000008e000000760000006300000066",
            INIT_1B => X"0000006f00000053000000470000002f0000003d00000062000000630000005d",
            INIT_1C => X"00000073000000600000002b000000400000006f000000750000007200000074",
            INIT_1D => X"00000077000000710000006d0000005e0000006e000000830000006a00000057",
            INIT_1E => X"0000005f000000580000004d00000076000000990000007c0000005d00000062",
            INIT_1F => X"0000005d000000510000003c000000350000002f000000530000006700000061",
            INIT_20 => X"000000a1000000690000003a000000790000007c00000071000000750000007a",
            INIT_21 => X"000000790000008700000059000000690000008d0000008f0000006f00000050",
            INIT_22 => X"00000051000000550000004e000000470000007d00000087000000670000004f",
            INIT_23 => X"0000004d000000520000004900000039000000230000003b0000006a00000067",
            INIT_24 => X"000000b00000008b000000640000009a00000095000000740000007400000076",
            INIT_25 => X"000000b4000000d6000000b40000008300000099000000830000006e00000055",
            INIT_26 => X"000000540000004a00000039000000440000007d000000850000007c00000062",
            INIT_27 => X"0000005100000055000000550000004c000000310000001e0000004b00000067",
            INIT_28 => X"000000b70000007400000097000000a90000009c000000700000007600000059",
            INIT_29 => X"000000c5000000e0000000bf000000870000009f000000890000006c0000006f",
            INIT_2A => X"0000004c000000500000002c00000055000000a5000000930000009300000064",
            INIT_2B => X"0000005300000066000000580000004f0000003b000000240000002e00000051",
            INIT_2C => X"000000bf0000006c00000090000000af000000a7000000780000007b0000005d",
            INIT_2D => X"0000005f000000b6000000ab0000008e000000a1000000ab000000770000006b",
            INIT_2E => X"00000062000000540000002600000079000000c9000000980000008b00000059",
            INIT_2F => X"000000500000005d00000068000000570000004b000000350000003700000038",
            INIT_30 => X"000000c20000006000000086000000b40000009c0000007b0000007b0000006d",
            INIT_31 => X"000000440000009a0000009000000072000000a6000000ca0000009500000071",
            INIT_32 => X"00000072000000720000003200000093000000bb000000950000007600000058",
            INIT_33 => X"00000053000000540000005f0000005700000057000000490000004a00000037",
            INIT_34 => X"000000c00000005f0000009a000000bc0000006e0000006a0000007c00000074",
            INIT_35 => X"00000048000000840000007d00000095000000ae000000d8000000ac00000083",
            INIT_36 => X"00000075000000720000004700000098000000b5000000900000006e00000055",
            INIT_37 => X"0000005000000049000000500000006400000065000000580000005900000049",
            INIT_38 => X"000000c40000006b000000a7000000ba0000006d00000059000000770000007a",
            INIT_39 => X"0000004a0000006a0000007b000000b9000000b4000000a50000008c0000008f",
            INIT_3A => X"00000088000000640000004700000098000000af00000085000000800000006d",
            INIT_3B => X"000000560000005d000000600000006e0000007400000060000000550000005f",
            INIT_3C => X"000000c500000081000000a7000000b20000008900000053000000780000007d",
            INIT_3D => X"0000005e0000007800000083000000dd000000ec0000008a0000008200000079",
            INIT_3E => X"000000700000006800000058000000860000009f000000930000006c00000055",
            INIT_3F => X"0000004800000058000000680000006d0000006e000000560000006000000068",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY2;


    MEM_IFMAP_LAYER0_ENTITY3 : if BRAM_NAME = "ifmap_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cb00000092000000a4000000b6000000aa000000560000007d0000007e",
            INIT_01 => X"00000079000000500000008f000000a300000098000000840000006a0000006a",
            INIT_02 => X"00000065000000650000005a0000008f0000008a0000008d0000008200000069",
            INIT_03 => X"0000004c0000004f0000005d0000005b00000053000000580000006c00000068",
            INIT_04 => X"000000d7000000a6000000a7000000b8000000b6000000660000006000000095",
            INIT_05 => X"000000890000005d000000740000006900000066000000690000005b0000006e",
            INIT_06 => X"0000005b00000067000000800000006000000038000000780000007e00000045",
            INIT_07 => X"0000003800000038000000460000005d0000005e00000070000000740000006e",
            INIT_08 => X"000000d3000000b8000000af000000b5000000b800000083000000580000008b",
            INIT_09 => X"00000094000000800000005a00000040000000790000006f000000750000008f",
            INIT_0A => X"0000005c000000600000008b000000750000006d00000063000000440000003b",
            INIT_0B => X"000000290000003e00000045000000690000007700000078000000730000006f",
            INIT_0C => X"000000c0000000bd000000b0000000b3000000b6000000950000005a00000079",
            INIT_0D => X"0000007c00000088000000860000003b000000760000006100000086000000b0",
            INIT_0E => X"000000760000004b000000770000007c00000081000000560000003100000033",
            INIT_0F => X"000000310000005a0000005b0000007600000079000000710000006f0000006b",
            INIT_10 => X"0000009c000000c1000000b2000000ad000000b50000009d0000006700000087",
            INIT_11 => X"000000af000000690000005a0000004d0000005a00000076000000ad000000b6",
            INIT_12 => X"00000094000000640000004e0000004d0000003d000000340000002e00000021",
            INIT_13 => X"0000003900000047000000640000007d0000007b0000006d0000007100000069",
            INIT_14 => X"00000078000000c8000000b2000000a9000000b3000000900000005700000099",
            INIT_15 => X"000000f7000000de0000008c0000008d0000009c000000b6000000c4000000c0",
            INIT_16 => X"000000ac000000850000006d0000003e00000031000000360000004600000051",
            INIT_17 => X"0000005500000054000000630000006500000068000000600000005c0000005a",
            INIT_18 => X"00000069000000c5000000b7000000ac000000b10000009200000070000000d3",
            INIT_19 => X"000000fc000000fd000000e00000008f000000840000008d0000008500000085",
            INIT_1A => X"0000007c0000005d00000057000000520000005400000054000000550000005d",
            INIT_1B => X"0000005e0000005b00000060000000680000006c00000061000000610000005f",
            INIT_1C => X"0000005900000089000000a8000000ae000000b6000000aa000000a6000000f5",
            INIT_1D => X"000000fb000000e70000008800000058000000500000004c0000004b00000048",
            INIT_1E => X"0000004f000000510000005100000052000000560000005a0000005900000057",
            INIT_1F => X"000000590000005d0000005e00000060000000600000005e0000005f0000005a",
            INIT_20 => X"0000005b000000570000006600000099000000b300000088000000bd000000fa",
            INIT_21 => X"000000f50000009f0000005e0000005400000054000000550000005300000054",
            INIT_22 => X"0000005600000054000000520000004f00000053000000560000005500000059",
            INIT_23 => X"0000005c00000067000000670000006500000066000000630000005e00000067",
            INIT_24 => X"0000006f0000005e000000550000006a0000009400000088000000d5000000fd",
            INIT_25 => X"000000c60000005d0000005b000000580000005a0000005a0000005300000052",
            INIT_26 => X"0000005200000051000000500000005300000056000000590000005c0000005f",
            INIT_27 => X"0000006c0000006e0000006d0000006c0000006c000000690000007b00000089",
            INIT_28 => X"000000720000006300000056000000530000005f00000091000000e5000000f5",
            INIT_29 => X"0000008f0000005c000000570000005e0000005c000000520000005200000053",
            INIT_2A => X"000000540000005300000056000000580000005a000000610000006a0000006e",
            INIT_2B => X"00000069000000610000005f0000005b0000006c000000820000008a0000007d",
            INIT_2C => X"0000006e000000620000005900000056000000530000006a000000db000000e4",
            INIT_2D => X"0000007e000000680000005e0000005700000061000000570000005000000052",
            INIT_2E => X"00000054000000570000005900000059000000610000005c0000005d00000066",
            INIT_2F => X"000000650000005d0000005500000065000000810000007e0000006200000060",
            INIT_30 => X"0000006c000000610000005c00000058000000580000005400000085000000c5",
            INIT_31 => X"00000064000000610000005e0000005f00000067000000640000006000000053",
            INIT_32 => X"0000004f00000050000000580000005c0000005c0000005f0000005d0000005c",
            INIT_33 => X"0000005a0000005d000000660000007d0000006e0000005a0000003c0000005d",
            INIT_34 => X"0000007c00000064000000580000005b00000057000000590000004f0000006b",
            INIT_35 => X"000000590000004d00000047000000520000005d00000064000000660000005c",
            INIT_36 => X"0000005e0000006300000063000000610000005f0000005e0000005800000053",
            INIT_37 => X"0000005b00000070000000840000008300000074000000610000004000000055",
            INIT_38 => X"0000007400000066000000550000005b0000005a0000005c0000005800000051",
            INIT_39 => X"0000005500000048000000430000004a00000047000000490000005000000056",
            INIT_3A => X"0000005f000000650000006d00000077000000710000005f0000005800000058",
            INIT_3B => X"00000069000000820000009c0000009100000073000000520000005200000040",
            INIT_3C => X"0000006b000000690000005900000056000000590000005c0000005700000051",
            INIT_3D => X"0000004f00000045000000420000004900000045000000490000003f0000003a",
            INIT_3E => X"000000460000005700000068000000770000006f000000600000005f00000057",
            INIT_3F => X"0000006d000000830000009200000087000000630000004d0000005400000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY3;


    MEM_IFMAP_LAYER0_ENTITY4 : if BRAM_NAME = "ifmap_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000310000002f00000033000000350000002e000000290000002f0000002d",
            INIT_01 => X"0000002c00000029000000290000003400000031000000290000002d0000002c",
            INIT_02 => X"0000002800000026000000270000002b0000002c0000002d0000002d0000002b",
            INIT_03 => X"0000002c000000270000002b0000002900000026000000240000002400000021",
            INIT_04 => X"00000033000000280000002d00000038000000310000002b0000002f0000002d",
            INIT_05 => X"0000002e00000026000000290000003600000034000000290000002800000021",
            INIT_06 => X"0000001e00000021000000290000003200000035000000370000003400000030",
            INIT_07 => X"000000320000002e0000002d00000026000000220000001f0000002000000022",
            INIT_08 => X"0000002f0000002100000024000000300000002a0000002c0000002d0000002d",
            INIT_09 => X"0000002b0000002b000000300000003900000033000000260000002500000023",
            INIT_0A => X"000000270000002f000000360000003100000034000000320000002f00000032",
            INIT_0B => X"0000003000000037000000330000002700000023000000220000002200000021",
            INIT_0C => X"00000028000000200000001f0000002c0000002b0000002e0000003000000030",
            INIT_0D => X"0000002c0000002d000000390000005f0000004b000000290000002f00000036",
            INIT_0E => X"0000003a000000430000002f000000410000004c000000540000004200000032",
            INIT_0F => X"00000034000000270000002d0000002e0000002b000000270000002700000024",
            INIT_10 => X"0000002900000030000000310000002f0000002b000000280000002f0000002c",
            INIT_11 => X"000000290000002a0000003b000000a40000006b000000380000003c00000047",
            INIT_12 => X"000000320000001f00000038000000620000006f00000076000000690000005d",
            INIT_13 => X"00000043000000460000002f0000002d000000300000002e0000002400000024",
            INIT_14 => X"000000360000004000000039000000350000002c000000270000002900000029",
            INIT_15 => X"00000025000000270000002a000000550000004e0000003a0000002b0000001f",
            INIT_16 => X"0000002b0000002d0000004c0000006e000000780000007a0000007400000060",
            INIT_17 => X"00000061000000560000002f00000025000000310000003a0000002c00000028",
            INIT_18 => X"0000003900000050000000110000001c000000300000002b000000280000002b",
            INIT_19 => X"0000002a0000002500000027000000340000003b0000004b0000004600000039",
            INIT_1A => X"00000048000000400000004a00000079000000840000006c0000005a0000005e",
            INIT_1B => X"000000670000004d0000004500000027000000240000003a0000003000000027",
            INIT_1C => X"0000005a0000005c0000002600000029000000380000002a0000002400000027",
            INIT_1D => X"000000310000003300000033000000310000004d0000006b0000005d0000004f",
            INIT_1E => X"0000005800000052000000450000006b0000008c000000700000005100000058",
            INIT_1F => X"000000540000004a0000003a0000003100000020000000320000003300000027",
            INIT_20 => X"00000090000000690000003b00000071000000520000002b0000002900000032",
            INIT_21 => X"000000420000005f0000003b0000004e0000007900000080000000650000004a",
            INIT_22 => X"0000004d00000052000000490000003d000000700000007b0000005d00000046",
            INIT_23 => X"000000450000004c00000043000000350000001b000000230000003b0000002d",
            INIT_24 => X"000000a30000008f000000690000009500000070000000330000002f0000003c",
            INIT_25 => X"00000092000000c6000000a600000077000000910000007d0000006b0000004f",
            INIT_26 => X"0000004f00000047000000350000003a000000700000007a0000007200000059",
            INIT_27 => X"0000004a0000004e0000004e000000470000002b0000000f0000002c00000039",
            INIT_28 => X"000000af0000007a0000009e000000a80000007a00000032000000330000002f",
            INIT_29 => X"000000b3000000e2000000bc000000830000009b000000840000006800000068",
            INIT_2A => X"000000450000004d000000280000004d0000009a000000890000008a0000005c",
            INIT_2B => X"0000004d000000600000004f000000490000003b000000210000001f0000002e",
            INIT_2C => X"000000bd0000007400000099000000b2000000880000003b000000370000002c",
            INIT_2D => X"00000050000000bc000000a400000085000000970000009f0000006a0000005f",
            INIT_2E => X"000000590000004f0000002200000071000000c00000008e0000008200000052",
            INIT_2F => X"0000004b000000580000005e000000510000004e00000037000000300000001a",
            INIT_30 => X"000000c20000006900000090000000b90000008500000044000000350000002f",
            INIT_31 => X"0000002c000000980000007e0000005e00000094000000b70000008100000062",
            INIT_32 => X"000000690000006d0000002f0000008c000000b20000008c0000006f00000053",
            INIT_33 => X"0000004f00000050000000550000005100000059000000490000004000000018",
            INIT_34 => X"000000c100000067000000a3000000c000000062000000420000003a00000032",
            INIT_35 => X"0000002700000078000000670000007f0000009b000000c80000009d00000075",
            INIT_36 => X"0000006b0000006d0000004400000093000000ae000000880000006800000050",
            INIT_37 => X"0000004c00000046000000480000005e00000063000000510000004500000022",
            INIT_38 => X"000000c400000070000000ac000000bc0000006d000000430000003e00000037",
            INIT_39 => X"000000220000005800000067000000a9000000a90000009f0000008c00000086",
            INIT_3A => X"0000007d0000005f0000004600000095000000aa0000007f0000007a00000069",
            INIT_3B => X"000000530000005b0000005a000000680000006f00000050000000350000002f",
            INIT_3C => X"000000c500000088000000ae000000b50000008e0000004d000000580000004d",
            INIT_3D => X"000000340000005d00000074000000d3000000e6000000890000008200000070",
            INIT_3E => X"000000650000005f0000004b00000076000000920000008a0000006500000050",
            INIT_3F => X"000000440000005700000063000000630000005d000000360000003000000030",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY4;


    MEM_IFMAP_LAYER0_ENTITY5 : if BRAM_NAME = "ifmap_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cc000000a0000000b2000000bc000000ac0000005a0000007e00000071",
            INIT_01 => X"0000005200000025000000850000009b0000008d00000075000000580000005a",
            INIT_02 => X"0000005c000000570000003a000000680000006d0000007e0000007600000061",
            INIT_03 => X"000000480000004d0000005e00000052000000370000002d000000370000002e",
            INIT_04 => X"000000d7000000b4000000b8000000c2000000ba000000690000006600000091",
            INIT_05 => X"0000006f0000003d000000690000005f00000059000000590000004900000062",
            INIT_06 => X"000000580000005f00000066000000400000002000000069000000730000003d",
            INIT_07 => X"0000003300000035000000410000004e00000040000000440000004000000036",
            INIT_08 => X"000000cd000000c0000000bd000000c1000000bc00000085000000600000008f",
            INIT_09 => X"0000008d0000006f00000050000000370000006c000000600000006400000085",
            INIT_0A => X"0000005d0000005d000000780000005d0000005c000000560000003a00000034",
            INIT_0B => X"000000270000003c000000280000003b0000003e000000360000002d0000002e",
            INIT_0C => X"000000b4000000bb000000b5000000b9000000b8000000980000006300000084",
            INIT_0D => X"00000082000000870000007e000000330000006c000000560000007b000000a8",
            INIT_0E => X"00000076000000490000006700000069000000760000004e0000002c00000032",
            INIT_0F => X"000000340000005d0000003c000000440000004000000034000000320000002e",
            INIT_10 => X"00000092000000bb000000af000000ac000000b4000000a00000006f00000092",
            INIT_11 => X"000000b90000006f00000057000000490000005600000074000000ad000000b1",
            INIT_12 => X"0000009400000065000000420000003f00000039000000360000003300000029",
            INIT_13 => X"00000045000000530000004b000000520000004c0000003d000000450000003f",
            INIT_14 => X"0000007c000000c8000000b0000000a8000000b3000000930000005b0000009f",
            INIT_15 => X"000000fa000000e10000009000000093000000a4000000c0000000d0000000c5",
            INIT_16 => X"000000b50000008f0000006d0000003e0000003a000000440000005700000066",
            INIT_17 => X"0000006e0000006f0000007a0000007700000078000000700000007000000073",
            INIT_18 => X"00000085000000d5000000c0000000b1000000b60000009600000071000000d1",
            INIT_19 => X"000000f7000000fc000000e80000009d00000095000000a20000009c00000098",
            INIT_1A => X"000000940000007700000068000000650000006f0000006e000000730000007d",
            INIT_1B => X"0000008300000082000000870000008d0000008e000000840000008900000084",
            INIT_1C => X"00000087000000a8000000bc000000bc000000c0000000ae000000a4000000ed",
            INIT_1D => X"000000f1000000e4000000990000006f00000069000000690000006b00000065",
            INIT_1E => X"000000730000007800000071000000740000007d0000007d0000007e00000080",
            INIT_1F => X"000000840000008b000000890000008900000087000000860000008b00000085",
            INIT_20 => X"0000008d0000008200000086000000b0000000bf00000089000000b5000000f2",
            INIT_21 => X"000000f5000000af0000007f0000007600000077000000790000007800000074",
            INIT_22 => X"00000075000000750000007300000071000000780000007d0000007d00000082",
            INIT_23 => X"00000086000000910000008e0000008e00000092000000900000008c00000095",
            INIT_24 => X"000000a20000008c0000007c00000088000000a70000008f000000d1000000f9",
            INIT_25 => X"000000cd00000076000000800000007d0000007f0000007f0000007900000073",
            INIT_26 => X"000000710000007000000071000000750000007b00000083000000860000008a",
            INIT_27 => X"000000960000009800000093000000950000009a00000098000000a7000000b6",
            INIT_28 => X"000000a500000093000000820000007a0000007e000000a4000000ea000000f7",
            INIT_29 => X"00000099000000720000007b0000008300000081000000770000007700000077",
            INIT_2A => X"00000077000000770000007b0000007f000000830000008d000000960000009a",
            INIT_2B => X"000000960000008d0000008c0000008a0000009e000000b2000000b6000000a9",
            INIT_2C => X"000000a2000000950000008a000000850000007e0000008a000000e9000000ea",
            INIT_2D => X"0000008c0000007e000000810000007c000000850000007b0000007400000077",
            INIT_2E => X"0000007a0000007e00000082000000840000008c0000008a0000008b00000094",
            INIT_2F => X"000000930000008b0000008500000099000000b6000000b00000008e0000008b",
            INIT_30 => X"000000a1000000930000008f0000008d0000008a0000007d0000009f000000d3",
            INIT_31 => X"000000770000007900000080000000820000008b000000870000008300000078",
            INIT_32 => X"00000076000000780000008200000087000000880000008b0000008a00000088",
            INIT_33 => X"000000870000008a00000097000000b2000000a40000008c0000006700000088",
            INIT_34 => X"000000b10000009400000089000000920000008b000000840000007100000085",
            INIT_35 => X"0000007200000069000000690000007500000080000000870000008900000080",
            INIT_36 => X"00000083000000890000008b0000008a0000008900000088000000830000007d",
            INIT_37 => X"000000850000009a000000b3000000b5000000a8000000920000006c0000007f",
            INIT_38 => X"000000a800000094000000840000008f0000008b000000860000007d00000070",
            INIT_39 => X"0000007300000068000000660000006d0000006a0000006c0000007300000078",
            INIT_3A => X"0000008000000087000000900000009c00000098000000860000007f0000007f",
            INIT_3B => X"00000090000000aa000000c5000000be000000a4000000820000007e0000006b",
            INIT_3C => X"000000a000000095000000840000008600000086000000840000007b00000073",
            INIT_3D => X"0000007200000069000000650000006c000000680000006c0000006200000059",
            INIT_3E => X"000000640000007600000089000000980000009100000083000000820000007b",
            INIT_3F => X"00000091000000a7000000b6000000af000000910000007c000000810000006e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY5;


    MEM_GOLD_LAYER0_ENTITY0 : if BRAM_NAME = "gold_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000012000000120000000f00000014000000170000000d0000000f0000001d",
            INIT_01 => X"0000001d0000000a0000000000000001000000060000000c0000001500000016",
            INIT_02 => X"000000120000000f000000130000001300000004000000080000000300000000",
            INIT_03 => X"00000004000000000000000000000000000000050000000b000000000000000b",
            INIT_04 => X"000000130000001b000000120000001b000000200000001e0000000000000000",
            INIT_05 => X"000000000000000000000000000000000000000100000001000000000000000c",
            INIT_06 => X"000000190000000b000000110000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000300000003",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000040000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0B => X"00000000000000000000000000000000000000040000001c0000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0E => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_10 => X"0000000000000000000000000000000b00000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000080000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_2C => X"0000000000000000000000000000000000000004000000070000000000000000",
            INIT_2D => X"0000000000000000000000000000000600000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000f0000001a0000000f0000003f0000000a",
            INIT_31 => X"000000000000000000000000000000320000003a000000380000002500000020",
            INIT_32 => X"00000022000000290000002500000027000000200000002c0000003a00000000",
            INIT_33 => X"000000000000001e0000001d0000001d00000020000000200000001f00000024",
            INIT_34 => X"0000001e000000220000002800000021000000300000002f0000002f0000000e",
            INIT_35 => X"0000000f00000021000000190000001d00000022000000230000002f00000033",
            INIT_36 => X"00000034000000280000003a000000290000003300000031000000410000002a",
            INIT_37 => X"000000300000002a0000001f000000170000001c000000210000002d0000001a",
            INIT_38 => X"0000001c00000029000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000003000000180000000e0000000600000000000000000000000000000000",
            INIT_3E => X"0000000b00000000000000000000000000000000000000020000000100000000",
            INIT_3F => X"0000001b0000000000000006000000000000000000000000000000000000001e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY0;


    MEM_GOLD_LAYER0_ENTITY1 : if BRAM_NAME = "gold_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000011000000140000000500000003000000000000001d",
            INIT_01 => X"00000010000000000000000800000000000000030000000f0000001700000000",
            INIT_02 => X"000000000000001a0000000a0000000600000004000000000000004400000003",
            INIT_03 => X"000000000000000b0000000000000002000000170000000b0000000000000000",
            INIT_04 => X"0000000c0000001e0000000b0000000000000000000000370000000000000004",
            INIT_05 => X"0000000a00000011000000020000002000000014000000060000000000000006",
            INIT_06 => X"0000002d00000000000000000000000000000020000000000000000000000011",
            INIT_07 => X"00000008000000000000001d0000002800000004000000110000000800000000",
            INIT_08 => X"000000000000000b0000000b0000000000000010000000000000000600000000",
            INIT_09 => X"00000000000000180000002400000000000000270000000e0000000900000012",
            INIT_0A => X"00000012000000150000000000000000000000000000000c0000000000000000",
            INIT_0B => X"0000002b0000002300000000000000580000000d000000280000002d00000011",
            INIT_0C => X"00000000000000000000001b000000220000001f0000000b0000000000000036",
            INIT_0D => X"00000023000000120000004500000000000000070000001f000000210000001a",
            INIT_0E => X"0000001e00000022000000280000002e0000002f0000002f0000002a00000038",
            INIT_0F => X"000000330000002500000000000000270000002500000024000000240000002a",
            INIT_10 => X"0000002f000000360000002f0000002e0000003a0000002c0000002e00000052",
            INIT_11 => X"00000000000000130000002b000000260000002a0000002a0000002f0000002e",
            INIT_12 => X"0000002f0000002a00000045000000280000002b000000330000002c00000019",
            INIT_13 => X"000000190000002800000023000000240000002e000000310000002d0000002e",
            INIT_14 => X"000000430000003a0000001f0000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000000000000020000000a0000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000100000000800000017000000000000001f0000001c0000000300000000",
            INIT_18 => X"000000000000002a00000000000000000000000000000000000000000000002b",
            INIT_19 => X"000000110000000000000000000000420000002d0000003f0000000000000000",
            INIT_1A => X"000000710000000000000000000000000000000e00000000000000280000002c",
            INIT_1B => X"00000025000000000000005a000000260000003b0000002a000000000000006c",
            INIT_1C => X"00000005000000230000000000000034000000240000005d000000480000003c",
            INIT_1D => X"000000000000002f000000520000001e0000003e000000000000005900000031",
            INIT_1E => X"0000003700000000000000000000002c000000610000003e0000006000000000",
            INIT_1F => X"000000730000005c000000120000003100000025000000480000007300000015",
            INIT_20 => X"0000003800000000000000000000005a0000004a0000006a0000000000000075",
            INIT_21 => X"00000047000000120000000c000000370000004d000000650000002800000031",
            INIT_22 => X"00000000000000060000008b0000003800000046000000000000004f00000050",
            INIT_23 => X"0000000600000025000000130000006800000042000000840000000b0000002a",
            INIT_24 => X"000000130000002e0000002c0000000000000029000000160000005b00000004",
            INIT_25 => X"00000000000000000000004a0000003a0000009f000000000000006400000018",
            INIT_26 => X"000000000000004d000000300000003b0000005a000000170000000000000000",
            INIT_27 => X"0000000c0000000f0000003c0000009400000000000000930000004c00000020",
            INIT_28 => X"0000007100000083000000410000001a0000001d000000230000002000000031",
            INIT_29 => X"0000001d0000002b0000004e00000000000000d8000000730000003a0000003c",
            INIT_2A => X"00000047000000380000003d0000003c0000003e000000400000004f0000005f",
            INIT_2B => X"000000120000000000000082000000af00000042000000490000003f0000003e",
            INIT_2C => X"00000039000000380000004000000050000000480000003d0000006a00000045",
            INIT_2D => X"00000000000000cb0000005a000000390000004d000000420000003c00000041",
            INIT_2E => X"000000480000004d0000004e000000380000007b000000760000004b0000003e",
            INIT_2F => X"0000005400000048000000350000004300000044000000380000004400000055",
            INIT_30 => X"0000003a0000001a0000006f0000008000000000000000000000000800000008",
            INIT_31 => X"0000000600000003000000050000000000000004000000000000000000000000",
            INIT_32 => X"000000000000000600000005000000070000000a0000000c000000070000000a",
            INIT_33 => X"000000490000001a000000000000000000000000000000240000000600000000",
            INIT_34 => X"0000000000000004000000000000000000000004000000040000000700000000",
            INIT_35 => X"00000000000000000000000d0000001a00000015000000070000001700000000",
            INIT_36 => X"00000000000000280000002500000009000000050000000d0000000000000037",
            INIT_37 => X"0000001b00000005000000000000000000000000000000000000000100000000",
            INIT_38 => X"000000260000005a000000130000000b0000008000000056000000060000000e",
            INIT_39 => X"000000000000000000000025000000250000000f000000180000000000000000",
            INIT_3A => X"00000000000000080000000000000000000000000000002a0000001a0000001f",
            INIT_3B => X"0000003a00000000000000000000000000000009000000270000000600000007",
            INIT_3C => X"00000000000000040000000000000021000000000000000a0000000900000011",
            INIT_3D => X"000000000000000b00000000000000170000001d00000015000000070000001c",
            INIT_3E => X"0000001000000019000000160000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000010000000040000000b00000004",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY1;


    MEM_GOLD_LAYER0_ENTITY2 : if BRAM_NAME = "gold_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000000000000000001a00000004000000000000000000000000",
            INIT_01 => X"00000000000000030000002f0000000000000000000000090000000400000011",
            INIT_02 => X"00000000000000000000004a0000000c0000000000000000000000000000001b",
            INIT_03 => X"0000001f00000000000000000000000000000000000000460000009c00000085",
            INIT_04 => X"0000002800000000000000000000000000000020000000410000001b00000000",
            INIT_05 => X"0000000000000000000000000000000f00000046000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000004000000070000001200000000000000000000001100000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000080000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001400000013",
            INIT_0C => X"00000004000000000000002800000022000000000000009d000000a3000000a2",
            INIT_0D => X"000000a5000000a40000009d000000ac000000b7000000ad000000940000007c",
            INIT_0E => X"0000007c000000840000009200000092000000a2000000ad000000a8000000ac",
            INIT_0F => X"000000a00000008c000000a9000000a00000007a0000003a0000002e0000003e",
            INIT_10 => X"0000004e0000006e0000008b000000890000006a000000ac000000b0000000af",
            INIT_11 => X"0000008e00000073000000480000002d000000070000001e0000000a00000027",
            INIT_12 => X"0000003a000000670000004d0000002b000000a4000000aa000000a200000059",
            INIT_13 => X"0000004d00000027000000150000000c000000330000002d0000001b00000025",
            INIT_14 => X"0000003a000000170000001f00000094000000600000004e0000004700000043",
            INIT_15 => X"0000002f0000001f000000000000003100000039000000170000001c0000002f",
            INIT_16 => X"00000016000000120000008e00000099000000250000003b0000004500000031",
            INIT_17 => X"0000002d000000000000003e0000002a0000001000000012000000170000000e",
            INIT_18 => X"0000002a000000620000009f0000002f000000320000003e0000002d0000002f",
            INIT_19 => X"000000000000003200000028000000100000000e000000260000001c0000000a",
            INIT_1A => X"0000002c0000006200000037000000260000002e00000027000000290000001e",
            INIT_1B => X"0000002f0000002d00000009000000220000004100000014000000000000002b",
            INIT_1C => X"0000000e000000550000002200000036000000300000000d0000005400000042",
            INIT_1D => X"000000260000000f0000002d0000007900000010000000050000002400000000",
            INIT_1E => X"000000350000002000000008000000280000002d000000340000001d00000006",
            INIT_1F => X"00000009000000620000008a0000000000000015000000230000000000000017",
            INIT_20 => X"0000001a00000000000000000000000600000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000060000003a00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000002200000023",
            INIT_29 => X"00000025000000200000001e0000002700000026000000240000001d00000017",
            INIT_2A => X"0000001a00000026000000240000001e00000018000000230000002c0000002a",
            INIT_2B => X"0000001f00000028000000200000000f0000001d0000000e0000001d00000000",
            INIT_2C => X"00000009000000200000002b0000001c00000006000000390000002800000021",
            INIT_2D => X"000000270000001a0000000000000006000000210000002e0000000000000000",
            INIT_2E => X"00000000000000250000002c000000000000004c00000021000000290000000f",
            INIT_2F => X"0000002400000004000000000000000000000048000000000000000900000000",
            INIT_30 => X"000000000000004a00000000000000260000000200000056000000090000000b",
            INIT_31 => X"0000000000000000000000000000005900000000000000000000000600000000",
            INIT_32 => X"0000002b000000000000000a000000000000001a0000003e0000001300000000",
            INIT_33 => X"00000000000000000000008e0000000000000000000000140000000000000000",
            INIT_34 => X"000000000000000000000020000000000000003f000000360000000000000000",
            INIT_35 => X"000000000000006600000000000000000000000a000000150000000000000000",
            INIT_36 => X"0000000000000000000000000000003800000042000000000000000000000000",
            INIT_37 => X"0000004200000000000000000000001d0000000f000000080000000000000002",
            INIT_38 => X"0000000000000021000000040000001100000000000000000000002400000000",
            INIT_39 => X"00000025000000000000001e0000002100000023000000000000000000000000",
            INIT_3A => X"0000002c000000000000000f0000002700000000000000020000000500000000",
            INIT_3B => X"0000000c0000003000000034000000140000002a000000040000000000000078",
            INIT_3C => X"0000000000000000000000220000000000000000000000000000000800000009",
            INIT_3D => X"0000000100000000000000000000002000000014000000000000004000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000002100000043000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY3 : if BRAM_NAME = "gold_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000005d00000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000400000000000000000000002b",
            INIT_05 => X"000000300000002d0000002c0000002f00000029000000300000003a00000037",
            INIT_06 => X"0000002a0000002500000026000000270000002a000000310000002c00000035",
            INIT_07 => X"000000300000002e0000002d000000000000001f000000290000003b0000000c",
            INIT_08 => X"00000000000000000000000e0000001f000000250000001c000000290000002e",
            INIT_09 => X"00000035000000320000003b0000002d00000023000000000000000000000000",
            INIT_0A => X"0000000000000000000000040000001a00000000000000000000002300000032",
            INIT_0B => X"0000002500000019000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000600000000000000110000000000000000000000120000001800000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000000000000500000000000000000000000b000000380000000300000003",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000070000003a000000070000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_14 => X"000000000000000000000000000000000000001a000000050000000000000000",
            INIT_15 => X"0000000f00000003000000180000000400000000000000080000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000008",
            INIT_17 => X"000000110000000a00000000000000000000001f000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000a000000110000000800000008000000040000000c0000000c0000000b",
            INIT_22 => X"0000000b000000210000002d0000002300000011000000080000000600000000",
            INIT_23 => X"0000000a0000000a0000000c0000000800000000000000050000002300000042",
            INIT_24 => X"0000000000000000000000000000000a000000170000000a0000003500000033",
            INIT_25 => X"0000000500000008000000050000003700000016000000090000000000000000",
            INIT_26 => X"0000000000000000000000000000000e0000000c000000000000000000000005",
            INIT_27 => X"0000000800000008000000000000000000000002000000000000001a00000004",
            INIT_28 => X"0000001000000006000000000000000e0000000100000000000000020000000e",
            INIT_29 => X"0000000000000000000000090000000000000007000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000f0000000000000006000000030000003e",
            INIT_2B => X"0000002800000000000000000000000000000000000000140000001500000007",
            INIT_2C => X"000000000000000000000000000000000000001c000000180000001200000000",
            INIT_2D => X"0000003100000000000000110000000000000011000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000020000003500000035",
            INIT_2F => X"000000210000000e000000000000000900000000000000050000000e00000000",
            INIT_30 => X"0000000000000001000000000000000000000000000000260000000000000000",
            INIT_31 => X"000000000000000000000026000000300000000000000000000000000000000c",
            INIT_32 => X"0000000000000004000000000000002300000009000000000000000000000000",
            INIT_33 => X"0000004e00000036000000110000000000000000000000180000000300000000",
            INIT_34 => X"000000070000000000000000000000000000001e000000510000003700000000",
            INIT_35 => X"000000000000000000000000000000050000000a00000035000000210000000c",
            INIT_36 => X"0000000000000056000000280000000400000005000000030000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000160000000000000018",
            INIT_38 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000180000004f0000000b",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000014000000000000000000000000000000220000000000000003",
            INIT_3C => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000d000000130000000a0000000e000000090000001500000008",
            INIT_3E => X"000000060000000c0000001c000000220000001b000000130000000600000002",
            INIT_3F => X"000000080000000b000000090000000d0000000f000000360000000f0000001a",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY3;


    MEM_GOLD_LAYER0_ENTITY4 : if BRAM_NAME = "gold_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f000000340000003500000024000000210000001a0000000a00000026",
            INIT_01 => X"000000240000000b0000000a0000000800000051000000330000002800000020",
            INIT_02 => X"000000530000005e0000004b0000002b000000190000001a0000003300000014",
            INIT_03 => X"0000000e00000012000000190000002e000000450000002f000000360000005b",
            INIT_04 => X"0000005d000000420000003b000000150000001b000000710000005e00000015",
            INIT_05 => X"000000350000007e00000044000000640000003b000000330000003b00000067",
            INIT_06 => X"000000380000003900000025000000010000007f0000009e0000002800000013",
            INIT_07 => X"000000bd0000007e0000007d0000004b0000002e0000005b0000007f00000050",
            INIT_08 => X"000000470000003c000000150000007a0000009400000043000000170000005a",
            INIT_09 => X"00000075000000a8000000650000004e0000007800000081000000460000003b",
            INIT_0A => X"0000004c000000330000008e000000a5000000400000003900000039000000a5",
            INIT_0B => X"000000850000006a000000500000005f000000780000004c000000480000004b",
            INIT_0C => X"00000026000000b0000000b80000006600000073000000380000006600000059",
            INIT_0D => X"0000004e000000510000003300000065000000410000002c0000002b0000000e",
            INIT_0E => X"000000c0000000b300000086000000750000006f000000330000005f00000079",
            INIT_0F => X"000000420000005a00000040000000250000002f0000002700000027000000c7",
            INIT_10 => X"000000ab0000008b000000a20000009e0000006500000091000000b900000079",
            INIT_11 => X"0000003c00000040000000470000005a0000007100000068000000c1000000cb",
            INIT_12 => X"0000009d000000c9000000e7000000a50000008a000000850000007c0000006f",
            INIT_13 => X"0000007800000080000000880000008a0000008e0000008c000000a1000000b1",
            INIT_14 => X"000000e5000000af0000007a0000007500000070000000710000007600000084",
            INIT_15 => X"0000008c000000950000009a000000a30000009d00000085000000a6000000ef",
            INIT_16 => X"0000008800000080000000790000007300000077000000820000008c0000009b",
            INIT_17 => X"00000093000000a3000000ab000000970000008f0000007f000000a700000074",
            INIT_18 => X"0000007f000000890000007e0000007c0000008800000086000000850000009a",
            INIT_19 => X"000000af0000008d000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000130000001c0000000b0000000000000000",
            INIT_1B => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_1C => X"00000014000000330000000000000000000000140000001e0000000000000000",
            INIT_1D => X"0000003f000000000000000000000000000000000000003e0000001c00000028",
            INIT_1E => X"00000000000000000000000000000000000000070000001e0000000000000019",
            INIT_1F => X"0000000000000000000000000000000c00000000000000000000000000000000",
            INIT_20 => X"00000000000000000000001a000000060000000e000000000000000000000000",
            INIT_21 => X"000000090000000000000000000000000000000f000000040000001d00000000",
            INIT_22 => X"00000000000000080000000000000000000000250000002f0000000000000002",
            INIT_23 => X"0000004f00000003000000000000000000000000000000060000000000000026",
            INIT_24 => X"0000001c00000000000000000000000000000000000000180000000d0000000d",
            INIT_25 => X"0000000000000000000000050000000000000009000000000000001800000008",
            INIT_26 => X"0000000000000000000000000000000200000000000000070000000000000000",
            INIT_27 => X"000000000000003d0000001e0000000000000000000000000000001c00000000",
            INIT_28 => X"000000100000000000000000000000000000002e000000000000002200000032",
            INIT_29 => X"00000003000000000000000000000036000000260000003a0000000d00000000",
            INIT_2A => X"0000000000000000000000000000000a00000000000000120000001500000000",
            INIT_2B => X"000000000000002e0000001f0000003100000001000000000000000000000008",
            INIT_2C => X"0000000000000000000000220000000000000000000000000000000000000019",
            INIT_2D => X"0000000f0000000d000000000000000000000000000000160000002100000041",
            INIT_2E => X"000000000000000000000000000000a2000000520000003f000000370000000c",
            INIT_2F => X"0000000600000000000000020000000000000000000000000000000d00000036",
            INIT_30 => X"0000000000000041000000560000000000000002000000000000000000000000",
            INIT_31 => X"0000000000000000000000030000000000000000000000020000000000000025",
            INIT_32 => X"0000003e00000006000000000000000000000001000000000000000000000007",
            INIT_33 => X"0000000a0000000000000000000000420000000c000000000000001800000036",
            INIT_34 => X"0000002400000013000000090000000000000000000000000000000500000000",
            INIT_35 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000040000001f0000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000050000002d000000000000000700000000000000020000000100000000",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000002",
            INIT_3E => X"0000003b00000000000000000000000300000000000000100000000100000006",
            INIT_3F => X"00000000000000000000002c000000000000000000000000000000000000005d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY4;


    MEM_GOLD_LAYER0_ENTITY5 : if BRAM_NAME = "gold_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_01 => X"000000000000001c0000000f0000000000000000000000000000005200000000",
            INIT_02 => X"0000000000000012000000130000000000000004000000000000000000000000",
            INIT_03 => X"0000000c000000170000000000000005000000000000002d0000000000000000",
            INIT_04 => X"0000001d00000003000000000000000000000016000000000000001100000000",
            INIT_05 => X"000000120000000000000000000000080000000000000011000000000000001b",
            INIT_06 => X"00000000000000000000000900000019000000000000003b0000000000000003",
            INIT_07 => X"0000001000000000000000050000000000000000000000120000001200000000",
            INIT_08 => X"00000000000000330000000d000000000000005800000000000000000000002d",
            INIT_09 => X"00000004000000000000000200000028000000330000003e0000002c0000001d",
            INIT_0A => X"0000007000000036000000000000003b000000000000002e0000004e0000004e",
            INIT_0B => X"00000044000000490000004f00000056000000580000005a000000530000005a",
            INIT_0C => X"0000006f00000048000000080000000000000049000000480000004a0000004c",
            INIT_0D => X"000000540000005b0000005b000000570000005d0000005e0000005a00000060",
            INIT_0E => X"0000008a000000000000003100000050000000450000004d0000005300000057",
            INIT_0F => X"000000610000006400000061000000740000005e000000500000006700000067",
            INIT_10 => X"00000041000000490000005f0000005500000049000000520000005200000052",
            INIT_11 => X"0000005e0000006b00000053000000450000002f0000002e000000330000002e",
            INIT_12 => X"0000002f0000002f000000310000002f0000002b000000230000001c00000027",
            INIT_13 => X"0000002600000027000000240000003200000032000000350000002d00000034",
            INIT_14 => X"0000005500000013000000250000000400000021000000130000001500000024",
            INIT_15 => X"0000002d000000280000001a0000003b000000340000002e000000380000002c",
            INIT_16 => X"00000000000000000000001a0000004f0000000a0000000b0000000400000027",
            INIT_17 => X"0000003900000000000000790000002c0000003600000025000000230000001a",
            INIT_18 => X"0000000800000018000000530000000000000012000000000000000e00000053",
            INIT_19 => X"00000000000000630000000a000000490000002c0000001a0000000000000000",
            INIT_1A => X"000000080000005f0000000b000000000000001e000000000000003900000000",
            INIT_1B => X"00000038000000000000002e0000004900000000000000000000000000000000",
            INIT_1C => X"000000bf000000000000000000000023000000040000000d0000000000000015",
            INIT_1D => X"0000000c0000000000000061000000500000000a0000000000000000000000a4",
            INIT_1E => X"00000000000000000000001e000000270000000d000000000000000000000001",
            INIT_1F => X"0000000000000045000000680000000000000008000000000000007c00000000",
            INIT_20 => X"000000000000002a00000022000000120000000000000017000000000000003c",
            INIT_21 => X"0000001100000003000000000000001c00000031000000060000002200000000",
            INIT_22 => X"000000260000003a000000440000000a00000018000000000000004a00000000",
            INIT_23 => X"000000190000002a0000000e000000170000000a000000000000000500000048",
            INIT_24 => X"000000560000001c000000510000001100000000000000a3000000000000000b",
            INIT_25 => X"0000005600000000000000000000000000000014000000280000002d0000001e",
            INIT_26 => X"0000000000000040000000280000000000000098000000000000000000000000",
            INIT_27 => X"00000000000000000000000900000010000000100000000e0000001100000000",
            INIT_28 => X"0000000300000041000000480000001f0000000000000009000000050000000a",
            INIT_29 => X"0000000800000010000000140000001700000010000000080000001700000000",
            INIT_2A => X"000000100000007400000000000000000000001100000000000000090000000d",
            INIT_2B => X"000000100000000d00000009000000000000002600000000000000000000000d",
            INIT_2C => X"000000190000000000000000000000160000000c000000090000001800000010",
            INIT_2D => X"000000000000000b000000310000000300000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000004000000000000000000000000000000000000000100000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000040000001200000000000000000000000000000000",
            INIT_34 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000001000000270000000000000000000000380000000800000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000014000000000000000000000000000000000000000f00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000001200000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY5;


    MEM_GOLD_LAYER0_ENTITY6 : if BRAM_NAME = "gold_layer0_entity6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001100000000000000000000000000000000000000000000001e00000030",
            INIT_01 => X"0000003e000000000000000000000000000000000000001c0000002400000001",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000001300000000000000000000002f00000036",
            INIT_0A => X"00000033000000350000003500000030000000390000003b000000360000002b",
            INIT_0B => X"0000002000000020000000250000002800000027000000300000003800000036",
            INIT_0C => X"0000003900000033000000420000003b00000039000000230000000200000002",
            INIT_0D => X"0000000600000006000000110000002700000030000000130000003600000039",
            INIT_0E => X"000000370000003d0000001e0000000000000000000000000000000400000000",
            INIT_0F => X"0000000100000000000000170000001500000000000000320000003700000040",
            INIT_10 => X"000000120000001e000000000000000000000000000000170000000000000000",
            INIT_11 => X"0000000000000000000000000000001200000034000000100000004400000033",
            INIT_12 => X"0000002500000006000000000000000000000010000000090000000000000000",
            INIT_13 => X"00000000000000000000000f00000031000000380000000b0000000d0000002b",
            INIT_14 => X"000000080000000b000000000000002a00000000000000000000000000000000",
            INIT_15 => X"000000000000002c000000070000003d0000000e000000110000002e00000017",
            INIT_16 => X"0000000800000003000000130000000000000000000000000000000000000004",
            INIT_17 => X"00000019000000000000002500000000000000220000002e0000000a00000000",
            INIT_18 => X"000000130000000f000000000000000000000002000000000000001500000011",
            INIT_19 => X"00000009000000000000001c00000000000000000000000c000000000000002c",
            INIT_1A => X"0000000000000000000000000000000000000021000000160000000e00000014",
            INIT_1B => X"000000000000000300000000000000000000001f000000060000000500000000",
            INIT_1C => X"00000000000000000000001e0000002800000005000000140000001500000000",
            INIT_1D => X"0000002c00000006000000110000001700000000000000000000000000000000",
            INIT_1E => X"000000000000000000000000000000000000000000000000000000320000003c",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000000000000000000000000000004f0000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000027",
            INIT_26 => X"0000002200000023000000290000002c00000020000000280000002b0000002f",
            INIT_27 => X"00000032000000290000001d0000001e000000290000002e0000002800000024",
            INIT_28 => X"000000240000002c000000210000000e00000043000000300000002e00000005",
            INIT_29 => X"000000210000002900000019000000150000002c0000003f0000000200000028",
            INIT_2A => X"000000290000002a00000020000000280000002400000010000000000000001c",
            INIT_2B => X"0000000c000000320000001a0000000b0000005c000000000000002e00000024",
            INIT_2C => X"000000380000000c000000270000002500000019000000000000002300000018",
            INIT_2D => X"0000001a00000026000000000000002c00000005000000410000000000000013",
            INIT_2E => X"000000270000002a000000240000002500000000000000140000003800000012",
            INIT_2F => X"0000002b0000001a0000002400000000000000370000002f0000000000000000",
            INIT_30 => X"00000016000000250000004300000000000000340000002a000000070000001d",
            INIT_31 => X"0000002000000011000000240000000e00000046000000000000000000000015",
            INIT_32 => X"0000001c00000039000000000000002b000000280000000d0000000000000025",
            INIT_33 => X"0000000b0000000600000029000000340000000200000000000000350000000b",
            INIT_34 => X"0000001800000000000000110000002c00000000000000110000000d0000000d",
            INIT_35 => X"000000000000003f0000000000000034000000000000000e0000001b00000000",
            INIT_36 => X"0000003f000000050000002b00000000000000000000001a0000000000000000",
            INIT_37 => X"00000039000000000000002a00000014000000000000001d0000002c0000000f",
            INIT_38 => X"0000002f0000000f00000000000000100000002f000000000000000000000038",
            INIT_39 => X"0000000000000029000000320000000000000005000000270000002b0000000f",
            INIT_3A => X"0000000800000008000000110000002100000000000000000000000000000000",
            INIT_3B => X"0000005200000005000000000000000000000000000000070000000300000000",
            INIT_3C => X"000000000000000000000003000000140000000000000000000000220000002e",
            INIT_3D => X"0000000000000006000000020000000500000001000000000000000000000002",
            INIT_3E => X"0000000000000000000000090000000000000000000000220000000d00000000",
            INIT_3F => X"0000000900000006000000000000000000000001000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY6;


    MEM_GOLD_LAYER0_ENTITY7 : if BRAM_NAME = "gold_layer0_entity7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001500000013000000000000000000000004000000140000000000000000",
            INIT_01 => X"0000000000000000000000000000000c0000000000000000000000120000001a",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY7;

    MEM_EMPTY_18Kb : if BRAM_NAME = "default" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate;


end a1;