library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    5, 0, 6, 10, 1, 0, 3, 3, 6, 7, 3, 0, 0, 0, 0, 4, 9, 16, 24, 37, 37, 32, 27, 21, 20, 20, 20, 21, 28, 32, 4, 0, 2, 6, 0, 0, 1, 3, 0, 0, 0, 7, 6, 2, 4, 10, 31, 38, 47, 52, 60, 58, 47, 48, 29, 24, 21, 19, 22, 27, 2, 0, 0, 4, 0, 0, 3, 2, 0, 0, 0, 21, 23, 9, 27, 50, 61, 56, 36, 40, 50, 60, 65, 57, 50, 30, 19, 17, 23, 26, 12, 5, 4, 5, 0, 0, 6, 2, 0, 0, 0, 56, 58, 50, 64, 90, 78, 24, 8, 23, 35, 52, 52, 58, 58, 55, 27, 12, 21, 28, 62, 41, 4, 0, 0, 0, 2, 1, 0, 0, 10, 57, 68, 84, 81, 76, 49, 0, 0, 17, 34, 44, 45, 46, 73, 88, 46, 6, 13, 29, 95, 86, 0, 0, 0, 0, 0, 1, 7, 15, 25, 24, 43, 74, 55, 43, 45, 0, 0, 10, 51, 49, 32, 49, 90, 88, 68, 14, 3, 27, 108, 58, 0, 0, 2, 0, 0, 0, 30, 39, 15, 0, 24, 70, 53, 42, 53, 25, 0, 0, 59, 61, 44, 60, 79, 88, 80, 39, 0, 15, 99, 18, 0, 0, 13, 1, 0, 0, 0, 43, 0, 0, 34, 77, 66, 54, 65, 51, 0, 0, 36, 63, 65, 55, 59, 69, 86, 74, 12, 0, 58, 0, 0, 20, 26, 19, 0, 0, 0, 28, 0, 0, 53, 65, 72, 56, 82, 60, 0, 0, 12, 55, 68, 46, 46, 59, 82, 93, 50, 8, 49, 0, 0, 31, 29, 28, 0, 0, 0, 48, 17, 0, 51, 57, 55, 69, 91, 39, 0, 0, 14, 57, 84, 46, 30, 57, 74, 94, 70, 35, 47, 0, 0, 30, 26, 24, 28, 0, 0, 51, 3, 0, 22, 58, 48, 44, 98, 9, 0, 0, 45, 74, 89, 47, 32, 48, 64, 76, 69, 52, 48, 0, 0, 49, 24, 16, 61, 0, 0, 31, 0, 0, 0, 57, 42, 29, 86, 0, 0, 0, 63, 85, 77, 55, 41, 40, 47, 56, 54, 54, 32, 0, 26, 90, 17, 3, 69, 10, 0, 0, 0, 0, 0, 49, 36, 39, 85, 0, 0, 6, 60, 70, 69, 53, 43, 28, 19, 42, 48, 40, 17, 0, 41, 103, 19, 0, 58, 26, 0, 0, 0, 0, 37, 47, 32, 47, 83, 0, 0, 6, 62, 60, 70, 55, 28, 17, 12, 40, 44, 27, 11, 0, 21, 98, 33, 0, 43, 42, 0, 0, 0, 21, 80, 37, 43, 54, 58, 0, 0, 0, 37, 66, 80, 57, 26, 23, 28, 40, 31, 4, 14, 0, 0, 86, 63, 0, 23, 51, 11, 0, 0, 63, 70, 43, 46, 43, 24, 0, 0, 11, 21, 66, 84, 71, 41, 29, 37, 30, 3, 0, 12, 0, 0, 69, 85, 0, 0, 50, 38, 21, 34, 39, 42, 20, 41, 47, 0, 2, 60, 44, 17, 78, 117, 78, 50, 17, 6, 3, 0, 10, 3, 0, 0, 41, 90, 15, 0, 29, 36, 82, 31, 7, 19, 0, 28, 73, 0, 3, 45, 32, 67, 105, 99, 59, 25, 0, 0, 0, 0, 11, 0, 0, 0, 18, 84, 31, 0, 33, 46, 82, 48, 0, 0, 0, 9, 82, 39, 19, 51, 71, 113, 109, 81, 47, 5, 0, 0, 9, 19, 22, 0, 0, 0, 13, 86, 24, 0, 0, 61, 66, 18, 0, 0, 0, 5, 68, 56, 68, 86, 104, 98, 83, 68, 39, 26, 15, 19, 47, 54, 50, 0, 0, 0, 17, 84, 0, 0, 0, 3, 51, 7, 0, 0, 0, 30, 75, 80, 85, 101, 82, 63, 52, 44, 49, 44, 42, 55, 71, 76, 74, 0, 0, 0, 11, 47, 0, 0, 0, 24, 78, 80, 44, 45, 61, 72, 95, 97, 92, 82, 61, 54, 52, 54, 60, 59, 54, 50, 60, 68, 64, 2, 0, 0, 13, 0, 0, 0, 0, 82, 147, 108, 73, 75, 75, 79, 81, 76, 75, 70, 61, 61, 60, 60, 55, 52, 49, 48, 57, 60, 54, 49, 14, 0, 14, 0, 0, 0, 61, 148, 125, 77, 63, 65, 66, 65, 63, 65, 67, 63, 56, 58, 59, 49, 42, 39, 46, 49, 54, 49, 39, 68, 39, 7, 6, 0, 0, 0, 132, 147, 73, 61, 61, 66, 67, 65, 65, 64, 62, 56, 53, 49, 47, 43, 42, 49, 58, 51, 41, 30, 19, 76, 62, 44, 19, 0, 0, 47, 153, 100, 58, 51, 64, 72, 65, 62, 62, 61, 57, 53, 56, 50, 44, 46, 59, 69, 64, 43, 25, 28, 38, 75, 69, 60, 40, 0, 0, 85, 137, 74, 56, 51, 55, 65, 66, 63, 63, 59, 57, 56, 56, 59, 54, 57, 65, 66, 49, 29, 33, 73, 73, 75, 65, 64, 57, 15, 0, 78, 133, 73, 61, 48, 48, 56, 61, 63, 58, 55, 53, 54, 60, 62, 61, 60, 52, 39, 22, 27, 68, 105, 75, 81, 65, 59, 64, 53, 40, 80, 101, 82, 68, 58, 58, 57, 61, 58, 47, 42, 41, 48, 58, 63, 66, 53, 25, 0, 4, 46, 81, 96, 79, 78, 67, 58, 62, 64, 62, 71, 81, 85, 68, 65, 69, 72, 72, 61, 48, 41, 31, 37, 59, 67, 64, 39, 6, 0, 8, 63, 96, 93, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 41, 44, 40, 25, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 31, 52, 69, 72, 65, 55, 49, 28, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 6, 1, 17, 29, 57, 61, 62, 90, 105, 102, 80, 62, 47, 30, 15, 0, 0, 0, 2, 17, 0, 0, 0, 0, 0, 0, 0, 0, 29, 96, 55, 48, 72, 75, 57, 45, 73, 114, 130, 127, 111, 93, 82, 65, 39, 10, 0, 0, 56, 59, 20, 0, 0, 0, 0, 0, 0, 0, 10, 48, 58, 66, 57, 53, 60, 66, 86, 108, 124, 126, 108, 101, 111, 90, 40, 14, 0, 0, 99, 72, 0, 0, 0, 0, 0, 0, 0, 7, 23, 36, 64, 88, 81, 78, 84, 71, 88, 110, 117, 104, 93, 103, 110, 95, 65, 19, 0, 0, 127, 99, 9, 0, 0, 0, 0, 0, 17, 43, 52, 46, 90, 110, 100, 96, 102, 80, 70, 106, 129, 101, 90, 98, 97, 86, 66, 36, 10, 0, 177, 100, 61, 53, 5, 0, 2, 13, 61, 70, 48, 72, 120, 124, 96, 91, 89, 91, 56, 62, 122, 117, 97, 78, 82, 93, 80, 47, 13, 12, 208, 147, 104, 94, 29, 0, 5, 65, 127, 171, 122, 103, 121, 120, 98, 89, 93, 79, 38, 63, 124, 125, 119, 94, 85, 92, 100, 79, 34, 2, 203, 153, 149, 114, 28, 0, 0, 61, 155, 190, 134, 102, 124, 118, 110, 100, 89, 83, 33, 98, 153, 151, 138, 98, 96, 105, 100, 88, 60, 13, 207, 141, 154, 139, 39, 0, 0, 14, 68, 152, 118, 114, 138, 143, 109, 103, 103, 72, 44, 143, 188, 157, 131, 92, 90, 106, 108, 100, 79, 34, 200, 122, 160, 160, 65, 0, 0, 8, 40, 120, 84, 98, 164, 171, 121, 107, 129, 93, 67, 160, 184, 146, 121, 103, 92, 101, 103, 97, 85, 47, 186, 126, 193, 169, 69, 13, 22, 23, 41, 99, 92, 133, 200, 195, 149, 117, 119, 96, 85, 157, 172, 145, 111, 95, 85, 80, 90, 96, 76, 34, 189, 138, 202, 184, 103, 43, 54, 39, 42, 59, 119, 168, 167, 151, 132, 137, 118, 66, 61, 146, 151, 134, 136, 118, 99, 95, 90, 84, 51, 3, 203, 163, 200, 200, 144, 86, 77, 65, 66, 76, 135, 219, 192, 127, 122, 120, 94, 55, 59, 109, 127, 129, 110, 83, 82, 89, 78, 60, 15, 0, 217, 187, 208, 223, 176, 121, 113, 102, 69, 70, 132, 133, 131, 107, 101, 117, 92, 50, 64, 107, 124, 131, 119, 101, 73, 72, 47, 10, 0, 0, 226, 205, 212, 229, 194, 126, 122, 147, 101, 80, 108, 74, 84, 76, 94, 122, 97, 85, 90, 48, 66, 127, 112, 73, 39, 23, 0, 0, 0, 0, 211, 210, 207, 216, 205, 150, 128, 159, 163, 114, 63, 71, 100, 93, 134, 141, 96, 102, 109, 100, 107, 100, 88, 69, 38, 9, 0, 0, 0, 0, 190, 203, 194, 203, 209, 166, 123, 141, 158, 182, 122, 95, 121, 111, 168, 184, 116, 94, 130, 146, 152, 115, 99, 102, 95, 92, 72, 77, 79, 77, 188, 211, 193, 197, 210, 174, 124, 181, 186, 140, 138, 115, 124, 161, 211, 212, 173, 125, 117, 129, 133, 133, 124, 130, 150, 158, 171, 182, 179, 175, 212, 231, 203, 203, 205, 146, 105, 202, 283, 255, 200, 207, 229, 248, 267, 264, 241, 215, 185, 155, 157, 171, 193, 209, 219, 228, 235, 234, 235, 232, 256, 275, 226, 212, 205, 129, 138, 239, 313, 331, 294, 237, 237, 240, 243, 249, 233, 212, 212, 213, 220, 222, 230, 242, 244, 244, 246, 253, 255, 251, 263, 270, 253, 226, 211, 164, 196, 285, 334, 300, 237, 204, 198, 196, 197, 201, 213, 218, 223, 229, 237, 242, 243, 242, 245, 246, 246, 253, 257, 258, 267, 235, 227, 242, 195, 157, 229, 324, 320, 257, 218, 214, 216, 212, 212, 213, 219, 221, 224, 230, 239, 244, 246, 249, 252, 260, 265, 269, 271, 268, 293, 255, 224, 226, 202, 181, 275, 334, 274, 218, 224, 219, 225, 221, 212, 211, 215, 219, 225, 236, 248, 255, 255, 263, 275, 281, 282, 286, 283, 280, 301, 274, 244, 214, 201, 236, 305, 322, 240, 216, 224, 229, 226, 217, 217, 216, 219, 224, 233, 245, 254, 269, 277, 279, 275, 276, 277, 285, 292, 301, 301, 281, 260, 239, 205, 245, 325, 303, 243, 232, 225, 227, 231, 220, 216, 217, 224, 233, 239, 250, 259, 258, 263, 269, 270, 268, 277, 302, 314, 288, 289, 277, 263, 254, 230, 221, 287, 289, 230, 232, 231, 237, 240, 233, 224, 213, 215, 224, 237, 248, 253, 254, 251, 248, 251, 262, 294, 312, 289, 240, 292, 265, 256, 255, 245, 226, 224, 236, 222, 212, 212, 225, 234, 239, 230, 218, 225, 236, 240, 244, 245, 241, 235, 228, 241, 272, 300, 306, 289, 247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 21, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 33, 29, 13, 11, 11, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 0, 4, 22, 29, 20, 12, 26, 24, 9, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 19, 20, 7, 0, 11, 16, 10, 16, 24, 28, 17, 0, 0, 0, 25, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 19, 22, 25, 20, 0, 3, 11, 11, 14, 13, 20, 15, 5, 0, 0, 53, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 13, 18, 20, 32, 14, 0, 0, 2, 12, 14, 6, 16, 15, 13, 0, 0, 83, 46, 2, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 10, 4, 20, 13, 39, 0, 0, 7, 3, 28, 22, 7, 18, 22, 19, 9, 0, 100, 50, 19, 0, 0, 0, 0, 0, 0, 20, 18, 0, 0, 11, 6, 14, 6, 47, 0, 0, 31, 21, 41, 25, 15, 17, 26, 21, 17, 0, 108, 43, 14, 4, 0, 0, 0, 0, 0, 16, 9, 0, 0, 13, 8, 5, 4, 49, 0, 0, 42, 32, 37, 22, 22, 22, 28, 20, 17, 0, 102, 24, 18, 41, 0, 0, 0, 0, 0, 6, 0, 0, 0, 29, 16, 6, 15, 54, 0, 10, 44, 33, 30, 26, 25, 21, 17, 14, 11, 0, 91, 17, 28, 53, 0, 0, 0, 0, 0, 1, 0, 0, 33, 43, 20, 12, 21, 40, 0, 14, 38, 25, 26, 30, 19, 14, 8, 2, 0, 0, 81, 24, 34, 46, 40, 0, 0, 0, 0, 0, 0, 9, 50, 34, 26, 22, 13, 14, 0, 3, 24, 30, 33, 37, 24, 17, 7, 0, 0, 0, 79, 42, 41, 41, 69, 0, 0, 0, 0, 0, 14, 45, 48, 30, 16, 23, 11, 0, 0, 6, 9, 13, 22, 28, 24, 18, 6, 0, 0, 0, 79, 61, 53, 48, 81, 43, 0, 0, 0, 0, 30, 16, 10, 12, 0, 30, 12, 0, 0, 9, 0, 18, 39, 34, 15, 2, 0, 0, 0, 0, 70, 69, 63, 55, 70, 63, 15, 18, 10, 0, 26, 0, 0, 0, 0, 36, 27, 0, 0, 0, 0, 33, 32, 29, 0, 0, 0, 0, 0, 0, 51, 63, 60, 52, 61, 76, 35, 31, 29, 13, 31, 0, 21, 0, 0, 40, 35, 0, 4, 9, 34, 40, 32, 32, 0, 0, 0, 0, 0, 0, 31, 55, 51, 42, 55, 83, 36, 17, 46, 43, 40, 10, 18, 0, 18, 43, 42, 17, 30, 50, 62, 55, 52, 51, 46, 21, 0, 0, 0, 0, 31, 63, 50, 39, 62, 87, 19, 0, 35, 39, 37, 34, 37, 48, 64, 70, 72, 49, 54, 61, 68, 67, 72, 78, 90, 77, 73, 68, 75, 75, 70, 90, 64, 45, 59, 62, 0, 21, 55, 88, 110, 104, 108, 119, 121, 123, 127, 102, 93, 90, 100, 107, 117, 128, 136, 138, 138, 132, 138, 138, 137, 131, 91, 56, 64, 44, 0, 45, 96, 155, 158, 131, 129, 131, 129, 130, 134, 124, 126, 133, 138, 141, 146, 152, 151, 155, 155, 155, 158, 160, 176, 159, 116, 80, 91, 34, 11, 67, 140, 159, 137, 122, 121, 120, 120, 125, 135, 137, 143, 149, 152, 156, 156, 157, 152, 155, 156, 158, 165, 166, 186, 168, 135, 105, 94, 20, 28, 108, 167, 144, 134, 131, 134, 135, 131, 132, 137, 140, 143, 149, 155, 158, 158, 157, 160, 163, 169, 172, 173, 162, 196, 180, 155, 128, 103, 39, 59, 141, 150, 131, 137, 136, 141, 138, 133, 132, 135, 139, 144, 151, 160, 165, 166, 170, 177, 180, 186, 178, 173, 175, 199, 188, 168, 148, 128, 80, 88, 159, 136, 135, 141, 136, 141, 138, 135, 135, 140, 143, 150, 155, 168, 175, 175, 178, 181, 185, 180, 180, 188, 200, 196, 191, 178, 163, 150, 124, 116, 172, 139, 144, 144, 138, 142, 138, 139, 138, 141, 144, 151, 158, 166, 170, 173, 176, 174, 173, 177, 198, 200, 198, 192, 189, 177, 171, 158, 148, 133, 160, 144, 150, 146, 146, 148, 144, 142, 133, 134, 141, 147, 152, 160, 165, 166, 161, 155, 158, 176, 193, 190, 178, 185, 179, 168, 169, 158, 149, 138, 138, 144, 144, 140, 149, 149, 148, 145, 138, 139, 142, 141, 148, 157, 153, 154, 145, 144, 150, 173, 192, 194, 169, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152, 163, 164, 157, 154, 159, 157, 158, 156, 154, 151, 150, 160, 170, 171, 168, 159, 148, 147, 144, 138, 138, 136, 141, 136, 133, 134, 139, 138, 130, 150, 160, 165, 156, 155, 160, 158, 161, 158, 154, 137, 131, 152, 166, 162, 160, 146, 143, 133, 112, 95, 92, 107, 118, 129, 138, 136, 137, 137, 130, 148, 150, 160, 157, 162, 164, 164, 163, 163, 165, 133, 118, 139, 153, 147, 147, 156, 137, 95, 72, 57, 51, 54, 69, 81, 103, 126, 134, 135, 134, 143, 145, 157, 161, 164, 167, 167, 164, 162, 161, 200, 184, 144, 142, 151, 136, 116, 80, 73, 67, 64, 51, 49, 51, 43, 72, 108, 126, 128, 129, 124, 135, 163, 165, 159, 166, 165, 160, 160, 148, 208, 178, 129, 103, 93, 72, 49, 59, 76, 68, 72, 77, 73, 50, 61, 51, 66, 105, 127, 126, 95, 78, 102, 137, 158, 167, 170, 163, 156, 148, 162, 138, 105, 77, 48, 46, 38, 57, 89, 87, 78, 82, 72, 78, 74, 50, 41, 72, 118, 127, 77, 38, 38, 92, 147, 164, 165, 163, 139, 137, 128, 97, 92, 79, 58, 66, 56, 46, 97, 127, 97, 68, 75, 92, 69, 50, 29, 47, 103, 124, 71, 19, 33, 86, 134, 157, 165, 144, 104, 68, 65, 86, 105, 89, 63, 61, 61, 56, 79, 110, 104, 71, 62, 65, 65, 46, 33, 24, 73, 123, 95, 27, 62, 103, 135, 150, 163, 145, 136, 91, 86, 105, 104, 91, 56, 55, 56, 59, 54, 75, 92, 76, 61, 61, 58, 53, 50, 27, 35, 95, 91, 60, 94, 115, 129, 145, 121, 177, 196, 157, 111, 122, 96, 82, 74, 60, 48, 49, 47, 72, 88, 96, 83, 67, 68, 60, 55, 38, 16, 47, 66, 85, 100, 123, 131, 155, 106, 149, 166, 155, 132, 140, 109, 76, 87, 61, 50, 26, 44, 111, 106, 113, 82, 57, 72, 71, 65, 47, 25, 29, 62, 67, 87, 129, 142, 161, 137, 98, 136, 142, 111, 118, 134, 93, 78, 76, 73, 22, 61, 131, 108, 104, 71, 57, 64, 80, 65, 51, 37, 47, 54, 64, 99, 100, 115, 151, 153, 94, 133, 131, 89, 104, 158, 139, 94, 74, 88, 36, 85, 122, 111, 86, 52, 51, 48, 54, 56, 56, 50, 75, 49, 78, 122, 65, 74, 122, 142, 95, 110, 102, 107, 84, 131, 126, 104, 103, 95, 41, 96, 134, 102, 85, 76, 70, 60, 53, 68, 78, 81, 93, 55, 88, 121, 63, 48, 89, 119, 80, 114, 101, 140, 169, 137, 107, 110, 108, 88, 59, 102, 136, 111, 86, 65, 51, 62, 65, 78, 104, 102, 95, 67, 85, 109, 89, 39, 88, 103, 74, 92, 93, 151, 184, 121, 106, 90, 83, 83, 53, 100, 160, 145, 91, 79, 65, 67, 81, 83, 94, 89, 108, 85, 81, 103, 113, 37, 66, 94, 99, 49, 95, 129, 112, 96, 79, 64, 60, 77, 72, 106, 83, 92, 117, 94, 62, 53, 71, 90, 93, 110, 141, 109, 92, 102, 116, 57, 42, 92, 110, 76, 68, 71, 84, 95, 81, 75, 42, 61, 111, 104, 49, 77, 99, 64, 46, 33, 46, 88, 108, 134, 145, 126, 101, 105, 115, 82, 41, 72, 65, 77, 97, 53, 93, 89, 69, 97, 56, 32, 95, 114, 116, 101, 57, 50, 29, 47, 64, 107, 132, 143, 139, 125, 104, 108, 111, 98, 64, 81, 59, 23, 48, 13, 46, 30, 58, 109, 78, 27, 47, 71, 88, 59, 22, 4, 0, 25, 41, 90, 110, 103, 101, 112, 102, 101, 109, 98, 56, 57, 111, 80, 29, 26, 58, 74, 117, 135, 117, 81, 63, 48, 15, 0, 2, 0, 2, 7, 28, 55, 62, 53, 52, 109, 112, 99, 108, 89, 33, 60, 139, 148, 111, 98, 87, 102, 111, 114, 105, 64, 49, 24, 5, 0, 0, 7, 10, 2, 6, 11, 21, 16, 5, 63, 104, 108, 104, 108, 69, 115, 138, 156, 141, 60, 33, 35, 29, 31, 33, 14, 10, 10, 7, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 34, 81, 108, 102, 86, 132, 150, 158, 75, 13, 4, 0, 2, 0, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 97, 73, 92, 134, 157, 93, 25, 3, 0, 4, 4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 8, 4, 0, 0, 0, 0, 0, 36, 57, 113, 146, 123, 34, 7, 4, 3, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 11, 0, 0, 0, 0, 20, 125, 162, 87, 33, 10, 4, 3, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 8, 28, 0, 0, 0, 0, 0, 75, 147, 70, 27, 21, 10, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 76, 26, 8, 4, 2, 13, 19, 20, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 0, 0, 7, 14, 21, 21, 15, 9, 5, 1, 0, 0, 0, 5, 21, 18, 7, 0, 0, 12, 11, 12, 17, 11, 7, 11, 6, 8, 8, 8, 10, 9, 9, 12, 10, 9, 6, 6, 9, 9, 10, 11, 9, 9, 4, 8, 8, 10, 11, 12, 8, 9, 17, 9, 8, 8, 12, 10, 4, 0, 0, 7, 9, 9, 5, 1, 0, 6, 2, 2, 6, 5, 13, 15, 12, 10, 7, 8, 6, 7, 4, 5, 10, 9, 9, 9, 12, 13, 19, 0, 0, 5, 5, 1, 7, 5, 26, 8, 0, 0, 0, 0, 0, 7, 11, 11, 7, 7, 8, 4, 2, 5, 5, 10, 9, 13, 13, 13, 31, 0, 21, 18, 8, 8, 9, 35, 23, 0, 0, 0, 1, 0, 0, 0, 0, 10, 10, 4, 8, 0, 19, 23, 13, 6, 9, 11, 11, 4, 0, 7, 52, 16, 0, 22, 21, 9, 0, 0, 0, 0, 4, 19, 0, 0, 2, 6, 12, 7, 9, 0, 21, 23, 7, 6, 11, 12, 7, 7, 0, 4, 25, 6, 3, 5, 0, 0, 0, 0, 0, 0, 17, 12, 0, 18, 5, 0, 5, 6, 9, 0, 13, 0, 0, 5, 11, 8, 3, 0, 0, 17, 0, 0, 3, 3, 0, 0, 0, 2, 6, 6, 6, 0, 14, 11, 12, 0, 0, 7, 9, 0, 23, 0, 0, 4, 9, 4, 0, 0, 0, 0, 0, 0, 7, 6, 3, 7, 0, 4, 9, 12, 0, 0, 10, 11, 1, 0, 0, 8, 8, 21, 0, 0, 0, 10, 6, 35, 0, 0, 0, 0, 0, 5, 16, 8, 0, 0, 16, 5, 0, 0, 3, 0, 0, 0, 3, 1, 0, 0, 7, 46, 0, 0, 0, 21, 0, 25, 0, 11, 21, 24, 0, 2, 18, 0, 8, 0, 24, 0, 0, 0, 0, 15, 16, 0, 0, 3, 3, 0, 0, 25, 0, 0, 7, 22, 4, 0, 7, 17, 43, 35, 15, 0, 0, 10, 1, 0, 26, 0, 0, 3, 5, 28, 5, 7, 4, 8, 4, 0, 0, 32, 0, 0, 21, 31, 14, 0, 3, 0, 22, 32, 0, 0, 1, 2, 5, 0, 17, 0, 0, 14, 21, 24, 0, 0, 7, 11, 1, 3, 0, 41, 0, 0, 31, 29, 11, 10, 5, 0, 40, 0, 0, 0, 27, 6, 0, 10, 15, 0, 0, 18, 14, 5, 0, 0, 5, 0, 0, 2, 5, 28, 0, 0, 20, 9, 2, 2, 0, 0, 20, 0, 0, 0, 46, 23, 0, 15, 13, 0, 0, 30, 16, 7, 15, 2, 0, 0, 0, 9, 21, 12, 0, 8, 3, 7, 0, 3, 4, 0, 9, 0, 0, 34, 16, 14, 26, 22, 0, 0, 17, 9, 3, 10, 13, 5, 0, 0, 8, 30, 9, 6, 0, 5, 0, 12, 0, 13, 0, 12, 0, 0, 61, 45, 21, 12, 12, 9, 0, 0, 22, 34, 16, 8, 9, 3, 3, 4, 20, 13, 0, 6, 0, 0, 6, 2, 7, 0, 0, 0, 0, 19, 28, 17, 17, 0, 2, 16, 0, 0, 28, 4, 6, 34, 18, 4, 13, 15, 16, 0, 4, 13, 0, 0, 15, 6, 0, 0, 21, 0, 0, 32, 0, 11, 4, 0, 0, 4, 3, 29, 0, 0, 33, 26, 16, 0, 0, 0, 0, 0, 11, 10, 0, 0, 11, 8, 1, 0, 2, 19, 0, 15, 0, 19, 0, 0, 0, 0, 3, 29, 5, 20, 24, 14, 13, 0, 0, 0, 0, 3, 1, 0, 0, 0, 3, 15, 24, 1, 0, 0, 9, 0, 0, 0, 0, 0, 6, 0, 0, 0, 25, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 31, 0, 0, 0, 0, 0, 0, 0, 0, 17, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 17, 16, 0, 0, 29, 0, 5, 2, 0, 20, 31, 31, 31, 29, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 25, 11, 4, 26, 0, 0, 0, 0, 49, 40, 0, 1, 2, 9, 18, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 0, 36, 0, 0, 0, 48, 63, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 26, 0, 0, 9, 75, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 55, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 59, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 24, 59, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 23, 32, 0, 1, 0, 1, 5, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 8, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 52, 55, 56, 51, 53, 52, 52, 52, 52, 51, 48, 47, 53, 60, 60, 60, 55, 51, 49, 52, 52, 53, 53, 51, 52, 49, 48, 53, 55, 53, 54, 58, 59, 49, 51, 51, 51, 50, 51, 45, 34, 22, 40, 55, 51, 50, 51, 48, 50, 35, 26, 25, 39, 48, 51, 59, 52, 50, 52, 52, 51, 51, 53, 53, 53, 55, 53, 55, 53, 35, 20, 0, 21, 44, 46, 50, 66, 54, 28, 1, 0, 0, 0, 14, 26, 31, 49, 52, 51, 52, 44, 49, 53, 56, 56, 58, 57, 56, 57, 42, 60, 42, 40, 52, 65, 68, 42, 26, 9, 0, 0, 0, 0, 0, 5, 18, 43, 52, 49, 44, 47, 46, 74, 67, 55, 55, 56, 54, 58, 64, 57, 46, 42, 34, 23, 24, 13, 13, 5, 0, 0, 0, 0, 0, 2, 14, 23, 44, 52, 44, 32, 19, 39, 53, 54, 57, 58, 55, 52, 57, 52, 35, 18, 5, 2, 7, 6, 4, 10, 0, 0, 0, 9, 13, 11, 18, 24, 29, 48, 48, 0, 0, 7, 8, 39, 55, 51, 43, 39, 32, 34, 11, 0, 0, 5, 14, 15, 11, 15, 26, 3, 0, 13, 21, 21, 11, 16, 25, 44, 51, 0, 0, 0, 0, 19, 49, 40, 13, 0, 0, 0, 0, 0, 2, 3, 10, 14, 26, 21, 15, 0, 0, 0, 5, 13, 10, 10, 15, 32, 57, 0, 0, 0, 0, 16, 50, 25, 14, 0, 0, 0, 0, 0, 0, 0, 1, 20, 11, 13, 0, 0, 0, 0, 4, 7, 2, 10, 17, 21, 41, 0, 0, 0, 0, 7, 48, 33, 37, 24, 0, 0, 0, 0, 0, 4, 0, 11, 1, 2, 0, 0, 0, 0, 9, 14, 6, 0, 6, 10, 24, 0, 0, 0, 0, 10, 47, 58, 26, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 9, 14, 7, 5, 0, 16, 0, 0, 0, 0, 28, 49, 56, 31, 33, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 4, 13, 14, 17, 10, 0, 0, 10, 0, 0, 0, 0, 11, 46, 55, 39, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 27, 40, 33, 20, 0, 0, 0, 0, 0, 0, 10, 7, 0, 4, 0, 0, 0, 11, 11, 11, 2, 0, 9, 13, 23, 0, 0, 0, 0, 0, 2, 11, 22, 19, 13, 0, 11, 1, 3, 13, 10, 14, 11, 16, 0, 1, 0, 0, 0, 9, 12, 15, 27, 28, 31, 0, 0, 0, 0, 0, 0, 3, 4, 0, 34, 26, 23, 26, 13, 14, 4, 8, 3, 23, 40, 42, 8, 9, 29, 27, 27, 24, 13, 19, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 24, 25, 0, 0, 0, 0, 0, 15, 10, 3, 13, 33, 36, 30, 33, 22, 25, 16, 26, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 16, 0, 8, 11, 22, 35, 18, 19, 4, 20, 26, 37, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 16, 0, 0, 0, 0, 0, 7, 34, 45, 41, 31, 25, 19, 11, 11, 23, 29, 35, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 27, 18, 9, 0, 0, 0, 0, 3, 16, 14, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 13, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 92, 86, 88, 92, 94, 95, 94, 97, 96, 93, 87, 89, 96, 97, 99, 103, 97, 93, 85, 82, 79, 80, 82, 83, 80, 81, 81, 83, 83, 92, 95, 87, 89, 93, 97, 96, 96, 100, 108, 98, 91, 95, 100, 102, 102, 91, 92, 88, 87, 81, 74, 73, 66, 75, 74, 82, 86, 88, 87, 98, 100, 91, 88, 94, 95, 94, 96, 101, 137, 102, 95, 99, 100, 87, 74, 71, 83, 89, 88, 80, 76, 70, 72, 71, 76, 83, 85, 85, 86, 96, 98, 90, 90, 95, 94, 93, 96, 98, 120, 77, 69, 78, 73, 64, 55, 72, 89, 80, 77, 70, 65, 67, 65, 61, 65, 77, 83, 81, 85, 69, 83, 85, 90, 98, 97, 96, 98, 100, 105, 78, 82, 77, 74, 78, 67, 78, 88, 77, 70, 63, 59, 64, 58, 52, 55, 71, 78, 72, 78, 58, 81, 97, 92, 95, 97, 98, 98, 101, 96, 94, 97, 81, 76, 81, 68, 69, 86, 83, 66, 61, 65, 63, 50, 46, 51, 56, 73, 69, 72, 57, 97, 96, 92, 96, 102, 104, 109, 92, 100, 110, 106, 80, 66, 70, 61, 60, 69, 79, 63, 59, 64, 59, 52, 52, 50, 48, 63, 71, 71, 67, 112, 92, 78, 96, 104, 129, 140, 118, 112, 124, 91, 69, 58, 64, 57, 50, 57, 82, 71, 69, 66, 62, 64, 59, 57, 46, 52, 71, 71, 89, 107, 85, 69, 92, 90, 146, 135, 102, 82, 97, 70, 61, 64, 55, 60, 40, 64, 101, 79, 85, 64, 63, 69, 60, 60, 48, 46, 63, 69, 99, 100, 81, 67, 95, 81, 113, 111, 66, 56, 86, 73, 58, 67, 57, 60, 39, 86, 116, 78, 87, 53, 59, 68, 64, 60, 58, 48, 59, 59, 102, 94, 78, 66, 90, 78, 82, 107, 61, 44, 85, 85, 65, 74, 71, 74, 39, 112, 111, 67, 74, 51, 61, 66, 64, 58, 61, 51, 57, 50, 108, 98, 59, 65, 83, 80, 67, 112, 56, 64, 100, 116, 78, 83, 82, 76, 42, 117, 100, 65, 71, 55, 62, 58, 61, 63, 68, 58, 60, 49, 116, 95, 46, 67, 89, 83, 64, 107, 66, 95, 108, 106, 74, 79, 81, 69, 47, 114, 89, 65, 75, 66, 66, 67, 68, 76, 77, 61, 60, 59, 116, 88, 51, 66, 96, 88, 74, 110, 87, 132, 119, 90, 82, 75, 70, 59, 50, 102, 83, 66, 68, 61, 51, 60, 67, 71, 70, 53, 61, 68, 111, 88, 68, 56, 102, 89, 86, 89, 101, 110, 83, 51, 55, 65, 58, 62, 57, 94, 72, 73, 72, 64, 59, 67, 66, 62, 55, 50, 67, 76, 104, 91, 80, 47, 86, 87, 80, 80, 104, 87, 56, 48, 58, 67, 62, 74, 77, 81, 56, 73, 64, 51, 48, 48, 52, 55, 56, 69, 83, 82, 97, 91, 85, 54, 75, 90, 76, 73, 94, 62, 68, 62, 75, 94, 68, 81, 89, 75, 73, 97, 69, 42, 38, 54, 50, 61, 62, 74, 79, 79, 92, 91, 87, 65, 62, 90, 65, 74, 83, 50, 91, 58, 81, 102, 65, 72, 88, 63, 81, 79, 48, 46, 47, 67, 61, 77, 73, 78, 80, 85, 89, 92, 91, 72, 58, 93, 85, 65, 70, 41, 75, 64, 101, 109, 73, 68, 75, 56, 53, 43, 37, 44, 51, 63, 63, 78, 83, 86, 95, 95, 87, 95, 95, 71, 49, 96, 112, 91, 87, 92, 110, 106, 127, 111, 82, 75, 79, 55, 57, 52, 60, 65, 71, 73, 76, 85, 92, 93, 101, 101, 88, 97, 98, 72, 59, 126, 131, 105, 99, 89, 99, 88, 79, 67, 59, 50, 56, 50, 62, 73, 74, 71, 70, 63, 71, 76, 88, 89, 95, 91, 78, 88, 96, 80, 83, 149, 129, 107, 72, 59, 53, 54, 47, 44, 45, 45, 56, 56, 68, 68, 65, 64, 61, 59, 62, 63, 67, 63, 66, 65, 64, 82, 85, 66, 95, 138, 116, 89, 57, 54, 66, 61, 56, 56, 55, 55, 57, 54, 60, 61, 58, 59, 58, 61, 60, 62, 63, 61, 61, 62, 64, 77, 82, 59, 115, 137, 100, 57, 54, 63, 63, 57, 53, 51, 50, 51, 51, 53, 58, 60, 59, 61, 65, 65, 62, 61, 62, 61, 68, 74, 59, 66, 66, 68, 127, 125, 72, 48, 65, 66, 55, 51, 49, 49, 52, 55, 58, 60, 62, 63, 65, 66, 66, 61, 57, 55, 63, 69, 77, 74, 58, 61, 60, 69, 126, 101, 52, 66, 75, 62, 57, 49, 50, 52, 52, 54, 57, 59, 61, 59, 61, 61, 59, 55, 55, 62, 76, 76, 64, 55, 57, 58, 57, 60, 94, 88, 29, 76, 69, 63, 61, 56, 57, 54, 52, 50, 53, 54, 56, 55, 57, 58, 55, 54, 59, 73, 73, 59, 36, 51, 56, 57, 52, 52, 64, 67, 30, 64, 61, 58, 57, 55, 59, 55, 57, 57, 58, 58, 56, 54, 54, 53, 54, 62, 72, 79, 67, 54, 40, 63, 50, 56, 49, 49, 53, 61, 46, 64, 58, 59, 53, 51, 51, 49, 55, 56, 59, 63, 62, 58, 55, 53, 61, 74, 83, 77, 61, 51, 46, 51, 49, 54, 48, 48, 49, 55, 53, 54, 54, 56, 49, 52, 49, 46, 48, 50, 57, 65, 60, 54, 56, 54, 67, 73, 79, 66, 50, 44, 50, 45, 451, 464, 459, 450, 460, 466, 465, 464, 463, 450, 441, 450, 476, 504, 507, 499, 476, 443, 406, 372, 355, 352, 367, 375, 381, 392, 404, 415, 408, 388, 461, 477, 472, 462, 468, 473, 471, 470, 461, 435, 426, 434, 460, 489, 484, 463, 427, 368, 325, 278, 259, 260, 281, 309, 333, 360, 389, 409, 408, 392, 458, 472, 475, 473, 477, 480, 477, 476, 469, 433, 416, 384, 414, 436, 419, 387, 333, 280, 230, 174, 143, 139, 175, 200, 255, 303, 351, 383, 396, 390, 421, 426, 450, 470, 485, 488, 484, 484, 485, 484, 433, 352, 359, 363, 321, 279, 244, 209, 166, 119, 93, 80, 88, 118, 160, 214, 288, 341, 371, 381, 350, 343, 402, 453, 482, 492, 488, 491, 493, 487, 457, 354, 302, 264, 225, 188, 162, 161, 149, 122, 107, 93, 98, 104, 104, 140, 215, 292, 345, 365, 232, 230, 338, 421, 470, 496, 494, 484, 471, 437, 388, 320, 250, 177, 141, 126, 121, 147, 160, 141, 126, 126, 133, 119, 100, 94, 145, 238, 320, 356, 132, 109, 252, 365, 446, 488, 482, 452, 420, 362, 319, 275, 210, 146, 121, 114, 106, 144, 184, 175, 142, 141, 149, 136, 105, 91, 108, 186, 286, 343, 73, 73, 190, 297, 407, 465, 432, 387, 309, 260, 243, 230, 176, 132, 117, 121, 111, 122, 180, 207, 157, 132, 136, 134, 112, 88, 90, 144, 244, 317, 50, 70, 172, 260, 371, 437, 395, 340, 231, 158, 175, 196, 157, 125, 116, 106, 107, 109, 157, 195, 158, 132, 111, 117, 121, 100, 84, 95, 181, 278, 67, 86, 158, 245, 355, 411, 396, 332, 243, 158, 174, 186, 153, 136, 120, 110, 97, 97, 167, 182, 147, 135, 108, 122, 120, 107, 88, 75, 109, 214, 51, 104, 158, 227, 345, 406, 366, 328, 272, 181, 194, 213, 170, 141, 140, 113, 90, 96, 190, 178, 140, 132, 107, 121, 131, 113, 90, 71, 78, 157, 36, 109, 152, 203, 333, 414, 358, 302, 277, 190, 229, 242, 196, 139, 145, 135, 87, 100, 194, 176, 132, 122, 105, 112, 125, 120, 105, 86, 89, 149, 42, 117, 115, 157, 299, 399, 369, 307, 275, 203, 226, 236, 199, 141, 138, 144, 103, 109, 186, 159, 116, 108, 99, 96, 110, 117, 112, 104, 121, 179, 57, 128, 90, 95, 215, 337, 338, 295, 271, 217, 218, 193, 165, 160, 150, 138, 118, 143, 199, 161, 130, 113, 96, 93, 102, 114, 133, 145, 172, 247, 60, 117, 85, 61, 121, 239, 265, 275, 249, 252, 234, 155, 137, 158, 160, 155, 146, 177, 244, 203, 148, 124, 111, 106, 116, 125, 154, 189, 241, 310, 57, 94, 83, 46, 70, 158, 203, 216, 243, 263, 231, 199, 160, 161, 159, 143, 152, 214, 259, 231, 195, 137, 102, 105, 122, 136, 170, 223, 293, 346, 58, 74, 83, 48, 36, 109, 154, 158, 190, 224, 186, 196, 177, 169, 151, 121, 156, 201, 225, 244, 223, 149, 120, 110, 137, 176, 231, 292, 356, 390, 89, 76, 85, 61, 28, 75, 136, 125, 128, 155, 160, 186, 161, 165, 130, 93, 146, 189, 172, 170, 160, 135, 104, 92, 135, 197, 294, 346, 385, 404, 132, 100, 102, 85, 40, 47, 94, 110, 107, 94, 132, 166, 153, 175, 120, 65, 124, 184, 186, 152, 103, 90, 73, 75, 125, 203, 321, 367, 380, 385, 155, 115, 121, 108, 58, 43, 84, 59, 59, 67, 83, 111, 118, 134, 100, 51, 62, 125, 139, 115, 61, 26, 18, 19, 64, 122, 198, 223, 225, 217, 126, 96, 115, 107, 60, 63, 142, 98, 11, 15, 32, 54, 71, 87, 67, 37, 18, 22, 26, 12, 0, 0, 0, 0, 0, 0, 40, 53, 42, 38, 55, 54, 83, 86, 52, 86, 172, 161, 97, 9, 3, 35, 40, 46, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 49, 76, 66, 131, 186, 155, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 50, 86, 171, 189, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 73, 161, 149, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 129, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 83, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 12, 0, 0, 0, 0, 6, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 4, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 8, 0, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 0, 0, 15, 14, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 8, 15, 0, 0, 0, 0, 0, 2, 8, 0, 0, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 13, 4, 0, 0, 0, 0, 1, 3, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 38, 38, 0, 21, 0, 29, 10, 0, 25, 9, 0, 0, 0, 0, 3, 7, 14, 0, 13, 8, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 24, 62, 36, 16, 0, 3, 0, 0, 2, 1, 0, 5, 8, 10, 19, 30, 20, 21, 16, 17, 20, 18, 10, 15, 29, 10, 1, 10, 18, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 2, 26, 21, 21, 22, 20, 21, 24, 21, 23, 23, 27, 24, 23, 11, 12, 14, 6, 9, 0, 6, 0, 0, 0, 0, 0, 0, 0, 4, 12, 12, 20, 16, 20, 24, 21, 23, 28, 28, 25, 27, 32, 25, 30, 5, 5, 9, 6, 4, 0, 0, 0, 0, 2, 16, 22, 20, 20, 16, 15, 18, 21, 21, 23, 28, 29, 31, 32, 32, 30, 30, 31, 34, 45, 27, 4, 1, 28, 8, 8, 0, 0, 0, 9, 21, 19, 18, 19, 20, 20, 22, 25, 26, 28, 34, 35, 33, 26, 26, 27, 27, 40, 46, 39, 36, 25, 8, 19, 2, 18, 0, 0, 0, 13, 20, 21, 18, 19, 23, 23, 25, 25, 28, 28, 26, 32, 28, 26, 23, 28, 38, 44, 25, 16, 37, 37, 30, 5, 0, 13, 26, 0, 6, 15, 24, 29, 23, 20, 19, 20, 22, 25, 26, 25, 22, 24, 27, 29, 33, 43, 36, 22, 10, 17, 31, 34, 37, 23, 0, 0, 28, 0, 4, 16, 18, 29, 29, 24, 22, 24, 24, 25, 22, 27, 24, 21, 25, 35, 47, 40, 29, 29, 27, 19, 29, 30, 33, 33, 9, 0, 36, 2, 8, 13, 12, 15, 17, 23, 25, 26, 25, 29, 31, 25, 21, 24, 30, 38, 45, 37, 37, 30, 38, 15, 31, 23, 30, 29, 32, 14, 25, 20, 17, 16, 16, 13, 12, 10, 10, 14, 22, 28, 29, 23, 23, 25, 25, 29, 29, 32, 24, 21, 36, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 119, 122, 120, 113, 117, 121, 121, 116, 117, 120, 120, 120, 123, 122, 118, 117, 118, 123, 120, 113, 104, 98, 100, 96, 95, 93, 88, 83, 79, 71, 110, 116, 115, 113, 119, 124, 125, 119, 119, 119, 132, 136, 126, 119, 121, 123, 128, 114, 105, 102, 97, 94, 88, 90, 89, 85, 88, 88, 84, 76, 106, 118, 117, 116, 120, 127, 125, 122, 126, 137, 171, 167, 135, 126, 131, 128, 97, 79, 94, 99, 91, 81, 80, 73, 80, 87, 88, 91, 91, 82, 115, 122, 122, 122, 124, 126, 123, 121, 133, 201, 201, 158, 134, 125, 98, 76, 59, 81, 111, 128, 115, 98, 74, 62, 71, 69, 74, 86, 94, 88, 123, 109, 99, 116, 127, 122, 119, 121, 131, 207, 194, 147, 116, 95, 64, 42, 54, 91, 136, 166, 153, 121, 94, 95, 63, 48, 58, 74, 86, 89, 92, 70, 85, 119, 129, 122, 118, 121, 127, 144, 132, 120, 106, 72, 53, 49, 72, 111, 153, 176, 160, 124, 118, 101, 65, 26, 28, 60, 80, 90, 71, 27, 82, 135, 133, 124, 128, 127, 141, 121, 115, 146, 145, 107, 85, 71, 74, 119, 158, 164, 146, 127, 113, 85, 62, 27, 14, 36, 62, 87, 100, 80, 120, 149, 139, 129, 131, 161, 175, 166, 167, 190, 171, 123, 95, 85, 73, 79, 128, 167, 151, 124, 100, 81, 59, 37, 11, 23, 49, 73, 140, 162, 189, 175, 144, 137, 159, 237, 249, 221, 205, 209, 182, 121, 97, 77, 59, 38, 95, 175, 180, 143, 101, 77, 76, 62, 21, 0, 31, 63, 199, 216, 229, 194, 153, 127, 211, 281, 307, 266, 236, 212, 191, 145, 99, 79, 47, 29, 122, 213, 221, 168, 109, 89, 85, 83, 49, 5, 9, 44, 218, 230, 253, 201, 158, 114, 173, 235, 279, 254, 225, 223, 213, 179, 118, 96, 51, 63, 190, 251, 241, 163, 105, 98, 96, 91, 66, 29, 14, 26, 201, 236, 271, 198, 150, 124, 106, 166, 207, 203, 224, 272, 255, 206, 157, 129, 64, 107, 230, 265, 230, 146, 97, 85, 93, 87, 86, 65, 47, 25, 205, 250, 250, 182, 143, 135, 101, 139, 152, 171, 240, 317, 289, 215, 178, 167, 93, 136, 230, 259, 203, 136, 105, 81, 83, 96, 108, 97, 82, 40, 233, 270, 226, 165, 131, 140, 112, 126, 139, 204, 275, 346, 291, 226, 192, 155, 96, 153, 226, 233, 201, 146, 98, 73, 77, 108, 128, 115, 84, 62, 259, 275, 240, 173, 133, 147, 129, 143, 134, 239, 320, 282, 225, 190, 169, 139, 98, 141, 209, 216, 187, 149, 109, 92, 95, 117, 129, 98, 72, 81, 281, 284, 274, 194, 160, 146, 151, 150, 159, 245, 286, 227, 179, 140, 136, 123, 97, 156, 191, 171, 156, 143, 86, 64, 79, 91, 98, 81, 91, 103, 296, 299, 302, 217, 177, 162, 171, 139, 174, 180, 155, 155, 136, 130, 138, 125, 112, 152, 141, 163, 174, 118, 62, 37, 50, 68, 73, 91, 113, 112, 308, 305, 308, 240, 176, 174, 187, 166, 153, 133, 113, 122, 119, 147, 155, 142, 139, 135, 110, 133, 124, 64, 22, 10, 30, 71, 93, 116, 119, 116, 307, 307, 303, 261, 186, 170, 181, 215, 179, 91, 107, 113, 144, 218, 202, 150, 151, 146, 144, 107, 51, 26, 0, 28, 42, 92, 128, 139, 130, 124, 302, 306, 299, 275, 197, 162, 186, 227, 228, 139, 134, 145, 219, 282, 258, 181, 142, 134, 119, 69, 29, 14, 24, 67, 85, 132, 155, 152, 148, 137, 301, 309, 304, 275, 193, 183, 288, 312, 260, 215, 194, 206, 266, 290, 274, 209, 138, 88, 54, 42, 45, 44, 64, 81, 109, 140, 163, 162, 154, 144, 283, 296, 303, 269, 196, 241, 376, 435, 389, 283, 220, 228, 242, 243, 230, 182, 142, 101, 77, 68, 82, 99, 110, 112, 125, 134, 145, 139, 132, 127, 254, 267, 287, 282, 229, 310, 414, 464, 385, 238, 171, 154, 149, 145, 144, 124, 108, 101, 102, 102, 108, 113, 118, 121, 127, 135, 139, 136, 135, 126, 190, 229, 265, 259, 262, 367, 447, 416, 257, 148, 111, 99, 97, 90, 93, 94, 92, 91, 98, 104, 109, 114, 117, 131, 138, 140, 140, 140, 136, 141, 131, 166, 216, 203, 269, 394, 442, 311, 177, 119, 109, 111, 103, 96, 96, 96, 94, 93, 100, 107, 113, 124, 138, 150, 149, 149, 146, 146, 161, 185, 128, 125, 155, 183, 279, 397, 387, 233, 145, 118, 114, 112, 105, 96, 94, 94, 97, 102, 108, 121, 129, 137, 148, 151, 148, 140, 149, 176, 203, 201, 132, 116, 115, 157, 274, 357, 312, 201, 131, 119, 120, 115, 108, 104, 102, 99, 102, 107, 118, 125, 133, 145, 146, 135, 126, 129, 169, 196, 184, 155, 140, 120, 113, 122, 216, 293, 231, 167, 127, 111, 118, 120, 117, 110, 104, 103, 112, 119, 126, 126, 125, 128, 125, 121, 128, 162, 188, 180, 137, 118, 138, 121, 117, 112, 134, 196, 157, 129, 102, 100, 114, 121, 121, 109, 106, 108, 118, 125, 133, 137, 126, 115, 111, 128, 162, 202, 199, 164, 96, 100, 136, 124, 115, 113, 106, 116, 107, 93, 75, 76, 86, 96, 106, 104, 104, 111, 126, 141, 151, 142, 122, 111, 116, 151, 203, 226, 207, 154, 98, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 23, 16, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 0, 5, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 13, 18, 5, 14, 14, 9, 2, 0, 0, 0, 0, 9, 11, 9, 3, 0, 0, 0, 0, 0, 0, 0, 16, 19, 0, 0, 0, 0, 0, 9, 23, 23, 16, 26, 25, 9, 7, 0, 0, 0, 0, 18, 19, 15, 0, 0, 0, 0, 0, 0, 0, 0, 33, 28, 14, 0, 0, 0, 0, 14, 39, 39, 30, 26, 31, 12, 2, 1, 0, 0, 0, 27, 27, 17, 2, 0, 0, 0, 0, 0, 0, 0, 39, 35, 25, 0, 0, 0, 0, 20, 35, 32, 16, 22, 32, 22, 5, 3, 0, 0, 7, 31, 35, 18, 5, 0, 0, 0, 0, 0, 0, 0, 36, 42, 39, 0, 0, 0, 0, 0, 10, 16, 24, 29, 37, 28, 13, 6, 0, 0, 20, 41, 37, 17, 2, 0, 0, 0, 2, 0, 0, 0, 34, 41, 46, 6, 0, 0, 0, 0, 0, 2, 26, 42, 37, 22, 17, 21, 3, 0, 24, 42, 30, 18, 10, 0, 0, 1, 4, 0, 0, 0, 41, 45, 47, 23, 0, 0, 0, 0, 0, 10, 41, 74, 53, 31, 16, 11, 4, 6, 20, 35, 32, 11, 0, 0, 0, 0, 1, 0, 0, 0, 49, 48, 52, 38, 0, 0, 0, 0, 0, 17, 33, 34, 33, 16, 15, 8, 0, 0, 14, 22, 23, 21, 13, 2, 0, 0, 0, 0, 0, 0, 61, 54, 56, 45, 17, 0, 2, 1, 0, 16, 36, 27, 15, 3, 11, 2, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 67, 63, 63, 52, 37, 10, 7, 3, 14, 8, 4, 15, 6, 6, 20, 7, 0, 0, 7, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 64, 64, 53, 39, 20, 19, 11, 12, 15, 0, 0, 0, 4, 27, 21, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 61, 58, 55, 42, 28, 32, 48, 16, 0, 0, 0, 7, 28, 34, 28, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 55, 53, 56, 39, 18, 26, 59, 68, 31, 24, 26, 40, 47, 52, 39, 17, 15, 13, 5, 0, 0, 5, 13, 0, 0, 0, 0, 0, 0, 58, 58, 56, 58, 42, 27, 49, 56, 58, 55, 30, 26, 41, 44, 50, 40, 13, 5, 12, 13, 12, 10, 16, 24, 28, 34, 40, 42, 43, 42, 51, 56, 60, 58, 41, 36, 65, 86, 87, 55, 42, 47, 53, 54, 57, 53, 40, 29, 26, 22, 27, 34, 40, 43, 50, 52, 51, 50, 53, 52, 59, 47, 54, 57, 28, 43, 76, 104, 98, 71, 57, 53, 54, 51, 55, 51, 41, 39, 41, 40, 43, 45, 49, 52, 54, 56, 55, 55, 55, 52, 67, 57, 50, 51, 40, 61, 93, 103, 77, 56, 42, 38, 38, 33, 35, 36, 35, 37, 42, 45, 47, 49, 50, 55, 53, 54, 56, 58, 58, 63, 56, 51, 49, 35, 41, 72, 104, 87, 65, 46, 43, 43, 40, 37, 38, 39, 39, 39, 42, 47, 49, 54, 57, 57, 54, 56, 57, 62, 67, 70, 59, 50, 50, 42, 40, 77, 101, 73, 54, 43, 41, 44, 43, 37, 37, 38, 41, 43, 46, 53, 53, 53, 58, 61, 62, 61, 67, 73, 72, 64, 63, 55, 49, 50, 53, 63, 86, 59, 44, 41, 45, 45, 44, 43, 40, 40, 42, 46, 50, 55, 59, 61, 60, 58, 60, 65, 75, 74, 67, 56, 67, 58, 54, 50, 61, 64, 60, 54, 41, 35, 39, 41, 43, 43, 42, 45, 50, 52, 53, 56, 56, 55, 54, 54, 61, 73, 80, 80, 67, 49, 65, 58, 56, 51, 50, 61, 53, 49, 40, 38, 41, 40, 39, 36, 37, 39, 45, 50, 57, 59, 54, 50, 49, 52, 63, 80, 84, 73, 49, 46, 62, 57, 53, 51, 44, 41, 41, 38, 34, 32, 36, 39, 43, 36, 31, 34, 41, 47, 52, 52, 49, 46, 43, 51, 64, 76, 80, 67, 49, 45, 19, 24, 31, 36, 32, 32, 33, 29, 25, 31, 37, 40, 34, 23, 21, 17, 17, 11, 8, 0, 0, 0, 0, 8, 17, 15, 7, 0, 0, 0, 10, 19, 27, 36, 35, 38, 37, 33, 36, 70, 80, 71, 45, 24, 29, 34, 16, 12, 0, 5, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 18, 29, 34, 37, 36, 35, 36, 31, 41, 129, 157, 157, 76, 35, 26, 4, 0, 0, 27, 67, 69, 54, 12, 0, 0, 0, 0, 0, 0, 0, 22, 32, 32, 34, 30, 29, 28, 25, 29, 86, 125, 132, 51, 0, 0, 0, 0, 9, 77, 126, 128, 106, 81, 44, 3, 0, 0, 0, 3, 2, 0, 0, 0, 10, 31, 30, 29, 26, 26, 53, 41, 57, 34, 0, 0, 0, 0, 49, 117, 158, 142, 114, 93, 71, 34, 0, 0, 0, 0, 12, 0, 0, 0, 0, 29, 27, 29, 32, 26, 24, 28, 53, 66, 53, 30, 14, 22, 59, 125, 174, 151, 100, 75, 64, 19, 0, 0, 0, 0, 9, 57, 34, 10, 43, 41, 29, 37, 63, 45, 46, 55, 106, 131, 98, 55, 28, 28, 32, 80, 134, 147, 98, 51, 31, 14, 0, 0, 0, 0, 0, 157, 135, 123, 126, 70, 32, 92, 175, 226, 200, 175, 172, 175, 117, 66, 23, 5, 6, 45, 96, 152, 126, 66, 32, 19, 11, 0, 0, 0, 0, 229, 215, 211, 172, 97, 21, 117, 243, 361, 343, 285, 221, 198, 141, 76, 44, 0, 0, 64, 139, 205, 156, 104, 60, 36, 34, 0, 0, 0, 0, 239, 232, 258, 202, 122, 35, 69, 189, 305, 334, 298, 259, 230, 169, 102, 60, 0, 18, 112, 211, 260, 165, 104, 52, 54, 53, 26, 0, 0, 0, 247, 217, 255, 219, 137, 58, 53, 116, 183, 248, 254, 264, 272, 222, 129, 102, 30, 74, 148, 252, 258, 147, 84, 42, 41, 48, 46, 18, 2, 0, 259, 228, 240, 196, 107, 61, 37, 92, 113, 205, 219, 287, 309, 277, 178, 128, 70, 122, 177, 253, 234, 127, 66, 28, 23, 35, 54, 52, 42, 0, 280, 254, 251, 170, 72, 51, 26, 60, 67, 184, 244, 302, 287, 265, 208, 151, 82, 130, 180, 246, 228, 143, 88, 54, 40, 56, 83, 84, 60, 14, 308, 275, 269, 181, 92, 54, 47, 66, 68, 217, 321, 353, 288, 200, 171, 141, 85, 114, 162, 227, 202, 132, 73, 46, 50, 81, 97, 79, 54, 10, 335, 304, 305, 216, 149, 85, 97, 63, 91, 175, 275, 303, 226, 148, 113, 92, 68, 114, 132, 190, 191, 144, 73, 39, 37, 63, 70, 48, 32, 17, 362, 330, 336, 254, 179, 125, 135, 113, 91, 113, 167, 143, 121, 99, 70, 80, 82, 89, 68, 98, 107, 110, 59, 1, 0, 22, 39, 41, 41, 41, 381, 351, 348, 282, 207, 147, 158, 166, 132, 66, 88, 79, 102, 116, 93, 95, 91, 111, 95, 57, 41, 44, 0, 0, 0, 0, 25, 53, 52, 41, 367, 355, 346, 298, 221, 170, 139, 179, 179, 89, 82, 56, 127, 170, 170, 137, 97, 92, 126, 104, 44, 0, 0, 0, 0, 43, 52, 74, 61, 39, 332, 348, 337, 304, 235, 201, 191, 190, 168, 90, 72, 63, 156, 227, 256, 205, 109, 49, 44, 25, 0, 0, 0, 0, 7, 62, 69, 69, 52, 31, 297, 349, 331, 294, 219, 206, 261, 351, 316, 199, 169, 186, 265, 331, 333, 271, 189, 72, 6, 0, 0, 0, 0, 21, 40, 64, 77, 70, 56, 40, 283, 358, 337, 295, 228, 248, 325, 457, 485, 362, 267, 240, 267, 285, 270, 217, 157, 88, 38, 9, 16, 36, 69, 82, 82, 86, 87, 79, 76, 59, 236, 324, 343, 320, 286, 338, 415, 504, 435, 333, 200, 131, 127, 124, 120, 104, 87, 59, 56, 62, 73, 79, 89, 100, 106, 107, 111, 111, 110, 101, 138, 218, 288, 293, 313, 378, 458, 471, 359, 204, 107, 80, 74, 74, 71, 64, 66, 60, 61, 67, 79, 89, 95, 111, 124, 133, 132, 128, 128, 127, 116, 126, 194, 237, 309, 387, 452, 389, 247, 120, 93, 89, 88, 82, 77, 70, 65, 65, 67, 76, 88, 99, 116, 135, 149, 154, 151, 148, 160, 173, 129, 109, 117, 167, 297, 409, 426, 316, 163, 96, 103, 99, 93, 83, 77, 72, 71, 73, 82, 95, 112, 130, 141, 145, 142, 134, 143, 164, 194, 213, 134, 109, 100, 116, 260, 382, 387, 269, 139, 99, 109, 103, 92, 79, 78, 82, 86, 91, 102, 107, 117, 131, 142, 139, 121, 119, 144, 177, 197, 193, 136, 113, 107, 111, 176, 283, 278, 225, 113, 105, 113, 114, 115, 96, 85, 80, 88, 99, 109, 116, 118, 116, 117, 119, 121, 139, 161, 177, 143, 123, 148, 122, 112, 115, 124, 143, 139, 130, 64, 67, 88, 106, 120, 116, 109, 104, 109, 117, 122, 118, 113, 106, 103, 116, 149, 187, 206, 182, 113, 87, 153, 125, 114, 116, 111, 99, 64, 64, 42, 35, 45, 60, 73, 85, 99, 112, 131, 148, 154, 143, 123, 103, 107, 139, 201, 246, 239, 182, 120, 77, 149, 128, 110, 112, 99, 90, 65, 47, 36, 30, 31, 40, 33, 31, 42, 65, 101, 139, 160, 155, 130, 103, 117, 154, 218, 252, 233, 167, 105, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 5, 12, 19, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 10, 0, 0, 0, 0, 13, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 15, 0, 0, 10, 18, 18, 20, 40, 30, 12, 0, 0, 0, 0, 0, 11, 22, 1, 0, 0, 1, 12, 9, 0, 0, 0, 0, 0, 0, 70, 64, 0, 0, 0, 12, 0, 12, 59, 52, 27, 19, 14, 4, 0, 0, 0, 30, 34, 0, 0, 0, 13, 46, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 0, 9, 69, 73, 22, 6, 21, 37, 17, 0, 0, 16, 53, 21, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 14, 10, 69, 112, 50, 0, 5, 41, 25, 1, 0, 0, 47, 45, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 7, 32, 21, 48, 115, 88, 0, 0, 5, 21, 2, 0, 0, 18, 64, 25, 0, 20, 12, 0, 0, 0, 38, 52, 0, 0, 0, 32, 0, 0, 0, 14, 16, 23, 87, 71, 1, 0, 0, 8, 9, 0, 0, 0, 48, 60, 7, 77, 24, 0, 0, 0, 105, 193, 88, 0, 22, 30, 0, 0, 0, 0, 0, 20, 100, 44, 0, 0, 0, 22, 19, 0, 0, 0, 0, 46, 35, 123, 47, 0, 0, 0, 59, 209, 164, 34, 57, 57, 0, 0, 0, 0, 0, 30, 142, 49, 4, 0, 0, 37, 38, 11, 0, 0, 0, 0, 24, 130, 58, 0, 0, 0, 0, 119, 140, 41, 69, 90, 0, 0, 0, 0, 0, 47, 161, 54, 0, 0, 0, 30, 48, 34, 16, 0, 0, 0, 17, 125, 27, 0, 2, 0, 0, 64, 102, 39, 56, 92, 34, 0, 0, 11, 0, 75, 148, 45, 0, 0, 0, 12, 28, 33, 26, 0, 0, 0, 28, 122, 0, 0, 7, 3, 0, 14, 69, 81, 62, 42, 41, 34, 23, 10, 0, 85, 144, 47, 0, 0, 0, 14, 23, 31, 32, 0, 0, 0, 33, 105, 3, 0, 0, 26, 0, 0, 54, 135, 116, 17, 8, 54, 58, 26, 0, 64, 121, 58, 10, 0, 0, 33, 56, 49, 39, 6, 0, 0, 32, 93, 37, 0, 0, 56, 0, 0, 49, 159, 160, 78, 33, 42, 44, 29, 1, 41, 81, 85, 47, 0, 0, 29, 69, 63, 32, 0, 0, 0, 32, 87, 70, 0, 0, 80, 42, 0, 6, 88, 89, 64, 14, 20, 13, 14, 25, 17, 2, 64, 84, 24, 9, 36, 51, 49, 14, 0, 0, 0, 45, 77, 80, 0, 0, 72, 92, 0, 0, 0, 44, 50, 5, 27, 0, 0, 64, 26, 0, 0, 30, 19, 10, 22, 10, 11, 7, 0, 0, 0, 63, 66, 79, 22, 0, 41, 90, 39, 4, 0, 38, 65, 43, 63, 0, 0, 40, 70, 50, 28, 0, 12, 20, 46, 19, 7, 3, 0, 0, 0, 81, 49, 73, 42, 0, 37, 84, 0, 0, 0, 7, 25, 48, 64, 0, 0, 0, 28, 60, 51, 20, 6, 17, 53, 56, 53, 29, 0, 1, 4, 103, 37, 65, 40, 0, 53, 138, 7, 0, 0, 0, 44, 95, 101, 66, 8, 0, 0, 0, 4, 15, 9, 18, 31, 54, 67, 55, 32, 31, 36, 148, 66, 67, 26, 0, 55, 150, 94, 6, 0, 56, 141, 166, 163, 149, 98, 64, 32, 13, 14, 31, 53, 63, 62, 69, 75, 75, 60, 56, 59, 192, 145, 108, 46, 4, 106, 136, 96, 66, 41, 76, 108, 112, 108, 107, 84, 65, 60, 64, 67, 66, 71, 77, 78, 72, 73, 81, 72, 70, 70, 140, 178, 170, 87, 76, 153, 126, 63, 23, 32, 48, 52, 52, 50, 56, 61, 62, 63, 69, 77, 74, 72, 73, 76, 70, 66, 71, 69, 66, 65, 60, 126, 177, 113, 122, 159, 93, 5, 21, 60, 61, 63, 62, 63, 63, 61, 60, 60, 64, 70, 69, 67, 72, 80, 81, 82, 86, 79, 71, 73, 53, 77, 123, 138, 193, 182, 40, 0, 23, 65, 70, 63, 60, 65, 64, 60, 59, 62, 67, 74, 80, 83, 85, 84, 88, 94, 101, 96, 93, 102, 62, 68, 77, 121, 234, 230, 34, 0, 39, 62, 72, 58, 46, 56, 66, 70, 73, 73, 76, 79, 86, 99, 97, 82, 77, 83, 102, 109, 103, 113, 61, 76, 78, 85, 186, 245, 89, 20, 70, 77, 86, 72, 52, 46, 54, 65, 72, 73, 77, 76, 75, 85, 90, 85, 74, 83, 93, 87, 65, 93, 55, 79, 86, 74, 96, 162, 101, 50, 68, 90, 102, 98, 89, 69, 61, 63, 64, 64, 61, 61, 65, 71, 78, 85, 85, 83, 64, 48, 29, 74, 53, 76, 87, 78, 63, 71, 69, 51, 48, 71, 83, 89, 97, 93, 96, 99, 92, 82, 65, 49, 52, 60, 77, 101, 112, 93, 61, 49, 48, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
