library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=3
    -7676, 60, -270, 3599, 7729, -6459, 4506, -5844, 5911, -1946,

    -- weights
    -- layer=3 filter=0 channel=0
    3, 13, 28, 3, 13, 26, 17, 15, -26, 17, -39, 21, -51, 1, 5, -9, -60, -8, -33, -34, 4, 32, -29, 28, -47, -19, 13, -8, 32, 19, 13, 17, 7, -63, 50, -13, 14, 2, 27, 0, -21, 4, 37, 46, -48, -3, -17, 16, 19, -41, -16, 20, 0, -24, -22, -17, -13, -37, 48, 26, 8, 0, -1, 1, -40, -25, 46, -19, 16, 26, 19, 0, -52, 2, 37, 6, 2, -16, -12, 31, 7, -34, -37, 24, 0, 14, 3, -41, -39, -43, 35, -4, 23, -39, -35, 14, 21, 29, -1, -53, -6, 38, -13, 9, -49, 0, -50, -36, 9, -27, 22, -15, 1, 38, -8, -31, 16, -79, 31, 34, -3, -8, -10, 9, -37, 40, -10, -36, -24, -17, -3, -56, 27, 16, -16, 24, -7, -76, 39, -13, 0, 22, 20, -52, -17, -26, -7, 25, 23, -15, 18, -14, 20, -24, -34, -2, -10, 7, -75, 8, -23, 26, -37, -27, 41, -14, 45, 15, 10, -46, -33, 23, 17, 5, 36, -54, -12, -39, -1, 43, -26, -47, -2, 12, 15, -4, -11, -29, -28, -18, 2, -5, -31, 20, -21, -31, 52, -41, 25, 52, -62, 56, -23, 15, -93, -69, -9, 35, 52, -30, 52, 27, 10, 12, -40, -43, 23, -39, -2, -8, 5, -26, 27, 12, -8, 31, -17, -33, -22, -42, 11, 26, -61, 24, -5, -9, 32, 11, 8, 40, 31, 1, 1, -18, -1, 24, 19, -11, 36, -13, 28, 21, -32, -2, 7, -25, 13, 7, 0, -14, 21, -26, 20, 15, -42, 21, -93, 29, -9, -41, -7, 4, 33, -15, 0, 15, -11, 22, -29, -6, 45, 10, -34, 28, 29, 32, -37, 21,
    -- layer=3 filter=0 channel=1
    25, 18, -22, -26, -35, 12, -4, -20, -56, 27, -8, 14, 3, 29, -9, 8, -13, -1, 21, 0, -47, -19, -1, -25, 66, 13, 10, 11, -20, -4, -7, 33, -58, -50, 4, -28, 0, 40, -21, -6, -6, 0, 13, 26, -12, 43, -9, -7, -20, 13, 59, -18, -32, -18, -29, 13, 37, -31, -60, 8, -32, 46, -74, -4, 9, 21, -22, -4, 19, 6, -19, -37, 43, 2, -53, 9, -11, 33, 43, -6, -17, 45, -10, -25, 3, 29, -1, -29, 15, -8, 22, -4, -6, 21, -9, -25, -41, 43, 0, -45, 10, 5, -6, 32, -83, -17, 8, -18, -20, -13, -25, 9, -86, -6, 43, -5, -2, -9, -46, 25, -7, 4, -76, 39, 27, 41, 61, -24, -66, -9, 26, -73, 34, -4, 65, 99, -67, -4, 0, -11, -11, -44, -3, 19, -76, -62, 24, 15, 61, 29, -20, 64, -9, 7, -79, -6, 3, -3, 49, 22, -41, -3, -32, -35, -27, 43, 22, -4, -63, -48, -5, 33, -96, -45, 33, -18, -50, -23, 20, 45, 37, -17, 19, 2, -8, 15, -59, 1, -28, 37, 25, -28, -14, -1, 39, -44, -54, 15, 60, -36, -73, -41, -27, -49, 0, 61, 43, -19, -105, 40, -11, 32, -41, -34, 26, 47, -7, -27, 19, -34, 6, 90, -13, 32, 20, 12, 54, -32, 33, 78, -17, -12, -42, -61, -42, -25, 40, 39, 28, -3, -46, -45, -11, 23, -34, 0, 31, -17, -7, 15, 30, 13, -19, 4, 36, -35, 12, 24, -14, -63, -64, 11, 23, 17, -35, -25, 37, 16, 60, -13, 45, 2, -40, -42, 39, 11, 5, -20, 28, -22, -16, 17, 11, -82, 3, 16, -14, 20,
    -- layer=3 filter=0 channel=2
    -25, -11, 2, 17, 8, -27, 54, 17, 38, 20, 44, 12, -1, 2, -32, 27, -2, 12, -10, -23, -3, -11, -39, -6, 19, -15, 15, -26, -33, 8, -14, 13, 3, 17, -7, 20, -6, 38, -28, -10, 24, 25, 40, 20, -3, -12, 2, 21, -39, -11, -4, 10, 19, -16, -1, -25, -8, -23, -37, 25, 10, -13, -57, 23, 33, -21, 15, -22, -26, -39, 30, 28, 46, -3, -50, 45, -10, 8, -46, 12, -40, -28, -25, 10, 6, 1, 9, -28, -58, 30, 8, -25, -3, -17, -14, -14, -16, -28, 43, 0, 7, -30, 19, -14, 3, -9, 17, 31, -39, 37, -20, 20, 19, 28, -37, 1, 46, -46, -16, 19, 35, 19, 46, 44, 9, -10, -12, 33, -38, 31, 35, 1, 5, 4, -40, -25, 62, 23, 25, -15, 15, 2, -6, -34, 34, -42, -18, -15, -66, 20, -40, 27, 23, 23, 22, -41, -11, 3, -40, 16, 35, -61, 9, -10, 42, -13, 62, 21, 48, 10, 36, -19, 47, 14, -11, -25, -3, -9, -9, 10, -34, -8, -44, -34, -35, 21, 32, -5, -31, -15, -23, -20, -32, -52, -35, -12, 30, -42, -11, 17, -28, -17, 11, 34, -34, 20, -62, 42, 9, -36, -19, -40, 45, 40, -47, -5, 13, 17, -32, 33, -28, -36, -44, 22, 0, -12, 1, -14, -52, -21, -12, 7, 49, 22, -4, -45, 24, 0, 1, 26, 18, -13, -39, -13, 0, 65, -21, -18, -16, 1, -52, 27, 7, -45, 1, -33, 37, -33, -7, 36, 50, -39, 27, 25, 43, -27, -82, 12, -35, -6, -4, 15, -1, -38, -30, 34, -36, 18, -29, 27, 12, -12, -33, 27, -25, 3, -64, 16,
    -- layer=3 filter=0 channel=3
    26, 7, -7, 24, -23, -9, -33, -31, 32, 6, 18, -47, 31, 14, 0, 15, 16, 18, -10, -16, 1, 31, 9, -50, -14, -31, 27, -5, 20, -1, 22, 22, 17, 0, -6, 5, -11, 3, 16, -3, 16, 17, 53, 20, 50, 13, 0, 0, -40, 9, -34, 1, 3, -34, -8, 0, 28, -19, -21, -5, -26, 4, 12, -19, -15, 0, -7, 41, 2, -8, -3, -24, -17, 27, -11, 2, 55, 28, -16, 8, -34, 7, -14, -5, 4, -20, 18, 11, 47, -14, 41, -2, -19, -10, 7, 1, 20, -21, 16, 20, -6, -42, -29, -1, 15, 8, 56, 23, 34, -38, -32, -16, -7, 2, 29, -10, -47, 14, -9, 0, -10, 39, -18, 8, -23, -16, -18, 15, 31, -47, 21, 41, -35, -33, -29, 3, 20, 6, 45, -9, 19, 8, -67, 4, -29, 4, -10, -35, -43, 21, -14, 28, 18, 11, 3, 5, 23, -17, -31, -32, 34, -11, 30, 34, -1, -12, 16, 37, -1, -10, -2, 17, -11, 14, -16, -7, 12, 28, -42, 7, -53, 15, -11, -19, -21, -28, 43, 21, -15, -7, -31, 1, 9, -37, -37, -9, 32, 5, -52, -28, 42, -12, 11, 23, 61, 20, 7, 8, -40, -21, 22, -39, 28, 22, 13, 8, -43, -13, 13, 12, -31, -12, -53, -34, -23, -6, -19, -3, 29, -50, -2, -27, 22, 15, -10, 21, 22, 14, -45, -7, -56, 35, -21, 12, 26, -38, -5, 2, -46, 9, -15, 9, -2, -3, -13, 24, -35, -39, 1, -13, 34, -19, -40, -13, 38, -14, -40, 20, -7, 8, -31, -31, 11, -6, -36, -39, -14, 6, 17, 17, -25, -5, 49, -13, 24, -12, -35, -23,
    -- layer=3 filter=0 channel=4
    8, 26, -37, 28, -3, -3, 19, 48, -34, -28, 5, -45, -54, 26, -4, -5, -47, -6, -1, -7, -54, -17, -1, 53, -6, 0, 1, -7, 4, -34, 31, 24, 24, -61, -8, -9, 18, 5, 32, 20, -51, 0, -13, -19, -39, 18, -3, 33, -4, 35, -33, 13, -32, -35, 6, -30, -14, 29, 2, 29, -14, -65, 29, 11, 2, -53, -2, -33, -26, -37, -21, 11, -83, 15, -13, -46, -30, -5, 4, 2, 7, -13, -1, -21, 26, -43, 2, 10, 41, 41, -17, -34, -5, -79, 15, 2, 3, 3, 9, 37, -13, -7, 17, 28, -20, -30, -5, 25, -67, -39, 2, 20, 22, -33, -37, 17, 6, -15, 25, -3, -29, -24, 0, 13, -33, 21, -25, 31, -12, -2, 1, 47, -46, -22, -8, -10, 10, 29, 3, -6, -7, -4, 34, -22, -24, 5, 3, -41, 6, 19, -12, 15, -16, -25, -28, -28, -3, 7, -53, -2, -18, -6, 15, 2, 26, -9, 4, 30, -63, -10, -6, 28, 7, -16, -59, 17, -5, -37, 14, -24, -7, 9, 8, -9, -33, -5, -28, 16, 0, -27, -11, 29, -28, -14, -1, -33, 54, -26, 11, -5, 0, 4, 9, 9, -15, 33, -10, 44, 4, 0, 13, 14, 26, 1, 20, 23, 23, 47, 20, 34, -8, -30, 14, -25, 29, -35, -14, 15, -60, 18, 2, -33, 36, 24, -10, -13, 30, 11, -95, 37, -43, 9, -19, -68, 23, 21, 2, -47, 20, 10, 73, -3, 0, 2, -27, 13, -1, 13, 23, 39, 38, -57, -13, 10, -35, 12, -91, -18, -34, -12, -54, 34, -33, 41, -3, 13, 55, 15, -39, 17, -4, 40, 21, 1, 0, 24, -19, -32,
    -- layer=3 filter=0 channel=5
    5, -31, -44, 29, -7, 5, 31, -34, 67, 11, 5, -35, 66, -17, 8, 5, 50, -25, -37, -7, 37, 5, -37, -17, 11, -36, 7, -51, -28, 23, -20, -1, -1, 41, 18, -14, 49, 8, -40, -10, 58, -5, 6, -11, 0, 0, -7, 35, 50, -19, 1, -21, 4, -3, -49, -12, 29, -10, -51, 18, 4, 40, -4, 35, 24, 13, -12, -38, -13, 7, 39, 1, 21, -52, -6, -29, 22, -26, -51, 13, -40, 23, 14, -42, -18, 43, 19, -38, -2, 17, 31, 24, 11, 10, 21, 5, 4, -18, -23, 25, 2, 8, -28, -42, 48, 29, -17, -1, 41, -9, -72, -5, -8, -6, -23, 1, -22, -20, 10, 12, 42, -15, 0, 15, 11, -68, 29, -32, 17, 4, 5, 8, -44, -17, -43, -7, 21, 27, -7, -2, 16, 44, -8, -46, -26, 29, 43, -40, -64, -22, -22, 8, 18, -48, 29, -17, -31, 9, -15, 3, 43, -4, 36, 30, -35, -22, -20, 0, 20, 29, 2, 8, 33, 36, -16, 18, 4, 69, -30, -25, -18, -3, -8, -34, -16, 8, 36, 3, 13, -36, 12, -31, 37, -72, -42, 30, 34, -64, 18, -27, 57, 2, -22, 39, 20, 5, -6, -17, 8, -39, 4, 13, -31, 6, -48, -31, -9, 11, -10, -13, -2, -16, -9, 33, 0, -12, 9, 12, -28, -20, -14, -24, 14, -10, -9, 28, -22, -28, -24, -33, -11, 34, 8, -1, 17, 46, -38, -27, -31, -7, 2, 43, -17, -8, -13, -31, -20, -29, 62, -3, -14, -44, -14, -10, 4, -9, 9, -22, -11, 10, 0, -37, -45, -2, -39, -61, -2, -2, -40, -53, -35, -8, 62, 57, -33, -29, -24, 27,
    -- layer=3 filter=0 channel=6
    0, 23, -24, 31, -15, 16, 7, -3, -26, -36, -11, -5, 13, -21, -18, 28, -72, 21, 6, -7, -9, -72, -11, -52, -38, 14, -16, 26, -12, 8, -49, -15, 24, 36, 8, 14, 41, -59, 21, -3, -99, -19, -12, 22, 10, -34, -1, 38, -86, -7, 20, 57, 74, -22, -36, -20, 33, 31, 10, -14, 1, -39, -1, 25, -25, -41, -57, 43, 7, -31, 23, -16, -58, 24, -34, 16, -18, 5, -5, 22, -8, -31, 42, -19, -14, -50, -37, -8, 74, -31, -54, 19, 27, -20, 20, 19, 35, 11, 35, 35, -28, -13, -29, 52, 31, -9, -45, -39, 75, 30, 8, -4, -7, -4, 23, -28, 18, -15, 25, -34, -51, 46, -7, 34, -21, 30, -63, -33, -6, 2, -20, 20, 5, -48, 82, -9, -60, 47, -52, 16, -4, -11, -36, 61, -61, 29, -54, 22, -24, 16, 4, -61, -16, 105, -20, -5, -6, -30, -9, 2, -33, 0, -47, 16, -12, -12, -30, -32, 0, 23, -57, 9, 31, 58, 4, 16, -51, -49, 6, -53, -33, -17, -45, -56, 88, 2, 21, -62, 0, -37, 10, 11, -6, -17, -35, -6, -50, 13, -62, 28, -3, 11, -45, 13, -50, 22, -31, 16, -61, 29, -25, -52, -1, -53, 22, 23, 11, -12, -16, 16, -4, -13, -35, -6, -5, 2, -38, 39, -41, 21, -48, -12, 0, 1, -80, 2, -24, 30, 41, 3, -28, 24, 2, -23, 28, -3, -25, -5, 20, -5, -11, -29, -29, -6, -26, -10, 21, -8, -37, 0, -25, 7, -44, 78, -31, -37, -81, -25, 26, 18, -55, 13, -54, -12, -31, -44, -17, 1, -7, -3, 5, 20, 8, -59, -30, -56, 8, -26,
    -- layer=3 filter=0 channel=7
    -12, 0, 12, -1, -13, 12, -13, 16, 0, -51, -48, -17, -17, -49, 19, -54, -13, -5, -33, -33, -8, 63, -36, 24, 46, 3, -48, -32, 17, -2, -30, 10, 51, -39, 31, 18, -43, 0, -13, 14, 49, -43, 14, 8, 45, -39, 15, -26, -44, -7, 30, -51, -38, 53, -35, -25, -21, -48, -19, -34, -3, -54, 2, -34, -22, 22, 37, -27, -19, 36, -13, -22, -1, -58, 21, 14, 8, -24, 35, -22, 6, -19, 36, 21, 24, -2, -38, 37, -73, -40, -41, 1, -23, -13, 5, 16, -13, 29, 21, 42, -11, -10, 36, -51, 4, -13, 16, -8, 0, -5, -26, -5, 15, -42, -27, -3, -38, -14, -24, -43, 38, -84, 43, -7, 3, -7, -13, -8, 53, 17, -4, -51, 0, 30, -66, 4, 4, 4, -46, -5, -81, 47, -39, -8, 33, 9, 9, -26, 10, -27, -27, -34, -13, -129, 13, 53, 24, 45, -81, 13, 58, 20, 9, -7, -33, 45, -5, 18, -3, 55, -44, -18, 24, 23, -13, -10, 27, 16, -25, -59, 6, 52, 1, -53, 15, 17, -1, 48, -14, -33, -38, -16, 11, 13, 3, -2, -67, -38, 30, -48, -4, 29, 19, -22, 19, 18, 51, 7, 91, 38, 28, 0, -36, -22, -20, -55, 39, 46, 12, -10, 8, -81, 44, -17, -26, -46, 3, 29, -77, -51, 33, 7, -18, 24, 24, 19, -17, 1, 4, 48, 36, -5, -36, 8, 13, -28, -46, -37, 33, 53, 11, -24, -3, -60, 3, 36, 6, 35, -24, 41, -7, 4, 4, -5, 22, -12, -51, 20, -15, 24, -11, 57, -33, 33, -25, 40, -33, 17, 17, -38, 51, 34, 50, 0, -10, -44, 14, 33,
    -- layer=3 filter=0 channel=8
    23, 12, 25, -49, 46, -12, -27, 22, -104, 24, 31, 20, -141, -25, 35, 0, -18, -17, 31, -24, 17, -23, -11, 14, 9, -24, 37, -6, -6, -39, -34, -23, 2, -10, 37, 25, 29, 10, -6, -35, -58, 49, -1, 20, -75, 15, 19, 10, -40, -14, 26, 1, 4, -21, -1, 57, -19, -24, 32, 18, 11, -31, -55, 1, -5, -45, 26, -34, 12, -11, 33, 35, -77, 28, 21, 2, -33, 7, -15, 20, -63, -74, -1, 18, -16, -26, -13, 37, -9, 3, -12, 35, 12, 13, -6, 6, -7, -29, -7, -26, 50, 26, 17, 6, -44, -7, 31, 17, 1, -28, 34, -52, -53, 1, -19, -20, 50, 18, 31, -8, -29, 44, -9, -19, 3, -6, -35, 26, -38, 32, 0, 13, 18, -19, -50, -7, -71, -16, 19, 32, -8, 9, 26, -58, 3, 4, 2, 2, 3, -19, 6, -48, 11, 12, 19, -12, -21, 66, -1, 29, -16, 8, 43, -2, 34, -6, -24, -46, -82, 17, 92, 9, -72, 0, 14, -29, -65, -26, 12, -13, 4, 1, -38, 1, -63, -50, -44, -3, -29, 42, -27, -18, 6, 3, -22, -7, 57, 1, -23, -9, 46, -18, 0, -21, 43, -90, 2, -77, -53, 0, 18, 54, -22, -18, 0, 12, -59, -19, 12, 3, 4, 30, -84, 5, -103, -25, 33, -46, 105, -3, 2, 42, -25, -10, 72, 13, -27, -100, 10, 68, -26, 9, 20, 72, 2, -19, 26, 8, -50, 37, -82, 40, 27, 64, -8, -1, -70, -53, 19, -18, 40, -28, -65, 35, 6, 20, 34, -26, -17, -31, 11, -41, -48, 17, 33, -15, -59, -16, -37, -7, -54, -49, -7, 4, -11, -11, -11, 3,
    -- layer=3 filter=0 channel=9
    31, -3, 49, -2, -12, 18, 0, 9, 45, 16, -25, 17, -26, 3, 18, -50, -2, 1, 25, 34, -20, 40, -5, 32, -24, 28, 5, 43, 31, -20, -34, -9, -9, 26, 18, -29, -15, -10, -31, 6, 16, 10, 11, -34, -14, -29, 11, 5, -33, 40, 41, 7, -8, 27, 2, 12, -26, 13, -32, 19, -20, -20, 3, -30, 41, 8, 54, -17, 32, 6, -36, 43, 26, 27, -44, -6, 10, -4, 60, -13, 16, 17, 27, 1, 0, 33, -6, -29, -56, 9, 3, 11, 32, 8, -24, -16, 19, -13, 17, -33, -3, 0, -3, -1, -40, 34, 10, -44, -35, 11, -12, -3, -20, -36, 7, 17, -5, 6, -7, -9, 1, -7, -50, -33, -11, -36, 31, -9, 16, -15, 29, -1, -1, 19, 46, 45, -6, 31, -67, 18, -4, -18, -35, 26, 25, 15, 12, 16, -20, -28, 23, -76, -2, 24, 19, 2, 24, -39, 37, 28, -22, -25, 32, 3, 11, 33, 1, -31, -11, -15, 1, 7, -71, 8, 44, 24, 24, 43, 19, 33, 38, 24, 7, 10, -10, -61, 3, -6, 24, 26, 13, 30, -20, 34, -20, -53, -49, 23, -4, -85, -85, -80, -1, -90, -27, 58, -22, -80, -54, 11, -7, 0, -43, 19, -30, 41, 58, -17, -53, -57, -26, 37, -5, -25, -35, 0, 28, -43, -23, 50, -22, 16, -56, -57, -3, 1, 46, 40, -2, -9, -52, -47, 38, 8, -34, 4, 14, -23, 10, 12, 28, 3, -8, -14, -28, 13, -35, 14, -11, -12, -16, 73, -28, -70, -28, -75, 30, -52, 39, -6, 16, -37, -73, -34, 51, -39, -17, -33, -23, -14, 58, 19, -36, -51, 28, 16, -7, -26,

    others => 0);
end iwght_package;
