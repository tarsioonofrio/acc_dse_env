library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=4
    -3455, -4615, 3456, 2032, 18894, -13794, 13410, -13876, 9478, -12687,

    -- weights
    -- layer=4 filter=0 channel=0
    21, -9, -59, 77, 7, 5, 67, 80, -24, 20, 105, 47, 39, -95, -48, 90, -102, 50, -17, 38, -38, -30, 10, -7, -83, -21, -59, -44, 7, 9, 101, -11, 59, 99, 38, -78, -5, -35, -65, 17, 79, -37, 25, -6, -90, 49, -62, -109, -41, -25, -126, 138, 39, -15, -25, -11, -43, 35, -26, 3, 74, -34, 0, -119,
    -- layer=4 filter=0 channel=1
    65, 119, -41, 38, -55, 104, -73, 42, 133, 133, -9, 92, -42, -93, 38, -67, -87, -92, -43, 66, 13, 36, 34, -27, -30, 18, -15, 135, -50, -99, -61, -76, -41, -61, 88, 37, -72, -90, -64, -35, 3, -81, 69, -8, 18, -29, -15, 8, 42, -38, -88, 137, 105, -89, 13, -56, -29, -64, 11, -7, -93, -130, 23, 21,
    -- layer=4 filter=0 channel=2
    -42, -69, -69, -20, 65, 14, 2, -22, 70, -52, -42, 30, 35, -12, -125, -15, 21, 35, -19, 28, -67, -6, 60, -17, 1, -29, 42, -96, 27, -44, 110, -8, 63, 14, 23, -56, 5, 18, -65, -28, -16, 82, 0, -7, -46, -33, -8, -49, 55, -59, 64, 25, -44, 101, -3, 2, -53, -67, -91, 115, -10, 24, 30, 89,
    -- layer=4 filter=0 channel=3
    -35, -1, -13, -61, -59, -42, -2, 0, 11, -106, -19, 2, 2, -5, -19, 16, 66, -27, -75, -44, 35, -33, 47, 0, -23, -51, 70, -11, -9, -18, 0, 101, -100, -71, -1, -66, 0, 22, -66, -4, 62, 70, -15, -46, -4, 30, 21, 102, 20, -1, 72, 10, 17, -44, 69, 59, -45, -51, 0, -37, 63, -9, -21, 25,
    -- layer=4 filter=0 channel=4
    -80, -51, 26, -113, 62, 16, 71, 66, -57, 15, -15, -1, -70, 37, -63, -32, -51, 36, -63, -63, -108, 90, -6, -39, -44, -14, 46, -64, -66, -61, -73, 46, 12, 19, -27, 83, -19, 14, 2, 35, -10, 6, -16, 82, 2, -25, 80, 69, 27, 73, -30, -40, -74, -8, -17, -12, -86, -16, 17, 28, 36, 52, -17, -139,
    -- layer=4 filter=0 channel=5
    -110, -1, -12, -5, 3, -35, 10, -40, 0, -95, 31, 26, 18, 60, -28, -52, 56, 21, -13, -41, -12, -29, -15, 47, -8, 40, 86, 13, 13, -23, 19, 41, -81, -38, -13, 47, -32, -40, -61, 62, 64, 87, 71, 13, -1, -68, 2, 21, -25, -58, 42, -69, 40, 48, -12, 1, 72, 25, 44, -30, 71, 26, -120, 120,
    -- layer=4 filter=0 channel=6
    -26, 8, -142, -147, -26, 9, 56, -84, -42, 19, 94, 106, -148, 47, -64, 31, 48, -38, -27, -89, 5, 20, 76, 34, 22, 11, -47, 2, -14, -87, -38, -77, -56, -16, -80, -66, 119, 64, 4, -43, -47, -108, -107, -103, 67, 41, -27, 95, 33, -112, 55, 8, 28, 26, -32, 107, 26, -38, -36, -109, -63, -100, -56, 16,
    -- layer=4 filter=0 channel=7
    22, -76, 138, -63, 131, -65, 26, 51, 52, 82, -23, -52, 2, 82, 67, -100, 36, 68, 46, 50, 18, 42, -60, 32, -92, -26, 95, -29, -115, 66, 15, 22, 0, 93, -33, 8, -32, -78, -65, -67, 75, 0, 100, 164, -24, -16, -99, 13, 19, -22, -45, -45, -83, -19, 66, -70, 3, 43, -33, -13, -22, 118, -108, -53,
    -- layer=4 filter=0 channel=8
    68, 116, -67, 6, -12, -85, -22, 24, 31, 19, -7, -50, 53, -51, -26, 55, -9, -154, 42, 84, 42, -97, -28, -40, 113, 54, -76, -86, 119, 2, -33, 26, 57, 85, -43, 5, -134, 60, -54, 5, -35, -51, -50, -75, 41, -46, 77, 9, -144, 37, -34, -48, 62, -94, -14, -74, 1, 3, 66, -6, 44, -53, 46, -56,
    -- layer=4 filter=0 channel=9
    33, 82, -42, 11, -89, 127, -69, -23, 47, 53, 67, -52, 34, -62, 57, -108, 14, -64, -1, -18, 42, 88, -55, -67, 4, -32, 47, 110, -80, 38, -44, -75, -57, -2, 86, -6, 31, 35, -78, -9, -68, 59, -75, -52, 13, 62, 57, -38, -13, 34, -47, 22, -16, -110, -27, -109, 60, 41, 82, -101, -85, -58, 5, -51,

    others => 0);
end iwght_package;
