library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    292, 
    
    -- channel=1
    555, 
    
    -- channel=2
    0, 
    
    -- channel=3
    277, 
    
    -- channel=4
    0, 
    
    -- channel=5
    94, 
    
    -- channel=6
    1015, 
    
    -- channel=7
    289, 
    
    -- channel=8
    0, 
    
    -- channel=9
    0, 
    
    -- channel=10
    151, 
    
    -- channel=11
    764, 
    
    -- channel=12
    307, 
    
    -- channel=13
    328, 
    
    -- channel=14
    315, 
    
    -- channel=15
    0, 
    
    -- channel=16
    79, 
    
    -- channel=17
    157, 
    
    -- channel=18
    0, 
    
    -- channel=19
    267, 
    
    -- channel=20
    303, 
    
    -- channel=21
    185, 
    
    -- channel=22
    172, 
    
    -- channel=23
    0, 
    
    -- channel=24
    358, 
    
    -- channel=25
    0, 
    
    -- channel=26
    519, 
    
    -- channel=27
    164, 
    
    -- channel=28
    200, 
    
    -- channel=29
    0, 
    
    -- channel=30
    53, 
    
    -- channel=31
    207, 
    
    -- channel=32
    0, 
    
    -- channel=33
    130, 
    
    -- channel=34
    668, 
    
    -- channel=35
    65, 
    
    -- channel=36
    421, 
    
    -- channel=37
    804, 
    
    -- channel=38
    0, 
    
    -- channel=39
    0, 
    
    -- channel=40
    384, 
    
    -- channel=41
    90, 
    
    -- channel=42
    83, 
    
    -- channel=43
    164, 
    
    -- channel=44
    0, 
    
    -- channel=45
    0, 
    
    -- channel=46
    315, 
    
    -- channel=47
    276, 
    
    -- channel=48
    383, 
    
    -- channel=49
    13, 
    
    -- channel=50
    562, 
    
    -- channel=51
    0, 
    
    -- channel=52
    436, 
    
    -- channel=53
    186, 
    
    -- channel=54
    0, 
    
    -- channel=55
    521, 
    
    -- channel=56
    448, 
    
    -- channel=57
    0, 
    
    -- channel=58
    417, 
    
    -- channel=59
    16, 
    
    -- channel=60
    279, 
    
    -- channel=61
    359, 
    
    -- channel=62
    0, 
    
    -- channel=63
    164, 
    
    
    others => 0);
end gold_package;
