library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 278, 0, 85, 
    407, 0, 183, 82, 0, 0, 0, 
    0, 0, 204, 71, 38, 242, 39, 
    0, 23, 0, 94, 0, 0, 36, 
    0, 127, 107, 0, 0, 452, 0, 
    0, 0, 381, 89, 55, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 144, 155, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 24, 
    0, 0, 0, 15, 0, 132, 0, 
    0, 0, 0, 0, 0, 210, 0, 
    116, 0, 0, 425, 204, 5, 24, 
    0, 563, 70, 39, 21, 18, 3, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 80, 0, 0, 
    135, 0, 306, 251, 136, 245, 163, 
    0, 317, 350, 245, 218, 211, 181, 
    
    -- channel=3
    219, 336, 63, 0, 0, 0, 109, 
    0, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 
    117, 0, 0, 101, 0, 0, 173, 
    0, 0, 0, 0, 0, 185, 0, 
    0, 0, 0, 27, 103, 45, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 193, 0, 0, 283, 
    0, 0, 0, 83, 0, 218, 46, 
    27, 88, 0, 0, 0, 170, 0, 
    0, 0, 0, 0, 0, 82, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    265, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 323, 0, 33, 0, 
    55, 0, 0, 0, 38, 0, 4, 
    0, 0, 0, 0, 0, 9, 0, 
    10, 0, 0, 46, 0, 30, 43, 
    0, 57, 0, 0, 395, 0, 0, 
    57, 0, 155, 158, 0, 0, 0, 
    0, 281, 0, 1, 0, 0, 0, 
    
    -- channel=6
    0, 0, 83, 600, 540, 484, 284, 
    167, 0, 131, 16, 0, 0, 127, 
    0, 0, 0, 0, 0, 87, 0, 
    0, 217, 124, 86, 0, 131, 0, 
    0, 0, 59, 38, 277, 284, 0, 
    7, 27, 527, 162, 11, 0, 0, 
    34, 247, 8, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    120, 0, 0, 0, 0, 0, 0, 
    66, 0, 0, 0, 110, 0, 18, 
    0, 0, 0, 0, 0, 0, 87, 
    0, 66, 25, 189, 0, 4, 66, 
    0, 443, 0, 0, 32, 1, 0, 
    0, 0, 0, 0, 0, 0, 73, 
    
    -- channel=8
    15, 0, 41, 66, 10, 151, 0, 
    79, 0, 274, 225, 0, 0, 20, 
    57, 0, 0, 0, 162, 0, 0, 
    0, 0, 0, 0, 97, 0, 0, 
    0, 204, 116, 238, 115, 0, 0, 
    0, 391, 273, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 
    99, 84, 21, 0, 145, 0, 0, 
    0, 0, 0, 0, 603, 0, 0, 
    0, 0, 0, 0, 216, 0, 0, 
    0, 418, 2, 0, 0, 0, 113, 
    0, 143, 0, 0, 32, 60, 0, 
    0, 0, 148, 0, 0, 0, 0, 
    
    -- channel=10
    0, 47, 295, 478, 325, 224, 47, 
    124, 166, 153, 278, 0, 155, 0, 
    89, 0, 0, 48, 39, 95, 0, 
    124, 0, 0, 110, 0, 0, 0, 
    0, 0, 46, 229, 209, 49, 151, 
    0, 489, 118, 249, 220, 204, 156, 
    0, 60, 95, 0, 44, 2, 242, 
    
    -- channel=11
    71, 105, 54, 106, 0, 159, 228, 
    159, 84, 0, 13, 54, 0, 0, 
    170, 244, 144, 0, 0, 0, 133, 
    106, 212, 163, 34, 229, 0, 173, 
    0, 0, 354, 251, 226, 60, 180, 
    201, 79, 0, 248, 123, 103, 57, 
    49, 142, 0, 5, 4, 0, 0, 
    
    -- channel=12
    0, 0, 0, 28, 67, 265, 104, 
    0, 0, 0, 227, 0, 155, 0, 
    170, 0, 0, 433, 0, 218, 78, 
    293, 95, 0, 280, 0, 139, 0, 
    169, 138, 0, 214, 76, 54, 0, 
    0, 0, 501, 0, 226, 0, 33, 
    0, 154, 78, 59, 26, 8, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    29, 0, 340, 0, 134, 0, 43, 
    26, 75, 0, 0, 126, 0, 0, 
    451, 0, 29, 0, 172, 0, 157, 
    315, 324, 391, 76, 249, 0, 168, 
    118, 0, 0, 328, 44, 0, 168, 
    50, 576, 0, 0, 47, 34, 0, 
    0, 763, 32, 12, 32, 54, 96, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 88, 110, 0, 
    0, 0, 0, 83, 226, 79, 126, 
    107, 153, 0, 31, 0, 0, 23, 
    152, 88, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 200, 258, 254, 
    0, 45, 71, 165, 301, 259, 180, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 72, 142, 
    289, 0, 0, 0, 0, 9, 30, 
    0, 0, 0, 113, 0, 0, 337, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 202, 119, 106, 0, 122, 
    240, 0, 0, 49, 29, 96, 115, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 53, 0, 0, 0, 0, 
    0, 111, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 175, 
    0, 0, 0, 0, 0, 0, 0, 
    103, 0, 0, 0, 0, 1, 79, 
    277, 0, 0, 137, 134, 177, 199, 
    
    -- channel=20
    121, 26, 128, 269, 162, 50, 126, 
    59, 279, 179, 0, 0, 40, 93, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 147, 0, 123, 0, 0, 0, 
    33, 0, 0, 0, 0, 67, 249, 
    0, 39, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 66, 0, 0, 0, 0, 121, 
    115, 42, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 134, 0, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 337, 230, 230, 188, 
    213, 0, 0, 0, 176, 166, 189, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 111, 0, 56, 70, 
    0, 264, 197, 20, 0, 51, 0, 
    0, 0, 142, 32, 57, 126, 102, 
    0, 0, 0, 0, 115, 0, 0, 
    199, 50, 26, 123, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 201, 0, 130, 0, 
    0, 0, 0, 0, 0, 0, 64, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 331, 160, 177, 
    18, 0, 0, 0, 191, 115, 0, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41, 0, 
    0, 0, 5, 0, 0, 0, 0, 
    0, 0, 82, 0, 0, 0, 0, 
    183, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 235, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 40, 0, 0, 
    80, 0, 0, 0, 15, 0, 0, 
    149, 0, 0, 0, 70, 0, 0, 
    21, 16, 0, 164, 115, 0, 0, 
    339, 385, 0, 387, 277, 325, 330, 
    453, 283, 208, 151, 193, 222, 303, 
    
    -- channel=27
    264, 0, 0, 160, 0, 8, 433, 
    12, 153, 0, 0, 251, 0, 64, 
    0, 0, 0, 0, 7, 0, 0, 
    0, 185, 46, 0, 0, 0, 143, 
    0, 0, 0, 0, 0, 62, 239, 
    283, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    271, 475, 529, 311, 60, 0, 56, 
    0, 330, 0, 0, 9, 90, 0, 
    0, 296, 0, 103, 125, 194, 0, 
    0, 0, 337, 136, 233, 219, 4, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 203, 0, 0, 0, 0, 
    0, 0, 48, 148, 0, 31, 0, 
    0, 380, 35, 231, 119, 46, 0, 
    0, 0, 61, 0, 124, 179, 0, 
    0, 0, 83, 83, 0, 0, 0, 
    0, 0, 264, 0, 0, 0, 0, 
    0, 0, 103, 0, 0, 0, 0, 
    
    -- channel=30
    93, 231, 0, 0, 0, 0, 0, 
    0, 80, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 
    0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    20, 18, 176, 92, 113, 80, 0, 
    44, 123, 78, 122, 8, 0, 0, 
    0, 102, 0, 7, 137, 0, 55, 
    134, 170, 0, 36, 67, 2, 77, 
    16, 208, 160, 98, 52, 42, 0, 
    0, 130, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
