library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    24, 47, 31, 33, 25, 40, 36, 44, 27, 0, 8, 25, 40, 42, 39, 
    28, 59, 29, 33, 25, 27, 19, 16, 19, 15, 0, 8, 11, 16, 27, 
    0, 0, 33, 43, 20, 34, 52, 44, 9, 0, 7, 18, 3, 0, 32, 
    48, 0, 27, 29, 18, 15, 12, 0, 0, 0, 50, 14, 48, 16, 0, 
    32, 0, 18, 0, 0, 0, 55, 42, 29, 0, 27, 28, 14, 33, 0, 
    0, 0, 50, 15, 47, 48, 65, 43, 52, 0, 5, 53, 0, 18, 21, 
    11, 2, 25, 92, 0, 0, 0, 25, 56, 0, 47, 37, 8, 4, 15, 
    0, 50, 0, 32, 0, 0, 25, 20, 59, 0, 38, 55, 0, 4, 61, 
    0, 0, 21, 0, 0, 40, 66, 15, 0, 25, 17, 66, 25, 39, 2, 
    12, 0, 59, 0, 12, 0, 6, 25, 0, 3, 35, 30, 0, 0, 16, 
    0, 0, 64, 0, 2, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 43, 8, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 
    30, 19, 0, 0, 1, 183, 14, 10, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 34, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 135, 167, 21, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 11, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 95, 90, 0, 72, 3, 2, 0, 35, 14, 
    0, 0, 0, 0, 0, 153, 0, 0, 0, 36, 62, 109, 58, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 63, 71, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    134, 0, 0, 0, 191, 117, 99, 80, 0, 0, 0, 0, 0, 0, 0, 
    0, 116, 0, 46, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 89, 95, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 89, 
    0, 0, 13, 110, 26, 33, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    46, 32, 54, 35, 37, 39, 40, 45, 37, 13, 17, 40, 36, 23, 19, 
    40, 36, 58, 28, 66, 0, 0, 0, 1, 21, 0, 0, 13, 37, 12, 
    0, 99, 43, 34, 59, 11, 0, 0, 33, 61, 0, 0, 0, 33, 27, 
    0, 98, 4, 54, 0, 72, 0, 0, 0, 151, 0, 0, 0, 0, 111, 
    0, 0, 0, 240, 0, 30, 0, 0, 0, 232, 0, 0, 0, 0, 81, 
    0, 0, 0, 112, 68, 84, 0, 0, 0, 302, 0, 0, 8, 0, 0, 
    43, 0, 6, 0, 91, 99, 0, 0, 0, 189, 0, 0, 0, 2, 0, 
    17, 0, 0, 0, 128, 67, 0, 0, 0, 135, 0, 0, 40, 0, 18, 
    0, 0, 0, 0, 7, 56, 0, 0, 44, 0, 0, 0, 47, 30, 31, 
    0, 0, 0, 61, 0, 106, 109, 0, 0, 3, 0, 0, 26, 45, 4, 
    0, 0, 0, 251, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 42, 0, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 63, 216, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 250, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    
    -- channel=3
    1, 0, 0, 0, 3, 0, 0, 4, 7, 0, 0, 0, 0, 0, 1, 
    6, 0, 0, 0, 0, 0, 5, 0, 0, 55, 28, 83, 86, 0, 0, 
    0, 0, 3, 5, 5, 80, 53, 167, 37, 0, 0, 0, 0, 44, 0, 
    15, 82, 12, 8, 3, 62, 0, 0, 0, 0, 0, 0, 8, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 35, 0, 0, 0, 42, 
    0, 0, 0, 1, 75, 0, 0, 12, 0, 0, 0, 8, 0, 0, 0, 
    21, 0, 57, 0, 11, 0, 0, 0, 0, 0, 7, 35, 50, 2, 0, 
    0, 6, 25, 16, 0, 0, 0, 0, 0, 0, 0, 74, 0, 0, 8, 
    0, 0, 0, 0, 0, 99, 113, 29, 0, 130, 59, 3, 49, 21, 0, 
    0, 0, 0, 85, 0, 0, 52, 0, 23, 0, 0, 10, 0, 0, 0, 
    9, 5, 31, 18, 0, 0, 0, 0, 0, 29, 52, 0, 0, 50, 51, 
    30, 0, 0, 0, 0, 156, 177, 170, 54, 0, 0, 0, 7, 9, 0, 
    0, 46, 23, 0, 98, 0, 0, 0, 6, 0, 0, 0, 0, 0, 1, 
    0, 0, 11, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 16, 156, 30, 7, 0, 0, 0, 2, 0, 18, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 51, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 6, 160, 0, 0, 0, 0, 0, 0, 
    74, 0, 0, 0, 0, 120, 9, 10, 0, 0, 12, 0, 80, 0, 0, 
    128, 0, 0, 0, 0, 0, 0, 20, 2, 0, 25, 38, 13, 0, 0, 
    79, 0, 29, 0, 0, 21, 50, 0, 42, 0, 0, 52, 0, 25, 0, 
    67, 0, 0, 25, 0, 0, 0, 10, 44, 0, 98, 61, 0, 15, 0, 
    0, 75, 0, 57, 0, 0, 94, 0, 104, 0, 82, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 189, 46, 0, 0, 11, 13, 0, 18, 0, 
    0, 0, 35, 0, 0, 86, 0, 0, 0, 100, 0, 129, 0, 0, 0, 
    0, 0, 68, 0, 41, 0, 0, 0, 0, 69, 189, 20, 0, 0, 21, 
    0, 0, 112, 0, 0, 0, 14, 136, 139, 56, 0, 0, 0, 0, 15, 
    53, 0, 1, 0, 376, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 89, 156, 0, 18, 0, 0, 0, 0, 0, 25, 18, 0, 
    15, 0, 0, 199, 15, 0, 0, 0, 0, 0, 3, 2, 0, 0, 152, 
    42, 0, 0, 85, 43, 0, 26, 0, 0, 0, 9, 0, 0, 10, 82, 
    
    -- channel=5
    66, 86, 79, 88, 88, 69, 84, 92, 95, 71, 62, 55, 73, 81, 90, 
    87, 80, 69, 94, 60, 151, 100, 104, 64, 30, 69, 50, 20, 35, 87, 
    126, 0, 86, 97, 72, 0, 141, 23, 0, 0, 29, 28, 83, 0, 49, 
    181, 0, 75, 71, 150, 5, 78, 39, 40, 0, 133, 0, 77, 69, 0, 
    102, 0, 112, 0, 105, 10, 95, 107, 71, 0, 22, 100, 30, 99, 0, 
    0, 12, 140, 67, 0, 0, 165, 50, 166, 0, 106, 101, 0, 46, 61, 
    0, 121, 22, 184, 0, 0, 31, 100, 114, 0, 109, 86, 1, 0, 59, 
    23, 64, 0, 110, 0, 0, 131, 16, 83, 0, 99, 88, 0, 0, 50, 
    59, 0, 161, 0, 73, 0, 39, 77, 0, 67, 0, 103, 0, 3, 48, 
    26, 0, 196, 0, 36, 0, 0, 82, 3, 26, 101, 0, 0, 13, 79, 
    0, 0, 152, 0, 248, 16, 0, 9, 110, 67, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 133, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 62, 109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 184, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 61, 51, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 95, 0, 0, 0, 0, 52, 0, 
    16, 168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 76, 
    0, 0, 0, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 90, 84, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 74, 0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 128, 43, 22, 7, 0, 0, 0, 8, 8, 0, 
    0, 0, 0, 34, 0, 38, 0, 0, 40, 0, 0, 41, 0, 0, 0, 
    0, 0, 0, 0, 27, 16, 0, 0, 0, 161, 85, 38, 48, 0, 0, 
    14, 0, 0, 0, 0, 0, 107, 181, 139, 0, 0, 0, 0, 23, 19, 
    133, 135, 67, 0, 0, 30, 0, 0, 3, 3, 1, 0, 0, 0, 0, 
    0, 53, 101, 0, 51, 0, 0, 0, 0, 0, 0, 0, 4, 26, 0, 
    0, 0, 114, 79, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 21, 0, 11, 72, 23, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 20, 36, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 22, 0, 30, 0, 26, 15, 0, 
    60, 18, 0, 0, 0, 0, 13, 23, 35, 0, 5, 19, 16, 39, 0, 
    24, 44, 0, 0, 0, 0, 47, 0, 77, 0, 25, 14, 0, 25, 20, 
    7, 122, 0, 0, 0, 0, 13, 13, 46, 0, 38, 35, 17, 16, 6, 
    34, 88, 0, 0, 0, 0, 21, 0, 0, 0, 32, 37, 0, 0, 0, 
    84, 68, 83, 13, 0, 0, 0, 39, 0, 0, 0, 6, 0, 0, 0, 
    56, 56, 121, 41, 16, 0, 0, 73, 1, 0, 19, 4, 0, 0, 0, 
    68, 36, 103, 0, 166, 64, 49, 61, 75, 65, 86, 115, 121, 80, 80, 
    106, 67, 32, 38, 141, 129, 132, 127, 155, 152, 177, 186, 204, 204, 204, 
    249, 105, 0, 120, 126, 174, 175, 168, 175, 186, 205, 211, 207, 202, 225, 
    260, 219, 34, 191, 150, 172, 191, 174, 176, 194, 218, 219, 231, 242, 252, 
    258, 241, 205, 145, 166, 166, 166, 171, 182, 210, 214, 200, 205, 275, 259, 
    
    -- channel=8
    213, 227, 225, 226, 225, 213, 235, 253, 225, 169, 136, 149, 174, 199, 196, 
    221, 242, 238, 234, 223, 232, 192, 181, 129, 61, 39, 48, 76, 132, 180, 
    132, 144, 234, 242, 243, 214, 111, 51, 23, 59, 28, 16, 44, 47, 150, 
    47, 102, 206, 230, 193, 110, 90, 28, 28, 42, 58, 47, 18, 25, 104, 
    0, 93, 167, 127, 110, 103, 64, 34, 34, 37, 55, 39, 34, 24, 58, 
    0, 43, 147, 212, 81, 53, 93, 47, 50, 61, 44, 4, 22, 15, 22, 
    0, 76, 72, 183, 142, 84, 61, 45, 25, 85, 15, 16, 27, 21, 40, 
    0, 14, 8, 89, 107, 66, 34, 42, 29, 130, 50, 21, 13, 52, 104, 
    0, 0, 0, 34, 63, 51, 45, 55, 18, 131, 38, 14, 37, 104, 185, 
    22, 13, 0, 32, 0, 27, 27, 61, 33, 20, 13, 0, 37, 163, 162, 
    5, 11, 0, 18, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    102, 118, 103, 99, 100, 97, 115, 143, 126, 112, 104, 101, 77, 78, 91, 
    98, 117, 116, 110, 102, 0, 34, 117, 147, 0, 0, 0, 20, 80, 71, 
    111, 154, 112, 121, 128, 194, 52, 12, 0, 0, 0, 0, 0, 0, 59, 
    0, 0, 75, 119, 75, 4, 0, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 109, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 74, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 62, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    35, 36, 25, 36, 35, 28, 33, 36, 37, 44, 24, 17, 18, 26, 42, 
    38, 38, 28, 40, 30, 80, 2, 29, 21, 28, 40, 28, 19, 39, 46, 
    47, 38, 39, 40, 45, 96, 15, 17, 2, 44, 20, 0, 40, 22, 56, 
    73, 46, 53, 35, 43, 6, 66, 0, 29, 13, 10, 15, 25, 28, 45, 
    0, 86, 0, 0, 53, 0, 0, 0, 41, 0, 24, 0, 38, 42, 0, 
    0, 52, 0, 0, 73, 0, 40, 7, 75, 13, 0, 0, 31, 17, 0, 
    0, 109, 0, 66, 78, 0, 68, 0, 54, 68, 0, 3, 17, 37, 17, 
    0, 43, 0, 75, 13, 64, 0, 4, 27, 56, 9, 21, 17, 26, 0, 
    0, 1, 0, 52, 0, 0, 24, 72, 7, 51, 83, 0, 21, 47, 41, 
    0, 0, 18, 25, 9, 0, 0, 99, 0, 3, 10, 19, 49, 52, 25, 
    102, 0, 23, 0, 0, 0, 0, 0, 0, 0, 34, 23, 11, 61, 52, 
    67, 0, 0, 64, 46, 0, 29, 22, 26, 35, 43, 35, 39, 35, 29, 
    39, 26, 0, 104, 0, 18, 25, 26, 37, 40, 40, 35, 33, 20, 24, 
    37, 31, 0, 139, 12, 20, 26, 29, 20, 23, 32, 49, 33, 40, 61, 
    24, 35, 25, 115, 47, 44, 35, 16, 24, 34, 38, 24, 29, 59, 40, 
    
    -- channel=11
    78, 89, 79, 82, 77, 84, 90, 86, 75, 78, 69, 65, 61, 63, 51, 
    73, 86, 83, 89, 75, 130, 89, 96, 60, 29, 41, 42, 46, 55, 61, 
    99, 60, 87, 84, 86, 145, 62, 13, 0, 63, 84, 33, 41, 24, 63, 
    57, 41, 93, 84, 98, 33, 90, 25, 29, 70, 87, 59, 19, 3, 37, 
    51, 140, 89, 33, 172, 98, 113, 45, 36, 0, 98, 51, 33, 8, 4, 
    64, 169, 96, 85, 187, 100, 147, 59, 46, 70, 138, 38, 41, 18, 0, 
    35, 202, 83, 76, 109, 116, 198, 85, 65, 126, 108, 44, 26, 39, 42, 
    95, 144, 46, 84, 47, 203, 123, 96, 49, 122, 102, 53, 33, 75, 30, 
    141, 168, 75, 103, 71, 70, 66, 78, 42, 87, 105, 23, 9, 40, 80, 
    160, 159, 112, 83, 106, 18, 35, 135, 72, 77, 26, 0, 32, 93, 82, 
    179, 155, 115, 111, 150, 94, 148, 161, 72, 0, 0, 0, 30, 62, 48, 
    132, 137, 100, 251, 251, 45, 51, 40, 21, 10, 22, 21, 26, 37, 29, 
    32, 96, 78, 302, 38, 21, 24, 16, 9, 8, 12, 30, 48, 30, 33, 
    23, 25, 101, 221, 22, 23, 20, 20, 13, 21, 27, 38, 17, 38, 87, 
    33, 22, 42, 72, 13, 21, 27, 15, 24, 33, 30, 7, 27, 81, 16, 
    
    -- channel=12
    0, 7, 8, 3, 0, 16, 0, 0, 11, 0, 0, 0, 0, 0, 1, 
    10, 26, 11, 0, 8, 172, 0, 33, 0, 30, 32, 14, 0, 0, 12, 
    21, 0, 11, 0, 14, 0, 0, 0, 31, 90, 0, 0, 0, 0, 30, 
    0, 163, 0, 20, 53, 0, 66, 0, 0, 18, 0, 0, 0, 0, 30, 
    0, 142, 0, 4, 133, 0, 0, 0, 0, 53, 0, 0, 22, 0, 17, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 300, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 60, 105, 0, 0, 0, 204, 0, 0, 0, 37, 0, 
    0, 0, 0, 0, 17, 131, 0, 0, 0, 112, 0, 0, 6, 0, 0, 
    0, 0, 0, 41, 13, 0, 0, 62, 0, 0, 39, 0, 0, 8, 63, 
    0, 0, 0, 32, 0, 0, 0, 44, 0, 0, 0, 0, 74, 85, 0, 
    71, 0, 0, 235, 0, 61, 97, 0, 0, 0, 46, 95, 37, 0, 0, 
    0, 0, 0, 186, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 28, 0, 
    0, 84, 0, 0, 0, 197, 0, 0, 0, 47, 0, 0, 0, 19, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 0, 0, 0, 0, 146, 
    0, 15, 0, 59, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 
    0, 45, 0, 0, 346, 0, 0, 0, 0, 146, 0, 0, 54, 0, 0, 
    0, 0, 4, 0, 215, 0, 89, 0, 0, 190, 0, 0, 0, 4, 0, 
    0, 25, 0, 0, 62, 212, 0, 7, 0, 135, 0, 0, 54, 7, 0, 
    0, 14, 0, 97, 0, 95, 17, 0, 45, 0, 182, 0, 29, 67, 0, 
    0, 0, 0, 77, 0, 0, 0, 0, 0, 42, 0, 34, 68, 2, 0, 
    180, 0, 0, 133, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    256, 58, 0, 81, 0, 0, 60, 61, 7, 0, 0, 0, 0, 0, 0, 
    0, 139, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 130, 67, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 256, 0, 50, 48, 0, 0, 0, 0, 0, 11, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    144, 139, 147, 151, 146, 131, 156, 171, 155, 116, 90, 102, 113, 121, 127, 
    154, 153, 154, 152, 158, 102, 118, 110, 57, 42, 0, 0, 32, 110, 125, 
    55, 124, 161, 160, 159, 77, 57, 21, 34, 0, 0, 0, 0, 38, 98, 
    0, 50, 145, 159, 102, 90, 20, 0, 0, 22, 0, 0, 0, 0, 70, 
    0, 0, 105, 159, 23, 0, 0, 0, 0, 34, 0, 0, 0, 0, 5, 
    0, 0, 110, 47, 6, 18, 0, 0, 0, 44, 0, 0, 0, 0, 0, 
    0, 0, 94, 98, 0, 37, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 55, 54, 17, 0, 0, 20, 0, 0, 0, 0, 0, 71, 
    0, 0, 0, 0, 17, 0, 18, 0, 32, 0, 47, 0, 0, 55, 94, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 26, 0, 0, 2, 75, 106, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
