library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    80, 84, 85, 85, 81, 81, 83, 87, 82, 64, 54, 60, 66, 66, 66, 
    80, 83, 85, 85, 88, 104, 62, 67, 40, 48, 26, 20, 35, 55, 66, 
    52, 66, 86, 87, 89, 84, 52, 24, 29, 56, 43, 37, 10, 25, 61, 
    6, 57, 72, 86, 72, 64, 51, 31, 28, 60, 46, 35, 25, 10, 45, 
    26, 58, 58, 91, 83, 57, 47, 34, 20, 60, 52, 23, 33, 10, 18, 
    44, 76, 66, 83, 109, 75, 66, 35, 11, 98, 55, 28, 36, 23, 10, 
    53, 46, 53, 56, 69, 97, 69, 54, 18, 86, 43, 29, 31, 42, 31, 
    65, 54, 24, 40, 59, 100, 56, 48, 42, 89, 60, 28, 37, 47, 57, 
    70, 68, 32, 58, 55, 46, 46, 46, 47, 29, 60, 20, 35, 59, 71, 
    93, 79, 32, 51, 32, 42, 60, 49, 40, 50, 8, 1, 26, 62, 61, 
    81, 73, 31, 120, 56, 30, 62, 50, 16, 0, 1, 3, 2, 8, 4, 
    28, 69, 54, 119, 42, 20, 12, 10, 6, 2, 2, 3, 9, 9, 6, 
    0, 29, 88, 87, 19, 8, 0, 2, 2, 4, 4, 8, 5, 5, 17, 
    0, 0, 58, 46, 19, 9, 2, 1, 4, 6, 4, 5, 0, 18, 0, 
    0, 0, 0, 4, 1, 9, 10, 8, 11, 11, 2, 6, 28, 12, 0, 
    
    -- channel=1
    54, 52, 56, 57, 56, 50, 57, 59, 55, 45, 37, 39, 46, 51, 52, 
    56, 55, 59, 57, 59, 45, 54, 41, 32, 24, 24, 17, 19, 42, 51, 
    24, 42, 58, 57, 58, 17, 22, 14, 29, 20, 20, 23, 23, 27, 40, 
    24, 37, 55, 55, 40, 38, 32, 32, 23, 22, 14, 17, 15, 23, 33, 
    33, 33, 55, 62, 46, 41, 12, 17, 9, 27, 23, 28, 20, 26, 24, 
    17, 8, 51, 27, 0, 18, 14, 26, 15, 30, 12, 14, 20, 23, 31, 
    27, 0, 32, 38, 12, 22, 11, 22, 18, 11, 11, 16, 16, 23, 31, 
    17, 2, 34, 35, 46, 20, 2, 2, 23, 14, 12, 10, 18, 20, 39, 
    5, 0, 11, 16, 27, 2, 14, 12, 32, 11, 9, 3, 14, 35, 53, 
    0, 4, 6, 4, 21, 22, 21, 21, 18, 15, 7, 17, 32, 40, 42, 
    0, 4, 0, 21, 37, 40, 14, 0, 12, 7, 14, 19, 5, 0, 2, 
    0, 0, 27, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=2
    35, 39, 40, 37, 36, 39, 43, 43, 39, 35, 27, 28, 29, 26, 23, 
    33, 44, 47, 41, 45, 27, 36, 37, 38, 7, 0, 0, 1, 22, 22, 
    16, 41, 39, 40, 45, 61, 3, 0, 0, 15, 0, 0, 0, 0, 19, 
    0, 0, 35, 45, 27, 30, 9, 0, 0, 39, 0, 0, 0, 0, 26, 
    0, 16, 22, 81, 44, 41, 3, 0, 0, 18, 8, 0, 0, 0, 0, 
    0, 6, 11, 34, 49, 36, 0, 0, 0, 48, 2, 0, 0, 0, 0, 
    0, 0, 14, 14, 50, 29, 40, 0, 0, 56, 0, 0, 0, 0, 0, 
    0, 2, 0, 10, 50, 72, 0, 2, 0, 39, 0, 0, 0, 0, 0, 
    1, 23, 0, 9, 0, 25, 0, 0, 3, 9, 11, 0, 0, 0, 23, 
    13, 20, 0, 21, 0, 0, 14, 6, 0, 5, 0, 0, 0, 27, 29, 
    30, 22, 0, 46, 0, 0, 37, 19, 0, 0, 0, 0, 0, 0, 0, 
    10, 14, 10, 78, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    47, 47, 44, 47, 49, 44, 48, 53, 54, 51, 43, 37, 36, 42, 45, 
    46, 47, 47, 50, 45, 30, 51, 50, 49, 24, 20, 26, 30, 36, 42, 
    52, 36, 50, 51, 52, 60, 49, 40, 16, 0, 10, 2, 19, 23, 29, 
    43, 1, 50, 49, 53, 29, 24, 10, 6, 0, 18, 17, 17, 16, 15, 
    16, 0, 45, 20, 7, 0, 22, 14, 16, 0, 17, 19, 7, 12, 12, 
    10, 6, 38, 39, 20, 12, 21, 19, 21, 0, 21, 22, 7, 7, 4, 
    0, 25, 35, 53, 15, 2, 29, 11, 27, 0, 28, 17, 7, 3, 10, 
    0, 12, 13, 37, 14, 3, 19, 19, 19, 0, 21, 25, 3, 8, 15, 
    4, 1, 17, 5, 17, 22, 28, 20, 2, 36, 35, 24, 6, 11, 28, 
    8, 2, 23, 0, 24, 0, 0, 15, 9, 21, 22, 9, 0, 19, 45, 
    1, 6, 28, 0, 0, 0, 0, 6, 10, 9, 0, 0, 0, 16, 26, 
    0, 0, 1, 0, 55, 21, 7, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 38, 0, 0, 0, 11, 1, 0, 
    31, 25, 0, 0, 0, 53, 21, 16, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 13, 6, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 14, 
    13, 0, 0, 41, 45, 14, 0, 0, 0, 0, 11, 14, 0, 0, 0, 
    0, 2, 9, 0, 15, 0, 2, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 49, 33, 0, 0, 6, 2, 0, 13, 0, 
    0, 0, 2, 0, 0, 53, 0, 0, 0, 18, 19, 50, 19, 0, 0, 
    3, 0, 0, 0, 0, 12, 0, 0, 2, 36, 47, 3, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 34, 10, 0, 0, 0, 0, 9, 7, 
    61, 19, 0, 0, 97, 66, 45, 40, 9, 4, 0, 3, 0, 0, 0, 
    0, 47, 0, 27, 64, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 
    0, 0, 36, 65, 10, 0, 0, 0, 0, 0, 6, 12, 3, 0, 49, 
    3, 0, 14, 48, 24, 20, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    11, 15, 12, 15, 13, 17, 15, 8, 11, 19, 18, 14, 16, 12, 7, 
    12, 15, 11, 18, 12, 62, 37, 28, 17, 23, 55, 37, 12, 9, 15, 
    31, 0, 15, 12, 9, 14, 27, 6, 14, 43, 66, 46, 50, 5, 14, 
    74, 18, 24, 14, 36, 20, 69, 42, 39, 16, 70, 33, 30, 19, 0, 
    94, 90, 45, 5, 139, 95, 82, 50, 32, 0, 74, 64, 36, 41, 0, 
    76, 91, 53, 16, 33, 52, 103, 57, 62, 21, 100, 48, 29, 43, 34, 
    72, 117, 26, 36, 18, 62, 105, 81, 65, 44, 87, 53, 30, 40, 46, 
    95, 109, 60, 62, 23, 84, 89, 44, 43, 31, 69, 48, 23, 40, 14, 
    118, 106, 93, 57, 61, 16, 37, 56, 35, 53, 23, 24, 1, 12, 25, 
    96, 95, 110, 53, 79, 30, 36, 109, 52, 31, 34, 6, 27, 35, 29, 
    91, 99, 101, 60, 183, 116, 101, 102, 88, 50, 40, 61, 63, 68, 69, 
    57, 85, 97, 125, 141, 46, 39, 36, 49, 53, 61, 62, 68, 70, 71, 
    86, 47, 56, 156, 68, 62, 62, 55, 54, 58, 65, 76, 79, 72, 85, 
    82, 71, 36, 134, 64, 61, 69, 59, 56, 64, 68, 67, 69, 79, 91, 
    89, 69, 65, 46, 49, 42, 51, 60, 68, 77, 72, 58, 76, 113, 85, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 5, 26, 4, 3, 0, 3, 0, 
    0, 25, 0, 0, 0, 3, 0, 0, 0, 36, 0, 8, 0, 0, 15, 
    0, 20, 0, 20, 0, 15, 1, 0, 0, 48, 9, 0, 3, 0, 12, 
    16, 29, 0, 15, 59, 32, 4, 0, 0, 76, 3, 0, 10, 0, 0, 
    22, 9, 6, 0, 31, 44, 8, 3, 0, 65, 0, 0, 11, 13, 0, 
    32, 11, 7, 0, 15, 42, 0, 14, 0, 45, 5, 0, 17, 10, 0, 
    27, 38, 0, 25, 9, 24, 6, 5, 16, 0, 18, 0, 15, 8, 0, 
    33, 39, 0, 45, 0, 19, 32, 0, 17, 4, 0, 0, 11, 8, 0, 
    50, 37, 0, 87, 0, 3, 39, 18, 0, 0, 7, 11, 21, 14, 2, 
    53, 49, 13, 72, 1, 19, 33, 32, 17, 14, 16, 22, 23, 25, 21, 
    16, 54, 72, 33, 0, 20, 16, 18, 15, 18, 23, 25, 23, 26, 32, 
    15, 24, 88, 0, 7, 23, 15, 18, 21, 24, 25, 25, 22, 38, 19, 
    13, 26, 33, 14, 10, 25, 20, 17, 23, 23, 17, 24, 40, 20, 0, 
    
    -- channel=9
    74, 83, 78, 80, 80, 76, 84, 91, 85, 76, 66, 63, 66, 67, 69, 
    75, 85, 85, 86, 82, 59, 76, 79, 81, 26, 7, 6, 22, 52, 66, 
    65, 68, 80, 86, 83, 101, 54, 28, 0, 0, 9, 5, 11, 9, 51, 
    35, 0, 74, 84, 76, 49, 33, 8, 0, 12, 26, 14, 8, 0, 27, 
    24, 2, 66, 65, 61, 32, 37, 7, 3, 0, 21, 14, 1, 3, 0, 
    0, 10, 60, 46, 40, 35, 33, 23, 8, 0, 33, 17, 6, 5, 0, 
    0, 24, 36, 84, 41, 7, 63, 22, 30, 0, 31, 0, 0, 0, 0, 
    0, 30, 0, 55, 33, 44, 46, 24, 18, 13, 26, 7, 0, 12, 27, 
    3, 10, 0, 10, 5, 32, 20, 8, 2, 38, 21, 24, 0, 11, 44, 
    21, 9, 16, 0, 19, 0, 4, 29, 0, 37, 30, 0, 0, 39, 69, 
    6, 11, 24, 0, 13, 0, 2, 36, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 12, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    52, 53, 58, 58, 59, 52, 59, 65, 65, 46, 35, 39, 48, 53, 56, 
    62, 62, 58, 58, 58, 66, 61, 53, 30, 32, 26, 23, 22, 39, 51, 
    30, 30, 61, 64, 58, 0, 47, 28, 27, 0, 0, 2, 9, 10, 36, 
    28, 22, 56, 63, 61, 42, 24, 10, 1, 0, 11, 0, 11, 16, 11, 
    16, 0, 51, 40, 28, 11, 5, 18, 0, 5, 9, 18, 6, 18, 6, 
    0, 0, 53, 32, 0, 5, 22, 14, 17, 0, 0, 12, 0, 7, 23, 
    6, 0, 30, 61, 0, 17, 0, 12, 7, 0, 2, 15, 2, 4, 9, 
    2, 0, 14, 39, 2, 0, 0, 0, 10, 0, 4, 9, 0, 0, 24, 
    0, 0, 11, 0, 24, 0, 15, 12, 2, 10, 0, 0, 0, 18, 40, 
    0, 0, 5, 0, 0, 4, 8, 3, 0, 0, 0, 7, 0, 28, 47, 
    0, 0, 0, 0, 31, 3, 0, 0, 0, 7, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    30, 30, 37, 33, 34, 34, 33, 34, 36, 25, 14, 21, 26, 26, 27, 
    37, 38, 40, 32, 41, 63, 13, 25, 2, 25, 11, 6, 14, 22, 27, 
    12, 25, 34, 33, 43, 33, 0, 0, 16, 56, 2, 0, 0, 16, 30, 
    0, 77, 26, 40, 29, 31, 22, 6, 11, 57, 0, 10, 0, 0, 47, 
    0, 61, 0, 65, 32, 28, 0, 0, 0, 69, 7, 0, 17, 0, 32, 
    0, 20, 0, 52, 41, 0, 0, 0, 0, 142, 0, 0, 20, 0, 1, 
    0, 0, 0, 0, 70, 58, 0, 0, 0, 120, 0, 0, 18, 27, 0, 
    0, 0, 0, 0, 58, 72, 0, 0, 0, 89, 0, 0, 25, 16, 1, 
    0, 7, 0, 29, 17, 0, 0, 21, 23, 5, 23, 0, 23, 28, 43, 
    2, 12, 0, 52, 0, 10, 27, 12, 13, 0, 0, 0, 39, 56, 18, 
    47, 7, 0, 123, 0, 10, 55, 0, 0, 0, 11, 25, 21, 1, 0, 
    24, 6, 0, 114, 0, 0, 0, 0, 0, 0, 0, 2, 1, 5, 0, 
    0, 29, 38, 16, 0, 0, 0, 0, 0, 6, 8, 9, 0, 0, 7, 
    0, 0, 71, 0, 0, 3, 0, 0, 2, 4, 2, 0, 0, 21, 0, 
    0, 0, 5, 0, 0, 6, 0, 0, 11, 5, 0, 1, 34, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 14, 15, 20, 6, 0, 
    29, 0, 0, 0, 0, 0, 0, 4, 10, 0, 14, 9, 20, 14, 0, 
    38, 0, 0, 0, 0, 0, 16, 9, 18, 0, 11, 13, 5, 14, 1, 
    46, 15, 0, 0, 7, 3, 0, 13, 19, 0, 23, 32, 11, 16, 9, 
    38, 32, 3, 0, 0, 0, 17, 10, 29, 0, 40, 22, 14, 5, 5, 
    26, 38, 29, 0, 0, 0, 36, 23, 12, 0, 18, 31, 11, 2, 0, 
    35, 33, 39, 6, 0, 30, 22, 6, 8, 15, 10, 35, 6, 0, 0, 
    23, 28, 47, 18, 33, 1, 5, 8, 15, 9, 35, 24, 0, 0, 0, 
    20, 27, 55, 0, 14, 15, 0, 45, 47, 42, 38, 27, 51, 68, 71, 
    82, 43, 33, 0, 89, 99, 81, 82, 75, 65, 67, 71, 69, 73, 74, 
    89, 69, 24, 34, 108, 62, 64, 63, 65, 65, 70, 70, 75, 79, 75, 
    98, 81, 44, 85, 64, 65, 66, 64, 63, 67, 77, 85, 87, 75, 94, 
    90, 81, 72, 104, 74, 68, 70, 63, 55, 65, 75, 74, 57, 83, 100, 
    
    -- channel=14
    57, 62, 56, 63, 64, 57, 64, 70, 70, 63, 54, 46, 48, 60, 63, 
    60, 64, 57, 67, 50, 47, 84, 73, 59, 17, 33, 48, 41, 34, 58, 
    87, 11, 63, 68, 62, 69, 79, 56, 11, 0, 31, 10, 47, 21, 28, 
    107, 0, 67, 58, 88, 17, 45, 26, 16, 0, 59, 28, 39, 39, 0, 
    44, 0, 79, 0, 20, 18, 69, 53, 45, 0, 34, 59, 17, 40, 12, 
    32, 7, 82, 64, 0, 9, 64, 46, 79, 0, 68, 61, 2, 21, 22, 
    14, 70, 42, 103, 0, 0, 45, 39, 74, 0, 71, 53, 11, 0, 35, 
    19, 39, 28, 67, 0, 0, 74, 32, 44, 0, 45, 68, 0, 17, 30, 
    30, 0, 78, 0, 49, 14, 48, 44, 0, 74, 35, 65, 3, 0, 33, 
    14, 0, 89, 0, 55, 5, 0, 41, 39, 29, 53, 7, 0, 17, 64, 
    0, 11, 90, 0, 46, 17, 0, 15, 40, 33, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 129, 43, 9, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 3, 9, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 25, 17, 0, 7, 
    40, 0, 0, 0, 0, 0, 26, 1, 11, 0, 31, 0, 22, 0, 0, 
    69, 18, 0, 0, 85, 0, 23, 7, 4, 0, 24, 12, 14, 30, 0, 
    0, 32, 0, 0, 19, 0, 54, 21, 31, 0, 12, 15, 9, 24, 5, 
    0, 42, 0, 20, 0, 0, 55, 27, 47, 0, 36, 7, 0, 16, 7, 
    0, 77, 0, 41, 0, 24, 19, 5, 31, 0, 31, 7, 1, 0, 2, 
    19, 35, 0, 40, 0, 0, 13, 12, 13, 0, 0, 10, 0, 8, 0, 
    36, 18, 60, 8, 27, 0, 3, 71, 0, 13, 30, 15, 18, 0, 0, 
    51, 14, 51, 0, 109, 20, 13, 58, 53, 21, 15, 27, 6, 17, 21, 
    0, 42, 58, 9, 39, 17, 0, 2, 26, 26, 32, 27, 36, 26, 33, 
    27, 0, 0, 30, 39, 31, 31, 26, 28, 29, 35, 31, 34, 39, 43, 
    47, 27, 0, 113, 40, 25, 32, 23, 31, 30, 26, 34, 40, 27, 32, 
    43, 38, 5, 48, 17, 14, 33, 38, 35, 35, 30, 29, 40, 48, 61, 
    
    -- channel=16
    84, 93, 87, 90, 87, 89, 92, 98, 96, 88, 78, 74, 77, 79, 81, 
    83, 98, 92, 95, 88, 75, 91, 97, 90, 41, 28, 34, 44, 61, 76, 
    88, 64, 91, 96, 93, 102, 76, 51, 26, 10, 26, 12, 24, 28, 57, 
    57, 0, 83, 93, 95, 57, 52, 26, 14, 13, 42, 34, 26, 14, 28, 
    31, 7, 76, 58, 63, 47, 57, 33, 25, 0, 37, 38, 17, 18, 15, 
    25, 15, 74, 93, 54, 55, 55, 37, 32, 0, 53, 38, 15, 18, 8, 
    14, 39, 51, 105, 42, 31, 64, 37, 43, 0, 48, 28, 9, 10, 19, 
    25, 31, 13, 65, 34, 44, 55, 37, 35, 19, 42, 34, 10, 26, 30, 
    31, 21, 30, 12, 47, 40, 39, 34, 4, 55, 50, 40, 14, 18, 56, 
    34, 19, 40, 0, 42, 20, 10, 39, 20, 49, 37, 12, 0, 45, 78, 
    12, 29, 43, 0, 21, 15, 11, 36, 24, 11, 0, 0, 0, 0, 5, 
    0, 0, 16, 11, 85, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 63, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 5, 0, 0, 0, 9, 0, 7, 4, 22, 16, 12, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 10, 46, 6, 23, 14, 3, 15, 
    0, 0, 0, 0, 0, 0, 9, 4, 15, 36, 3, 0, 7, 0, 16, 
    38, 30, 0, 8, 75, 45, 0, 0, 0, 38, 18, 15, 21, 5, 0, 
    31, 23, 11, 0, 34, 17, 22, 7, 0, 51, 18, 6, 18, 13, 3, 
    32, 22, 4, 0, 10, 41, 34, 38, 12, 39, 21, 10, 26, 27, 0, 
    34, 49, 14, 23, 0, 57, 16, 2, 14, 6, 29, 24, 34, 8, 0, 
    44, 49, 6, 45, 12, 24, 24, 0, 20, 27, 20, 17, 11, 0, 0, 
    54, 42, 19, 44, 0, 0, 45, 54, 21, 11, 12, 15, 33, 38, 28, 
    102, 75, 28, 46, 64, 73, 74, 74, 53, 50, 50, 58, 58, 57, 56, 
    56, 93, 70, 50, 55, 50, 51, 51, 47, 48, 53, 52, 60, 66, 56, 
    61, 60, 109, 55, 43, 54, 45, 50, 55, 56, 64, 70, 65, 64, 83, 
    59, 65, 70, 73, 53, 66, 65, 53, 50, 50, 55, 60, 56, 53, 51, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 0, 0, 24, 28, 0, 
    0, 78, 0, 0, 0, 48, 0, 0, 0, 44, 0, 0, 0, 32, 34, 
    0, 64, 0, 0, 0, 9, 0, 0, 0, 96, 0, 0, 0, 0, 94, 
    0, 10, 0, 51, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 29, 
    0, 27, 0, 0, 148, 0, 0, 0, 0, 160, 0, 0, 19, 0, 0, 
    0, 0, 18, 0, 96, 29, 0, 0, 0, 147, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 27, 87, 0, 9, 0, 91, 0, 0, 30, 10, 0, 
    0, 0, 0, 51, 0, 43, 0, 0, 31, 0, 45, 0, 38, 29, 0, 
    0, 0, 0, 58, 0, 0, 28, 0, 0, 21, 0, 9, 45, 28, 0, 
    96, 0, 0, 124, 0, 0, 39, 9, 0, 0, 0, 0, 10, 37, 2, 
    135, 76, 0, 79, 0, 0, 34, 32, 3, 6, 9, 10, 3, 1, 0, 
    0, 108, 94, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 10, 2, 
    0, 7, 158, 0, 0, 4, 0, 0, 8, 4, 2, 17, 0, 20, 1, 
    0, 7, 14, 50, 0, 37, 29, 3, 0, 0, 0, 5, 21, 0, 0, 
    
    -- channel=19
    1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 27, 6, 0, 0, 26, 19, 0, 
    20, 45, 0, 0, 0, 51, 19, 26, 0, 0, 0, 0, 0, 26, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 6, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 0, 0, 0, 0, 18, 
    0, 0, 0, 8, 93, 12, 0, 0, 0, 1, 0, 0, 2, 0, 0, 
    0, 0, 31, 0, 33, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 24, 0, 12, 0, 0, 8, 1, 0, 
    0, 0, 0, 5, 0, 52, 10, 0, 0, 0, 46, 22, 23, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 15, 12, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 22, 16, 
    76, 31, 0, 0, 25, 63, 51, 49, 19, 0, 0, 0, 0, 0, 0, 
    0, 57, 22, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 64, 31, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 10, 
    0, 0, 6, 57, 9, 21, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 19, 2, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 5, 1, 4, 38, 0, 12, 0, 0, 0, 
    0, 31, 0, 4, 16, 5, 3, 0, 0, 21, 15, 0, 4, 0, 0, 
    26, 41, 0, 0, 58, 13, 6, 0, 0, 69, 14, 0, 14, 0, 0, 
    20, 36, 0, 0, 25, 37, 40, 0, 0, 67, 7, 2, 7, 19, 0, 
    36, 26, 8, 0, 16, 75, 0, 15, 0, 40, 11, 1, 21, 10, 0, 
    43, 56, 9, 30, 9, 10, 3, 18, 14, 0, 40, 0, 0, 0, 0, 
    46, 54, 10, 42, 27, 0, 13, 23, 18, 17, 0, 0, 9, 0, 0, 
    72, 50, 7, 86, 17, 43, 70, 48, 13, 0, 25, 36, 46, 43, 36, 
    98, 62, 27, 97, 58, 37, 50, 48, 46, 47, 54, 56, 59, 65, 63, 
    64, 86, 64, 83, 17, 49, 48, 46, 48, 55, 61, 68, 68, 68, 72, 
    67, 63, 109, 44, 42, 54, 46, 52, 54, 60, 65, 72, 62, 91, 74, 
    60, 68, 62, 54, 46, 62, 59, 48, 55, 57, 60, 59, 78, 78, 49, 
    
    -- channel=21
    1, 8, 1, 9, 10, 4, 3, 8, 17, 20, 13, 0, 3, 10, 19, 
    3, 5, 0, 12, 0, 3, 39, 25, 29, 0, 28, 23, 0, 0, 13, 
    45, 0, 4, 11, 0, 0, 57, 31, 0, 0, 26, 11, 43, 0, 0, 
    123, 0, 8, 1, 42, 0, 34, 26, 8, 0, 58, 6, 39, 26, 0, 
    88, 0, 41, 0, 28, 7, 62, 51, 32, 0, 24, 65, 5, 47, 0, 
    49, 0, 49, 11, 0, 0, 64, 45, 83, 0, 68, 69, 0, 27, 22, 
    39, 47, 0, 82, 0, 0, 30, 42, 84, 0, 82, 54, 0, 0, 25, 
    33, 45, 17, 49, 0, 0, 79, 9, 42, 0, 46, 64, 0, 0, 1, 
    48, 0, 100, 0, 31, 0, 30, 30, 0, 37, 0, 63, 0, 0, 0, 
    10, 0, 120, 0, 57, 0, 0, 44, 10, 14, 56, 4, 0, 0, 18, 
    0, 0, 108, 0, 108, 39, 0, 19, 69, 46, 4, 0, 0, 0, 28, 
    0, 0, 18, 0, 138, 61, 0, 3, 15, 0, 0, 0, 0, 0, 4, 
    11, 0, 0, 39, 132, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 105, 35, 0, 12, 0, 0, 0, 0, 0, 0, 0, 11, 
    30, 0, 0, 10, 13, 0, 0, 0, 0, 0, 10, 0, 0, 22, 48, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 12, 0, 0, 
    19, 25, 0, 0, 0, 0, 9, 6, 1, 0, 0, 0, 0, 9, 0, 
    4, 31, 0, 0, 29, 28, 0, 5, 0, 0, 3, 12, 6, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 15, 0, 0, 0, 4, 30, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 6, 5, 
    7, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 14, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 17, 14, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 22, 66, 68, 3, 0, 0, 20, 48, 61, 47, 17, 18, 
    0, 0, 0, 1, 0, 0, 0, 0, 9, 24, 30, 28, 34, 34, 31, 
    49, 0, 0, 0, 0, 28, 27, 26, 29, 37, 42, 48, 28, 21, 49, 
    38, 43, 0, 0, 1, 28, 37, 32, 26, 34, 31, 20, 29, 54, 5, 
    39, 37, 31, 0, 12, 8, 0, 20, 37, 45, 36, 31, 53, 55, 37, 
    
    -- channel=23
    0, 0, 5, 8, 9, 6, 4, 1, 9, 0, 0, 0, 2, 10, 7, 
    10, 10, 6, 7, 5, 58, 38, 11, 0, 1, 45, 28, 0, 0, 8, 
    0, 0, 5, 6, 1, 0, 0, 0, 13, 3, 13, 12, 30, 0, 0, 
    62, 27, 12, 7, 27, 3, 46, 23, 7, 0, 13, 0, 0, 11, 0, 
    52, 56, 35, 0, 104, 80, 24, 23, 0, 0, 34, 45, 12, 31, 0, 
    9, 0, 31, 0, 0, 0, 41, 30, 47, 0, 20, 0, 0, 17, 44, 
    28, 12, 0, 18, 0, 10, 0, 27, 22, 0, 8, 25, 3, 9, 26, 
    34, 16, 49, 37, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    29, 0, 43, 0, 40, 0, 0, 21, 0, 16, 0, 0, 0, 0, 24, 
    0, 0, 37, 0, 19, 6, 0, 54, 23, 0, 0, 0, 7, 15, 7, 
    0, 0, 16, 3, 142, 104, 8, 0, 11, 27, 33, 48, 27, 2, 9, 
    0, 0, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 9, 23, 6, 
    
    -- channel=24
    5, 14, 7, 12, 7, 10, 10, 4, 6, 13, 14, 8, 11, 10, 7, 
    5, 8, 6, 14, 5, 42, 31, 21, 18, 14, 44, 24, 0, 1, 11, 
    31, 0, 5, 9, 0, 6, 41, 4, 9, 21, 79, 58, 58, 0, 7, 
    93, 0, 13, 3, 29, 0, 65, 51, 42, 0, 91, 41, 51, 32, 0, 
    121, 58, 45, 0, 122, 76, 97, 69, 45, 0, 76, 80, 39, 57, 0, 
    93, 87, 65, 8, 38, 71, 121, 71, 79, 0, 115, 76, 30, 53, 39, 
    93, 123, 28, 52, 0, 45, 116, 89, 94, 0, 114, 69, 27, 39, 58, 
    107, 125, 54, 54, 3, 69, 117, 57, 68, 6, 93, 70, 24, 44, 32, 
    132, 103, 120, 53, 52, 21, 54, 59, 27, 34, 34, 56, 2, 18, 20, 
    109, 99, 150, 25, 103, 27, 22, 111, 49, 56, 57, 15, 15, 14, 25, 
    67, 96, 133, 14, 202, 111, 77, 118, 116, 48, 33, 49, 46, 36, 47, 
    34, 77, 113, 72, 179, 82, 43, 44, 65, 54, 63, 62, 71, 74, 81, 
    90, 26, 34, 150, 127, 70, 71, 62, 62, 62, 66, 76, 83, 77, 83, 
    100, 70, 0, 172, 86, 64, 78, 67, 64, 70, 72, 77, 78, 76, 103, 
    108, 79, 62, 60, 58, 49, 65, 71, 71, 80, 84, 65, 69, 121, 112, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 16, 6, 0, 
    20, 26, 0, 0, 0, 48, 13, 23, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 7, 3, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 3, 49, 1, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 4, 19, 0, 8, 0, 7, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 25, 1, 0, 0, 3, 0, 5, 0, 
    0, 0, 0, 0, 0, 45, 6, 0, 0, 7, 34, 36, 10, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 31, 32, 7, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 28, 3, 0, 0, 0, 0, 22, 25, 
    66, 15, 0, 0, 78, 64, 46, 45, 19, 6, 0, 1, 0, 0, 0, 
    0, 44, 0, 19, 55, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 27, 68, 3, 0, 0, 0, 0, 0, 0, 12, 2, 0, 37, 
    0, 0, 7, 70, 18, 18, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    48, 48, 49, 54, 53, 45, 52, 56, 55, 46, 32, 27, 35, 46, 50, 
    48, 50, 51, 56, 48, 48, 67, 47, 32, 10, 25, 23, 11, 20, 46, 
    46, 1, 53, 55, 53, 34, 42, 20, 12, 0, 35, 19, 34, 3, 17, 
    75, 0, 51, 48, 60, 20, 46, 34, 16, 0, 43, 19, 23, 18, 0, 
    56, 14, 67, 5, 57, 50, 51, 39, 22, 0, 37, 52, 17, 31, 0, 
    42, 7, 67, 50, 0, 18, 54, 44, 52, 0, 59, 40, 6, 23, 21, 
    38, 39, 16, 74, 0, 5, 41, 41, 52, 0, 53, 39, 8, 7, 35, 
    37, 35, 30, 48, 9, 2, 56, 15, 32, 0, 36, 41, 0, 15, 28, 
    42, 14, 62, 0, 46, 0, 26, 32, 0, 42, 13, 28, 0, 6, 40, 
    22, 18, 65, 0, 44, 14, 0, 48, 32, 18, 23, 0, 0, 18, 44, 
    0, 21, 59, 0, 83, 54, 0, 14, 32, 19, 0, 0, 0, 0, 4, 
    0, 0, 28, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 
    
    -- channel=27
    12, 0, 6, 5, 5, 1, 8, 6, 2, 7, 15, 11, 7, 10, 3, 
    6, 0, 2, 4, 3, 0, 33, 3, 14, 0, 0, 9, 11, 11, 3, 
    0, 12, 8, 3, 3, 0, 23, 16, 23, 0, 1, 6, 3, 27, 0, 
    0, 0, 12, 0, 0, 4, 0, 27, 3, 0, 6, 8, 7, 24, 0, 
    43, 0, 48, 20, 0, 35, 4, 17, 0, 8, 0, 31, 0, 4, 30, 
    104, 0, 67, 27, 0, 64, 0, 7, 0, 0, 36, 48, 0, 6, 25, 
    123, 0, 57, 0, 0, 0, 0, 25, 0, 0, 37, 23, 1, 0, 20, 
    92, 0, 82, 0, 0, 0, 46, 6, 16, 0, 11, 16, 0, 0, 25, 
    44, 0, 87, 0, 52, 16, 9, 0, 8, 0, 0, 33, 0, 0, 0, 
    0, 0, 23, 0, 33, 65, 13, 0, 45, 16, 20, 11, 0, 0, 16, 
    0, 9, 16, 0, 5, 30, 0, 0, 50, 14, 0, 0, 2, 0, 17, 
    0, 0, 38, 0, 14, 60, 0, 3, 14, 1, 0, 0, 0, 0, 0, 
    12, 0, 40, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 3, 17, 0, 25, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 8, 0, 6, 0, 0, 4, 0, 0, 0, 0, 0, 0, 17, 
    
    -- channel=28
    34, 41, 34, 38, 35, 34, 40, 36, 31, 38, 39, 35, 34, 32, 28, 
    34, 32, 34, 42, 32, 54, 48, 43, 40, 21, 39, 27, 19, 29, 35, 
    52, 30, 35, 37, 30, 48, 51, 12, 6, 27, 71, 57, 56, 14, 35, 
    76, 0, 42, 31, 47, 16, 59, 44, 44, 22, 87, 43, 47, 30, 6, 
    99, 68, 66, 0, 113, 65, 89, 57, 46, 0, 68, 65, 39, 49, 0, 
    76, 102, 81, 12, 64, 70, 108, 63, 67, 0, 110, 70, 37, 48, 30, 
    67, 124, 54, 57, 24, 46, 123, 84, 83, 17, 106, 56, 28, 34, 55, 
    82, 117, 53, 66, 13, 86, 124, 69, 67, 29, 90, 60, 28, 55, 48, 
    110, 101, 93, 66, 43, 41, 54, 51, 39, 46, 39, 62, 12, 33, 37, 
    107, 98, 126, 31, 90, 30, 30, 97, 46, 68, 67, 14, 27, 38, 48, 
    82, 92, 118, 17, 161, 80, 81, 126, 110, 42, 16, 30, 39, 49, 50, 
    60, 92, 106, 86, 173, 74, 39, 38, 52, 43, 52, 49, 55, 59, 62, 
    73, 43, 46, 152, 109, 54, 56, 50, 48, 46, 50, 57, 70, 63, 64, 
    79, 55, 16, 184, 70, 51, 58, 50, 49, 54, 57, 64, 62, 54, 96, 
    85, 60, 51, 71, 49, 43, 60, 59, 54, 60, 63, 50, 49, 95, 88, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 3, 4, 10, 2, 0, 
    4, 1, 0, 0, 0, 0, 0, 0, 12, 12, 0, 0, 8, 2, 0, 
    22, 32, 0, 0, 33, 0, 0, 0, 0, 21, 5, 7, 15, 9, 0, 
    19, 24, 0, 0, 0, 0, 8, 0, 3, 29, 10, 5, 12, 12, 3, 
    17, 29, 0, 0, 0, 17, 19, 18, 6, 16, 10, 8, 20, 13, 0, 
    27, 40, 14, 19, 0, 15, 1, 1, 10, 0, 6, 14, 14, 0, 0, 
    37, 41, 21, 31, 8, 1, 9, 1, 7, 9, 12, 12, 8, 0, 0, 
    48, 28, 23, 43, 3, 1, 33, 47, 27, 14, 30, 36, 43, 36, 25, 
    102, 68, 28, 32, 42, 75, 73, 73, 73, 71, 82, 86, 93, 94, 92, 
    103, 94, 59, 36, 67, 79, 78, 79, 80, 85, 92, 95, 97, 99, 104, 
    113, 96, 90, 76, 69, 84, 78, 79, 84, 91, 100, 108, 105, 113, 116, 
    109, 108, 91, 94, 80, 92, 94, 86, 81, 88, 92, 99, 100, 107, 103, 
    
    -- channel=30
    35, 38, 30, 31, 30, 31, 34, 39, 29, 25, 22, 24, 17, 17, 17, 
    26, 32, 32, 33, 32, 18, 5, 23, 25, 5, 0, 0, 14, 23, 16, 
    23, 51, 35, 36, 39, 104, 24, 13, 0, 8, 0, 0, 0, 4, 26, 
    0, 0, 29, 35, 18, 14, 0, 0, 0, 38, 0, 6, 0, 0, 31, 
    0, 0, 3, 22, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 40, 2, 34, 136, 30, 5, 0, 0, 22, 3, 0, 1, 0, 0, 
    0, 33, 30, 12, 66, 22, 45, 0, 0, 52, 6, 0, 0, 0, 0, 
    0, 17, 0, 0, 12, 59, 20, 37, 0, 61, 20, 0, 2, 12, 9, 
    0, 30, 0, 22, 0, 60, 22, 0, 0, 18, 53, 6, 10, 20, 12, 
    49, 37, 0, 23, 0, 0, 4, 0, 0, 24, 0, 0, 0, 11, 17, 
    67, 27, 1, 28, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 
    66, 50, 0, 61, 68, 32, 29, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 43, 30, 74, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    3, 0, 0, 1, 7, 0, 0, 4, 9, 1, 0, 0, 0, 3, 7, 
    8, 2, 0, 0, 1, 6, 13, 0, 0, 17, 26, 25, 12, 2, 3, 
    0, 0, 6, 5, 6, 0, 19, 35, 15, 0, 0, 0, 8, 6, 0, 
    24, 19, 13, 7, 8, 21, 4, 0, 0, 0, 0, 0, 5, 8, 0, 
    10, 0, 11, 0, 0, 0, 0, 0, 0, 8, 7, 5, 0, 4, 5, 
    2, 0, 5, 7, 0, 0, 0, 4, 12, 0, 0, 3, 0, 0, 12, 
    9, 0, 6, 5, 0, 0, 0, 0, 0, 0, 4, 13, 12, 3, 0, 
    0, 0, 20, 19, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 14, 0, 12, 0, 18, 9, 0, 41, 0, 0, 0, 0, 0, 
    0, 0, 2, 9, 0, 0, 5, 0, 0, 0, 0, 5, 0, 0, 4, 
    0, 0, 9, 0, 8, 0, 0, 0, 0, 24, 25, 4, 5, 22, 33, 
    0, 0, 0, 0, 0, 20, 19, 18, 8, 2, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 6, 0, 0, 0, 3, 2, 2, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 8, 1, 7, 0, 0, 0, 0, 3, 0, 1, 0, 0, 4, 
    
    
    others => 0);
end ifmap_package;
