library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    113, 9432, 5516, -364, -7354, 8721, -12605, 2341, -3759, -5175, 3397, -8637, -4899, 5114, -5064, 4018, -4891, -5353, -25189, -1254, 14621, -10862, -9102, -2929, 14904, 5953, 16902, 3147, 19864, 1889, -3451, -2593,

    -- weights
    -- filter=0 channel=0
    1, -7, 11, -13, -8, -14, -10, 7, -9,
    -- filter=0 channel=1
    -16, -9, 6, 16, -15, 20, 18, -9, 14,
    -- filter=0 channel=2
    -1, 2, 18, 0, -11, -10, -1, 5, -10,
    -- filter=0 channel=3
    1, 11, 5, 3, 4, 6, 19, 11, -5,
    -- filter=0 channel=4
    -3, 15, 7, 13, 16, 17, 12, 3, -13,
    -- filter=0 channel=5
    17, 14, -13, 20, 0, 12, -5, -7, 16,
    -- filter=0 channel=6
    -3, -1, 9, -10, 5, 3, 4, -13, 19,
    -- filter=0 channel=7
    -17, 6, -2, 3, 1, -2, -11, -14, -13,
    -- filter=0 channel=8
    14, -2, -7, 5, -10, -14, -15, -8, 1,
    -- filter=0 channel=9
    -13, 0, 12, -5, -13, -19, 14, 20, 19,
    -- filter=0 channel=10
    15, 4, 16, 12, 10, 8, 17, -6, -8,
    -- filter=0 channel=11
    4, 0, -5, 6, 1, 7, 3, 3, -7,
    -- filter=0 channel=12
    -3, -3, 0, -19, 17, -18, -21, -5, -10,
    -- filter=0 channel=13
    4, -10, -10, 8, -16, -9, 0, 16, 20,
    -- filter=0 channel=14
    10, -10, 6, -1, 15, -6, -9, -1, -3,
    -- filter=0 channel=15
    2, -18, 4, 10, -7, -20, 16, -17, -10,
    -- filter=1 channel=0
    19, 15, -7, -19, -3, 3, 4, 10, 2,
    -- filter=1 channel=1
    21, 4, -1, 25, 18, 7, 23, 0, 1,
    -- filter=1 channel=2
    0, -28, -36, 23, -25, -29, 20, 0, 5,
    -- filter=1 channel=3
    5, 14, 5, -6, 15, 21, -17, -7, -17,
    -- filter=1 channel=4
    4, -3, -16, 14, -9, -9, -15, -22, 5,
    -- filter=1 channel=5
    1, -17, 12, -10, -4, 7, -19, -6, 4,
    -- filter=1 channel=6
    -8, -8, 19, -9, 14, 15, 10, -9, 17,
    -- filter=1 channel=7
    -1, 15, 3, -8, 9, 18, -5, 14, 15,
    -- filter=1 channel=8
    15, 32, 25, -11, -3, 27, 18, -6, 16,
    -- filter=1 channel=9
    14, 11, 17, 14, 23, 35, 21, -4, 32,
    -- filter=1 channel=10
    29, -5, -8, 32, 24, 14, 27, 11, 0,
    -- filter=1 channel=11
    1, 23, 29, -6, 7, -8, -6, -12, -1,
    -- filter=1 channel=12
    7, -14, 4, 13, -9, 9, 0, 14, -30,
    -- filter=1 channel=13
    5, -13, 3, -3, 3, 3, 1, -17, -37,
    -- filter=1 channel=14
    -14, -22, -37, 5, 0, -14, 14, -18, -9,
    -- filter=1 channel=15
    0, -1, -27, 5, -16, 4, -23, -23, 5,
    -- filter=2 channel=0
    -4, 6, 16, 11, -7, 9, -15, -3, 17,
    -- filter=2 channel=1
    7, -15, 1, 3, -14, -7, -14, 0, 13,
    -- filter=2 channel=2
    9, 10, 1, -10, 23, 25, 17, 34, 12,
    -- filter=2 channel=3
    -1, 20, -11, 12, -4, -19, 8, -14, 0,
    -- filter=2 channel=4
    -33, -40, -44, -15, -6, -22, -39, -17, -28,
    -- filter=2 channel=5
    -10, -21, 2, -18, -17, -21, 1, -26, 11,
    -- filter=2 channel=6
    -8, 2, -16, -2, -1, 11, -8, -10, 6,
    -- filter=2 channel=7
    -18, 1, -22, -18, 2, 8, 0, -12, -19,
    -- filter=2 channel=8
    19, 12, 5, 0, 21, 17, 22, 13, 21,
    -- filter=2 channel=9
    6, 9, -17, -2, 0, -6, 9, -8, 10,
    -- filter=2 channel=10
    -7, 7, 11, -20, -4, -22, 5, -26, 12,
    -- filter=2 channel=11
    39, 9, 41, 31, 13, 39, 10, 39, 21,
    -- filter=2 channel=12
    -17, 6, 4, 12, 7, -10, 8, -2, 25,
    -- filter=2 channel=13
    -27, -27, -32, -13, 2, -16, -9, -13, -11,
    -- filter=2 channel=14
    -10, -22, 2, 17, 0, 14, -15, -18, 17,
    -- filter=2 channel=15
    -5, -20, -17, -5, -32, -28, -8, -14, -1,
    -- filter=3 channel=0
    6, -17, 13, -15, -5, 11, -13, 17, -14,
    -- filter=3 channel=1
    15, 0, -18, -12, 17, -6, 8, 3, -4,
    -- filter=3 channel=2
    25, -3, -16, 23, -14, -9, 25, -11, -4,
    -- filter=3 channel=3
    -8, 12, 2, 5, 4, 10, 8, 16, 7,
    -- filter=3 channel=4
    3, 19, 2, 25, 15, -7, 21, 28, -2,
    -- filter=3 channel=5
    0, -18, 15, 14, 17, 18, -10, 21, 12,
    -- filter=3 channel=6
    1, 17, -10, -9, -18, 18, 14, 4, 0,
    -- filter=3 channel=7
    12, 16, -6, -19, -11, -7, -15, 17, -1,
    -- filter=3 channel=8
    25, 22, -7, -16, 18, 15, -13, 18, -11,
    -- filter=3 channel=9
    -14, -17, -13, 3, -13, -14, 3, 0, 5,
    -- filter=3 channel=10
    15, 0, 0, -9, 15, 7, 11, 0, 17,
    -- filter=3 channel=11
    9, -4, 16, -6, 3, 14, -14, -12, 5,
    -- filter=3 channel=12
    19, -12, -12, 23, 6, 6, 16, -11, -23,
    -- filter=3 channel=13
    6, 3, -35, -16, -23, -7, 14, -6, 3,
    -- filter=3 channel=14
    12, -9, -23, 22, -10, -11, 15, -12, -10,
    -- filter=3 channel=15
    9, 2, -8, 12, -19, -11, -1, -7, -26,
    -- filter=4 channel=0
    -19, 19, -19, 1, -11, 0, 9, 11, 11,
    -- filter=4 channel=1
    -7, -11, 0, -10, 20, -15, 23, 0, -4,
    -- filter=4 channel=2
    22, -2, 0, -8, 18, 20, 26, -1, -9,
    -- filter=4 channel=3
    -14, 6, -18, -3, -17, 8, 16, 11, 16,
    -- filter=4 channel=4
    0, 0, -28, 5, -4, -5, -25, -31, -11,
    -- filter=4 channel=5
    1, -1, -3, -20, -24, -4, -9, 12, 14,
    -- filter=4 channel=6
    8, -21, 3, 14, 17, -15, 6, -14, 0,
    -- filter=4 channel=7
    -4, 4, -1, 7, -1, 16, -22, 20, 0,
    -- filter=4 channel=8
    -5, 12, 3, -8, 20, -5, 12, -5, 22,
    -- filter=4 channel=9
    -4, -8, -15, -5, 16, -6, -9, 4, 2,
    -- filter=4 channel=10
    -9, 12, -8, 11, 20, 8, 11, -10, 11,
    -- filter=4 channel=11
    19, 22, 22, 8, 36, 22, 19, 13, 12,
    -- filter=4 channel=12
    -13, -3, -20, -3, 7, 7, 0, 23, 23,
    -- filter=4 channel=13
    -11, -6, -23, -6, -4, -19, 1, 0, 15,
    -- filter=4 channel=14
    -17, 12, 0, -3, 19, 1, -4, 10, 6,
    -- filter=4 channel=15
    3, 11, 8, -24, -23, -14, 1, 10, -11,
    -- filter=5 channel=0
    14, 18, 7, 18, -16, 10, 4, -8, 9,
    -- filter=5 channel=1
    -12, -23, -7, -5, -17, -17, 10, -19, -23,
    -- filter=5 channel=2
    -1, 6, 19, 5, 14, -5, 22, 2, 22,
    -- filter=5 channel=3
    -5, -9, 5, 0, 7, 14, 8, 4, -3,
    -- filter=5 channel=4
    -16, 3, 6, -27, -15, 3, -20, -18, -3,
    -- filter=5 channel=5
    16, 0, 9, -24, 13, 4, -18, -15, -12,
    -- filter=5 channel=6
    -15, 11, -2, -14, 0, -5, 6, -6, -5,
    -- filter=5 channel=7
    -14, 2, -15, 12, -5, 16, 1, 1, 7,
    -- filter=5 channel=8
    -12, 2, 2, -24, 7, 14, -14, -17, 8,
    -- filter=5 channel=9
    -2, -29, -7, -45, -18, -24, -30, -44, -5,
    -- filter=5 channel=10
    -14, -3, -8, -16, 2, -21, -19, -2, -24,
    -- filter=5 channel=11
    11, 10, 25, -20, -12, -13, -16, -6, 2,
    -- filter=5 channel=12
    22, 32, 11, 18, 11, -6, -12, -13, -10,
    -- filter=5 channel=13
    0, 30, 17, 4, 26, -17, 2, 6, 1,
    -- filter=5 channel=14
    18, 0, 1, 26, 11, 14, -13, 1, 2,
    -- filter=5 channel=15
    5, -12, 26, 6, 20, 11, -11, 25, 6,
    -- filter=6 channel=0
    -2, -12, -14, -5, 7, -17, 14, -12, 1,
    -- filter=6 channel=1
    3, 8, 8, 26, 11, 7, -13, -11, 7,
    -- filter=6 channel=2
    -16, -13, 4, 13, -14, -7, -3, 6, 0,
    -- filter=6 channel=3
    0, -16, -6, -4, -19, 5, 1, -1, -5,
    -- filter=6 channel=4
    -17, -8, -9, -39, -1, -25, -16, -24, -26,
    -- filter=6 channel=5
    -6, 15, 14, 2, -26, -1, 0, -9, -17,
    -- filter=6 channel=6
    0, -18, -8, -8, 17, -13, 20, 18, 9,
    -- filter=6 channel=7
    -13, -8, 3, -6, 6, 16, -14, -11, -1,
    -- filter=6 channel=8
    11, 24, 15, 23, 4, -14, -2, 9, -25,
    -- filter=6 channel=9
    23, 0, 15, -6, 11, -4, 4, 12, -20,
    -- filter=6 channel=10
    31, 13, 13, 13, 29, 20, 19, -1, -15,
    -- filter=6 channel=11
    14, 17, 33, -15, 16, 0, -27, -2, 8,
    -- filter=6 channel=12
    21, 46, 30, 20, 37, 1, 5, 8, -18,
    -- filter=6 channel=13
    45, -1, 12, 26, 20, 1, 6, -12, -19,
    -- filter=6 channel=14
    24, 18, -2, 17, 17, 10, 20, -12, -5,
    -- filter=6 channel=15
    -3, 13, -5, 2, 0, 17, -10, -14, 5,
    -- filter=7 channel=0
    12, -14, 20, -13, -19, -15, -1, -17, 20,
    -- filter=7 channel=1
    17, 5, 10, -22, -21, 1, 2, -9, -23,
    -- filter=7 channel=2
    -4, 7, 13, -23, -10, 22, -14, 9, 23,
    -- filter=7 channel=3
    -14, 8, 11, -16, 8, 12, -18, -18, 10,
    -- filter=7 channel=4
    -25, -10, 2, -25, -6, -6, 12, -25, 8,
    -- filter=7 channel=5
    -9, -14, -3, -3, -16, -16, 14, -2, -5,
    -- filter=7 channel=6
    4, 2, -18, -17, 0, 3, 4, -10, 14,
    -- filter=7 channel=7
    17, 13, 4, -21, -9, 8, 10, 16, 16,
    -- filter=7 channel=8
    -16, -8, -16, 23, 21, -9, 7, 23, 0,
    -- filter=7 channel=9
    12, -25, -14, 2, -14, -12, -10, 0, -28,
    -- filter=7 channel=10
    -2, -28, 6, -6, -6, 11, 0, -20, -18,
    -- filter=7 channel=11
    19, -11, -6, 21, 7, 27, 0, -3, 8,
    -- filter=7 channel=12
    -14, -20, -2, -11, 4, 26, 8, 29, 27,
    -- filter=7 channel=13
    16, 12, 9, -18, 16, 11, 3, -8, 21,
    -- filter=7 channel=14
    -14, -9, -14, 3, -1, 9, -8, -9, 20,
    -- filter=7 channel=15
    0, -4, -1, 20, 18, 27, 17, -16, 27,
    -- filter=8 channel=0
    -5, 4, 19, -7, 13, 0, -19, -1, 0,
    -- filter=8 channel=1
    -18, 2, -13, 2, -4, 9, 1, 9, 9,
    -- filter=8 channel=2
    20, -17, -18, 6, -16, 3, -5, -3, -4,
    -- filter=8 channel=3
    -17, 7, 3, -7, 16, 16, 1, -4, 18,
    -- filter=8 channel=4
    16, 10, 33, -9, 18, 23, 19, 1, 21,
    -- filter=8 channel=5
    2, 21, -1, 21, 2, -19, -14, -14, 10,
    -- filter=8 channel=6
    -16, 3, -10, -10, -18, -12, 8, 1, 6,
    -- filter=8 channel=7
    -6, 5, 17, -11, 5, 15, -2, -14, -9,
    -- filter=8 channel=8
    16, 1, -7, -18, 6, 10, -24, 4, 11,
    -- filter=8 channel=9
    19, 10, 25, -23, 7, -4, 8, 5, -17,
    -- filter=8 channel=10
    -10, -12, -16, -18, 7, -16, -19, -10, 12,
    -- filter=8 channel=11
    21, 21, -2, 7, 19, 13, 12, -21, -20,
    -- filter=8 channel=12
    25, 16, 10, -14, 7, -14, 13, -22, -24,
    -- filter=8 channel=13
    21, -4, -3, 5, -8, -7, 7, -2, -15,
    -- filter=8 channel=14
    2, -4, -13, -1, 16, 0, 4, 12, 11,
    -- filter=8 channel=15
    7, -8, -9, 22, -7, 16, -10, 9, 14,
    -- filter=9 channel=0
    -15, -11, -1, 18, 20, 13, 13, -16, 5,
    -- filter=9 channel=1
    -21, -13, 7, 0, -18, -2, 2, -24, -22,
    -- filter=9 channel=2
    5, 25, 19, -11, 0, 0, 16, -7, -9,
    -- filter=9 channel=3
    4, -6, 11, 19, 4, -11, 1, -1, 6,
    -- filter=9 channel=4
    0, -15, -26, 7, -12, -18, -11, 4, 10,
    -- filter=9 channel=5
    -23, -18, 0, 12, 16, 12, 11, 4, 6,
    -- filter=9 channel=6
    0, -15, -11, -9, -19, -5, -1, 11, -18,
    -- filter=9 channel=7
    -10, 17, -17, -15, 11, 13, 0, -3, 6,
    -- filter=9 channel=8
    -17, -7, 5, -1, -8, 11, -1, -16, 6,
    -- filter=9 channel=9
    -27, -3, -6, -24, -21, -6, -9, 4, 3,
    -- filter=9 channel=10
    -8, -24, -1, -10, 7, -19, -8, 0, -11,
    -- filter=9 channel=11
    17, 2, 31, 32, 29, 4, 0, 12, -13,
    -- filter=9 channel=12
    3, 9, 23, 9, -11, 10, 8, 22, 9,
    -- filter=9 channel=13
    3, -2, 7, -2, 20, 20, 5, -19, -17,
    -- filter=9 channel=14
    -20, 10, 17, -4, 18, -14, 4, 27, 6,
    -- filter=9 channel=15
    -1, 6, 11, -18, -18, 6, -21, 2, 0,
    -- filter=10 channel=0
    -3, -3, -2, 7, -15, 15, 9, -11, 1,
    -- filter=10 channel=1
    -13, 3, -2, 0, -15, -8, -11, 18, -19,
    -- filter=10 channel=2
    0, 7, 23, -7, -3, 18, -3, -10, 9,
    -- filter=10 channel=3
    17, 2, 19, 17, -13, 0, 21, -20, -3,
    -- filter=10 channel=4
    17, -15, -13, -14, -6, 4, -15, -15, -16,
    -- filter=10 channel=5
    -13, 10, 20, 5, 11, 8, 2, -12, -2,
    -- filter=10 channel=6
    1, 17, -9, -6, 6, 4, 7, 6, -9,
    -- filter=10 channel=7
    -5, 16, -19, 0, 13, 8, -13, -11, -3,
    -- filter=10 channel=8
    12, -5, 4, -12, 10, -10, 10, -10, -6,
    -- filter=10 channel=9
    7, 14, -5, -1, 1, 5, -11, 3, 18,
    -- filter=10 channel=10
    19, -16, 11, -20, -8, -2, -2, 13, 2,
    -- filter=10 channel=11
    18, 15, -3, -10, -5, 18, 1, 3, -6,
    -- filter=10 channel=12
    -12, -8, 1, -3, -18, 8, -21, -10, 2,
    -- filter=10 channel=13
    0, 11, -16, -3, -20, -12, 20, -20, -12,
    -- filter=10 channel=14
    17, -14, -15, -17, -1, -18, -3, -13, 8,
    -- filter=10 channel=15
    -1, 0, 10, -12, 6, -10, -9, 12, -3,
    -- filter=11 channel=0
    -2, 13, -5, -3, 16, 8, 4, 1, 15,
    -- filter=11 channel=1
    -13, 24, 2, -15, 15, 7, -9, 0, 17,
    -- filter=11 channel=2
    12, -19, -6, 12, -19, 5, -7, -21, -6,
    -- filter=11 channel=3
    6, 20, 15, -13, -6, 3, -7, 3, -10,
    -- filter=11 channel=4
    -12, 2, 44, 6, 25, 30, -21, -11, 16,
    -- filter=11 channel=5
    -16, -1, 12, 4, 2, -15, 2, -8, -7,
    -- filter=11 channel=6
    0, 20, 16, -4, -20, -2, 16, -16, 13,
    -- filter=11 channel=7
    -21, 11, 13, -12, -12, -12, -5, 16, 18,
    -- filter=11 channel=8
    -18, 0, -20, -7, 7, 16, -6, -8, 0,
    -- filter=11 channel=9
    -6, -4, -12, -21, -25, 2, 5, -35, -31,
    -- filter=11 channel=10
    15, 11, -9, 21, -10, -3, -1, -1, -18,
    -- filter=11 channel=11
    -14, 17, 14, -15, 2, 17, -19, -8, -15,
    -- filter=11 channel=12
    35, 13, 17, 26, 17, 9, 21, 30, -11,
    -- filter=11 channel=13
    30, 18, -10, 37, 33, -8, 37, 30, -5,
    -- filter=11 channel=14
    15, 9, -16, 14, -1, -9, 24, 34, 22,
    -- filter=11 channel=15
    -4, 16, 3, 37, 3, -1, 35, 35, 6,
    -- filter=12 channel=0
    9, 11, -18, 8, 13, 3, 9, 16, 2,
    -- filter=12 channel=1
    17, -17, -10, -20, 9, -17, 2, -6, 18,
    -- filter=12 channel=2
    25, -3, 16, 0, -3, 2, 5, 20, 22,
    -- filter=12 channel=3
    -13, 10, -17, 13, -17, 4, -10, 10, 14,
    -- filter=12 channel=4
    13, 9, -11, -13, 15, 25, -8, 20, 22,
    -- filter=12 channel=5
    -8, 20, 12, 20, 0, 22, 16, 4, -1,
    -- filter=12 channel=6
    -9, -17, -4, 15, -3, -1, 10, -11, -8,
    -- filter=12 channel=7
    3, 22, 19, 12, -2, 2, 11, 2, -3,
    -- filter=12 channel=8
    -1, 7, -12, -9, 6, -18, -10, 1, 8,
    -- filter=12 channel=9
    3, 5, -7, 7, -16, -19, 0, 19, 19,
    -- filter=12 channel=10
    -7, -6, 19, -12, -3, -10, -12, 19, 4,
    -- filter=12 channel=11
    -11, 15, -15, -8, 0, 0, 19, 17, -12,
    -- filter=12 channel=12
    2, -11, 0, -27, 10, -7, 4, -20, 12,
    -- filter=12 channel=13
    -20, -23, 11, -11, -18, -14, -18, -11, 21,
    -- filter=12 channel=14
    23, -13, 10, 17, 18, 10, -11, -4, 7,
    -- filter=12 channel=15
    6, -1, 4, 15, -5, 10, 7, 14, 3,
    -- filter=13 channel=0
    7, -20, 4, 6, -16, 9, -20, 13, -8,
    -- filter=13 channel=1
    17, 15, 7, 14, 18, 14, 9, -12, 15,
    -- filter=13 channel=2
    -16, -19, 7, -11, -23, -10, 18, -21, -11,
    -- filter=13 channel=3
    -15, 15, 9, 20, -12, -20, -15, 0, 18,
    -- filter=13 channel=4
    37, 3, 7, 47, 37, 10, 13, 37, 30,
    -- filter=13 channel=5
    13, -9, 11, -17, 11, 0, 3, 5, 14,
    -- filter=13 channel=6
    3, 3, 19, 18, -2, -19, -10, -11, -16,
    -- filter=13 channel=7
    -11, -3, 23, -6, 0, -13, -6, 19, -14,
    -- filter=13 channel=8
    31, 20, -2, 3, -2, -14, 30, 24, -8,
    -- filter=13 channel=9
    -13, -18, -22, -1, 1, 9, -18, 12, -6,
    -- filter=13 channel=10
    30, -15, -20, 12, 14, -9, -8, 5, -25,
    -- filter=13 channel=11
    19, -6, -28, 10, 5, -1, 9, 23, 4,
    -- filter=13 channel=12
    18, -9, -37, 36, -11, -19, 31, 4, -43,
    -- filter=13 channel=13
    4, -20, -23, 21, -39, -15, 8, -29, -38,
    -- filter=13 channel=14
    13, 8, 1, -9, -7, 0, 23, -29, -1,
    -- filter=13 channel=15
    22, -15, 17, 19, -14, -5, 27, -11, 3,
    -- filter=14 channel=0
    9, -19, 19, 12, 15, -20, -9, 2, -3,
    -- filter=14 channel=1
    -19, 20, -15, 4, 3, -20, -17, -15, 3,
    -- filter=14 channel=2
    16, -19, -9, 14, 9, 19, -14, 1, 15,
    -- filter=14 channel=3
    -18, -20, -20, 8, 19, -16, 0, -6, 20,
    -- filter=14 channel=4
    9, -16, -21, 8, 13, 19, 9, -5, 8,
    -- filter=14 channel=5
    -9, 9, 9, 17, -6, 3, -4, 0, 2,
    -- filter=14 channel=6
    4, 0, -3, -8, 18, 19, 5, -19, -3,
    -- filter=14 channel=7
    -3, 1, 19, -4, 19, 2, -12, 14, -18,
    -- filter=14 channel=8
    15, -6, -4, -7, 4, 1, 0, 20, -14,
    -- filter=14 channel=9
    6, 11, 20, -17, -5, -18, -20, 6, 10,
    -- filter=14 channel=10
    19, 6, -11, -20, -3, 2, 8, 0, -15,
    -- filter=14 channel=11
    -21, 0, 0, 19, -18, 0, 4, -6, 18,
    -- filter=14 channel=12
    5, -14, -10, -12, -12, -20, 1, 0, 4,
    -- filter=14 channel=13
    -3, 3, -15, -11, -5, -5, 4, -7, -5,
    -- filter=14 channel=14
    9, -15, -8, -4, -10, -19, -16, -13, -3,
    -- filter=14 channel=15
    -6, 19, 17, -5, -11, -8, -11, -8, 3,
    -- filter=15 channel=0
    0, 2, 1, -10, -18, 18, -8, 20, 10,
    -- filter=15 channel=1
    -4, 13, -6, 0, 14, 13, -20, 0, 7,
    -- filter=15 channel=2
    20, -21, -5, 15, 2, -14, 0, 16, -6,
    -- filter=15 channel=3
    0, -3, 9, 10, 11, -5, -10, 2, 14,
    -- filter=15 channel=4
    28, 16, -8, 6, -11, 6, 6, 6, -14,
    -- filter=15 channel=5
    11, -5, 12, -19, -7, 20, -19, -4, 16,
    -- filter=15 channel=6
    20, 8, 9, -10, -19, -18, -15, -16, 11,
    -- filter=15 channel=7
    -16, -17, 4, -13, 19, -15, 14, -17, 8,
    -- filter=15 channel=8
    29, -1, -9, 16, 12, -9, 9, 11, 11,
    -- filter=15 channel=9
    10, 20, -2, -4, 11, 16, -7, 23, -8,
    -- filter=15 channel=10
    -7, 5, 5, 11, 0, 17, 22, -13, -7,
    -- filter=15 channel=11
    23, 19, 7, 28, 28, 8, 30, 34, 17,
    -- filter=15 channel=12
    2, -12, -30, 25, -21, -4, 4, 13, -13,
    -- filter=15 channel=13
    -25, -30, 3, -26, -34, -26, -13, -17, 0,
    -- filter=15 channel=14
    -2, 0, -18, 2, 10, -13, 23, -20, -17,
    -- filter=15 channel=15
    6, -21, -2, 7, -19, -29, 14, -19, -12,
    -- filter=16 channel=0
    -17, 4, 17, -14, 4, -10, -21, -9, -1,
    -- filter=16 channel=1
    -20, 11, 11, -16, 15, -13, 9, 8, -18,
    -- filter=16 channel=2
    -7, 14, 17, 21, 13, -18, -2, -18, -12,
    -- filter=16 channel=3
    5, 6, -12, -9, -9, 3, 11, -21, 13,
    -- filter=16 channel=4
    0, -14, 4, -7, 15, 2, 24, 20, 18,
    -- filter=16 channel=5
    6, 10, -12, -12, 17, 3, 4, 13, 19,
    -- filter=16 channel=6
    -12, -3, 14, 18, 20, 3, -19, 10, 18,
    -- filter=16 channel=7
    -4, -12, 14, 17, 22, -15, 16, 12, -4,
    -- filter=16 channel=8
    -3, -10, 12, -16, -4, 3, -10, 23, 13,
    -- filter=16 channel=9
    -11, -18, 2, 19, 15, 16, 26, 22, 9,
    -- filter=16 channel=10
    -5, 10, -10, -12, 17, -10, 12, -6, 19,
    -- filter=16 channel=11
    0, -6, -20, 1, -5, -7, 6, 21, 23,
    -- filter=16 channel=12
    -23, -12, 8, -28, -7, -6, 16, 22, -9,
    -- filter=16 channel=13
    -26, 9, 6, -5, -18, -21, -3, -3, 7,
    -- filter=16 channel=14
    21, 23, 9, 15, -24, -14, 12, 1, 14,
    -- filter=16 channel=15
    13, -14, 9, 11, -8, -11, -18, -3, 11,
    -- filter=17 channel=0
    -8, -8, 17, -15, -8, -20, 13, 5, 4,
    -- filter=17 channel=1
    -6, 4, -1, -10, 13, -5, 17, 2, 11,
    -- filter=17 channel=2
    0, 4, 14, 2, -8, 9, -3, -18, -12,
    -- filter=17 channel=3
    -16, -19, 20, -10, -9, 16, 4, 10, 1,
    -- filter=17 channel=4
    37, 15, 34, 15, 37, 34, 2, 31, 25,
    -- filter=17 channel=5
    16, -3, 20, 19, -6, 27, 7, 23, 5,
    -- filter=17 channel=6
    20, -3, 17, -5, -19, 20, -1, -12, -6,
    -- filter=17 channel=7
    9, -6, 21, 11, 15, 2, 21, -15, -2,
    -- filter=17 channel=8
    -29, -37, -3, -20, 0, 18, -20, 12, 13,
    -- filter=17 channel=9
    19, 17, 8, 21, 22, 37, 19, 18, 14,
    -- filter=17 channel=10
    -18, 19, -8, 11, -7, -12, 15, 23, -1,
    -- filter=17 channel=11
    2, -14, 13, -6, -8, 13, 13, 4, 11,
    -- filter=17 channel=12
    -21, -15, -12, -13, -12, 17, 25, 33, 30,
    -- filter=17 channel=13
    -18, 0, -6, -12, -13, 14, 24, 17, 32,
    -- filter=17 channel=14
    -5, 5, 9, -6, -25, -20, -12, 14, -8,
    -- filter=17 channel=15
    -6, -14, -13, 9, 7, 1, -12, -15, -2,
    -- filter=18 channel=0
    -15, 20, -6, 6, 18, 16, -20, -6, 5,
    -- filter=18 channel=1
    2, 25, 12, -10, 8, 16, 25, -4, 0,
    -- filter=18 channel=2
    -15, -11, -8, 14, -17, -11, 14, 2, -9,
    -- filter=18 channel=3
    -1, -18, -4, -18, -8, 13, 3, -2, -3,
    -- filter=18 channel=4
    -1, 1, 20, -15, 34, 41, 12, 28, 24,
    -- filter=18 channel=5
    15, 19, -4, 9, -20, 6, 15, 1, 12,
    -- filter=18 channel=6
    6, 8, -6, 14, 0, -17, 11, -8, 0,
    -- filter=18 channel=7
    -20, 13, -3, 9, 8, 0, -1, 19, 8,
    -- filter=18 channel=8
    -22, -6, -8, -13, 4, -1, 0, -1, -8,
    -- filter=18 channel=9
    12, 21, -13, 11, 16, -8, 9, 4, -16,
    -- filter=18 channel=10
    15, 9, 6, 25, -7, 10, 21, 28, -19,
    -- filter=18 channel=11
    -11, 17, 25, -23, 17, -1, -41, -23, -21,
    -- filter=18 channel=12
    18, 30, -6, 9, 47, -4, 33, 26, -12,
    -- filter=18 channel=13
    26, 5, 1, 37, 34, -2, 36, 3, 0,
    -- filter=18 channel=14
    -13, 3, 2, 11, 15, 0, 38, 16, 5,
    -- filter=18 channel=15
    -3, -1, 22, 19, 2, 8, 27, 32, 21,
    -- filter=19 channel=0
    8, -8, -1, -14, 13, 1, -11, 10, -19,
    -- filter=19 channel=1
    6, 5, 0, 14, -17, -4, 5, -13, 7,
    -- filter=19 channel=2
    -4, 18, 16, -17, 19, -6, 9, -11, 15,
    -- filter=19 channel=3
    9, 3, -3, 14, 3, 11, 1, 0, -10,
    -- filter=19 channel=4
    -6, 15, 7, 9, 17, 0, 6, 11, -18,
    -- filter=19 channel=5
    6, -17, -4, -20, 12, -16, 8, 14, 19,
    -- filter=19 channel=6
    -8, -8, 1, 1, 6, -11, -14, -20, -17,
    -- filter=19 channel=7
    11, 5, 10, 8, -8, 6, -19, 0, 17,
    -- filter=19 channel=8
    4, -4, 0, 18, 8, -4, -19, -18, 17,
    -- filter=19 channel=9
    -8, -15, -9, 6, -9, 19, -6, -7, -16,
    -- filter=19 channel=10
    -2, -14, 4, 2, -3, -10, -4, 15, -12,
    -- filter=19 channel=11
    2, 10, 1, 14, 5, 18, -5, -18, 0,
    -- filter=19 channel=12
    13, 15, 18, 7, -20, -8, -4, -14, 19,
    -- filter=19 channel=13
    0, -8, -5, -16, -21, 7, -14, -3, 4,
    -- filter=19 channel=14
    16, -3, 7, 5, -16, -14, 20, -2, 5,
    -- filter=19 channel=15
    -15, 7, 19, -5, -20, -8, 0, -18, -16,
    -- filter=20 channel=0
    8, 6, -18, 19, -16, 17, 11, -14, 2,
    -- filter=20 channel=1
    -17, 2, -4, 0, -12, -14, 4, 9, 17,
    -- filter=20 channel=2
    4, 14, -1, 28, 19, 23, 9, 34, -5,
    -- filter=20 channel=3
    -3, -18, -10, 4, -18, -10, -9, 19, 16,
    -- filter=20 channel=4
    2, -24, -3, -20, -26, -19, -17, -30, -14,
    -- filter=20 channel=5
    17, -11, -20, 5, 2, 0, 15, 0, -7,
    -- filter=20 channel=6
    -7, -20, -2, -11, 9, -5, 10, 20, -6,
    -- filter=20 channel=7
    -12, 0, -7, -19, 9, 0, -15, 15, 1,
    -- filter=20 channel=8
    -1, -25, -12, -23, -20, -13, 9, 6, 9,
    -- filter=20 channel=9
    -21, -4, 14, -3, -23, 5, -15, -19, 10,
    -- filter=20 channel=10
    -18, -29, -3, -3, -26, -4, 0, 3, -3,
    -- filter=20 channel=11
    -16, 11, 0, 11, 23, 26, -4, 26, 13,
    -- filter=20 channel=12
    -26, -15, -6, 19, 8, 19, 18, 19, 25,
    -- filter=20 channel=13
    -21, -1, -23, 0, 10, 2, 5, 19, -9,
    -- filter=20 channel=14
    17, -6, 0, -20, 22, -8, -9, 8, 5,
    -- filter=20 channel=15
    -1, 7, -4, -3, 9, -2, 17, 25, 13,
    -- filter=21 channel=0
    -3, -18, -17, -12, -5, -10, 1, 12, -6,
    -- filter=21 channel=1
    19, 26, 20, 24, 9, -12, -1, -12, 10,
    -- filter=21 channel=2
    27, -10, -37, 10, 0, -4, 21, 21, -9,
    -- filter=21 channel=3
    12, 11, 19, 9, -6, 10, 7, -9, -17,
    -- filter=21 channel=4
    0, -9, 6, 2, 4, 25, -21, -16, 22,
    -- filter=21 channel=5
    12, -13, -2, 18, -17, 8, -11, -25, -18,
    -- filter=21 channel=6
    -16, -9, 16, 12, -7, -20, -10, 0, 11,
    -- filter=21 channel=7
    8, -6, -4, -21, 2, -3, -21, -10, 3,
    -- filter=21 channel=8
    16, 20, 30, 6, 35, 20, 9, 2, 0,
    -- filter=21 channel=9
    15, 1, 26, 10, -3, -8, 3, 6, -17,
    -- filter=21 channel=10
    7, 33, -13, 5, 36, 1, 26, 32, -19,
    -- filter=21 channel=11
    -6, 25, 24, 0, 23, 19, -21, -24, -7,
    -- filter=21 channel=12
    17, 47, 16, 35, 31, 18, 18, -6, -18,
    -- filter=21 channel=13
    25, 30, -35, 46, 20, -34, 10, 5, -56,
    -- filter=21 channel=14
    0, 18, -28, 21, 23, -12, 20, 0, -10,
    -- filter=21 channel=15
    -10, 17, 0, 19, -4, -21, 14, 13, 0,
    -- filter=22 channel=0
    -19, 4, -15, 10, 12, 5, -9, -18, 19,
    -- filter=22 channel=1
    -8, 18, 15, -10, 10, 0, -3, -9, 10,
    -- filter=22 channel=2
    4, -4, -33, 0, -17, -7, -3, -3, -32,
    -- filter=22 channel=3
    14, -9, 0, -2, -13, 17, 15, -11, 6,
    -- filter=22 channel=4
    -11, -5, -6, -14, 13, -23, -20, -17, -20,
    -- filter=22 channel=5
    22, -15, 7, 20, -8, 11, -1, 11, -16,
    -- filter=22 channel=6
    4, 16, 15, 0, 6, -20, 14, 17, -2,
    -- filter=22 channel=7
    0, -21, -2, -5, -4, 13, -13, -5, -18,
    -- filter=22 channel=8
    -7, 0, -3, 21, 27, 15, 17, 27, 0,
    -- filter=22 channel=9
    21, 13, 7, 29, 10, 9, 15, -2, -4,
    -- filter=22 channel=10
    29, 31, -1, 25, 17, 5, -6, 16, 14,
    -- filter=22 channel=11
    -4, 13, -13, -26, -16, -9, -33, -13, -29,
    -- filter=22 channel=12
    21, 8, -3, 23, 35, 8, -10, 3, 7,
    -- filter=22 channel=13
    36, 0, 13, 34, 22, -1, 33, 2, 13,
    -- filter=22 channel=14
    6, -12, 0, 0, -9, -5, 0, 12, 0,
    -- filter=22 channel=15
    15, -2, -10, 1, 20, -9, -10, 19, -5,
    -- filter=23 channel=0
    5, 4, 1, -7, -18, -11, -16, 7, -20,
    -- filter=23 channel=1
    18, 15, -4, 11, 6, -8, -21, 18, -16,
    -- filter=23 channel=2
    -7, -18, -12, -7, -18, 12, 15, -14, 12,
    -- filter=23 channel=3
    -15, -3, 18, -17, -17, 12, 2, 11, 9,
    -- filter=23 channel=4
    -19, 12, -12, -18, 3, -5, 8, -6, -2,
    -- filter=23 channel=5
    -12, 9, -19, -8, 19, 2, 10, 4, 10,
    -- filter=23 channel=6
    5, -9, 0, 0, -13, -17, 2, 11, -6,
    -- filter=23 channel=7
    0, -19, -18, -1, 17, -12, 15, 11, 2,
    -- filter=23 channel=8
    -9, -11, -11, 14, -5, -12, -6, -15, -5,
    -- filter=23 channel=9
    -8, 20, -8, 7, 11, 8, -10, -5, -4,
    -- filter=23 channel=10
    2, -1, 2, -1, 9, 15, -21, -2, -6,
    -- filter=23 channel=11
    19, -3, -8, -9, -2, -16, 10, 0, -13,
    -- filter=23 channel=12
    -12, 17, -3, 12, 7, -12, 9, -15, 3,
    -- filter=23 channel=13
    3, -4, -15, 12, -5, -16, -17, 14, -3,
    -- filter=23 channel=14
    -2, -18, 12, 11, 6, 3, 15, -7, 8,
    -- filter=23 channel=15
    -11, -20, -17, 0, -7, 11, 11, -19, -8,
    -- filter=24 channel=0
    -19, 13, -1, -10, 8, 16, 5, 0, 21,
    -- filter=24 channel=1
    4, -27, -1, -17, -27, -10, -16, 10, -3,
    -- filter=24 channel=2
    26, 31, 30, 12, 35, 24, 5, 23, 10,
    -- filter=24 channel=3
    11, -19, 7, 14, -2, -15, 10, 12, 10,
    -- filter=24 channel=4
    -19, 1, -24, -31, -16, 0, -13, 3, 0,
    -- filter=24 channel=5
    -21, -11, -3, 0, -9, 3, 17, 0, 17,
    -- filter=24 channel=6
    -17, 0, 18, 13, 10, -15, 16, -6, 8,
    -- filter=24 channel=7
    4, -4, -3, -16, -17, -13, 19, -13, 3,
    -- filter=24 channel=8
    -6, -4, 1, 7, -5, -20, -26, -28, -20,
    -- filter=24 channel=9
    -24, -35, -15, -34, -34, -42, -28, -16, -24,
    -- filter=24 channel=10
    12, -26, -17, 0, 7, -2, -10, 2, -3,
    -- filter=24 channel=11
    16, -16, -11, -14, -2, -12, -18, -11, -22,
    -- filter=24 channel=12
    17, 19, 8, -1, -9, 8, -29, -10, 16,
    -- filter=24 channel=13
    -1, 23, 17, -7, -18, 10, -18, 13, 6,
    -- filter=24 channel=14
    -4, 2, 25, 13, 20, -8, 0, 17, -13,
    -- filter=24 channel=15
    23, 24, -7, -12, 19, 14, -17, 12, 27,
    -- filter=25 channel=0
    17, 10, -2, -7, 4, 7, 21, -10, 16,
    -- filter=25 channel=1
    -26, 1, 0, -20, -26, -18, 11, 13, -1,
    -- filter=25 channel=2
    -8, 39, 24, 33, 35, 26, 22, 40, 25,
    -- filter=25 channel=3
    -10, 14, 6, 12, 0, 18, 12, 8, 13,
    -- filter=25 channel=4
    -32, -42, -6, -37, -37, -18, -44, -43, -15,
    -- filter=25 channel=5
    9, 14, -18, -18, -26, -28, -9, -13, -11,
    -- filter=25 channel=6
    21, -5, -3, -1, 11, -19, 10, -19, -5,
    -- filter=25 channel=7
    -23, -10, 13, -23, 10, -24, 0, -10, -1,
    -- filter=25 channel=8
    -8, -9, -1, -15, 15, 23, -11, -19, 11,
    -- filter=25 channel=9
    3, -38, -34, -10, -15, -8, -28, -10, -22,
    -- filter=25 channel=10
    -15, -19, -4, -1, 6, -24, -16, 0, -8,
    -- filter=25 channel=11
    17, 19, 3, -8, 11, 21, -19, -12, 12,
    -- filter=25 channel=12
    11, 27, 30, -2, 34, 40, 5, -3, 1,
    -- filter=25 channel=13
    -15, 10, -7, -2, 10, 9, 4, 0, -14,
    -- filter=25 channel=14
    1, 18, 1, 7, 27, 15, 21, 21, -6,
    -- filter=25 channel=15
    -14, -16, 17, 4, 9, 22, 14, -5, -5,
    -- filter=26 channel=0
    -17, -14, -13, 0, -17, -1, 16, 8, -7,
    -- filter=26 channel=1
    1, -14, -23, -10, 4, -22, -6, 0, -4,
    -- filter=26 channel=2
    -10, 17, 35, 12, -7, 30, -7, 9, 34,
    -- filter=26 channel=3
    19, 14, 12, -12, 17, 1, 19, 8, 1,
    -- filter=26 channel=4
    -7, 7, 4, 15, -11, -10, 0, 22, 21,
    -- filter=26 channel=5
    0, 12, -6, -21, -9, -13, -1, 2, -12,
    -- filter=26 channel=6
    13, 15, 0, -19, 14, 5, 20, 5, -19,
    -- filter=26 channel=7
    13, 15, -17, -14, -11, 17, -4, -4, -19,
    -- filter=26 channel=8
    -11, -6, -6, -2, -15, 14, 18, 11, -9,
    -- filter=26 channel=9
    -15, -27, -29, 10, -10, -29, 18, -10, 0,
    -- filter=26 channel=10
    7, -18, -21, 0, -31, -8, -16, -16, -3,
    -- filter=26 channel=11
    0, 10, -8, 19, 0, -3, 23, 28, 33,
    -- filter=26 channel=12
    -18, 0, 4, -12, -26, -23, 17, 10, 12,
    -- filter=26 channel=13
    3, -19, -9, -2, 6, -1, -5, -14, 13,
    -- filter=26 channel=14
    11, 18, 20, -7, 7, 19, -17, -20, -12,
    -- filter=26 channel=15
    -13, -11, 11, -17, 10, 17, -13, 11, 0,
    -- filter=27 channel=0
    16, -13, -7, -12, -15, 16, 19, -21, 9,
    -- filter=27 channel=1
    -7, 15, 20, -5, 19, 17, -5, -12, -7,
    -- filter=27 channel=2
    -15, 0, -8, -1, -26, -9, 10, -5, -17,
    -- filter=27 channel=3
    8, -8, -19, -17, -14, 20, -9, -1, -15,
    -- filter=27 channel=4
    -27, -14, -9, -31, 1, 6, -20, -24, 17,
    -- filter=27 channel=5
    19, -9, -1, -3, -2, 6, -11, 8, -19,
    -- filter=27 channel=6
    -14, 4, -11, 0, -4, -15, 2, 10, -11,
    -- filter=27 channel=7
    -16, 18, -13, -14, -14, 3, 1, 19, 8,
    -- filter=27 channel=8
    22, -6, 7, 28, 1, 23, 9, -8, 22,
    -- filter=27 channel=9
    35, 36, 44, 16, 39, 33, 4, 23, 34,
    -- filter=27 channel=10
    30, 14, 7, 16, 41, 37, 24, 13, 0,
    -- filter=27 channel=11
    -3, -8, 4, -4, 20, -2, 16, -15, -4,
    -- filter=27 channel=12
    23, 0, 8, 25, 20, -13, 12, -20, -27,
    -- filter=27 channel=13
    -6, -14, 4, -1, -1, -1, 20, -23, -3,
    -- filter=27 channel=14
    -11, -28, 0, -16, -11, -27, -12, -18, -27,
    -- filter=27 channel=15
    17, 11, 4, -14, 0, -12, 6, -29, -28,
    -- filter=28 channel=0
    -21, 15, 9, -8, -5, -14, 4, 11, 0,
    -- filter=28 channel=1
    16, 8, 0, 2, 7, -10, 12, -21, -15,
    -- filter=28 channel=2
    13, 32, 55, 13, 0, 37, -40, -4, 43,
    -- filter=28 channel=3
    16, -8, 16, -14, 13, -6, -6, 12, -6,
    -- filter=28 channel=4
    34, 29, 37, 54, 18, 28, 74, 40, 8,
    -- filter=28 channel=5
    -1, 28, 15, 17, 30, 16, -11, 3, 6,
    -- filter=28 channel=6
    -7, -13, -11, 17, -20, -8, 8, 1, 10,
    -- filter=28 channel=7
    0, -18, -4, 21, -10, -7, 11, 14, 10,
    -- filter=28 channel=8
    -33, -20, 13, -14, -40, -8, 5, -15, -37,
    -- filter=28 channel=9
    15, -22, 18, -4, -3, -16, 28, 13, 13,
    -- filter=28 channel=10
    0, 26, 24, -8, 2, 30, 21, -13, -5,
    -- filter=28 channel=11
    -18, -33, -24, -39, -49, -49, -26, -36, -45,
    -- filter=28 channel=12
    -14, -5, 28, -53, -20, 8, -25, -50, -13,
    -- filter=28 channel=13
    -16, 20, 41, -22, 3, 19, -32, 2, 32,
    -- filter=28 channel=14
    1, 34, 17, -10, -12, 39, -32, -31, -3,
    -- filter=28 channel=15
    35, 8, 12, 2, 17, 39, 7, 14, 23,
    -- filter=29 channel=0
    -12, -1, -2, -7, -7, -6, 0, 4, 13,
    -- filter=29 channel=1
    -20, -15, 15, -5, -4, 17, -3, -3, 15,
    -- filter=29 channel=2
    6, -2, 1, 0, -2, -19, -9, 0, -1,
    -- filter=29 channel=3
    -4, 1, 16, 15, -8, 5, -6, 7, 7,
    -- filter=29 channel=4
    -14, 0, 9, 9, -7, -2, -16, 16, 0,
    -- filter=29 channel=5
    -14, 10, 2, -6, 0, 19, -18, 5, -16,
    -- filter=29 channel=6
    -8, 18, 11, 18, 6, 18, -18, 3, -1,
    -- filter=29 channel=7
    -11, -18, 13, -5, -8, 13, 20, 9, -15,
    -- filter=29 channel=8
    0, -18, 0, -4, 13, 16, -8, 0, -9,
    -- filter=29 channel=9
    -11, 5, 15, -7, -3, -12, -8, -7, 8,
    -- filter=29 channel=10
    -19, -5, -5, 20, -7, -9, 19, -12, 5,
    -- filter=29 channel=11
    -15, -9, 8, 5, 12, -7, 20, -13, 12,
    -- filter=29 channel=12
    5, 0, -1, -8, 0, 9, -1, -2, -9,
    -- filter=29 channel=13
    -10, -6, 20, -5, -12, -19, -7, -18, -3,
    -- filter=29 channel=14
    -16, -5, -11, 8, -8, -20, -16, -8, -6,
    -- filter=29 channel=15
    4, -5, -7, -8, 17, 13, 18, -19, 3,
    -- filter=30 channel=0
    -18, 17, 8, -5, 16, -13, -16, -3, -20,
    -- filter=30 channel=1
    -3, -16, -3, -18, 0, -11, -21, 4, 8,
    -- filter=30 channel=2
    17, 4, 2, 1, 28, 15, -6, 9, -1,
    -- filter=30 channel=3
    -4, -7, -4, -4, 7, 19, 13, 18, -18,
    -- filter=30 channel=4
    7, 15, 36, 18, 20, 35, -7, -1, 30,
    -- filter=30 channel=5
    -6, 13, -16, 0, 24, 6, -16, -7, -14,
    -- filter=30 channel=6
    -17, -20, -13, 19, -2, 17, 19, 0, 5,
    -- filter=30 channel=7
    -19, -12, 5, -7, -7, -10, 10, -5, -6,
    -- filter=30 channel=8
    3, 4, -16, -14, -21, 0, -18, 2, -24,
    -- filter=30 channel=9
    3, 9, 7, -26, -17, -16, 11, -7, -13,
    -- filter=30 channel=10
    6, 10, -16, 18, -3, 9, -15, -13, 16,
    -- filter=30 channel=11
    -17, -11, -13, -14, -20, -22, -41, -34, -36,
    -- filter=30 channel=12
    9, -5, 29, 0, 27, 17, -10, -23, -1,
    -- filter=30 channel=13
    34, 14, 37, -10, 16, 12, -12, -13, -4,
    -- filter=30 channel=14
    7, 17, -3, -13, 1, 23, 9, 21, 5,
    -- filter=30 channel=15
    12, 33, 20, 27, 18, 35, 19, 16, 31,
    -- filter=31 channel=0
    12, 2, -9, 0, 16, -17, -13, -19, 10,
    -- filter=31 channel=1
    8, -4, -15, -20, 20, 8, 10, -13, -10,
    -- filter=31 channel=2
    4, -1, -6, -1, -13, -14, 12, 3, 11,
    -- filter=31 channel=3
    -5, 13, -2, 16, -5, 17, 10, -1, -21,
    -- filter=31 channel=4
    18, -6, 19, 18, -14, 20, -2, 13, 5,
    -- filter=31 channel=5
    -1, -9, -6, 1, 15, -15, 20, 20, -2,
    -- filter=31 channel=6
    -2, 6, 5, 9, 8, 1, -2, 3, -18,
    -- filter=31 channel=7
    -8, 9, 1, -16, 10, -14, -16, 15, 12,
    -- filter=31 channel=8
    16, -18, 10, -14, -9, -12, 4, -14, 11,
    -- filter=31 channel=9
    -17, 20, 2, 2, -15, 15, 3, 12, 6,
    -- filter=31 channel=10
    -14, 3, 7, 18, 18, 8, 8, 0, -18,
    -- filter=31 channel=11
    -1, -1, 4, 2, 1, 17, 9, 7, -12,
    -- filter=31 channel=12
    8, -12, 5, 0, -12, -12, 4, -11, -18,
    -- filter=31 channel=13
    14, -16, 7, -5, -2, 3, -16, -19, 16,
    -- filter=31 channel=14
    -15, 6, -7, -20, -5, 5, 19, -14, 4,
    -- filter=31 channel=15
    -2, -7, -9, -12, 1, -17, 15, -15, 5,

    others => 0);
end iwght_package;
