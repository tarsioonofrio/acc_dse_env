LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias
					-- layer=2
					2953, -1047, -839, -6929, -1616, 14488, -3568, -855, -2211, 4138, -824, -1779, 15116, 375, 2552, 1444, -6669, -3510, -1104, -1222, 3411, -2554, 364, 2180, 10655, 6091, 11296, 9406, -748, 12319, 15754, -219, -735, -403, -2710, -4734, -947, -1357, 3249, 889, 10558, 669, -878, 9416, 3357, -5295, -1163, -549, -3667, 5391, -2917, 12526, 5142, -693, -1758, -879, -4568, -806, -568, 1103, -522, 13102, -503, 9675, -2939, -677, 3290, 5241, -4315, -1779, 6977, -9406, -846, -651, -2471, -2822, -1126, 3920, -813, -554, -8572, 6953, -1016, -7336, -1648, 2967, -1122, -2408, -1618, 4417, 4791, -1335, -2777, -1749, 2474, 4433, -2031, -1991, 3803, -1615, -647, 3682, -2621, -4703, -2741, -4490, -1246, -880, 8790, -4554, 4340, -1196, 2777, -424, -3421, 2498, -7792, 4011, -5285, 8226, 860, 13158, -2211, -839, -858, -4281, 5009, 7277, -740, 14634, 10075, 2826, -1352, -1114, 1683, -751, 7673, 11180, -2190, -472, 288, -4708, 3271, 3981, -570, 1412, 8983, 2762, 2854, -1804, 1525, -480, -2627, 5817, -349, -573, 6814, -746, 891, -1710, 13578, 11082, -486, 4235, -2315, -1722, -1654, -2271, -2331, -6803, -1628, -2813, 12652, -564, -1697, -319, -2396, -1134, -2572, -1989, -999, -4849, -2820, -3308, 1032, -1163, -483, -3760, 1050, 15390, -989, -4873, 1548, 13155, 11152, -8700, -599, -4367, 2169, -1150, -6324, -2437, -1849, -1223, -1603, 256, 7583, -2216, 9480, -1198, -3253, 3316, 4067, -8431, 2210, -1573, 5829, 7101, 10221, -605, 4106, -3290, -3061, -4057, -2326, -855, 12351, -3236, -986, 5092, -700, -558, 3856, -9954, 2212, 4845, 7765, -5791, 822, 1345, 13187, -762, -3594, -1011, 7416, -5802, 10027, 1227, -4332, 7272, -2767, -518, 5589, 2467, -4864, -1145,

					-- weights
					-- layer=2 filter=0 channel=0
					-33, -8, -18, 7, -2, 11, 7, -21, -44,
					-- layer=2 filter=0 channel=1
					-31, -13, -10, 4, 4, -2, -16, 27, 14,
					-- layer=2 filter=0 channel=2
					-2, 3, 0, 3, 4, 6, -1, -6, 9,
					-- layer=2 filter=0 channel=3
					-41, -17, -13, 37, -8, 0, -4, 19, 23,
					-- layer=2 filter=0 channel=4
					-24, 15, 18, 11, -4, 33, -9, 1, 2,
					-- layer=2 filter=0 channel=5
					22, 17, 4, 19, 3, 25, -29, -28, 0,
					-- layer=2 filter=0 channel=6
					8, 8, -2, -34, -21, 20, -9, 30, 37,
					-- layer=2 filter=0 channel=7
					-5, 40, 34, 2, 32, 30, 40, 9, 0,
					-- layer=2 filter=0 channel=8
					5, 0, -4, 4, -9, -4, -4, 2, 1,
					-- layer=2 filter=0 channel=9
					-59, -39, -27, -64, -26, -82, 16, 0, -7,
					-- layer=2 filter=0 channel=10
					-60, -48, -3, -6, -10, -9, 31, 18, -10,
					-- layer=2 filter=0 channel=11
					24, 13, 15, -14, 9, -16, -21, -26, -53,
					-- layer=2 filter=0 channel=12
					-8, -6, -1, 20, 25, 3, 0, 28, 6,
					-- layer=2 filter=0 channel=13
					4, 5, 0, -4, 10, -5, 12, -7, 6,
					-- layer=2 filter=0 channel=14
					-24, -9, 8, -7, 16, -5, -5, 23, -13,
					-- layer=2 filter=0 channel=15
					-36, -38, -29, -47, -30, 7, -50, 30, 51,
					-- layer=2 filter=0 channel=16
					-16, 23, -7, -16, 23, -6, -15, 0, -30,
					-- layer=2 filter=0 channel=17
					-8, 10, 10, -8, -8, 0, 3, -7, -6,
					-- layer=2 filter=0 channel=18
					-3, -6, -28, 23, 4, -32, -48, 0, -12,
					-- layer=2 filter=0 channel=19
					39, -3, -33, 1, 5, 13, 2, 32, 40,
					-- layer=2 filter=0 channel=20
					-2, -9, 8, 0, -5, 0, 10, 4, 5,
					-- layer=2 filter=0 channel=21
					3, 0, -5, -10, 2, -3, 1, -4, 10,
					-- layer=2 filter=0 channel=22
					-3, 3, -4, -1, 2, -7, -7, 3, -1,
					-- layer=2 filter=0 channel=23
					27, 19, -11, -18, -1, 9, 7, 13, -5,
					-- layer=2 filter=0 channel=24
					-35, -25, 1, 10, -6, 3, 4, -20, -47,
					-- layer=2 filter=0 channel=25
					-6, 14, 38, 17, -2, 19, -4, -40, -50,
					-- layer=2 filter=0 channel=26
					-1, 9, 5, -3, 8, 1, -9, -1, 2,
					-- layer=2 filter=0 channel=27
					-1, 11, 15, 6, 6, 7, -48, -20, -22,
					-- layer=2 filter=0 channel=28
					14, 24, -25, 5, 34, -1, 25, 20, -19,
					-- layer=2 filter=0 channel=29
					0, 0, 10, 1, 0, -2, 5, -8, 1,
					-- layer=2 filter=0 channel=30
					-42, -35, -17, -47, -35, -35, 4, -12, 26,
					-- layer=2 filter=0 channel=31
					-28, -51, -3, 8, 95, -20, -17, -24, -20,
					-- layer=2 filter=0 channel=32
					-6, 4, 7, 12, 9, -3, 2, -4, 3,
					-- layer=2 filter=0 channel=33
					-18, 36, -36, 0, 29, 26, -29, 13, -14,
					-- layer=2 filter=0 channel=34
					29, 9, -10, -37, -27, -45, -101, 3, 17,
					-- layer=2 filter=0 channel=35
					-1, 26, -6, -15, 15, 23, -33, -13, -13,
					-- layer=2 filter=0 channel=36
					-4, -1, 5, 0, -13, 3, -4, 0, -4,
					-- layer=2 filter=0 channel=37
					15, 41, 32, 3, -3, 12, -50, -8, -9,
					-- layer=2 filter=0 channel=38
					0, -5, 15, -20, -19, 20, -38, -5, -10,
					-- layer=2 filter=0 channel=39
					-15, -13, -18, -19, 5, 16, 8, 20, 28,
					-- layer=2 filter=0 channel=40
					-7, 14, -21, -15, -17, -6, -67, 14, -17,
					-- layer=2 filter=0 channel=41
					11, 0, -3, 6, -5, -5, -5, -5, 2,
					-- layer=2 filter=0 channel=42
					0, 8, 13, -4, -12, 0, 21, 28, 27,
					-- layer=2 filter=0 channel=43
					-21, -10, -85, 31, -13, 4, 0, -29, 67,
					-- layer=2 filter=0 channel=44
					3, -5, -6, -5, 2, -14, 5, 5, -8,
					-- layer=2 filter=0 channel=45
					12, 51, 19, 33, 55, 52, 0, -35, -21,
					-- layer=2 filter=0 channel=46
					-66, -42, -18, -52, -15, 29, -33, -23, 24,
					-- layer=2 filter=0 channel=47
					-8, 10, -11, -4, 0, -8, 23, -6, -38,
					-- layer=2 filter=0 channel=48
					-8, -5, 6, 9, -5, 2, -2, -9, -2,
					-- layer=2 filter=0 channel=49
					-22, -29, -45, 7, -5, -64, 28, 33, -15,
					-- layer=2 filter=0 channel=50
					5, -1, -9, -9, -11, 4, 23, 8, 31,
					-- layer=2 filter=0 channel=51
					-12, 0, 20, -14, -21, 1, 1, -7, -11,
					-- layer=2 filter=0 channel=52
					-2, 14, 3, -20, -28, -3, -29, 0, 44,
					-- layer=2 filter=0 channel=53
					-80, -57, -39, -9, -93, -45, 9, 5, 32,
					-- layer=2 filter=0 channel=54
					21, -5, -6, 21, 0, 14, 23, 9, 3,
					-- layer=2 filter=0 channel=55
					13, 14, 1, 4, 0, -8, -8, -14, -2,
					-- layer=2 filter=0 channel=56
					14, 21, 11, -15, 5, 1, -25, -31, -35,
					-- layer=2 filter=0 channel=57
					13, 5, -8, 6, -7, -10, 12, -5, 6,
					-- layer=2 filter=0 channel=58
					-7, 19, 40, 29, 32, 35, 6, 23, 19,
					-- layer=2 filter=0 channel=59
					15, 13, -4, 31, 47, 29, -16, 21, 38,
					-- layer=2 filter=0 channel=60
					21, -9, -2, 25, -17, 34, 7, 61, -11,
					-- layer=2 filter=0 channel=61
					-22, -35, -50, -23, -64, -15, 34, -7, -33,
					-- layer=2 filter=0 channel=62
					16, 23, 10, -11, -27, -25, -28, 48, 25,
					-- layer=2 filter=0 channel=63
					10, -9, -45, 0, -19, -8, 26, 2, -1,
					-- layer=2 filter=0 channel=64
					-20, -9, -5, -13, -21, 14, 12, 19, 9,
					-- layer=2 filter=0 channel=65
					-5, -8, -11, -24, -32, -27, -17, -13, 12,
					-- layer=2 filter=0 channel=66
					-18, 32, -8, 54, -47, 1, 49, 8, -25,
					-- layer=2 filter=0 channel=67
					-41, -36, -38, -74, -42, -8, -22, -34, 14,
					-- layer=2 filter=0 channel=68
					10, 8, 7, 8, -3, -6, -6, 10, -1,
					-- layer=2 filter=0 channel=69
					-34, -23, 8, -7, 5, 19, 13, 23, 4,
					-- layer=2 filter=0 channel=70
					31, 31, -27, 6, 27, 24, -24, -42, -22,
					-- layer=2 filter=0 channel=71
					18, 16, 10, 7, 15, 25, -6, -27, 2,
					-- layer=2 filter=0 channel=72
					16, 33, 21, 8, 42, 32, 37, 51, 14,
					-- layer=2 filter=0 channel=73
					-81, -62, -68, 49, -11, -9, 37, -20, 6,
					-- layer=2 filter=0 channel=74
					-53, -37, -27, -47, 15, 0, -24, 8, -14,
					-- layer=2 filter=0 channel=75
					34, 28, -6, 10, 59, -1, -9, 3, -5,
					-- layer=2 filter=0 channel=76
					-61, -48, -53, -62, -71, -34, -27, 12, -16,
					-- layer=2 filter=0 channel=77
					0, -7, -10, -3, 2, -2, -6, 7, -8,
					-- layer=2 filter=0 channel=78
					-7, 6, -7, -1, -31, -24, -32, -16, -12,
					-- layer=2 filter=0 channel=79
					-6, 6, 7, 3, -4, -5, 8, 9, 6,
					-- layer=2 filter=0 channel=80
					-25, -36, -15, -8, -13, -14, -13, -9, 20,
					-- layer=2 filter=0 channel=81
					8, 16, 0, 13, 11, 7, 17, 5, 10,
					-- layer=2 filter=0 channel=82
					11, 4, -6, 4, 1, 11, 6, 1, -7,
					-- layer=2 filter=0 channel=83
					-14, 5, -20, -8, 17, 0, 3, 23, 20,
					-- layer=2 filter=0 channel=84
					-1, -9, -8, 0, 1, 3, -7, 3, 0,
					-- layer=2 filter=0 channel=85
					10, -2, -3, 0, 0, 11, 6, -2, -8,
					-- layer=2 filter=0 channel=86
					-3, -4, -4, -11, 18, -3, 4, 4, -1,
					-- layer=2 filter=0 channel=87
					20, -23, 11, -14, -68, 16, -37, -8, 22,
					-- layer=2 filter=0 channel=88
					-31, -16, -19, -20, -10, -1, 0, 12, 19,
					-- layer=2 filter=0 channel=89
					-21, -18, 24, 6, 32, 5, 0, 20, 0,
					-- layer=2 filter=0 channel=90
					-7, 0, -9, -5, -9, 2, -4, -2, -3,
					-- layer=2 filter=0 channel=91
					-4, 0, 39, 15, 56, 22, 3, 54, 17,
					-- layer=2 filter=0 channel=92
					-16, 8, 17, 10, 27, 2, 8, 43, 8,
					-- layer=2 filter=0 channel=93
					-18, 55, -10, 12, 0, 32, -18, 30, 77,
					-- layer=2 filter=0 channel=94
					1, -33, -83, -34, -81, -66, 27, 20, 17,
					-- layer=2 filter=0 channel=95
					12, 11, 8, -13, -1, 14, -6, 14, 9,
					-- layer=2 filter=0 channel=96
					26, 51, -4, 7, -21, 6, 4, 49, 73,
					-- layer=2 filter=0 channel=97
					-6, -11, 4, 9, -12, -22, -9, 6, 2,
					-- layer=2 filter=0 channel=98
					14, 19, -14, -24, 27, 9, 5, -23, -52,
					-- layer=2 filter=0 channel=99
					20, -42, -19, -9, -40, 1, -3, 48, 17,
					-- layer=2 filter=0 channel=100
					11, -16, 5, 8, 9, 29, -27, 17, 27,
					-- layer=2 filter=0 channel=101
					27, 51, 30, -11, 0, 15, -4, -26, -56,
					-- layer=2 filter=0 channel=102
					-8, -16, -33, -1, -29, 1, -12, 37, 40,
					-- layer=2 filter=0 channel=103
					2, -6, 15, -30, 32, 8, 11, 16, -45,
					-- layer=2 filter=0 channel=104
					-15, -14, -1, -59, -64, -36, 5, 26, -14,
					-- layer=2 filter=0 channel=105
					-1, 37, -22, 22, -30, -15, -24, 37, -74,
					-- layer=2 filter=0 channel=106
					-35, 0, 23, 9, 29, 27, 4, 13, -39,
					-- layer=2 filter=0 channel=107
					-16, -8, 29, 3, 16, -22, 24, -43, 0,
					-- layer=2 filter=0 channel=108
					1, -13, 6, 11, 12, 5, 5, 0, 15,
					-- layer=2 filter=0 channel=109
					2, -3, 10, -2, -3, 14, 4, -6, 0,
					-- layer=2 filter=0 channel=110
					8, 16, 2, -16, 36, 5, 31, 14, -14,
					-- layer=2 filter=0 channel=111
					7, -1, 0, -1, 0, -3, -4, 7, -5,
					-- layer=2 filter=0 channel=112
					-31, -6, 5, -80, -56, -16, 16, -29, -84,
					-- layer=2 filter=0 channel=113
					-13, -6, -1, -33, -22, -39, 18, -15, -6,
					-- layer=2 filter=0 channel=114
					-5, 0, -4, -7, -11, -11, -13, 0, -13,
					-- layer=2 filter=0 channel=115
					0, -5, 5, 7, -2, -3, -12, 3, -6,
					-- layer=2 filter=0 channel=116
					9, -13, 28, -16, -22, 31, -42, 51, 25,
					-- layer=2 filter=0 channel=117
					-45, -40, -19, -48, 0, -17, 44, 28, -7,
					-- layer=2 filter=0 channel=118
					12, 38, 25, 23, -26, -29, -26, -6, 13,
					-- layer=2 filter=0 channel=119
					1, 15, 39, 16, 33, 30, -17, 20, -22,
					-- layer=2 filter=0 channel=120
					5, -6, 9, 8, 5, 10, 4, 6, 5,
					-- layer=2 filter=0 channel=121
					0, 1, -2, -4, 6, 4, -6, -1, 5,
					-- layer=2 filter=0 channel=122
					-9, -16, 8, -3, -10, 5, -10, 0, 3,
					-- layer=2 filter=0 channel=123
					11, 29, -14, -7, 22, 2, 4, 13, 21,
					-- layer=2 filter=0 channel=124
					-38, 14, -36, -1, -14, 13, 8, 19, 5,
					-- layer=2 filter=0 channel=125
					-10, -4, 7, 5, -4, -1, -9, 11, 10,
					-- layer=2 filter=0 channel=126
					-20, 11, -17, -9, -12, 18, -13, 57, 48,
					-- layer=2 filter=0 channel=127
					-15, 2, 5, 4, -18, -23, 20, 14, 16,
					-- layer=2 filter=1 channel=0
					0, 27, 3, 0, 32, 1, 52, 22, 28,
					-- layer=2 filter=1 channel=1
					4, 5, -21, 10, -4, -53, -2, -36, 5,
					-- layer=2 filter=1 channel=2
					9, 2, -4, -1, -2, 6, -4, 0, 8,
					-- layer=2 filter=1 channel=3
					1, -7, -4, 47, 24, -11, 38, 44, 22,
					-- layer=2 filter=1 channel=4
					-9, -76, -28, -35, 0, 14, 7, -9, -14,
					-- layer=2 filter=1 channel=5
					-12, 33, 5, -9, -18, 12, -3, -18, -4,
					-- layer=2 filter=1 channel=6
					-17, -25, 19, -9, 50, 23, -16, 31, -16,
					-- layer=2 filter=1 channel=7
					-13, -16, 5, 17, 8, 8, 24, 2, 8,
					-- layer=2 filter=1 channel=8
					2, -2, -3, -5, 2, -10, 8, -10, 4,
					-- layer=2 filter=1 channel=9
					-3, -12, -12, -16, 19, 4, 29, -7, 12,
					-- layer=2 filter=1 channel=10
					1, 24, -1, 21, 48, 15, 41, 46, 48,
					-- layer=2 filter=1 channel=11
					-2, -16, 28, 4, -22, 0, 5, -17, -9,
					-- layer=2 filter=1 channel=12
					11, 0, -8, 5, -38, -62, 9, -59, -9,
					-- layer=2 filter=1 channel=13
					11, -8, -8, 3, 5, 0, 11, -8, 3,
					-- layer=2 filter=1 channel=14
					17, 6, 15, 1, -15, -41, 9, -49, -16,
					-- layer=2 filter=1 channel=15
					35, -27, 18, -26, 2, 21, 12, -16, 2,
					-- layer=2 filter=1 channel=16
					42, -22, 14, -27, -31, 26, -7, 36, 51,
					-- layer=2 filter=1 channel=17
					-11, -6, 5, -8, 9, -3, 10, 2, -5,
					-- layer=2 filter=1 channel=18
					31, -64, -23, 3, -13, 22, 6, -10, -5,
					-- layer=2 filter=1 channel=19
					27, 41, 6, 29, 36, 18, -4, 37, 2,
					-- layer=2 filter=1 channel=20
					-1, 1, 4, 3, -8, 7, -8, 8, 10,
					-- layer=2 filter=1 channel=21
					20, 20, 0, 16, 7, 16, 12, 5, 8,
					-- layer=2 filter=1 channel=22
					-9, 1, -4, -9, -1, 8, -3, 0, -3,
					-- layer=2 filter=1 channel=23
					-16, -19, -2, -49, 16, -24, 14, 48, -5,
					-- layer=2 filter=1 channel=24
					22, 8, 23, 9, -4, -6, 6, 11, 9,
					-- layer=2 filter=1 channel=25
					11, 29, 11, 2, -17, -47, 7, -9, -24,
					-- layer=2 filter=1 channel=26
					-7, -3, -9, -1, 4, 8, 5, -3, 6,
					-- layer=2 filter=1 channel=27
					-23, -12, 26, -17, -10, -8, -4, -45, -15,
					-- layer=2 filter=1 channel=28
					17, -36, -51, -26, -58, -30, -8, 22, 29,
					-- layer=2 filter=1 channel=29
					-7, 7, 9, 0, -9, -3, -7, -10, 8,
					-- layer=2 filter=1 channel=30
					-33, 22, -53, -21, -70, -6, -1, -9, -13,
					-- layer=2 filter=1 channel=31
					44, -20, -53, -43, -20, -5, -20, 3, -29,
					-- layer=2 filter=1 channel=32
					0, 0, 10, -2, 9, -7, 6, 1, -4,
					-- layer=2 filter=1 channel=33
					13, 32, 15, 26, 41, 13, -10, -22, 2,
					-- layer=2 filter=1 channel=34
					21, 48, 0, 8, -11, 23, -33, 19, 28,
					-- layer=2 filter=1 channel=35
					-1, -42, 1, 0, -18, 28, -9, 9, 20,
					-- layer=2 filter=1 channel=36
					-12, -4, -6, 8, 3, -13, -9, 0, -2,
					-- layer=2 filter=1 channel=37
					-11, -15, -10, 5, -5, 7, -3, -18, -30,
					-- layer=2 filter=1 channel=38
					-35, 26, -18, 9, 10, 17, -11, -24, 11,
					-- layer=2 filter=1 channel=39
					2, -3, 3, 28, 29, 24, 36, 8, 29,
					-- layer=2 filter=1 channel=40
					44, -26, -5, -20, 30, -3, -36, -1, -31,
					-- layer=2 filter=1 channel=41
					-7, 0, -5, -8, 5, -8, -7, 6, -3,
					-- layer=2 filter=1 channel=42
					11, -21, 32, -34, 26, 38, 24, 16, 13,
					-- layer=2 filter=1 channel=43
					4, -23, -10, 9, -2, 0, 32, 15, 13,
					-- layer=2 filter=1 channel=44
					7, -8, 1, 3, 0, -5, 9, -8, 5,
					-- layer=2 filter=1 channel=45
					-50, -24, -28, -38, -50, -8, -12, -70, -14,
					-- layer=2 filter=1 channel=46
					-24, 33, -47, 7, -8, 19, 42, 41, -3,
					-- layer=2 filter=1 channel=47
					18, 7, -10, 8, -33, -33, 7, 18, 24,
					-- layer=2 filter=1 channel=48
					-7, -1, 2, 11, 1, 5, 4, -1, 0,
					-- layer=2 filter=1 channel=49
					17, -61, -24, -44, 16, -17, 5, -25, 20,
					-- layer=2 filter=1 channel=50
					7, 0, -17, 15, -16, 6, 0, -4, 1,
					-- layer=2 filter=1 channel=51
					-16, -4, -5, -11, -2, -2, 13, 6, -12,
					-- layer=2 filter=1 channel=52
					9, -82, -22, 5, -17, 23, -12, -32, 6,
					-- layer=2 filter=1 channel=53
					-10, -90, -15, -20, 12, 32, -10, 38, 48,
					-- layer=2 filter=1 channel=54
					6, -20, -38, -22, 7, -9, 3, 19, 15,
					-- layer=2 filter=1 channel=55
					0, -5, 14, -11, 9, -5, -2, 0, 4,
					-- layer=2 filter=1 channel=56
					11, -16, 46, 0, -29, 7, -1, -13, -10,
					-- layer=2 filter=1 channel=57
					2, 8, -6, -7, -6, -7, -7, -1, 5,
					-- layer=2 filter=1 channel=58
					8, -3, -4, -23, -37, -23, -10, -55, -16,
					-- layer=2 filter=1 channel=59
					-14, 34, 17, -10, 54, -5, -33, -24, -2,
					-- layer=2 filter=1 channel=60
					3, 49, -23, 38, 28, 13, 37, 5, -31,
					-- layer=2 filter=1 channel=61
					-27, -9, -20, -5, 45, -51, 23, 13, 15,
					-- layer=2 filter=1 channel=62
					19, -41, -6, -24, -13, 20, -7, 5, 15,
					-- layer=2 filter=1 channel=63
					-24, -8, -32, -14, -23, -48, 33, 3, 26,
					-- layer=2 filter=1 channel=64
					2, 0, -17, -9, -17, -2, -20, 18, -3,
					-- layer=2 filter=1 channel=65
					-49, 19, -42, 13, 26, 16, -8, -3, -16,
					-- layer=2 filter=1 channel=66
					-26, -12, -1, -43, -11, -5, 27, -7, 7,
					-- layer=2 filter=1 channel=67
					-61, 36, 18, 16, 2, 14, 34, 6, 20,
					-- layer=2 filter=1 channel=68
					-9, 5, 1, -1, 8, 5, -5, 8, -8,
					-- layer=2 filter=1 channel=69
					17, -10, 9, -16, 0, -22, 13, 16, 37,
					-- layer=2 filter=1 channel=70
					-17, -31, -46, -9, -4, 19, -10, 20, 22,
					-- layer=2 filter=1 channel=71
					-50, -12, 52, -52, -11, -1, 18, -26, -15,
					-- layer=2 filter=1 channel=72
					23, 61, -1, 26, 42, 12, -23, -18, -50,
					-- layer=2 filter=1 channel=73
					-1, 7, 66, -57, 23, 38, 16, 5, 0,
					-- layer=2 filter=1 channel=74
					-16, 36, -7, 16, 18, -22, -4, 18, 28,
					-- layer=2 filter=1 channel=75
					24, 6, -9, 21, -39, -72, 29, 30, 21,
					-- layer=2 filter=1 channel=76
					-1, -20, -26, -26, 54, 27, 29, 41, 13,
					-- layer=2 filter=1 channel=77
					-10, -5, -11, -2, -4, 6, 0, -1, 0,
					-- layer=2 filter=1 channel=78
					7, -33, 23, -10, -31, 8, -16, -9, 1,
					-- layer=2 filter=1 channel=79
					10, 9, -1, 10, 2, -8, -8, 11, 9,
					-- layer=2 filter=1 channel=80
					-10, -34, -20, 9, 0, 38, -12, 14, 37,
					-- layer=2 filter=1 channel=81
					-3, 0, -7, -4, -4, 8, -4, -8, 6,
					-- layer=2 filter=1 channel=82
					-2, 3, -3, 3, 2, -10, -2, 6, 11,
					-- layer=2 filter=1 channel=83
					18, -42, -29, -34, -58, -42, -56, -2, -7,
					-- layer=2 filter=1 channel=84
					-10, 0, -3, 1, 5, -1, 8, 3, 5,
					-- layer=2 filter=1 channel=85
					-13, -10, -11, -3, -4, -8, 6, -5, 1,
					-- layer=2 filter=1 channel=86
					6, 9, 1, 1, -11, 4, -2, -3, -9,
					-- layer=2 filter=1 channel=87
					21, -46, 12, -29, 45, 35, -30, 38, -5,
					-- layer=2 filter=1 channel=88
					-3, 34, -46, -40, -40, -33, -25, 14, -16,
					-- layer=2 filter=1 channel=89
					7, 22, 20, 2, 35, -25, -26, -62, 11,
					-- layer=2 filter=1 channel=90
					-3, 7, 7, -7, -5, 0, -5, 2, 9,
					-- layer=2 filter=1 channel=91
					28, 22, 3, 14, 14, -19, -2, -21, -38,
					-- layer=2 filter=1 channel=92
					1, 0, -25, 22, 17, -44, 2, -68, -14,
					-- layer=2 filter=1 channel=93
					30, 51, -11, 43, -26, 67, -30, 15, 10,
					-- layer=2 filter=1 channel=94
					-50, -35, 16, -50, 39, -53, 6, 30, 0,
					-- layer=2 filter=1 channel=95
					6, 4, -10, -14, 3, 0, -11, 4, 5,
					-- layer=2 filter=1 channel=96
					-16, 9, 10, -57, 36, 37, -12, 25, 0,
					-- layer=2 filter=1 channel=97
					37, 10, 7, 30, 11, -25, 8, 23, 43,
					-- layer=2 filter=1 channel=98
					-2, -73, -11, 17, -15, 0, 6, 6, 2,
					-- layer=2 filter=1 channel=99
					-7, -39, -21, -18, 18, 39, -19, 5, -41,
					-- layer=2 filter=1 channel=100
					-20, 43, -11, -10, 4, 29, -8, -25, 30,
					-- layer=2 filter=1 channel=101
					5, 8, 27, -19, -30, -6, 48, -7, -21,
					-- layer=2 filter=1 channel=102
					1, -27, -12, 12, 3, 40, 14, -15, 2,
					-- layer=2 filter=1 channel=103
					51, 14, -29, 18, 44, 82, 22, -33, 53,
					-- layer=2 filter=1 channel=104
					5, -85, 14, -39, 8, -1, -21, -2, -2,
					-- layer=2 filter=1 channel=105
					-18, 1, 15, -24, -22, -11, 12, 13, 53,
					-- layer=2 filter=1 channel=106
					24, 56, 4, 11, -16, -35, 31, 17, -1,
					-- layer=2 filter=1 channel=107
					-32, -16, 46, -26, 23, 25, 52, 2, 26,
					-- layer=2 filter=1 channel=108
					-10, -8, 12, -41, -12, -32, -18, -31, -26,
					-- layer=2 filter=1 channel=109
					1, 18, 8, -12, 21, 6, -6, 8, -11,
					-- layer=2 filter=1 channel=110
					25, 38, 26, 6, 40, 39, -9, 2, 22,
					-- layer=2 filter=1 channel=111
					0, 4, -2, -2, -5, 7, -7, 10, -5,
					-- layer=2 filter=1 channel=112
					-41, 10, 10, -3, -4, -11, 40, 5, -5,
					-- layer=2 filter=1 channel=113
					-54, -12, -60, -9, -65, -67, -18, -28, -8,
					-- layer=2 filter=1 channel=114
					-9, -4, -14, -3, -14, -17, -10, -18, -21,
					-- layer=2 filter=1 channel=115
					3, 8, -4, 4, -3, -7, -4, 4, -5,
					-- layer=2 filter=1 channel=116
					38, 14, 26, 22, 46, 45, -42, 15, -17,
					-- layer=2 filter=1 channel=117
					0, 5, 20, 23, 0, -14, -5, 16, 20,
					-- layer=2 filter=1 channel=118
					-14, -57, -1, -13, 9, 39, -29, 30, 4,
					-- layer=2 filter=1 channel=119
					58, -55, -61, -23, -36, -6, -16, -20, 0,
					-- layer=2 filter=1 channel=120
					-9, 9, -4, 1, -6, 6, 5, 6, -5,
					-- layer=2 filter=1 channel=121
					-8, 6, 3, -6, 5, 0, 3, 0, 12,
					-- layer=2 filter=1 channel=122
					2, 2, -3, 4, -2, 15, -9, 1, 9,
					-- layer=2 filter=1 channel=123
					-1, 33, 12, 22, 18, 2, 6, 1, -15,
					-- layer=2 filter=1 channel=124
					22, 21, 9, -14, 7, 23, 15, 13, 0,
					-- layer=2 filter=1 channel=125
					3, -5, -8, -8, 5, 2, 7, 0, -7,
					-- layer=2 filter=1 channel=126
					16, 40, -11, 21, 24, -9, 55, -20, -8,
					-- layer=2 filter=1 channel=127
					14, 13, -34, -9, -29, -20, -2, -23, -14,
					-- layer=2 filter=2 channel=0
					-3, 0, 0, 8, -4, -7, 3, 7, 3,
					-- layer=2 filter=2 channel=1
					-1, -7, -9, 0, -2, -7, -3, -6, 6,
					-- layer=2 filter=2 channel=2
					-9, 0, 1, -5, -8, 6, -3, -7, -5,
					-- layer=2 filter=2 channel=3
					-6, -1, -10, 4, -12, 6, -3, 5, 7,
					-- layer=2 filter=2 channel=4
					-4, 2, -13, -8, -8, 3, -7, -8, -7,
					-- layer=2 filter=2 channel=5
					-7, -6, -9, 6, -8, 6, -12, -10, -2,
					-- layer=2 filter=2 channel=6
					-5, -8, -2, 3, 1, -11, -10, -4, 8,
					-- layer=2 filter=2 channel=7
					3, 1, 6, -5, 3, -8, -11, -12, -15,
					-- layer=2 filter=2 channel=8
					9, 3, 3, 6, -3, 9, 1, -2, 7,
					-- layer=2 filter=2 channel=9
					1, 3, -4, 3, -10, -7, -4, 0, -11,
					-- layer=2 filter=2 channel=10
					-9, -5, -3, 5, -7, -11, -7, -1, -3,
					-- layer=2 filter=2 channel=11
					-2, -11, 6, -9, 4, -12, -3, 7, 4,
					-- layer=2 filter=2 channel=12
					7, 5, 3, 7, -1, 1, -11, -15, -12,
					-- layer=2 filter=2 channel=13
					-5, -6, -3, 8, -2, 0, 1, 5, -7,
					-- layer=2 filter=2 channel=14
					-1, 3, -7, 0, -12, 0, 4, 5, 6,
					-- layer=2 filter=2 channel=15
					2, 3, -7, -4, 4, -10, -7, 5, -13,
					-- layer=2 filter=2 channel=16
					6, -13, -8, -9, -9, -10, 8, 3, 3,
					-- layer=2 filter=2 channel=17
					8, -7, 5, 4, 0, -6, 8, -2, 3,
					-- layer=2 filter=2 channel=18
					-4, -2, -14, -3, -1, -11, 6, -2, 0,
					-- layer=2 filter=2 channel=19
					7, 7, -1, 8, 1, -8, -3, 0, -9,
					-- layer=2 filter=2 channel=20
					-4, 0, 1, -10, 3, 4, 0, -2, -8,
					-- layer=2 filter=2 channel=21
					-4, 3, 6, -1, -1, 5, 3, 0, 10,
					-- layer=2 filter=2 channel=22
					-5, -4, 1, -3, -1, 5, -8, 4, -4,
					-- layer=2 filter=2 channel=23
					-9, -8, -8, 8, 7, 8, -5, 0, 6,
					-- layer=2 filter=2 channel=24
					1, -5, -6, 0, 6, -1, -3, 7, 3,
					-- layer=2 filter=2 channel=25
					6, 0, 1, -3, 4, -1, -1, -4, -3,
					-- layer=2 filter=2 channel=26
					-2, 0, 2, 5, -5, 7, 1, -5, -2,
					-- layer=2 filter=2 channel=27
					0, -6, 1, 4, -12, 5, 5, 0, 6,
					-- layer=2 filter=2 channel=28
					-5, -13, -5, -6, 2, -6, 8, -8, 0,
					-- layer=2 filter=2 channel=29
					6, -10, 1, 6, -5, 8, 0, -6, -9,
					-- layer=2 filter=2 channel=30
					1, 7, -11, 0, -1, -7, -10, -9, 0,
					-- layer=2 filter=2 channel=31
					-2, 1, -11, -2, -3, -9, 4, 1, 8,
					-- layer=2 filter=2 channel=32
					4, 2, 10, -6, -7, 3, 8, 0, 7,
					-- layer=2 filter=2 channel=33
					1, -8, -8, -8, 5, 2, -14, -2, 6,
					-- layer=2 filter=2 channel=34
					-7, 0, -6, 0, 6, 8, -7, -7, -5,
					-- layer=2 filter=2 channel=35
					1, -1, -8, -4, -13, -9, 3, 0, 6,
					-- layer=2 filter=2 channel=36
					-7, 10, -3, -8, -3, 4, 9, -10, 0,
					-- layer=2 filter=2 channel=37
					4, 2, -2, 7, -3, -7, 0, -11, -11,
					-- layer=2 filter=2 channel=38
					5, -1, 1, 6, 5, -13, -5, 1, -11,
					-- layer=2 filter=2 channel=39
					0, 0, -2, -7, -2, 5, -13, 0, -10,
					-- layer=2 filter=2 channel=40
					5, -6, 9, 6, -8, 3, -9, -2, 9,
					-- layer=2 filter=2 channel=41
					-9, 4, 0, 3, 2, 6, 9, -3, 8,
					-- layer=2 filter=2 channel=42
					0, 8, 10, -2, 7, 5, 2, -7, 4,
					-- layer=2 filter=2 channel=43
					4, 4, -14, -2, 1, 2, 1, -6, -3,
					-- layer=2 filter=2 channel=44
					-1, 10, 10, 8, 0, -8, 10, 9, -2,
					-- layer=2 filter=2 channel=45
					6, 3, 6, 4, 1, -2, 4, 4, -7,
					-- layer=2 filter=2 channel=46
					-11, -8, 0, -8, -4, -5, -4, -8, 0,
					-- layer=2 filter=2 channel=47
					-6, -15, -5, -5, -11, -3, -7, 2, 0,
					-- layer=2 filter=2 channel=48
					-1, -9, 2, -8, 2, -8, 0, -2, 5,
					-- layer=2 filter=2 channel=49
					-5, -3, -6, 4, -7, 10, -6, -2, -1,
					-- layer=2 filter=2 channel=50
					-2, -9, 4, 0, 7, -8, 8, -7, 9,
					-- layer=2 filter=2 channel=51
					6, 6, -6, 3, -12, -8, 3, 0, 6,
					-- layer=2 filter=2 channel=52
					0, -4, -4, -3, 7, -10, -3, -5, -5,
					-- layer=2 filter=2 channel=53
					-2, 2, 2, 6, 3, -9, 7, 2, -9,
					-- layer=2 filter=2 channel=54
					4, -11, 2, -6, -3, 0, -1, -9, 1,
					-- layer=2 filter=2 channel=55
					-4, 3, 3, -8, 8, -4, -6, 7, 3,
					-- layer=2 filter=2 channel=56
					-12, 3, 3, 3, 5, -2, 2, -2, -5,
					-- layer=2 filter=2 channel=57
					-4, 10, -7, -6, 7, 0, 1, 7, -11,
					-- layer=2 filter=2 channel=58
					3, -9, -9, 0, 7, 3, -13, -6, -1,
					-- layer=2 filter=2 channel=59
					-8, 2, 6, -10, 2, 4, 3, 4, -13,
					-- layer=2 filter=2 channel=60
					3, -8, 1, -3, 3, -6, -7, -9, -1,
					-- layer=2 filter=2 channel=61
					-8, -12, -9, -3, 3, -7, 6, -8, -7,
					-- layer=2 filter=2 channel=62
					-3, 3, -10, -3, 3, 3, 3, 4, -9,
					-- layer=2 filter=2 channel=63
					5, 9, 9, -4, 0, -8, -5, 7, -6,
					-- layer=2 filter=2 channel=64
					0, -5, 6, 6, 1, 0, 1, -2, -5,
					-- layer=2 filter=2 channel=65
					9, -8, -10, -8, -4, 2, -5, 4, -4,
					-- layer=2 filter=2 channel=66
					-6, -4, 8, 0, -4, 2, -6, 6, 5,
					-- layer=2 filter=2 channel=67
					-12, -10, -8, -4, -8, -9, -5, 0, -9,
					-- layer=2 filter=2 channel=68
					2, 6, 2, -11, 0, 4, -12, -6, 0,
					-- layer=2 filter=2 channel=69
					-9, -4, 5, 0, 8, 0, -10, -5, -3,
					-- layer=2 filter=2 channel=70
					2, 4, -14, 0, 1, -8, 8, 5, -9,
					-- layer=2 filter=2 channel=71
					-6, 2, 3, 7, -12, -13, 2, -11, 6,
					-- layer=2 filter=2 channel=72
					0, 6, -8, -6, -1, 1, -13, -6, -5,
					-- layer=2 filter=2 channel=73
					-5, -11, 7, 0, -7, 5, -8, -4, 4,
					-- layer=2 filter=2 channel=74
					4, 4, -8, -10, -9, 0, -3, 1, 7,
					-- layer=2 filter=2 channel=75
					-11, -1, 6, 4, 1, -6, -1, 2, 0,
					-- layer=2 filter=2 channel=76
					-3, -7, -3, -1, -11, -6, -8, 3, -12,
					-- layer=2 filter=2 channel=77
					6, -8, 7, 0, 3, -5, 1, -3, -3,
					-- layer=2 filter=2 channel=78
					-4, -12, -6, 5, -11, -7, -7, 3, -8,
					-- layer=2 filter=2 channel=79
					7, -4, -9, 4, -5, -4, 0, 3, 3,
					-- layer=2 filter=2 channel=80
					-5, -12, 7, -6, 2, -1, -1, -8, -5,
					-- layer=2 filter=2 channel=81
					-10, -2, -9, -11, 7, 7, -7, 8, 3,
					-- layer=2 filter=2 channel=82
					0, 4, -8, 6, 10, 1, -9, -2, 0,
					-- layer=2 filter=2 channel=83
					-10, 6, 5, -2, -5, 5, -6, -9, -4,
					-- layer=2 filter=2 channel=84
					7, -7, 5, -1, 2, -7, 5, 2, -5,
					-- layer=2 filter=2 channel=85
					6, 0, 0, 3, 0, 8, -3, 8, 0,
					-- layer=2 filter=2 channel=86
					8, 3, -5, -2, -1, 4, 6, 0, 3,
					-- layer=2 filter=2 channel=87
					-4, -7, -3, 7, -7, -11, -10, 8, -10,
					-- layer=2 filter=2 channel=88
					7, 0, 5, 0, 3, 2, -8, -7, 5,
					-- layer=2 filter=2 channel=89
					2, 8, -7, 1, -8, -2, -14, -5, -6,
					-- layer=2 filter=2 channel=90
					0, -4, -4, 8, -10, -7, 1, -6, 9,
					-- layer=2 filter=2 channel=91
					-1, 1, 2, -4, -6, -2, 5, -5, -2,
					-- layer=2 filter=2 channel=92
					3, -2, -3, -1, 3, 5, -15, 0, 5,
					-- layer=2 filter=2 channel=93
					6, -8, 4, -1, -2, 6, -4, -12, 3,
					-- layer=2 filter=2 channel=94
					2, -7, -2, -4, 0, 0, 8, 7, -3,
					-- layer=2 filter=2 channel=95
					8, -1, -6, -8, 3, -6, 0, -1, -6,
					-- layer=2 filter=2 channel=96
					8, -9, -2, 3, 3, -4, 5, -10, -5,
					-- layer=2 filter=2 channel=97
					-12, 3, -11, -2, 0, -4, -4, -12, -9,
					-- layer=2 filter=2 channel=98
					4, 1, -17, -3, -12, -2, -11, -6, 4,
					-- layer=2 filter=2 channel=99
					-11, -10, -1, 8, 8, 1, 6, 5, -7,
					-- layer=2 filter=2 channel=100
					-4, -2, -3, -8, 3, 7, -7, 3, 4,
					-- layer=2 filter=2 channel=101
					-3, 4, -5, -12, -4, -1, -7, -5, -8,
					-- layer=2 filter=2 channel=102
					13, -4, 1, 10, -3, -2, -7, 0, 2,
					-- layer=2 filter=2 channel=103
					-11, 5, -1, 5, -8, 4, 8, 5, -9,
					-- layer=2 filter=2 channel=104
					-3, -10, -16, -9, 1, -4, 0, -6, -4,
					-- layer=2 filter=2 channel=105
					4, 0, -2, -9, 3, -7, -10, -4, 3,
					-- layer=2 filter=2 channel=106
					2, 6, 1, 1, 4, -3, -6, 0, 2,
					-- layer=2 filter=2 channel=107
					7, -10, -6, 5, 3, 1, 7, 3, 0,
					-- layer=2 filter=2 channel=108
					-11, 1, -11, -7, -2, -15, 4, -10, -12,
					-- layer=2 filter=2 channel=109
					7, 5, 2, 8, -11, 8, -10, -10, -10,
					-- layer=2 filter=2 channel=110
					-5, 0, -1, 8, -9, 0, -12, -9, -1,
					-- layer=2 filter=2 channel=111
					-5, -1, -7, 5, 1, -11, -1, 3, -5,
					-- layer=2 filter=2 channel=112
					4, -12, 2, 5, 6, 1, -2, -9, 0,
					-- layer=2 filter=2 channel=113
					-1, 10, 5, -8, -6, 2, -10, 1, -7,
					-- layer=2 filter=2 channel=114
					-1, -4, 1, -8, 8, 9, 0, 0, -1,
					-- layer=2 filter=2 channel=115
					-7, -7, 1, 10, 6, -9, 9, 6, 5,
					-- layer=2 filter=2 channel=116
					-10, -4, -5, -3, -11, -2, 5, 2, -11,
					-- layer=2 filter=2 channel=117
					-8, 2, -11, -8, 7, -7, -4, -11, -7,
					-- layer=2 filter=2 channel=118
					0, 0, -9, -6, -4, -5, -1, 2, -4,
					-- layer=2 filter=2 channel=119
					7, -2, 0, -12, -8, 3, 8, 1, -2,
					-- layer=2 filter=2 channel=120
					-3, 7, -1, -2, -6, 9, -2, 0, 5,
					-- layer=2 filter=2 channel=121
					-8, 3, -3, -7, -8, 8, 1, 3, 0,
					-- layer=2 filter=2 channel=122
					0, -2, -1, -6, -5, 8, 6, 3, -8,
					-- layer=2 filter=2 channel=123
					5, -14, 1, 9, 0, -6, 5, 0, 0,
					-- layer=2 filter=2 channel=124
					-12, -8, 4, -11, 0, -10, -8, -7, -7,
					-- layer=2 filter=2 channel=125
					-4, -2, -2, 6, 8, 10, 1, 4, -6,
					-- layer=2 filter=2 channel=126
					-9, 1, -2, -11, -1, -1, 6, 4, 2,
					-- layer=2 filter=2 channel=127
					-1, -5, -3, -9, 0, 9, -7, -1, 7,
					-- layer=2 filter=3 channel=0
					21, 31, 10, 21, 27, 33, -10, -13, -11,
					-- layer=2 filter=3 channel=1
					-7, -6, 20, -6, -27, 12, -15, -5, 7,
					-- layer=2 filter=3 channel=2
					-8, -3, -4, 6, -9, 0, 1, -1, 1,
					-- layer=2 filter=3 channel=3
					9, 30, 14, -32, 28, 21, -54, -18, -5,
					-- layer=2 filter=3 channel=4
					26, -11, -14, 2, -6, 17, -49, 0, 21,
					-- layer=2 filter=3 channel=5
					-11, -26, -17, 21, 51, 28, 0, 9, 0,
					-- layer=2 filter=3 channel=6
					-28, -15, -45, 11, 4, -7, 21, 79, 39,
					-- layer=2 filter=3 channel=7
					33, 75, 48, -22, 23, 7, -31, 9, -8,
					-- layer=2 filter=3 channel=8
					8, 9, -1, -3, -5, -3, 9, -3, 0,
					-- layer=2 filter=3 channel=9
					1, 11, 22, -15, -4, -14, 12, -20, 16,
					-- layer=2 filter=3 channel=10
					26, 23, 21, 6, 22, 7, -15, -34, -25,
					-- layer=2 filter=3 channel=11
					-26, -12, -24, -5, 11, -15, 4, -14, -28,
					-- layer=2 filter=3 channel=12
					-7, -7, 19, 13, 25, 28, -5, 14, 25,
					-- layer=2 filter=3 channel=13
					2, -7, -6, 7, 10, -7, -4, -8, 9,
					-- layer=2 filter=3 channel=14
					13, 4, 24, 7, 8, -4, -14, 7, 29,
					-- layer=2 filter=3 channel=15
					30, -1, -26, 56, 32, -2, 18, -21, -6,
					-- layer=2 filter=3 channel=16
					20, 22, 11, 2, 17, -9, -31, -28, -17,
					-- layer=2 filter=3 channel=17
					-1, -9, 0, -9, -2, -3, -4, -5, 5,
					-- layer=2 filter=3 channel=18
					-13, 15, -7, 34, -22, -29, 21, 28, 0,
					-- layer=2 filter=3 channel=19
					0, -33, -9, -25, -19, 7, 0, 3, 33,
					-- layer=2 filter=3 channel=20
					5, -10, 1, -5, 2, -1, -7, -6, 0,
					-- layer=2 filter=3 channel=21
					-32, -11, -24, -16, 2, -2, -14, -21, -27,
					-- layer=2 filter=3 channel=22
					-7, 2, 3, 3, 6, -3, 0, -8, -1,
					-- layer=2 filter=3 channel=23
					4, -10, 2, 9, -1, 19, -13, -12, 22,
					-- layer=2 filter=3 channel=24
					-39, 3, 7, -31, 5, 0, -10, -2, -4,
					-- layer=2 filter=3 channel=25
					-43, -27, -22, -30, -9, 0, -40, 3, 10,
					-- layer=2 filter=3 channel=26
					-8, -7, -2, -8, -4, -4, -12, 0, 3,
					-- layer=2 filter=3 channel=27
					-18, -49, -30, 0, 30, 12, 13, 20, 3,
					-- layer=2 filter=3 channel=28
					18, 22, -10, 55, 16, 21, -92, -53, -38,
					-- layer=2 filter=3 channel=29
					5, -2, -1, 8, -8, 3, -5, 3, -3,
					-- layer=2 filter=3 channel=30
					-8, -1, 7, 8, -13, 2, -7, -26, 7,
					-- layer=2 filter=3 channel=31
					68, -25, -96, 23, -45, -42, 12, -42, 1,
					-- layer=2 filter=3 channel=32
					-11, 8, -1, 5, -3, -12, 8, -5, 0,
					-- layer=2 filter=3 channel=33
					65, 24, 28, 5, 18, 3, -61, 8, -16,
					-- layer=2 filter=3 channel=34
					17, 6, -7, -6, -42, -32, 28, -24, -46,
					-- layer=2 filter=3 channel=35
					26, -1, -16, 23, 11, 15, -81, -19, -47,
					-- layer=2 filter=3 channel=36
					1, 10, 2, 11, 7, -6, -5, -12, 0,
					-- layer=2 filter=3 channel=37
					-16, -14, -14, 31, 6, -1, 3, 7, -2,
					-- layer=2 filter=3 channel=38
					0, -18, -29, 27, 9, -17, 4, 8, 0,
					-- layer=2 filter=3 channel=39
					14, 6, 13, 4, -12, -5, -5, -23, -16,
					-- layer=2 filter=3 channel=40
					-59, 75, -61, 21, -5, -8, -3, -33, -23,
					-- layer=2 filter=3 channel=41
					-7, 0, -8, 10, 3, 5, -8, 8, 0,
					-- layer=2 filter=3 channel=42
					-3, 16, 0, 9, 28, 2, -17, -1, 0,
					-- layer=2 filter=3 channel=43
					-13, 6, 4, 2, 2, 7, -53, -23, -19,
					-- layer=2 filter=3 channel=44
					-11, -10, -8, 6, 4, -8, 6, 3, 4,
					-- layer=2 filter=3 channel=45
					0, -40, -5, -34, 9, 9, -48, 26, 18,
					-- layer=2 filter=3 channel=46
					24, 9, 9, 11, 6, 1, -8, -3, -35,
					-- layer=2 filter=3 channel=47
					39, 48, 15, 21, 18, 33, -69, -6, -19,
					-- layer=2 filter=3 channel=48
					2, 2, -3, -5, 1, -3, -10, -3, -7,
					-- layer=2 filter=3 channel=49
					-44, -12, 14, 15, -9, -3, 16, 51, 23,
					-- layer=2 filter=3 channel=50
					12, -15, 0, -27, -4, -9, -27, -7, -3,
					-- layer=2 filter=3 channel=51
					-25, -8, -21, 11, -1, -15, -1, -10, -27,
					-- layer=2 filter=3 channel=52
					-43, -6, -6, -4, -23, -10, 27, 18, 3,
					-- layer=2 filter=3 channel=53
					5, -54, -69, 31, -37, 58, 10, -17, 12,
					-- layer=2 filter=3 channel=54
					-5, 0, -24, -21, -12, -24, -46, -23, -20,
					-- layer=2 filter=3 channel=55
					4, 0, 3, 4, -4, 6, 6, 8, 6,
					-- layer=2 filter=3 channel=56
					4, -16, -42, 25, 25, 12, 10, 17, 4,
					-- layer=2 filter=3 channel=57
					0, -4, -10, 9, -12, -1, 0, 5, 17,
					-- layer=2 filter=3 channel=58
					-1, -1, -20, 26, 2, 42, 13, 15, 23,
					-- layer=2 filter=3 channel=59
					25, 13, 20, 11, -23, -28, -8, 45, -20,
					-- layer=2 filter=3 channel=60
					8, 0, -11, 11, 14, -38, 10, 5, 22,
					-- layer=2 filter=3 channel=61
					-5, -24, -35, 18, 12, -41, -10, 46, 7,
					-- layer=2 filter=3 channel=62
					-12, -17, -39, -16, -9, -41, 26, 20, 5,
					-- layer=2 filter=3 channel=63
					-2, 19, 16, 12, 28, 22, -3, -3, -9,
					-- layer=2 filter=3 channel=64
					-5, -5, 17, 11, 12, 7, 7, 4, 0,
					-- layer=2 filter=3 channel=65
					-9, -19, -17, 21, -7, -29, 7, 24, 0,
					-- layer=2 filter=3 channel=66
					-7, 25, 1, -34, 49, -14, -24, -22, 9,
					-- layer=2 filter=3 channel=67
					23, 16, 20, -6, 15, -43, -1, -30, -13,
					-- layer=2 filter=3 channel=68
					0, 4, 7, 6, 4, 9, 9, 4, -1,
					-- layer=2 filter=3 channel=69
					-2, -10, 23, 17, 6, 1, -3, 1, 5,
					-- layer=2 filter=3 channel=70
					6, -13, -34, 38, 21, 18, -72, -33, -36,
					-- layer=2 filter=3 channel=71
					-41, -64, -36, -14, -18, -11, 1, 40, 7,
					-- layer=2 filter=3 channel=72
					43, 18, 7, 8, 9, -14, -50, 5, -12,
					-- layer=2 filter=3 channel=73
					23, -29, -64, 21, -6, 21, 31, -24, 10,
					-- layer=2 filter=3 channel=74
					23, 30, 14, 23, -4, -17, -9, -30, -14,
					-- layer=2 filter=3 channel=75
					-12, 49, -15, 47, 45, 54, 8, -9, 25,
					-- layer=2 filter=3 channel=76
					26, -31, -42, 54, -78, -25, 44, 9, 31,
					-- layer=2 filter=3 channel=77
					-4, 0, -8, 0, 0, 0, 3, 5, 2,
					-- layer=2 filter=3 channel=78
					-34, 1, -9, 10, -2, -13, -5, -19, -41,
					-- layer=2 filter=3 channel=79
					-7, -3, 7, -5, 2, -7, -6, -4, -8,
					-- layer=2 filter=3 channel=80
					19, 1, 7, 10, -6, 18, -40, -27, -2,
					-- layer=2 filter=3 channel=81
					2, -5, -9, -4, 1, -5, -5, 10, -7,
					-- layer=2 filter=3 channel=82
					4, 8, -5, 4, 12, -1, -6, 6, 3,
					-- layer=2 filter=3 channel=83
					16, -4, 9, 19, 7, 19, -37, -45, -38,
					-- layer=2 filter=3 channel=84
					2, -5, 7, 1, 9, 10, 4, 4, -6,
					-- layer=2 filter=3 channel=85
					4, 3, 8, 12, 7, -13, -5, -6, 9,
					-- layer=2 filter=3 channel=86
					10, -7, 3, 3, 0, -1, -8, -7, 1,
					-- layer=2 filter=3 channel=87
					16, -14, -47, -7, -73, -39, -2, -1, 18,
					-- layer=2 filter=3 channel=88
					15, 23, 8, 39, 1, 1, 10, 8, -10,
					-- layer=2 filter=3 channel=89
					-2, -2, 18, 32, -19, 3, 4, 20, 13,
					-- layer=2 filter=3 channel=90
					-1, 3, 2, -2, 9, -8, -5, -1, -1,
					-- layer=2 filter=3 channel=91
					-4, 17, -19, 31, -11, 31, -6, 12, 24,
					-- layer=2 filter=3 channel=92
					4, -4, 17, 8, 11, 17, -18, 12, 6,
					-- layer=2 filter=3 channel=93
					-12, -33, -6, 7, -49, 15, 32, 23, 35,
					-- layer=2 filter=3 channel=94
					15, -11, -19, -36, 51, -7, 40, 65, 25,
					-- layer=2 filter=3 channel=95
					-14, -7, 4, 2, 11, 9, 5, 5, 9,
					-- layer=2 filter=3 channel=96
					-26, -74, 3, 21, -48, -26, 58, 29, 32,
					-- layer=2 filter=3 channel=97
					-17, 5, 16, -9, 7, 45, 9, 10, 3,
					-- layer=2 filter=3 channel=98
					23, 24, -10, 20, 19, 6, -83, -41, -26,
					-- layer=2 filter=3 channel=99
					-17, -16, -15, -29, 22, -20, 34, 32, 14,
					-- layer=2 filter=3 channel=100
					14, -23, -13, 12, 12, 8, -21, -53, -10,
					-- layer=2 filter=3 channel=101
					-16, -14, -13, 13, 16, 21, -33, 1, 28,
					-- layer=2 filter=3 channel=102
					-49, -64, -7, 22, -32, -59, 29, 24, 10,
					-- layer=2 filter=3 channel=103
					-9, -17, -33, 14, -30, -21, -56, -7, -2,
					-- layer=2 filter=3 channel=104
					7, -47, -40, 0, 3, 0, 9, 35, 7,
					-- layer=2 filter=3 channel=105
					19, -15, -28, 7, -12, -37, 26, 33, -10,
					-- layer=2 filter=3 channel=106
					-5, 1, -33, 7, 5, 15, -8, 17, 20,
					-- layer=2 filter=3 channel=107
					18, 10, 18, -30, 39, 27, -1, -11, -24,
					-- layer=2 filter=3 channel=108
					-56, -72, -12, -7, 0, -4, 4, 23, 20,
					-- layer=2 filter=3 channel=109
					1, 0, 7, 8, 12, 3, 19, -4, 8,
					-- layer=2 filter=3 channel=110
					6, 10, 20, 13, 4, 15, 5, 7, 30,
					-- layer=2 filter=3 channel=111
					-10, 11, -7, -8, 6, 0, 5, 11, -9,
					-- layer=2 filter=3 channel=112
					-6, -4, -6, 25, 24, 25, 0, 5, -5,
					-- layer=2 filter=3 channel=113
					-9, 7, 7, 23, -14, 37, -14, -30, -36,
					-- layer=2 filter=3 channel=114
					-4, 16, 13, -1, -1, 5, 7, 7, 0,
					-- layer=2 filter=3 channel=115
					0, 1, -5, 3, 1, 8, -3, -1, 6,
					-- layer=2 filter=3 channel=116
					7, 9, -25, 20, -43, -28, 14, -5, 18,
					-- layer=2 filter=3 channel=117
					7, 40, -16, -43, 8, -47, -70, -57, -32,
					-- layer=2 filter=3 channel=118
					15, 26, -8, 7, -11, 21, -17, -8, -8,
					-- layer=2 filter=3 channel=119
					-15, -22, -11, 10, 29, -8, -23, -13, 8,
					-- layer=2 filter=3 channel=120
					-9, 3, -1, -2, -8, -9, 4, 2, 6,
					-- layer=2 filter=3 channel=121
					2, 0, -8, 11, 5, 3, 4, 3, 0,
					-- layer=2 filter=3 channel=122
					-2, 4, 1, -2, 15, 0, -1, -14, -2,
					-- layer=2 filter=3 channel=123
					33, 25, 20, -23, -24, -13, -13, 17, -36,
					-- layer=2 filter=3 channel=124
					23, -8, 4, 3, 18, 17, 29, 14, -30,
					-- layer=2 filter=3 channel=125
					8, 5, -4, -9, 3, 2, 12, 7, 7,
					-- layer=2 filter=3 channel=126
					-34, 1, 30, -38, 18, 34, -26, 20, 64,
					-- layer=2 filter=3 channel=127
					-6, -8, 23, 14, -3, -1, -23, -1, -30,
					-- layer=2 filter=4 channel=0
					-4, 3, -3, 0, -9, 1, 8, 5, -5,
					-- layer=2 filter=4 channel=1
					-19, -11, 3, -8, 0, -3, -13, -5, -1,
					-- layer=2 filter=4 channel=2
					-1, 12, -2, 3, 10, -8, -5, -3, 11,
					-- layer=2 filter=4 channel=3
					-3, -2, -6, 2, -3, -14, -12, -1, -8,
					-- layer=2 filter=4 channel=4
					-4, -13, -2, -2, -2, -17, 5, 0, -7,
					-- layer=2 filter=4 channel=5
					4, -1, -3, -9, 1, 5, 0, -2, -5,
					-- layer=2 filter=4 channel=6
					-14, 0, -20, -7, -9, 12, 8, -1, 12,
					-- layer=2 filter=4 channel=7
					-23, -20, -15, 0, 2, -15, 1, -15, -13,
					-- layer=2 filter=4 channel=8
					10, 1, -2, 6, 5, -8, 4, 0, 8,
					-- layer=2 filter=4 channel=9
					-2, 2, 7, -8, -8, -6, -5, 2, 5,
					-- layer=2 filter=4 channel=10
					-8, -7, -7, 3, -5, -14, 4, 5, -5,
					-- layer=2 filter=4 channel=11
					-4, -2, -11, 0, 0, -3, -2, -13, -5,
					-- layer=2 filter=4 channel=12
					-6, -3, -9, -7, -6, -21, 0, -3, -9,
					-- layer=2 filter=4 channel=13
					9, 11, 11, 8, 7, -11, 8, -10, 7,
					-- layer=2 filter=4 channel=14
					-21, -20, 0, -11, -9, -19, -15, 3, -6,
					-- layer=2 filter=4 channel=15
					-8, 0, -3, -6, -13, -16, -13, -20, -7,
					-- layer=2 filter=4 channel=16
					6, -1, 0, -1, -6, 7, 3, -6, -2,
					-- layer=2 filter=4 channel=17
					10, -1, -5, -3, 1, 6, -2, -9, -2,
					-- layer=2 filter=4 channel=18
					-9, -8, -11, -10, 8, -5, -2, -7, -16,
					-- layer=2 filter=4 channel=19
					-17, -20, -16, -12, -6, -8, -11, -4, 3,
					-- layer=2 filter=4 channel=20
					-3, 3, 8, 9, 10, 7, 8, 9, 2,
					-- layer=2 filter=4 channel=21
					5, -1, -2, 0, 1, -1, 0, 10, 9,
					-- layer=2 filter=4 channel=22
					-9, 4, 0, -8, 1, 3, 2, 7, 6,
					-- layer=2 filter=4 channel=23
					0, 3, -9, -6, 0, -10, 3, 1, -6,
					-- layer=2 filter=4 channel=24
					0, 1, -11, -7, 0, -14, -8, -7, -4,
					-- layer=2 filter=4 channel=25
					-13, -8, -6, -5, -18, -11, -7, -1, -19,
					-- layer=2 filter=4 channel=26
					6, -10, -4, 0, 0, 0, -2, -9, 0,
					-- layer=2 filter=4 channel=27
					-7, -13, 1, -8, 15, 12, 12, 20, 24,
					-- layer=2 filter=4 channel=28
					-12, -27, -20, 0, 4, -19, -6, -4, -8,
					-- layer=2 filter=4 channel=29
					5, 10, 8, 11, 8, -2, -3, 3, 7,
					-- layer=2 filter=4 channel=30
					11, -8, -7, -4, -3, 5, -4, -11, -11,
					-- layer=2 filter=4 channel=31
					-1, -9, 0, -1, 3, 13, 6, -11, 1,
					-- layer=2 filter=4 channel=32
					7, 12, 11, 11, -5, 0, -7, 7, 7,
					-- layer=2 filter=4 channel=33
					-9, -12, -16, 15, 11, 8, 11, -13, 10,
					-- layer=2 filter=4 channel=34
					-10, -23, 5, -9, -6, -14, 19, 15, 14,
					-- layer=2 filter=4 channel=35
					-18, -13, -25, -6, -10, -17, -7, -16, -15,
					-- layer=2 filter=4 channel=36
					4, -1, -6, -4, -8, 1, 5, -7, 9,
					-- layer=2 filter=4 channel=37
					4, -9, -5, -11, -12, -6, -4, -4, 4,
					-- layer=2 filter=4 channel=38
					-2, 1, 0, -16, 0, 3, -5, 4, 7,
					-- layer=2 filter=4 channel=39
					1, 4, 0, -4, -6, 2, 2, -11, -11,
					-- layer=2 filter=4 channel=40
					-32, -25, 4, 1, 2, -14, 17, -5, 2,
					-- layer=2 filter=4 channel=41
					8, -8, -10, -2, 8, -2, 9, 5, 5,
					-- layer=2 filter=4 channel=42
					-9, -6, -5, -1, 0, -10, -8, 3, -6,
					-- layer=2 filter=4 channel=43
					6, -11, -16, 0, 5, -1, -7, -8, 6,
					-- layer=2 filter=4 channel=44
					6, 3, -3, -10, -9, -4, 1, 5, 0,
					-- layer=2 filter=4 channel=45
					-16, -9, 0, -11, -9, -14, 7, -8, -3,
					-- layer=2 filter=4 channel=46
					-4, -4, -7, 1, -10, -13, 6, 2, 7,
					-- layer=2 filter=4 channel=47
					0, -12, -4, 10, 3, -7, 12, -17, -8,
					-- layer=2 filter=4 channel=48
					7, 2, -4, -5, -3, 4, 2, 9, 9,
					-- layer=2 filter=4 channel=49
					-13, -15, -5, -2, -19, -13, -9, -21, -13,
					-- layer=2 filter=4 channel=50
					-7, 5, 11, -9, 10, 1, 5, -12, -8,
					-- layer=2 filter=4 channel=51
					-1, -2, -9, -9, 7, 9, -7, 2, 0,
					-- layer=2 filter=4 channel=52
					5, -3, 8, -15, -5, -6, -11, 6, 2,
					-- layer=2 filter=4 channel=53
					-8, -3, -12, -13, -12, -7, 11, -11, 5,
					-- layer=2 filter=4 channel=54
					-21, -22, -4, -22, -16, -7, -12, -8, -13,
					-- layer=2 filter=4 channel=55
					-7, 0, -8, -1, 4, -4, -8, 6, -4,
					-- layer=2 filter=4 channel=56
					7, -3, -7, 0, -12, 0, 3, 7, -6,
					-- layer=2 filter=4 channel=57
					-5, 5, 11, -3, 4, 8, 4, 2, 7,
					-- layer=2 filter=4 channel=58
					-8, 3, -16, -9, -11, -14, 1, -11, -17,
					-- layer=2 filter=4 channel=59
					-16, 7, 4, -12, -4, 0, -1, -4, -6,
					-- layer=2 filter=4 channel=60
					-20, -1, -6, -17, -18, 2, -22, 2, -10,
					-- layer=2 filter=4 channel=61
					2, -5, -10, 0, -9, 4, -31, -1, 0,
					-- layer=2 filter=4 channel=62
					-4, -12, -10, -5, -17, -4, -5, 1, 0,
					-- layer=2 filter=4 channel=63
					7, 9, -6, -2, 6, -11, 9, 1, -5,
					-- layer=2 filter=4 channel=64
					-3, -14, -4, 7, 0, -9, 0, -9, -5,
					-- layer=2 filter=4 channel=65
					-18, -4, -2, -7, 0, 2, -1, 8, -5,
					-- layer=2 filter=4 channel=66
					4, -2, -2, 1, -9, 4, -5, 2, 3,
					-- layer=2 filter=4 channel=67
					-6, 7, -3, 5, -1, -4, 0, -9, 6,
					-- layer=2 filter=4 channel=68
					12, 0, -2, 3, -7, 1, 6, -8, -4,
					-- layer=2 filter=4 channel=69
					4, 5, -9, 3, 2, -6, -7, 0, -15,
					-- layer=2 filter=4 channel=70
					-26, -11, -10, -13, -7, -6, -3, -17, -1,
					-- layer=2 filter=4 channel=71
					-13, -11, 7, -19, -16, -5, -4, -4, -12,
					-- layer=2 filter=4 channel=72
					-18, -11, -5, -4, -9, 8, -8, 4, 10,
					-- layer=2 filter=4 channel=73
					-10, 1, -5, -12, -13, 2, -8, -15, -9,
					-- layer=2 filter=4 channel=74
					-2, -4, -12, 0, -1, 4, -4, 2, -1,
					-- layer=2 filter=4 channel=75
					-8, -15, 5, -7, 4, 2, 9, -2, -5,
					-- layer=2 filter=4 channel=76
					-19, 5, -18, -2, 4, -8, 19, -14, 1,
					-- layer=2 filter=4 channel=77
					-9, -9, -3, -4, 6, 7, 2, 8, -4,
					-- layer=2 filter=4 channel=78
					-8, -14, -8, -8, 0, -1, -10, 0, -3,
					-- layer=2 filter=4 channel=79
					8, 4, -2, 2, -1, 4, 2, -3, -3,
					-- layer=2 filter=4 channel=80
					-8, 6, -2, 3, -1, -4, -8, -9, -3,
					-- layer=2 filter=4 channel=81
					4, 5, -9, 3, -3, 6, -9, -2, -2,
					-- layer=2 filter=4 channel=82
					-1, -9, 5, 6, -6, 7, 0, 2, -8,
					-- layer=2 filter=4 channel=83
					2, 2, -3, 6, -2, -8, -2, -11, -9,
					-- layer=2 filter=4 channel=84
					7, -1, -8, 3, -4, -6, 2, -9, -6,
					-- layer=2 filter=4 channel=85
					-1, -4, 0, 4, 5, -8, -4, 5, 2,
					-- layer=2 filter=4 channel=86
					-10, -5, 3, 9, 0, -6, 6, -7, 2,
					-- layer=2 filter=4 channel=87
					-16, -3, -12, 3, -1, -17, -2, -16, 2,
					-- layer=2 filter=4 channel=88
					5, 8, 6, -7, 0, -5, 9, -5, 2,
					-- layer=2 filter=4 channel=89
					-28, -22, -24, -13, -13, -7, -18, -1, -5,
					-- layer=2 filter=4 channel=90
					-5, -8, 2, 7, -4, -6, -6, 7, -9,
					-- layer=2 filter=4 channel=91
					-1, -4, -1, -2, -13, -5, -14, -14, -3,
					-- layer=2 filter=4 channel=92
					-14, -18, -3, -14, -13, -15, -4, 3, -3,
					-- layer=2 filter=4 channel=93
					1, -12, -13, -11, 8, -6, -2, 13, -7,
					-- layer=2 filter=4 channel=94
					-2, -23, -31, -34, -12, 3, -13, -12, 7,
					-- layer=2 filter=4 channel=95
					-5, 5, -6, 3, 5, 9, 5, 0, 3,
					-- layer=2 filter=4 channel=96
					15, -1, 9, -2, 0, 8, 2, 17, 13,
					-- layer=2 filter=4 channel=97
					0, -1, -11, 0, -12, -10, -4, -16, 2,
					-- layer=2 filter=4 channel=98
					-24, -19, 1, 7, 12, 5, 5, -14, -11,
					-- layer=2 filter=4 channel=99
					-14, 0, 0, -16, -11, 0, -3, -10, 6,
					-- layer=2 filter=4 channel=100
					-4, -9, 6, 5, -1, -10, 1, -2, -10,
					-- layer=2 filter=4 channel=101
					0, 0, -5, 2, -10, 5, -9, -8, 3,
					-- layer=2 filter=4 channel=102
					3, -17, -19, 8, 4, -16, 16, -3, -18,
					-- layer=2 filter=4 channel=103
					-5, 0, 3, -6, -8, 7, -8, -1, -4,
					-- layer=2 filter=4 channel=104
					-9, -6, -16, 5, -22, -3, 4, -6, -2,
					-- layer=2 filter=4 channel=105
					-5, 3, -3, -6, 0, -11, -4, 4, 4,
					-- layer=2 filter=4 channel=106
					-1, 5, -13, -13, 3, 3, -3, -13, -9,
					-- layer=2 filter=4 channel=107
					9, -3, -10, 0, -8, -5, -2, -9, -2,
					-- layer=2 filter=4 channel=108
					-8, -1, -6, -13, -3, 0, 2, -2, -8,
					-- layer=2 filter=4 channel=109
					11, -2, 1, 0, -5, 0, 2, 1, -7,
					-- layer=2 filter=4 channel=110
					-14, -5, -12, -4, -13, -12, 0, -16, -15,
					-- layer=2 filter=4 channel=111
					6, -9, -2, 0, 0, -5, 2, 6, -4,
					-- layer=2 filter=4 channel=112
					-2, -7, 4, -13, -2, 0, -8, 0, 4,
					-- layer=2 filter=4 channel=113
					6, -7, 3, -10, 0, 4, 7, -9, 2,
					-- layer=2 filter=4 channel=114
					-6, -6, -7, 8, -6, 9, -7, -8, 8,
					-- layer=2 filter=4 channel=115
					8, 8, 11, 1, 2, -6, 2, 8, 7,
					-- layer=2 filter=4 channel=116
					-6, -7, -2, 3, 18, -14, -6, -17, -9,
					-- layer=2 filter=4 channel=117
					-9, -15, -22, -4, -14, -4, -23, -7, -7,
					-- layer=2 filter=4 channel=118
					-8, -10, -12, 0, -15, -14, -12, 0, -8,
					-- layer=2 filter=4 channel=119
					-10, -12, -7, 0, -9, -7, -10, -12, -4,
					-- layer=2 filter=4 channel=120
					6, 6, 8, 2, -7, -6, 0, -9, 3,
					-- layer=2 filter=4 channel=121
					4, 2, 9, -1, -6, 1, -1, 1, -7,
					-- layer=2 filter=4 channel=122
					-1, 8, 8, 4, 0, 5, -6, -6, -4,
					-- layer=2 filter=4 channel=123
					-8, -10, -1, -8, -9, -11, -13, -14, -9,
					-- layer=2 filter=4 channel=124
					-26, -14, -24, -8, -12, -8, -18, -2, 14,
					-- layer=2 filter=4 channel=125
					7, -8, -5, -2, -6, 10, 7, -4, -4,
					-- layer=2 filter=4 channel=126
					6, 0, 0, -1, 1, 6, -29, -11, 12,
					-- layer=2 filter=4 channel=127
					-7, -5, -5, 8, -11, -4, 8, -1, -1,
					-- layer=2 filter=5 channel=0
					14, 21, 0, 14, 16, 18, -17, 21, -8,
					-- layer=2 filter=5 channel=1
					44, -31, 1, -38, -22, -37, -28, -22, -6,
					-- layer=2 filter=5 channel=2
					-5, 9, 9, 8, 1, 3, -8, -5, 3,
					-- layer=2 filter=5 channel=3
					16, 8, 10, 11, 10, -1, -28, -18, -2,
					-- layer=2 filter=5 channel=4
					-53, -26, -30, -8, 13, 11, 2, -3, 8,
					-- layer=2 filter=5 channel=5
					12, 22, 1, -19, 15, 4, 9, 15, 30,
					-- layer=2 filter=5 channel=6
					27, -14, 27, 28, -14, 6, 20, 0, 27,
					-- layer=2 filter=5 channel=7
					-35, -40, -24, 2, -56, 37, -40, -32, -47,
					-- layer=2 filter=5 channel=8
					2, -7, -1, -6, -4, -10, 4, -1, 7,
					-- layer=2 filter=5 channel=9
					24, 2, -3, -34, 12, 0, -18, -12, -6,
					-- layer=2 filter=5 channel=10
					3, 35, 22, 7, 19, 44, -2, 17, -2,
					-- layer=2 filter=5 channel=11
					7, 7, -10, 10, 6, 5, -2, 20, 14,
					-- layer=2 filter=5 channel=12
					10, -5, -55, -53, -27, -46, -40, -40, -9,
					-- layer=2 filter=5 channel=13
					-8, -6, -1, 5, 0, -8, 8, -1, 6,
					-- layer=2 filter=5 channel=14
					28, -23, -60, -44, -8, -49, -28, -33, 14,
					-- layer=2 filter=5 channel=15
					26, -59, 46, -27, 13, 10, -2, 3, 47,
					-- layer=2 filter=5 channel=16
					-25, -28, -38, 0, 3, -9, 15, 18, 20,
					-- layer=2 filter=5 channel=17
					1, 6, -4, 6, 0, 4, 2, 10, -6,
					-- layer=2 filter=5 channel=18
					1, -29, 1, 34, 12, -24, -7, -20, -7,
					-- layer=2 filter=5 channel=19
					-15, 2, 36, -14, -38, 17, -10, -10, -10,
					-- layer=2 filter=5 channel=20
					1, 4, -5, -6, 5, 6, -3, 2, 5,
					-- layer=2 filter=5 channel=21
					17, 17, 1, 7, 13, 9, 7, 0, 0,
					-- layer=2 filter=5 channel=22
					10, 10, 2, -3, 6, 1, 2, 5, 0,
					-- layer=2 filter=5 channel=23
					-10, 28, 14, 0, -6, 7, 11, -28, 8,
					-- layer=2 filter=5 channel=24
					5, 9, -14, 36, -5, 7, 8, -3, -15,
					-- layer=2 filter=5 channel=25
					6, 0, -9, 26, -19, -14, 1, -8, -25,
					-- layer=2 filter=5 channel=26
					-10, -7, -3, -7, -7, -9, 10, -7, -4,
					-- layer=2 filter=5 channel=27
					-18, -10, -39, -47, -4, 4, -51, -14, 18,
					-- layer=2 filter=5 channel=28
					-21, -16, -30, -4, -28, -28, -43, -15, -22,
					-- layer=2 filter=5 channel=29
					-8, 6, 0, -1, 12, 0, 4, 7, 7,
					-- layer=2 filter=5 channel=30
					-13, -6, -14, -17, 6, 4, 0, 0, -9,
					-- layer=2 filter=5 channel=31
					-29, -11, 33, -22, 11, 43, -1, 35, 1,
					-- layer=2 filter=5 channel=32
					-1, -1, 11, -9, -4, -4, 1, 2, -1,
					-- layer=2 filter=5 channel=33
					-10, 6, 5, -64, -45, -25, -65, -69, -4,
					-- layer=2 filter=5 channel=34
					-41, 23, -7, -4, -4, 18, 4, 28, 43,
					-- layer=2 filter=5 channel=35
					-22, 1, -3, -33, -31, -11, -23, -52, -14,
					-- layer=2 filter=5 channel=36
					11, 0, -1, 7, 8, 14, -5, 9, 5,
					-- layer=2 filter=5 channel=37
					-5, -1, 0, 3, 37, 8, -2, 25, 26,
					-- layer=2 filter=5 channel=38
					-25, -27, 13, -41, -2, -3, -1, 1, 19,
					-- layer=2 filter=5 channel=39
					-30, -50, -30, -72, -37, 19, -40, -46, 15,
					-- layer=2 filter=5 channel=40
					-28, -44, -10, 2, -10, -27, -33, 0, 6,
					-- layer=2 filter=5 channel=41
					-9, 0, 0, -1, -8, -3, 9, -4, 4,
					-- layer=2 filter=5 channel=42
					14, 11, -10, -6, -3, -4, -8, -14, 8,
					-- layer=2 filter=5 channel=43
					5, 18, -24, 19, 12, -22, -13, 10, -13,
					-- layer=2 filter=5 channel=44
					1, -8, -7, 9, -9, 5, -3, -5, -3,
					-- layer=2 filter=5 channel=45
					-55, -80, -60, -90, -41, -48, -113, -30, 7,
					-- layer=2 filter=5 channel=46
					-11, 0, -13, -26, 12, -6, -13, 0, -9,
					-- layer=2 filter=5 channel=47
					-48, -17, -38, -30, -40, -8, -97, -74, 13,
					-- layer=2 filter=5 channel=48
					-4, -9, -7, 5, -9, 0, 0, -4, 0,
					-- layer=2 filter=5 channel=49
					32, -33, -25, 62, 17, -5, 23, -29, 34,
					-- layer=2 filter=5 channel=50
					0, -6, -11, -11, 12, -17, 4, 10, 5,
					-- layer=2 filter=5 channel=51
					19, 2, 11, 4, 26, 1, 8, 25, 19,
					-- layer=2 filter=5 channel=52
					9, -18, 35, 25, 16, 5, 29, 22, 24,
					-- layer=2 filter=5 channel=53
					-33, -51, -32, 2, 0, 52, -28, 18, 60,
					-- layer=2 filter=5 channel=54
					4, 18, 0, 8, -21, 38, -18, 7, -2,
					-- layer=2 filter=5 channel=55
					4, -8, -6, -3, 4, 0, -1, -4, 9,
					-- layer=2 filter=5 channel=56
					-15, 9, -5, -2, 0, -5, -20, 2, 10,
					-- layer=2 filter=5 channel=57
					4, -5, -7, 5, -3, -4, 4, 9, -7,
					-- layer=2 filter=5 channel=58
					-9, -2, 14, -101, -52, -29, -58, -35, -6,
					-- layer=2 filter=5 channel=59
					-43, -15, 1, -68, -40, 11, -47, 31, 22,
					-- layer=2 filter=5 channel=60
					11, -13, 37, 9, -3, 50, -4, 34, 17,
					-- layer=2 filter=5 channel=61
					0, 2, 14, 21, -50, 10, -28, 16, -28,
					-- layer=2 filter=5 channel=62
					9, -5, 18, 34, 2, -19, 22, 10, 4,
					-- layer=2 filter=5 channel=63
					-48, -7, -14, 0, -41, 33, -30, 0, -27,
					-- layer=2 filter=5 channel=64
					8, -5, 9, 3, -18, 29, 42, -12, 4,
					-- layer=2 filter=5 channel=65
					-12, 9, 39, 22, -15, -3, 4, 17, 6,
					-- layer=2 filter=5 channel=66
					19, 0, 20, 25, -16, 11, -38, -14, 0,
					-- layer=2 filter=5 channel=67
					-26, 0, 14, -47, -8, -6, -18, -1, -21,
					-- layer=2 filter=5 channel=68
					-10, 10, -9, 4, 7, 8, -4, -7, 4,
					-- layer=2 filter=5 channel=69
					14, -14, -25, -10, -3, 15, -7, -33, 27,
					-- layer=2 filter=5 channel=70
					-25, 15, 5, -35, -16, 26, 18, -21, 33,
					-- layer=2 filter=5 channel=71
					-13, -20, -44, -1, -59, -68, -24, -48, -35,
					-- layer=2 filter=5 channel=72
					16, -12, 11, 0, -15, 23, 0, 32, 30,
					-- layer=2 filter=5 channel=73
					0, 33, 31, 42, 51, 26, -24, 61, 21,
					-- layer=2 filter=5 channel=74
					-39, 0, -6, -32, -47, -12, -19, 31, 1,
					-- layer=2 filter=5 channel=75
					-38, -8, -64, -65, -43, -64, -3, -5, -23,
					-- layer=2 filter=5 channel=76
					-35, -25, -4, 19, 8, 25, -22, 17, 30,
					-- layer=2 filter=5 channel=77
					0, 6, 3, -6, 10, 11, -1, 5, -6,
					-- layer=2 filter=5 channel=78
					8, 23, 9, 51, 11, 15, 19, 28, -2,
					-- layer=2 filter=5 channel=79
					-6, -4, 3, -4, -1, 2, 4, -1, -1,
					-- layer=2 filter=5 channel=80
					-39, -7, -23, -21, 7, 8, 30, -29, -8,
					-- layer=2 filter=5 channel=81
					-1, 1, 3, 13, 7, 3, 1, 0, -5,
					-- layer=2 filter=5 channel=82
					-9, -3, 4, -5, -1, 8, -1, -5, 4,
					-- layer=2 filter=5 channel=83
					-36, -2, 18, -11, -19, 15, 26, -25, 6,
					-- layer=2 filter=5 channel=84
					4, -4, 0, 3, -8, -3, -7, 0, 10,
					-- layer=2 filter=5 channel=85
					4, 0, 8, -3, -12, 8, -6, -8, 11,
					-- layer=2 filter=5 channel=86
					11, 2, -10, 1, -3, -6, 0, -8, 5,
					-- layer=2 filter=5 channel=87
					-19, 15, 24, 10, 6, 21, -37, 34, 30,
					-- layer=2 filter=5 channel=88
					-22, -40, -30, -53, -38, -31, -61, -2, -11,
					-- layer=2 filter=5 channel=89
					21, -16, -6, -68, -19, -19, -20, 5, 29,
					-- layer=2 filter=5 channel=90
					-7, -5, -9, 5, 6, -9, 0, -9, 8,
					-- layer=2 filter=5 channel=91
					0, -11, 0, -85, -21, -9, -48, 18, 24,
					-- layer=2 filter=5 channel=92
					43, -10, -24, -60, -19, -62, -50, -17, 10,
					-- layer=2 filter=5 channel=93
					-12, 61, 71, 21, 26, 3, 13, 18, -5,
					-- layer=2 filter=5 channel=94
					15, -20, -12, 32, -38, 12, -25, 26, -2,
					-- layer=2 filter=5 channel=95
					-12, -3, -14, -13, -9, -10, -16, 0, -6,
					-- layer=2 filter=5 channel=96
					18, 49, 32, 7, 49, 1, -17, 13, 25,
					-- layer=2 filter=5 channel=97
					-11, -15, -40, 20, -8, -7, -11, -18, -12,
					-- layer=2 filter=5 channel=98
					-48, 0, -4, -3, -19, 28, -34, 11, -16,
					-- layer=2 filter=5 channel=99
					13, 3, 40, 7, -23, 7, 2, 10, 20,
					-- layer=2 filter=5 channel=100
					-33, -6, 33, -34, -8, 16, -30, 16, 23,
					-- layer=2 filter=5 channel=101
					0, -10, -30, -13, -21, -59, -21, -26, -42,
					-- layer=2 filter=5 channel=102
					27, 28, 20, 12, 17, -10, 16, 8, 18,
					-- layer=2 filter=5 channel=103
					-56, -8, 8, -1, -3, -60, 16, 1, -11,
					-- layer=2 filter=5 channel=104
					7, -30, -4, 32, 41, -1, 7, 45, 19,
					-- layer=2 filter=5 channel=105
					-42, -43, -29, -21, -72, -51, 11, 1, -17,
					-- layer=2 filter=5 channel=106
					-8, -20, -27, -18, -27, -34, -18, -14, -12,
					-- layer=2 filter=5 channel=107
					32, -10, 46, 1, 48, -9, -54, 36, 59,
					-- layer=2 filter=5 channel=108
					35, -4, -26, -32, 22, -15, 0, -11, 14,
					-- layer=2 filter=5 channel=109
					13, 0, -7, 13, 12, 2, 18, 6, -13,
					-- layer=2 filter=5 channel=110
					0, 24, 14, -19, -11, -14, -9, -17, -17,
					-- layer=2 filter=5 channel=111
					4, 4, 5, 7, -5, -6, -6, -10, 5,
					-- layer=2 filter=5 channel=112
					-30, -5, -11, -9, -15, 9, -23, -9, -13,
					-- layer=2 filter=5 channel=113
					-43, -17, 9, -12, 9, 7, -25, -1, -30,
					-- layer=2 filter=5 channel=114
					-2, -5, -17, 0, -7, -6, -3, -7, -12,
					-- layer=2 filter=5 channel=115
					-2, -8, -2, -4, 0, -12, 1, 4, -6,
					-- layer=2 filter=5 channel=116
					-11, -17, 31, -20, 1, -13, -36, 16, 61,
					-- layer=2 filter=5 channel=117
					-26, -1, 13, 32, -67, 37, -45, 0, -39,
					-- layer=2 filter=5 channel=118
					17, 35, 8, 54, 32, 1, 11, -3, 5,
					-- layer=2 filter=5 channel=119
					-16, -30, -40, -5, -35, -57, -60, -52, -44,
					-- layer=2 filter=5 channel=120
					4, 2, -4, 9, 4, 0, -5, 6, 0,
					-- layer=2 filter=5 channel=121
					-5, 7, 5, 10, -3, -1, 0, -1, 1,
					-- layer=2 filter=5 channel=122
					3, 14, 8, -5, 4, 9, 1, 12, -1,
					-- layer=2 filter=5 channel=123
					-44, -19, 19, 4, -27, 45, -49, -22, -30,
					-- layer=2 filter=5 channel=124
					30, -32, -6, 8, -15, 7, -33, 4, 19,
					-- layer=2 filter=5 channel=125
					9, 3, -4, -5, 6, 3, 6, -6, -8,
					-- layer=2 filter=5 channel=126
					-12, 96, 34, -18, 17, 26, -33, 48, -5,
					-- layer=2 filter=5 channel=127
					-25, -4, 5, -41, 0, 17, -26, -47, 7,
					-- layer=2 filter=6 channel=0
					3, -28, -7, 4, -6, -1, -21, -6, -1,
					-- layer=2 filter=6 channel=1
					2, -5, -18, 0, -5, -30, -21, -1, -13,
					-- layer=2 filter=6 channel=2
					1, 7, -6, -8, -7, -4, 0, 11, -4,
					-- layer=2 filter=6 channel=3
					-8, -22, 5, -12, -31, -17, 2, -11, -5,
					-- layer=2 filter=6 channel=4
					-20, -4, -1, -1, 6, -5, 17, 5, 12,
					-- layer=2 filter=6 channel=5
					-6, -28, -7, -13, -18, -5, -9, 0, 1,
					-- layer=2 filter=6 channel=6
					-10, -10, -28, -19, 1, -25, -9, -1, -29,
					-- layer=2 filter=6 channel=7
					0, 10, 20, -9, -22, -12, -11, -16, -5,
					-- layer=2 filter=6 channel=8
					-3, -4, 4, 4, 7, -6, -8, -4, -9,
					-- layer=2 filter=6 channel=9
					1, 0, -12, -16, -12, 16, -5, -3, 7,
					-- layer=2 filter=6 channel=10
					-6, -26, 0, -6, -5, 0, -15, 2, 7,
					-- layer=2 filter=6 channel=11
					-23, -5, -12, -26, -30, -19, -5, -23, -5,
					-- layer=2 filter=6 channel=12
					1, -3, -16, 5, -17, -24, -7, -13, -13,
					-- layer=2 filter=6 channel=13
					-8, -6, -8, 8, 4, -7, -3, 4, 5,
					-- layer=2 filter=6 channel=14
					-24, -24, -21, -4, -15, -22, -9, -17, -15,
					-- layer=2 filter=6 channel=15
					-29, 8, -20, 26, -1, -5, 6, 0, -14,
					-- layer=2 filter=6 channel=16
					-14, -18, -21, 3, -6, -22, 6, -16, -6,
					-- layer=2 filter=6 channel=17
					0, -4, -8, -11, 0, -1, 0, -4, 9,
					-- layer=2 filter=6 channel=18
					-21, -1, -6, -6, 6, -13, 7, -4, -6,
					-- layer=2 filter=6 channel=19
					17, -1, 10, 10, -13, -24, -9, -11, -24,
					-- layer=2 filter=6 channel=20
					-1, -11, 3, -6, -3, 0, 4, -7, 2,
					-- layer=2 filter=6 channel=21
					5, -8, 5, 7, 8, 5, -7, -6, -3,
					-- layer=2 filter=6 channel=22
					-5, -3, -1, 10, -3, 0, 6, 2, -7,
					-- layer=2 filter=6 channel=23
					-2, 4, -19, 0, -4, -15, 16, 0, 4,
					-- layer=2 filter=6 channel=24
					-14, -8, -2, -23, -16, -6, -19, -24, -27,
					-- layer=2 filter=6 channel=25
					-24, -4, -8, -18, -19, -20, -26, -14, -33,
					-- layer=2 filter=6 channel=26
					-4, 7, -2, -8, -9, -2, 5, 7, 2,
					-- layer=2 filter=6 channel=27
					3, -20, 3, -16, -30, 5, -14, -2, 0,
					-- layer=2 filter=6 channel=28
					-12, -1, 5, 0, 0, -17, -3, -15, -8,
					-- layer=2 filter=6 channel=29
					-12, 1, -7, 3, -4, -1, -4, -6, 1,
					-- layer=2 filter=6 channel=30
					-9, -5, -7, -13, 11, -1, -21, -12, -15,
					-- layer=2 filter=6 channel=31
					-25, 1, -1, 16, 7, 5, 9, -8, -10,
					-- layer=2 filter=6 channel=32
					-8, -6, 1, 0, 2, 2, 1, 4, 8,
					-- layer=2 filter=6 channel=33
					-8, 15, 3, 2, 2, -18, 0, -7, 4,
					-- layer=2 filter=6 channel=34
					-10, -24, -3, 5, 8, -7, -15, -1, -25,
					-- layer=2 filter=6 channel=35
					10, -1, 2, 2, -9, -8, -11, -1, -11,
					-- layer=2 filter=6 channel=36
					-12, -2, -2, -3, -1, -2, 8, -10, -8,
					-- layer=2 filter=6 channel=37
					-4, -4, -10, -20, -20, -4, -16, -17, -6,
					-- layer=2 filter=6 channel=38
					-14, -10, -14, -16, -16, -7, -20, -20, -16,
					-- layer=2 filter=6 channel=39
					-10, -2, -16, -6, -27, -12, -7, 4, -1,
					-- layer=2 filter=6 channel=40
					-37, -6, 0, -3, 13, 17, 10, -13, -7,
					-- layer=2 filter=6 channel=41
					-1, -9, 2, 9, 3, -9, 4, -4, 8,
					-- layer=2 filter=6 channel=42
					-12, -31, -13, -9, -10, -8, 11, -7, -3,
					-- layer=2 filter=6 channel=43
					-21, -14, 20, -11, 0, 7, 12, -7, 14,
					-- layer=2 filter=6 channel=44
					8, 9, -9, 0, 2, 8, 11, 9, -10,
					-- layer=2 filter=6 channel=45
					-4, -9, -1, 15, -11, -8, 12, 32, 18,
					-- layer=2 filter=6 channel=46
					-8, -11, -5, -13, -12, -9, -21, 9, 1,
					-- layer=2 filter=6 channel=47
					-6, -10, -3, -4, -1, -8, -23, -15, 9,
					-- layer=2 filter=6 channel=48
					6, -4, -3, 0, 10, 6, -7, -1, 7,
					-- layer=2 filter=6 channel=49
					-13, 6, -8, -5, -10, -19, 15, -15, -1,
					-- layer=2 filter=6 channel=50
					-8, -9, -4, -8, -11, 12, -7, 13, 4,
					-- layer=2 filter=6 channel=51
					-12, -14, -17, -31, -26, -18, -12, -19, -6,
					-- layer=2 filter=6 channel=52
					23, 1, -6, -6, -14, -1, 7, -5, -11,
					-- layer=2 filter=6 channel=53
					-30, -10, -5, -1, -12, -9, -2, -6, -13,
					-- layer=2 filter=6 channel=54
					-3, -8, 9, 12, -6, -7, -7, -25, -29,
					-- layer=2 filter=6 channel=55
					-7, -4, -3, 6, -6, -4, 8, -9, 4,
					-- layer=2 filter=6 channel=56
					-21, -26, -15, -12, -15, -32, -1, -3, -15,
					-- layer=2 filter=6 channel=57
					-7, 9, 12, 0, 0, 7, 2, -8, -1,
					-- layer=2 filter=6 channel=58
					27, -9, -16, 9, -6, -20, -2, -19, -13,
					-- layer=2 filter=6 channel=59
					-6, 22, 12, 2, -5, -17, -34, -9, -25,
					-- layer=2 filter=6 channel=60
					-13, -9, -29, -21, -12, -9, -33, -16, -5,
					-- layer=2 filter=6 channel=61
					-7, -3, -8, -12, -5, -10, -35, -11, 2,
					-- layer=2 filter=6 channel=62
					3, -7, -4, -13, 18, -9, -15, -15, -14,
					-- layer=2 filter=6 channel=63
					-16, -9, -15, 2, -9, -8, -13, -14, 3,
					-- layer=2 filter=6 channel=64
					-6, -10, -18, 1, -2, -1, -1, -16, -14,
					-- layer=2 filter=6 channel=65
					-17, 3, -15, -27, -10, -17, -21, -1, -17,
					-- layer=2 filter=6 channel=66
					-13, -4, -18, -11, -3, -19, 15, -9, -17,
					-- layer=2 filter=6 channel=67
					-9, -6, 17, -15, -14, 14, -4, -4, -9,
					-- layer=2 filter=6 channel=68
					0, -6, -11, -10, -4, 2, -3, -10, 6,
					-- layer=2 filter=6 channel=69
					-13, -5, -27, 1, -16, -4, 0, -20, -6,
					-- layer=2 filter=6 channel=70
					0, -17, -15, -2, -10, -8, 0, -9, -7,
					-- layer=2 filter=6 channel=71
					15, -18, -8, -12, -33, -7, -22, -4, 0,
					-- layer=2 filter=6 channel=72
					-15, -8, -13, -22, -19, -27, -2, -14, -15,
					-- layer=2 filter=6 channel=73
					-6, 6, -18, 3, -18, -21, 2, 8, -10,
					-- layer=2 filter=6 channel=74
					-11, -12, 6, -9, -7, 4, -1, 0, -6,
					-- layer=2 filter=6 channel=75
					7, -20, -30, 3, -2, -23, -3, -26, -13,
					-- layer=2 filter=6 channel=76
					-12, 25, 0, 2, -24, -7, -2, 8, -11,
					-- layer=2 filter=6 channel=77
					-10, 7, 7, 0, 6, -7, 6, -3, -5,
					-- layer=2 filter=6 channel=78
					-17, -9, -21, -38, -17, -10, -10, -19, -40,
					-- layer=2 filter=6 channel=79
					-5, 2, 0, -1, -3, -3, 6, -4, 8,
					-- layer=2 filter=6 channel=80
					-17, -4, -4, 2, -11, 5, 4, -2, 6,
					-- layer=2 filter=6 channel=81
					-2, -12, 5, -5, 5, -12, -8, -5, -10,
					-- layer=2 filter=6 channel=82
					-8, 10, 1, 5, 9, 1, 0, -6, -6,
					-- layer=2 filter=6 channel=83
					13, -3, -9, -3, -1, 0, 6, 15, 9,
					-- layer=2 filter=6 channel=84
					0, 4, 6, 7, 9, 0, -2, -6, -6,
					-- layer=2 filter=6 channel=85
					-9, 0, 3, -9, 0, -2, -8, 9, -10,
					-- layer=2 filter=6 channel=86
					-5, -9, -10, 0, -2, -2, -4, -11, -8,
					-- layer=2 filter=6 channel=87
					-20, 20, -17, -9, -1, -6, 12, -15, 3,
					-- layer=2 filter=6 channel=88
					-5, -8, -3, -7, -17, 1, -13, -7, -12,
					-- layer=2 filter=6 channel=89
					11, -5, -14, 0, -14, -26, -2, -5, -20,
					-- layer=2 filter=6 channel=90
					6, 0, 6, 6, -4, 1, 4, 3, -5,
					-- layer=2 filter=6 channel=91
					1, -4, -17, -2, -37, -23, -1, -6, -1,
					-- layer=2 filter=6 channel=92
					-2, 5, -9, 3, -21, -22, -10, 11, -12,
					-- layer=2 filter=6 channel=93
					-1, -7, -17, -18, 3, 0, -14, -9, -38,
					-- layer=2 filter=6 channel=94
					-8, -1, -12, -15, -16, -18, -7, -6, -8,
					-- layer=2 filter=6 channel=95
					4, -1, -10, 4, 6, 0, -2, 7, 0,
					-- layer=2 filter=6 channel=96
					-7, 6, -8, 2, 6, 2, 0, -18, -13,
					-- layer=2 filter=6 channel=97
					0, -11, 6, -9, -18, -5, -16, -27, -14,
					-- layer=2 filter=6 channel=98
					-12, -11, 0, -3, -6, -26, -1, -25, -18,
					-- layer=2 filter=6 channel=99
					14, 12, -5, -12, -27, -23, -17, -21, -10,
					-- layer=2 filter=6 channel=100
					10, -25, -2, -5, 6, 8, -5, 14, -1,
					-- layer=2 filter=6 channel=101
					-12, 0, -15, -12, -27, -2, -36, -36, -14,
					-- layer=2 filter=6 channel=102
					0, 5, -14, 0, 4, -13, 4, -6, -10,
					-- layer=2 filter=6 channel=103
					0, 19, -3, -28, -2, -3, -1, 0, -3,
					-- layer=2 filter=6 channel=104
					-16, 9, -27, 3, -5, -8, 11, -20, -23,
					-- layer=2 filter=6 channel=105
					-5, 7, 15, -16, -5, -19, -1, 0, -9,
					-- layer=2 filter=6 channel=106
					-10, -15, 1, -6, -16, -14, -18, -15, -13,
					-- layer=2 filter=6 channel=107
					6, -19, 0, 8, -19, -27, 1, -1, -12,
					-- layer=2 filter=6 channel=108
					14, -8, -34, -1, -10, -10, 13, 1, 5,
					-- layer=2 filter=6 channel=109
					-3, 9, -8, -4, -2, -9, 0, 6, -11,
					-- layer=2 filter=6 channel=110
					-14, -10, -14, -1, -33, -34, 3, -26, -26,
					-- layer=2 filter=6 channel=111
					-2, 9, 3, 2, 0, -6, 6, 1, -3,
					-- layer=2 filter=6 channel=112
					-7, -7, -17, -12, -21, -37, -25, -10, -25,
					-- layer=2 filter=6 channel=113
					-8, 3, -11, -1, -9, -8, -19, -1, 1,
					-- layer=2 filter=6 channel=114
					3, -7, -3, -5, 3, 1, 0, -8, 1,
					-- layer=2 filter=6 channel=115
					4, 1, 4, 3, 0, -1, 9, -3, -3,
					-- layer=2 filter=6 channel=116
					-7, 8, -15, 15, -2, -9, 6, -9, 0,
					-- layer=2 filter=6 channel=117
					-14, 4, 13, -7, -28, -9, -29, -19, -10,
					-- layer=2 filter=6 channel=118
					-16, -9, 2, -20, 3, 5, 7, 2, 9,
					-- layer=2 filter=6 channel=119
					-2, -16, 4, -6, 8, 2, -21, -10, 2,
					-- layer=2 filter=6 channel=120
					-9, -2, -5, 4, -5, 0, 0, -5, -6,
					-- layer=2 filter=6 channel=121
					-3, 10, 10, 4, -6, -9, -5, 8, 1,
					-- layer=2 filter=6 channel=122
					0, 1, -5, 1, 0, 10, -1, -8, 9,
					-- layer=2 filter=6 channel=123
					-3, -4, 1, -5, -1, -28, -9, -37, -5,
					-- layer=2 filter=6 channel=124
					-16, 26, -1, 6, 9, -24, 7, -6, -31,
					-- layer=2 filter=6 channel=125
					-3, 0, -2, -8, 4, -7, -7, 5, -3,
					-- layer=2 filter=6 channel=126
					13, -25, 0, -1, -12, 0, -13, -2, 0,
					-- layer=2 filter=6 channel=127
					0, -5, -7, -4, -6, -7, -1, -3, -11,
					-- layer=2 filter=7 channel=0
					0, -15, -8, 8, 13, 19, 1, -4, 1,
					-- layer=2 filter=7 channel=1
					14, 12, -9, 12, 5, -21, -3, 13, 22,
					-- layer=2 filter=7 channel=2
					-2, 5, 10, 12, 11, -6, -1, 4, 1,
					-- layer=2 filter=7 channel=3
					-13, -24, 18, -54, -4, -13, 3, 15, 3,
					-- layer=2 filter=7 channel=4
					-18, 16, 0, -36, -16, -10, 11, -2, 8,
					-- layer=2 filter=7 channel=5
					-19, -13, -31, 11, -3, 1, 4, -18, 1,
					-- layer=2 filter=7 channel=6
					13, 24, 69, 9, 2, 3, -13, -18, -36,
					-- layer=2 filter=7 channel=7
					-43, 5, 3, -45, -10, 1, 6, 57, -25,
					-- layer=2 filter=7 channel=8
					3, -9, 6, -7, 1, 2, -3, 8, 5,
					-- layer=2 filter=7 channel=9
					-39, -35, 3, -6, -18, 1, -13, -5, 20,
					-- layer=2 filter=7 channel=10
					-2, -8, 4, -17, -6, 23, -11, 6, 18,
					-- layer=2 filter=7 channel=11
					-15, -13, -21, 6, -8, -4, 1, 0, -26,
					-- layer=2 filter=7 channel=12
					10, 2, -29, -12, 2, -2, 22, 19, 19,
					-- layer=2 filter=7 channel=13
					-7, -6, -4, 6, 6, -4, 7, 6, -3,
					-- layer=2 filter=7 channel=14
					-1, 15, -8, 14, -2, -23, 7, 4, 0,
					-- layer=2 filter=7 channel=15
					-12, -11, -1, 26, 59, 20, -34, -57, -9,
					-- layer=2 filter=7 channel=16
					-28, -12, -17, -40, -36, -29, -5, 16, 7,
					-- layer=2 filter=7 channel=17
					4, -8, -3, -6, 0, 10, -6, 6, -9,
					-- layer=2 filter=7 channel=18
					-3, 5, 13, 27, 24, 12, 8, 20, 8,
					-- layer=2 filter=7 channel=19
					13, -9, -8, 23, 25, -16, 21, 20, 23,
					-- layer=2 filter=7 channel=20
					1, -1, -1, 0, -5, -7, -2, 5, -4,
					-- layer=2 filter=7 channel=21
					-3, 14, 7, 7, 5, -2, -2, 3, -7,
					-- layer=2 filter=7 channel=22
					3, -12, 1, 4, 0, 3, 2, -1, -2,
					-- layer=2 filter=7 channel=23
					-19, -6, -19, 2, -25, -21, 13, 15, 9,
					-- layer=2 filter=7 channel=24
					12, 44, 60, -41, -5, -2, -14, -2, 1,
					-- layer=2 filter=7 channel=25
					10, 44, 34, -29, -13, -15, -11, -1, -9,
					-- layer=2 filter=7 channel=26
					-2, 3, -3, -3, -8, -10, 5, 2, 0,
					-- layer=2 filter=7 channel=27
					-7, -18, -44, 6, 28, 36, -33, -12, 2,
					-- layer=2 filter=7 channel=28
					-9, -14, -5, -27, -3, 2, 16, -15, -18,
					-- layer=2 filter=7 channel=29
					-3, 2, 1, 0, -10, -1, -5, -1, 10,
					-- layer=2 filter=7 channel=30
					-4, -5, -14, 18, 6, 14, -17, -17, 15,
					-- layer=2 filter=7 channel=31
					-29, -68, -37, -23, -42, -26, -28, -54, -20,
					-- layer=2 filter=7 channel=32
					-5, 6, 9, 6, 9, -4, 10, -1, 4,
					-- layer=2 filter=7 channel=33
					-19, 11, 0, -19, 7, -6, 26, 22, -8,
					-- layer=2 filter=7 channel=34
					-6, -5, -31, -15, 18, 4, -20, 24, -10,
					-- layer=2 filter=7 channel=35
					-19, 17, -3, -30, 18, 15, 26, 14, 11,
					-- layer=2 filter=7 channel=36
					-7, 0, 4, -6, 4, -1, 8, -5, 5,
					-- layer=2 filter=7 channel=37
					14, -5, -7, 3, 10, 3, -9, -11, -10,
					-- layer=2 filter=7 channel=38
					13, -6, -21, 1, -5, 26, -42, -41, -5,
					-- layer=2 filter=7 channel=39
					-1, -24, -6, -40, -34, -13, 21, 35, 15,
					-- layer=2 filter=7 channel=40
					10, 15, -4, 29, -18, 34, -24, 34, -13,
					-- layer=2 filter=7 channel=41
					0, -8, -8, -5, -3, 2, 0, -6, 0,
					-- layer=2 filter=7 channel=42
					6, -14, -26, 3, 3, -4, 4, 21, -12,
					-- layer=2 filter=7 channel=43
					-45, -15, -9, 14, 23, 33, 0, 41, 23,
					-- layer=2 filter=7 channel=44
					3, 1, -3, 8, -1, 3, 6, -6, 0,
					-- layer=2 filter=7 channel=45
					-7, 9, 1, -3, -8, 25, -22, 2, 0,
					-- layer=2 filter=7 channel=46
					-27, -29, 6, 11, 0, 29, -25, 9, 26,
					-- layer=2 filter=7 channel=47
					-15, 25, 33, -5, -3, 31, 6, -1, -23,
					-- layer=2 filter=7 channel=48
					2, -9, -6, 8, -1, 6, 6, 3, 8,
					-- layer=2 filter=7 channel=49
					-21, 25, 29, 0, 45, 12, 8, 13, 36,
					-- layer=2 filter=7 channel=50
					-2, 18, 17, -7, 25, -1, 28, 29, 14,
					-- layer=2 filter=7 channel=51
					-15, -17, 2, -4, -3, -10, -21, -13, -26,
					-- layer=2 filter=7 channel=52
					0, -9, -1, 21, 1, -23, 17, -4, 0,
					-- layer=2 filter=7 channel=53
					0, 1, 2, 8, -3, -19, 6, -50, -19,
					-- layer=2 filter=7 channel=54
					7, 20, -1, -6, -34, -12, 19, -4, -8,
					-- layer=2 filter=7 channel=55
					8, 10, 5, -12, 11, 2, 0, -9, 3,
					-- layer=2 filter=7 channel=56
					-13, -24, -27, 9, 25, 1, 17, 1, -11,
					-- layer=2 filter=7 channel=57
					0, 9, 14, -6, 12, 16, -2, -10, 0,
					-- layer=2 filter=7 channel=58
					5, 0, -15, 18, -6, -28, 11, 24, 19,
					-- layer=2 filter=7 channel=59
					19, 27, 9, 0, 5, -5, 37, 15, 35,
					-- layer=2 filter=7 channel=60
					31, 25, 18, 23, -10, -8, -18, -7, -25,
					-- layer=2 filter=7 channel=61
					-32, 10, 17, -35, -12, -14, -9, -13, -49,
					-- layer=2 filter=7 channel=62
					18, -4, 29, 29, 14, -22, 18, 21, 4,
					-- layer=2 filter=7 channel=63
					-7, 3, 23, -3, -33, 19, 3, -23, -26,
					-- layer=2 filter=7 channel=64
					10, 21, -10, -14, -8, -1, -11, 0, 24,
					-- layer=2 filter=7 channel=65
					0, -15, 33, -20, -33, -28, -25, -18, -37,
					-- layer=2 filter=7 channel=66
					-2, -35, -37, 0, 1, 8, 23, 23, -6,
					-- layer=2 filter=7 channel=67
					-55, -58, -16, -27, -25, -13, -11, 20, 20,
					-- layer=2 filter=7 channel=68
					1, -6, -1, 1, -3, -2, 9, 8, 6,
					-- layer=2 filter=7 channel=69
					6, 8, 0, 0, -10, 2, -18, 18, 24,
					-- layer=2 filter=7 channel=70
					1, -2, -20, -7, 12, 4, 16, -3, 1,
					-- layer=2 filter=7 channel=71
					-11, -1, -42, 4, 36, 12, 8, 1, 5,
					-- layer=2 filter=7 channel=72
					-10, 12, -3, -4, -1, -13, 30, 21, -9,
					-- layer=2 filter=7 channel=73
					13, -26, -9, 41, -21, -8, -23, -14, 3,
					-- layer=2 filter=7 channel=74
					-10, -17, -2, -10, 3, 6, -17, 35, 4,
					-- layer=2 filter=7 channel=75
					2, 6, 2, 1, 28, -9, 88, 63, -4,
					-- layer=2 filter=7 channel=76
					-30, -37, -14, -4, -30, -22, 0, -56, -16,
					-- layer=2 filter=7 channel=77
					-7, -4, 4, 5, 4, 4, 0, -9, -4,
					-- layer=2 filter=7 channel=78
					-20, 8, 38, -11, -4, -7, -4, -6, 6,
					-- layer=2 filter=7 channel=79
					-9, 12, -8, 6, -8, 9, -4, -2, -5,
					-- layer=2 filter=7 channel=80
					-16, -19, 7, -24, -8, -2, -18, 33, 22,
					-- layer=2 filter=7 channel=81
					-7, -5, -9, -9, -18, -12, -13, -14, 0,
					-- layer=2 filter=7 channel=82
					0, -6, -8, -6, -9, 3, -7, -11, 0,
					-- layer=2 filter=7 channel=83
					-14, -10, 3, -2, 11, -9, -33, -4, -18,
					-- layer=2 filter=7 channel=84
					-5, 7, 4, -2, -8, -11, 1, -1, 7,
					-- layer=2 filter=7 channel=85
					-1, -6, 0, -4, 4, 0, 0, 6, 5,
					-- layer=2 filter=7 channel=86
					-5, 8, 16, -4, 14, 12, 0, -5, 7,
					-- layer=2 filter=7 channel=87
					17, 19, 1, 37, -25, -12, -16, -6, -13,
					-- layer=2 filter=7 channel=88
					-16, -24, -17, -12, -23, 7, -8, -12, -10,
					-- layer=2 filter=7 channel=89
					8, 19, 3, 15, 17, 0, 45, 40, 28,
					-- layer=2 filter=7 channel=90
					1, 8, -3, -4, -6, 6, -5, 4, -5,
					-- layer=2 filter=7 channel=91
					16, 0, -9, -8, 3, 5, 30, 13, 28,
					-- layer=2 filter=7 channel=92
					9, 38, 7, 16, 17, 13, 19, 19, 18,
					-- layer=2 filter=7 channel=93
					24, 19, 31, 0, -23, -26, 38, -10, 9,
					-- layer=2 filter=7 channel=94
					-47, -8, -7, -6, -19, -14, -10, 0, 0,
					-- layer=2 filter=7 channel=95
					4, 5, 15, 9, 0, 5, 20, 14, 0,
					-- layer=2 filter=7 channel=96
					33, 18, 9, 37, 8, 9, 26, -42, -13,
					-- layer=2 filter=7 channel=97
					-8, 12, 50, -23, 13, -2, -32, 12, 0,
					-- layer=2 filter=7 channel=98
					-5, -10, 14, -28, 8, 11, 5, 22, -16,
					-- layer=2 filter=7 channel=99
					-42, -18, -27, 8, 39, -25, 19, -34, -8,
					-- layer=2 filter=7 channel=100
					-2, -29, -49, -21, 31, 0, -9, -11, 7,
					-- layer=2 filter=7 channel=101
					-12, -12, -13, 0, -16, 2, 30, 0, 19,
					-- layer=2 filter=7 channel=102
					-7, 30, -23, -12, 16, -32, 6, -53, 1,
					-- layer=2 filter=7 channel=103
					-41, 15, 33, 8, 9, 5, -20, 7, -14,
					-- layer=2 filter=7 channel=104
					2, 6, -10, -3, 26, -12, -17, 39, 36,
					-- layer=2 filter=7 channel=105
					-59, -19, -9, -1, -39, -76, 2, 0, -18,
					-- layer=2 filter=7 channel=106
					-6, 40, 33, -24, -12, -2, -5, -17, -10,
					-- layer=2 filter=7 channel=107
					-41, 17, 18, 49, 33, 29, -16, 41, -2,
					-- layer=2 filter=7 channel=108
					2, 5, -10, 22, 32, 4, -38, -31, 8,
					-- layer=2 filter=7 channel=109
					-3, 0, 10, -9, 13, -6, -6, 4, -2,
					-- layer=2 filter=7 channel=110
					13, 16, 28, -16, 5, 33, 13, 7, -18,
					-- layer=2 filter=7 channel=111
					-1, 6, -3, 4, 11, 8, -5, 8, -2,
					-- layer=2 filter=7 channel=112
					-29, -11, -16, -31, -3, 2, -25, -8, -15,
					-- layer=2 filter=7 channel=113
					21, -24, -8, 2, -20, 10, -32, -29, 16,
					-- layer=2 filter=7 channel=114
					8, 17, 7, 0, 11, -4, 5, 3, -6,
					-- layer=2 filter=7 channel=115
					4, -4, 4, 12, 9, 6, -3, -7, -5,
					-- layer=2 filter=7 channel=116
					12, 22, -13, 22, -21, -4, -14, 0, -13,
					-- layer=2 filter=7 channel=117
					-75, -17, -27, -31, -14, 3, 38, 38, -16,
					-- layer=2 filter=7 channel=118
					-10, -15, 22, -5, 14, 24, -12, 26, 30,
					-- layer=2 filter=7 channel=119
					1, 12, 10, -29, 0, 5, 3, -1, -35,
					-- layer=2 filter=7 channel=120
					-6, 4, 8, -6, 7, 6, 4, 9, -4,
					-- layer=2 filter=7 channel=121
					10, -2, 9, -3, 1, 1, 6, 5, -5,
					-- layer=2 filter=7 channel=122
					11, 2, 10, 4, -1, 8, -12, -12, -6,
					-- layer=2 filter=7 channel=123
					-26, -1, 40, -11, -11, -8, 53, 27, 10,
					-- layer=2 filter=7 channel=124
					-43, -13, -4, -1, -5, 0, 6, 1, 22,
					-- layer=2 filter=7 channel=125
					3, 8, -8, 3, 5, 0, 5, -3, 4,
					-- layer=2 filter=7 channel=126
					24, 13, -8, -9, -46, 59, -21, -53, 28,
					-- layer=2 filter=7 channel=127
					3, 8, 13, -4, -29, -10, -17, -41, -16,
					-- layer=2 filter=8 channel=0
					-29, -22, -37, -12, -16, -23, 12, 11, 4,
					-- layer=2 filter=8 channel=1
					38, -12, -15, -42, -45, 10, -11, 0, 59,
					-- layer=2 filter=8 channel=2
					10, 1, 9, 0, 5, 4, 2, 5, -6,
					-- layer=2 filter=8 channel=3
					-28, -7, -40, 21, 14, -52, 9, -30, -45,
					-- layer=2 filter=8 channel=4
					-53, -41, 3, -31, 4, -3, 19, -21, 5,
					-- layer=2 filter=8 channel=5
					-24, -19, 1, 8, 8, -14, 8, -4, 5,
					-- layer=2 filter=8 channel=6
					5, -5, -16, 18, 7, 0, 11, -22, 26,
					-- layer=2 filter=8 channel=7
					21, 4, -32, -4, -15, 5, 7, 49, 9,
					-- layer=2 filter=8 channel=8
					2, -1, 5, 2, 8, 0, 7, 1, 6,
					-- layer=2 filter=8 channel=9
					-23, -19, -54, -9, -49, -41, 6, -26, -16,
					-- layer=2 filter=8 channel=10
					3, -10, -3, 6, 12, -33, 3, 0, -41,
					-- layer=2 filter=8 channel=11
					-31, -8, 2, 19, 5, 18, 29, -3, 16,
					-- layer=2 filter=8 channel=12
					-2, -38, -30, -78, -71, -24, 11, 14, 54,
					-- layer=2 filter=8 channel=13
					0, 2, 7, 0, 2, 0, 0, 3, -2,
					-- layer=2 filter=8 channel=14
					-5, -34, -17, -32, -42, -17, -7, -7, 31,
					-- layer=2 filter=8 channel=15
					-12, 34, -5, 4, -6, -6, 11, -24, -8,
					-- layer=2 filter=8 channel=16
					3, 15, 5, -38, 23, 10, -11, 13, -83,
					-- layer=2 filter=8 channel=17
					2, 3, 8, 4, -10, -6, 7, -2, -5,
					-- layer=2 filter=8 channel=18
					-13, -72, 8, -5, -5, -3, 31, 13, -5,
					-- layer=2 filter=8 channel=19
					24, 28, -15, 3, 1, 21, -3, 6, 10,
					-- layer=2 filter=8 channel=20
					5, -9, 5, -3, 2, 4, -8, -7, -7,
					-- layer=2 filter=8 channel=21
					-5, 0, 8, 6, -4, 3, 8, -3, -8,
					-- layer=2 filter=8 channel=22
					-10, 10, 2, -3, -1, 4, -6, 4, 8,
					-- layer=2 filter=8 channel=23
					-32, -25, -4, -7, 34, 0, -53, -15, -6,
					-- layer=2 filter=8 channel=24
					-20, -41, 2, 1, -21, -18, 17, -17, -23,
					-- layer=2 filter=8 channel=25
					-33, -40, 10, -23, -24, -4, 17, 18, 1,
					-- layer=2 filter=8 channel=26
					4, 3, -5, -7, 10, 1, -9, 0, 5,
					-- layer=2 filter=8 channel=27
					8, -2, -27, 24, -4, -11, 23, -7, -24,
					-- layer=2 filter=8 channel=28
					-5, -14, -17, -25, 10, -38, -3, 14, 9,
					-- layer=2 filter=8 channel=29
					-7, -7, -1, -11, -6, 7, -3, -1, -8,
					-- layer=2 filter=8 channel=30
					-43, -64, 11, -50, -65, -6, 7, 10, 17,
					-- layer=2 filter=8 channel=31
					-26, 11, -16, -55, 29, 11, -1, 26, -41,
					-- layer=2 filter=8 channel=32
					-5, -5, -1, 6, -3, -1, -8, 9, -6,
					-- layer=2 filter=8 channel=33
					-13, 10, -28, -11, -6, -14, 32, 16, -9,
					-- layer=2 filter=8 channel=34
					9, -36, 14, -50, 31, 49, -10, 62, -17,
					-- layer=2 filter=8 channel=35
					-14, -30, -19, -21, -20, -9, 10, 7, 22,
					-- layer=2 filter=8 channel=36
					3, 1, -9, 6, 3, -6, 6, 0, -6,
					-- layer=2 filter=8 channel=37
					-14, 0, 11, 2, -1, 16, 11, -19, -14,
					-- layer=2 filter=8 channel=38
					-15, 11, -62, -10, -14, -23, -30, -17, -19,
					-- layer=2 filter=8 channel=39
					2, -31, 8, 17, 10, -30, 2, -39, -50,
					-- layer=2 filter=8 channel=40
					-23, -8, 25, -24, -18, 9, 15, 32, -6,
					-- layer=2 filter=8 channel=41
					3, -6, -2, 8, -5, 10, -7, 4, -9,
					-- layer=2 filter=8 channel=42
					-42, -11, -47, -36, -16, -87, -26, -5, -7,
					-- layer=2 filter=8 channel=43
					-47, -87, 0, -17, 13, -14, -5, -18, -35,
					-- layer=2 filter=8 channel=44
					-8, -3, 11, 9, -7, -8, 8, 4, 7,
					-- layer=2 filter=8 channel=45
					-2, -21, -70, -2, 3, 9, 45, 42, 13,
					-- layer=2 filter=8 channel=46
					-24, -47, -34, -32, -43, -25, 13, -41, -25,
					-- layer=2 filter=8 channel=47
					-25, -36, 0, -8, 18, -2, 25, 46, -10,
					-- layer=2 filter=8 channel=48
					3, -4, -7, 2, -5, -8, -9, 2, -6,
					-- layer=2 filter=8 channel=49
					9, -49, 13, 21, -48, -1, 37, 7, 2,
					-- layer=2 filter=8 channel=50
					-16, 0, 17, 3, -5, 9, -9, -13, 4,
					-- layer=2 filter=8 channel=51
					-34, -26, 17, -12, -1, 23, 4, 12, 26,
					-- layer=2 filter=8 channel=52
					1, -21, 21, 3, 3, 28, 28, 0, 47,
					-- layer=2 filter=8 channel=53
					-21, -16, -23, -34, -66, 8, 13, -33, 33,
					-- layer=2 filter=8 channel=54
					3, 7, -1, 17, -10, 57, -6, 11, 36,
					-- layer=2 filter=8 channel=55
					8, -11, 7, 0, 9, -4, 5, 4, -3,
					-- layer=2 filter=8 channel=56
					-34, -36, 11, 11, -11, 15, 28, -20, 14,
					-- layer=2 filter=8 channel=57
					0, -9, 11, -2, -1, 4, -7, -3, 4,
					-- layer=2 filter=8 channel=58
					-11, -17, -26, -50, -48, -7, -5, -32, 35,
					-- layer=2 filter=8 channel=59
					27, -3, -61, -21, -19, -29, 14, -72, -23,
					-- layer=2 filter=8 channel=60
					8, -8, -15, 15, -23, -30, -70, 12, -21,
					-- layer=2 filter=8 channel=61
					-19, -11, -12, 34, -23, -35, -17, 29, -25,
					-- layer=2 filter=8 channel=62
					10, -1, -34, 30, 19, 11, 22, -6, 2,
					-- layer=2 filter=8 channel=63
					-15, -55, -6, 6, -49, -24, -41, -21, -53,
					-- layer=2 filter=8 channel=64
					-36, -9, -9, -14, 20, -7, -17, 5, -13,
					-- layer=2 filter=8 channel=65
					-17, 15, -52, 17, 6, 19, 10, 24, -1,
					-- layer=2 filter=8 channel=66
					30, -19, -50, -19, 12, 6, 13, -13, -7,
					-- layer=2 filter=8 channel=67
					-9, -7, -21, -18, -30, -46, -12, -23, 4,
					-- layer=2 filter=8 channel=68
					3, 3, -1, -11, -3, 4, 6, 2, 1,
					-- layer=2 filter=8 channel=69
					-25, 0, -35, -14, 27, -29, -6, -15, -47,
					-- layer=2 filter=8 channel=70
					-11, -7, -3, -33, -21, -18, 17, 12, 13,
					-- layer=2 filter=8 channel=71
					30, -12, -4, 16, -30, -10, 19, 31, 10,
					-- layer=2 filter=8 channel=72
					1, 17, -7, -8, -5, 14, -34, 21, 0,
					-- layer=2 filter=8 channel=73
					-42, 0, 2, -37, 4, -12, 3, -27, -18,
					-- layer=2 filter=8 channel=74
					13, 6, -48, -5, -41, -15, -42, -40, -25,
					-- layer=2 filter=8 channel=75
					46, 31, -43, -68, 2, -65, -50, -48, 8,
					-- layer=2 filter=8 channel=76
					-75, -24, -38, -41, 36, 26, 42, -14, 19,
					-- layer=2 filter=8 channel=77
					-2, 2, 2, -6, 6, -1, -4, 8, 2,
					-- layer=2 filter=8 channel=78
					4, -24, 3, 26, 28, 15, 18, -13, -7,
					-- layer=2 filter=8 channel=79
					-9, 11, 5, 4, 3, 0, -5, 0, 0,
					-- layer=2 filter=8 channel=80
					-37, 11, -2, -25, 35, -22, 27, 6, -89,
					-- layer=2 filter=8 channel=81
					3, 9, -3, -4, -1, 1, -3, 0, -11,
					-- layer=2 filter=8 channel=82
					4, 6, -4, 2, 3, -1, -4, -6, -2,
					-- layer=2 filter=8 channel=83
					-46, -47, -27, -53, -29, -61, 4, 21, -12,
					-- layer=2 filter=8 channel=84
					2, -9, -7, 8, 7, 7, -3, -5, 1,
					-- layer=2 filter=8 channel=85
					-4, 9, 0, 5, -2, -2, 9, 8, 5,
					-- layer=2 filter=8 channel=86
					11, 0, 2, 11, -8, -10, -5, -6, 0,
					-- layer=2 filter=8 channel=87
					-1, 2, -55, -24, -18, 10, 50, -14, 38,
					-- layer=2 filter=8 channel=88
					-29, -63, -58, -30, -26, -25, -27, -37, 3,
					-- layer=2 filter=8 channel=89
					-8, -4, -35, -41, -28, -20, 4, -29, 46,
					-- layer=2 filter=8 channel=90
					3, 3, 0, -1, -6, -9, 5, -1, 4,
					-- layer=2 filter=8 channel=91
					9, 23, -14, -63, -40, -40, -31, -37, -23,
					-- layer=2 filter=8 channel=92
					20, 0, -38, -36, -52, -41, -19, 1, 48,
					-- layer=2 filter=8 channel=93
					38, 3, -55, 32, 6, -10, 1, 35, -37,
					-- layer=2 filter=8 channel=94
					-6, -32, -18, 65, -19, 11, -15, -10, 5,
					-- layer=2 filter=8 channel=95
					-1, 1, 5, 3, 0, 0, -4, -1, -8,
					-- layer=2 filter=8 channel=96
					3, -26, -9, -5, -59, 5, -39, -57, 52,
					-- layer=2 filter=8 channel=97
					-24, 0, -17, 5, 23, -1, 44, 11, -51,
					-- layer=2 filter=8 channel=98
					-2, -23, 15, -2, 21, 15, 0, 34, -12,
					-- layer=2 filter=8 channel=99
					4, 14, 4, 20, 22, 34, 25, 7, 4,
					-- layer=2 filter=8 channel=100
					16, 5, -60, -35, -30, -58, -28, -39, -47,
					-- layer=2 filter=8 channel=101
					38, -8, 14, -3, -36, -19, 31, 14, 19,
					-- layer=2 filter=8 channel=102
					-26, -27, 18, -10, -44, 2, 1, -19, 31,
					-- layer=2 filter=8 channel=103
					0, 12, 33, 34, 16, 16, 3, -8, 33,
					-- layer=2 filter=8 channel=104
					-14, -49, -15, -7, -29, 20, 11, -17, 22,
					-- layer=2 filter=8 channel=105
					-49, -21, -25, 32, 4, -27, 44, 8, -7,
					-- layer=2 filter=8 channel=106
					-5, 0, -7, -39, -15, -53, 27, 19, -7,
					-- layer=2 filter=8 channel=107
					-4, 4, -36, 19, 29, -17, 20, 8, 15,
					-- layer=2 filter=8 channel=108
					21, -41, 0, -3, -56, -12, 9, -1, 10,
					-- layer=2 filter=8 channel=109
					-10, -6, -5, 6, 9, -9, 4, 3, 11,
					-- layer=2 filter=8 channel=110
					-14, -24, 24, -48, -17, -23, -17, 30, 7,
					-- layer=2 filter=8 channel=111
					5, -3, -12, -3, 6, -6, -8, -7, -6,
					-- layer=2 filter=8 channel=112
					-29, -53, -38, 43, -7, -9, 42, 35, -37,
					-- layer=2 filter=8 channel=113
					-27, -48, -9, -27, -60, 8, 3, -14, -8,
					-- layer=2 filter=8 channel=114
					3, 6, 10, 9, -6, -11, -9, -10, 10,
					-- layer=2 filter=8 channel=115
					5, 6, 10, 2, 2, 7, -8, 8, 8,
					-- layer=2 filter=8 channel=116
					-14, -2, -21, -22, -44, 1, 20, -13, 36,
					-- layer=2 filter=8 channel=117
					-9, -17, 18, 11, -11, 36, -9, 73, 18,
					-- layer=2 filter=8 channel=118
					-30, -9, -19, 21, 23, -1, 37, -9, -19,
					-- layer=2 filter=8 channel=119
					-5, -27, -16, 12, 1, -17, 45, 11, 30,
					-- layer=2 filter=8 channel=120
					2, 3, -9, -9, 9, 6, -4, -6, 0,
					-- layer=2 filter=8 channel=121
					0, -6, -12, -3, 0, 3, 1, -5, 1,
					-- layer=2 filter=8 channel=122
					10, -3, -1, 9, -1, -8, 5, -8, -7,
					-- layer=2 filter=8 channel=123
					11, 24, -6, -20, 21, 37, 6, 37, -36,
					-- layer=2 filter=8 channel=124
					-7, 1, -21, -19, 60, 7, 59, 21, -14,
					-- layer=2 filter=8 channel=125
					-10, 1, 10, -9, 10, 1, 1, -6, 3,
					-- layer=2 filter=8 channel=126
					7, -18, 15, -23, -36, -52, -49, -27, -15,
					-- layer=2 filter=8 channel=127
					6, -41, -35, -57, -58, -35, 42, -25, 1,
					-- layer=2 filter=9 channel=0
					2, -16, -9, 3, -4, -21, -7, -4, -5,
					-- layer=2 filter=9 channel=1
					0, 22, 14, 5, 3, 11, 9, -16, 19,
					-- layer=2 filter=9 channel=2
					2, -2, 7, -6, -7, 0, -10, -5, 1,
					-- layer=2 filter=9 channel=3
					19, -6, -53, 16, 17, -10, -19, -3, -26,
					-- layer=2 filter=9 channel=4
					-50, -50, -7, -38, -40, -25, -58, -61, 0,
					-- layer=2 filter=9 channel=5
					0, -26, 9, 6, -11, -18, -2, -5, 3,
					-- layer=2 filter=9 channel=6
					7, 14, 23, 2, -22, -42, 7, 8, 17,
					-- layer=2 filter=9 channel=7
					30, 32, 11, -9, 16, -23, -33, -16, -17,
					-- layer=2 filter=9 channel=8
					-5, -2, 6, 7, 1, -5, -3, -3, -4,
					-- layer=2 filter=9 channel=9
					-25, -32, -65, -63, -71, -65, -80, -44, -51,
					-- layer=2 filter=9 channel=10
					2, -20, -61, -9, -5, -13, -28, -12, -47,
					-- layer=2 filter=9 channel=11
					-3, -7, 14, 8, 0, -3, 21, 16, 23,
					-- layer=2 filter=9 channel=12
					3, 15, -11, -23, 1, 0, 6, 5, 2,
					-- layer=2 filter=9 channel=13
					0, -2, 6, 4, -8, -4, -4, 4, 6,
					-- layer=2 filter=9 channel=14
					14, 12, 10, 14, 5, 5, 25, -3, 30,
					-- layer=2 filter=9 channel=15
					6, 19, 0, 10, 7, -1, -15, 18, -13,
					-- layer=2 filter=9 channel=16
					-8, 34, 2, 74, 58, 24, -33, -15, -9,
					-- layer=2 filter=9 channel=17
					6, 6, 10, 3, 8, -2, -4, -11, 5,
					-- layer=2 filter=9 channel=18
					0, -15, 3, 27, -40, -34, -14, -18, 6,
					-- layer=2 filter=9 channel=19
					9, 7, 45, 26, 28, 10, 9, -12, 9,
					-- layer=2 filter=9 channel=20
					9, -3, 5, -4, -5, -4, 8, -4, -3,
					-- layer=2 filter=9 channel=21
					1, 1, -4, -7, -3, -13, -24, -16, -7,
					-- layer=2 filter=9 channel=22
					0, -1, 4, 5, -3, 5, 8, 7, 0,
					-- layer=2 filter=9 channel=23
					-71, -16, -50, -17, -12, -3, -29, -68, -43,
					-- layer=2 filter=9 channel=24
					-35, -73, -63, -13, 5, -3, -8, 4, 19,
					-- layer=2 filter=9 channel=25
					-10, -38, -29, -5, 25, 17, 22, 44, 30,
					-- layer=2 filter=9 channel=26
					2, 7, -6, 6, -10, -8, -9, -5, -3,
					-- layer=2 filter=9 channel=27
					18, -5, 21, 19, 15, 23, 0, -6, 16,
					-- layer=2 filter=9 channel=28
					0, 3, -17, 32, 41, 1, -35, 1, -51,
					-- layer=2 filter=9 channel=29
					6, -11, -2, 7, 5, 0, -10, 0, 6,
					-- layer=2 filter=9 channel=30
					-33, -19, 1, 18, -30, -40, -70, -31, -55,
					-- layer=2 filter=9 channel=31
					-16, 14, 12, 27, -5, -7, -25, -11, -24,
					-- layer=2 filter=9 channel=32
					-6, -6, -2, 8, 7, -1, 10, 1, -7,
					-- layer=2 filter=9 channel=33
					9, 9, 8, -21, -10, -34, 22, 12, -27,
					-- layer=2 filter=9 channel=34
					-8, 16, 15, 53, -12, 16, 15, 10, 44,
					-- layer=2 filter=9 channel=35
					-4, 3, -17, 47, 28, 14, -16, -14, -32,
					-- layer=2 filter=9 channel=36
					10, 2, -11, 5, -2, 1, -4, 2, -11,
					-- layer=2 filter=9 channel=37
					3, -11, 2, 16, -16, 0, 12, -3, 19,
					-- layer=2 filter=9 channel=38
					4, 8, 18, 13, 1, 33, -12, -15, 25,
					-- layer=2 filter=9 channel=39
					-15, -30, -50, 10, -8, -45, -26, -19, -62,
					-- layer=2 filter=9 channel=40
					35, 13, -10, 13, -9, -32, -16, 46, 42,
					-- layer=2 filter=9 channel=41
					8, 0, 3, 0, 6, 0, -5, 3, -9,
					-- layer=2 filter=9 channel=42
					18, 21, -39, 3, 5, 8, -24, 2, -14,
					-- layer=2 filter=9 channel=43
					-29, -39, -15, -7, -20, -20, -37, -24, -21,
					-- layer=2 filter=9 channel=44
					-7, 1, 4, 4, 6, -1, -8, -2, -9,
					-- layer=2 filter=9 channel=45
					-9, 12, -1, -1, -43, -10, 15, -20, -6,
					-- layer=2 filter=9 channel=46
					1, -34, -19, -27, -42, -41, -46, -3, -55,
					-- layer=2 filter=9 channel=47
					17, 35, 8, 1, 11, 25, 1, -8, -38,
					-- layer=2 filter=9 channel=48
					0, 7, 2, 1, 0, 2, 11, -6, 4,
					-- layer=2 filter=9 channel=49
					19, 17, 42, 5, -37, -3, 0, 6, -29,
					-- layer=2 filter=9 channel=50
					-22, -15, -14, -4, -14, -10, 6, 0, 10,
					-- layer=2 filter=9 channel=51
					-13, -6, -1, 4, -8, 5, 14, 13, 20,
					-- layer=2 filter=9 channel=52
					4, 15, 36, 7, -5, -5, -6, 10, 14,
					-- layer=2 filter=9 channel=53
					-32, 71, 4, 9, -18, 27, -26, 7, 2,
					-- layer=2 filter=9 channel=54
					0, 27, 25, 13, 11, 0, 16, 17, 12,
					-- layer=2 filter=9 channel=55
					8, 7, 0, 12, -4, -8, -1, 3, 9,
					-- layer=2 filter=9 channel=56
					2, 0, -10, 27, 9, -3, 11, 4, 12,
					-- layer=2 filter=9 channel=57
					3, 10, 1, -7, -1, -2, -7, -3, 5,
					-- layer=2 filter=9 channel=58
					11, 39, 11, 4, 10, -3, 11, -22, 27,
					-- layer=2 filter=9 channel=59
					5, 32, 5, 16, 8, 12, 18, 16, 37,
					-- layer=2 filter=9 channel=60
					-13, -40, 0, 5, 0, -12, 15, 6, 44,
					-- layer=2 filter=9 channel=61
					0, 1, 3, 12, -31, -26, 0, -14, 7,
					-- layer=2 filter=9 channel=62
					-8, 3, 19, 15, -35, -15, 20, -6, 12,
					-- layer=2 filter=9 channel=63
					-50, -14, -107, 1, -12, -84, -59, -48, -89,
					-- layer=2 filter=9 channel=64
					11, 4, -41, 28, 26, 21, 26, 24, 33,
					-- layer=2 filter=9 channel=65
					-29, -7, 32, -21, -30, -49, -16, -12, -15,
					-- layer=2 filter=9 channel=66
					18, 11, 12, -39, -8, 1, 3, 34, -23,
					-- layer=2 filter=9 channel=67
					-25, -88, -48, -22, -3, -51, -59, -62, -44,
					-- layer=2 filter=9 channel=68
					1, 7, -11, 7, 5, 7, 2, -10, -4,
					-- layer=2 filter=9 channel=69
					37, 16, -46, 38, 8, 18, 48, 30, 44,
					-- layer=2 filter=9 channel=70
					8, 4, -19, 11, 6, 2, -14, -14, -25,
					-- layer=2 filter=9 channel=71
					12, -16, -2, 25, 26, 38, 15, 13, 49,
					-- layer=2 filter=9 channel=72
					14, 11, 6, 24, 47, -23, 9, 29, 0,
					-- layer=2 filter=9 channel=73
					26, 52, 46, 42, 6, 2, -2, 15, -30,
					-- layer=2 filter=9 channel=74
					-4, -34, -62, 49, -40, -44, -19, -53, -30,
					-- layer=2 filter=9 channel=75
					23, -2, 1, 32, 11, -16, -28, 20, 14,
					-- layer=2 filter=9 channel=76
					16, 56, 17, -1, 21, 24, -33, -10, 13,
					-- layer=2 filter=9 channel=77
					-4, 7, -6, 6, -11, 0, 6, -8, 6,
					-- layer=2 filter=9 channel=78
					-20, -29, 18, 6, -4, -11, 10, 15, 31,
					-- layer=2 filter=9 channel=79
					4, 4, -1, -6, -5, 0, 1, 2, -5,
					-- layer=2 filter=9 channel=80
					-47, -36, -42, -20, 0, -18, -81, -96, -17,
					-- layer=2 filter=9 channel=81
					-4, 0, 8, 9, 13, 12, 3, 7, 6,
					-- layer=2 filter=9 channel=82
					-9, -5, 4, 10, 2, 10, -13, 0, 6,
					-- layer=2 filter=9 channel=83
					-60, -73, -25, -19, -24, 4, -51, -50, -28,
					-- layer=2 filter=9 channel=84
					6, -2, 7, -11, 3, 8, -1, -11, 2,
					-- layer=2 filter=9 channel=85
					7, 0, -1, 5, -14, -16, 4, -4, -8,
					-- layer=2 filter=9 channel=86
					1, -2, 9, 5, -10, -2, 2, -11, 6,
					-- layer=2 filter=9 channel=87
					-40, 24, 3, 9, 0, 5, -11, 6, 25,
					-- layer=2 filter=9 channel=88
					-33, -28, -28, -5, -26, -37, -10, -5, -12,
					-- layer=2 filter=9 channel=89
					24, 6, 20, -14, 18, -6, 8, 13, 25,
					-- layer=2 filter=9 channel=90
					0, 7, -4, 7, -8, 0, 0, 3, 5,
					-- layer=2 filter=9 channel=91
					26, 20, 0, -13, 31, -7, 2, 2, 34,
					-- layer=2 filter=9 channel=92
					-5, 18, 6, -6, 19, 4, 35, 5, 21,
					-- layer=2 filter=9 channel=93
					-5, 13, 44, -24, -7, -32, 12, -52, -32,
					-- layer=2 filter=9 channel=94
					-7, 30, 45, -13, -7, -51, -33, -30, 17,
					-- layer=2 filter=9 channel=95
					9, -23, -5, 1, -6, 1, 2, -2, 2,
					-- layer=2 filter=9 channel=96
					-49, -34, 22, -26, 14, 19, -12, -44, -14,
					-- layer=2 filter=9 channel=97
					-34, -85, -80, -48, -12, -61, -57, -42, -43,
					-- layer=2 filter=9 channel=98
					12, 37, -6, 31, 32, 24, 14, 9, 7,
					-- layer=2 filter=9 channel=99
					14, 24, 35, -9, -21, -2, 23, -7, 28,
					-- layer=2 filter=9 channel=100
					-15, -26, 15, -60, -13, -21, -36, -55, -27,
					-- layer=2 filter=9 channel=101
					17, -18, -30, 36, 21, 35, 24, 33, 26,
					-- layer=2 filter=9 channel=102
					-42, -45, 18, -16, -14, -24, -35, -69, -33,
					-- layer=2 filter=9 channel=103
					16, 11, -21, 11, -49, 48, 66, -2, -9,
					-- layer=2 filter=9 channel=104
					-25, -5, 16, 35, 2, 0, -14, -29, 6,
					-- layer=2 filter=9 channel=105
					-52, 39, 59, -4, 73, 46, 21, -12, 7,
					-- layer=2 filter=9 channel=106
					-15, -32, -26, 11, 29, 14, 25, 15, 46,
					-- layer=2 filter=9 channel=107
					-17, 7, -52, 17, 8, -3, 19, -3, -32,
					-- layer=2 filter=9 channel=108
					-1, -18, 22, 10, -2, 24, -15, -31, 25,
					-- layer=2 filter=9 channel=109
					-5, 5, -9, -5, -4, 0, -25, 4, -3,
					-- layer=2 filter=9 channel=110
					-22, 12, -36, 6, 12, 24, -27, 11, -2,
					-- layer=2 filter=9 channel=111
					-7, -3, -9, 8, 9, 6, -8, -2, 0,
					-- layer=2 filter=9 channel=112
					-19, -13, -29, 11, 24, 11, 24, 19, 5,
					-- layer=2 filter=9 channel=113
					-55, -30, -45, 19, -74, -39, -63, -19, -77,
					-- layer=2 filter=9 channel=114
					25, 15, 14, 5, 10, 3, 19, 10, 2,
					-- layer=2 filter=9 channel=115
					-5, 1, -6, 5, 3, -7, 1, -2, -3,
					-- layer=2 filter=9 channel=116
					-22, 21, -10, 3, 9, -1, -21, 7, -1,
					-- layer=2 filter=9 channel=117
					40, 61, 38, 8, 29, 49, 15, 7, -5,
					-- layer=2 filter=9 channel=118
					-25, -29, -6, -15, -19, -9, -26, 9, -22,
					-- layer=2 filter=9 channel=119
					-30, -33, -20, -52, -86, -45, -26, -78, -44,
					-- layer=2 filter=9 channel=120
					-10, -9, 7, 2, -5, 3, 4, -8, -3,
					-- layer=2 filter=9 channel=121
					10, 0, 5, 6, 4, -10, 0, 0, 9,
					-- layer=2 filter=9 channel=122
					9, 9, -7, 7, 5, 3, 0, 3, 3,
					-- layer=2 filter=9 channel=123
					6, 26, 12, -3, 27, 2, -12, 5, -33,
					-- layer=2 filter=9 channel=124
					-13, 0, 19, 22, 21, -6, -32, -2, -17,
					-- layer=2 filter=9 channel=125
					5, -8, -7, -9, 1, 2, -4, -7, 6,
					-- layer=2 filter=9 channel=126
					12, -44, -54, -17, -4, -80, -9, -61, -33,
					-- layer=2 filter=9 channel=127
					-33, -26, -11, -2, -14, -31, -24, -57, -16,
					-- layer=2 filter=10 channel=0
					2, 1, -11, -8, 2, 3, -7, -1, 3,
					-- layer=2 filter=10 channel=1
					0, -9, -11, -14, -13, 0, -7, 3, -15,
					-- layer=2 filter=10 channel=2
					-2, 4, 5, 2, -10, -8, 0, 0, 7,
					-- layer=2 filter=10 channel=3
					3, -9, 7, 0, -9, -1, 6, -12, -9,
					-- layer=2 filter=10 channel=4
					-2, 2, 6, 0, -7, 5, -11, -2, 0,
					-- layer=2 filter=10 channel=5
					-1, 7, 5, -5, 1, 5, 0, -10, -6,
					-- layer=2 filter=10 channel=6
					-2, -8, -5, -12, -4, 0, 1, 2, -6,
					-- layer=2 filter=10 channel=7
					-4, -4, -2, -4, -5, -10, -3, -7, -5,
					-- layer=2 filter=10 channel=8
					-3, -6, 1, 4, -1, 7, 2, -5, -7,
					-- layer=2 filter=10 channel=9
					2, -9, -10, 2, -11, -4, 1, -4, -1,
					-- layer=2 filter=10 channel=10
					-6, -9, -12, 9, -7, 6, -8, 2, 0,
					-- layer=2 filter=10 channel=11
					-9, -12, 1, -10, -4, -12, -1, -3, -8,
					-- layer=2 filter=10 channel=12
					-7, -2, -6, 1, -13, -4, -9, 1, 0,
					-- layer=2 filter=10 channel=13
					3, -1, 7, 1, 3, -2, -8, 0, 7,
					-- layer=2 filter=10 channel=14
					6, -12, 2, -11, -12, -8, -8, 5, -4,
					-- layer=2 filter=10 channel=15
					-8, -13, 7, 7, 2, 7, -4, 0, -12,
					-- layer=2 filter=10 channel=16
					4, 3, 6, 5, -3, -11, -5, 0, 0,
					-- layer=2 filter=10 channel=17
					-8, 5, 4, 5, -9, 0, 3, 8, -8,
					-- layer=2 filter=10 channel=18
					0, -13, -8, -10, -1, 5, 0, -16, -4,
					-- layer=2 filter=10 channel=19
					-17, 2, 4, -5, -20, 0, -7, -1, -1,
					-- layer=2 filter=10 channel=20
					-2, 9, -8, -4, 5, 9, 3, -2, 7,
					-- layer=2 filter=10 channel=21
					4, -10, 3, 5, -12, 0, -7, 4, 8,
					-- layer=2 filter=10 channel=22
					-2, 6, -5, 3, 8, -1, 4, -9, 9,
					-- layer=2 filter=10 channel=23
					-1, 2, -4, 3, -2, 0, -3, -3, 6,
					-- layer=2 filter=10 channel=24
					5, 0, -5, 6, -4, 7, -6, 4, -7,
					-- layer=2 filter=10 channel=25
					1, -15, 2, -5, -5, 0, -9, 7, -8,
					-- layer=2 filter=10 channel=26
					9, 7, 5, -2, 1, -1, 8, -6, -7,
					-- layer=2 filter=10 channel=27
					-5, 0, -8, -11, -5, -3, 0, -2, -3,
					-- layer=2 filter=10 channel=28
					2, -8, -17, -7, -14, 6, -1, 2, -4,
					-- layer=2 filter=10 channel=29
					-5, -7, 7, 7, 6, -3, -9, -8, -2,
					-- layer=2 filter=10 channel=30
					5, -5, 0, -10, 0, 3, -2, 4, -9,
					-- layer=2 filter=10 channel=31
					1, 2, -2, -12, -7, 7, -1, -11, -5,
					-- layer=2 filter=10 channel=32
					1, -1, -8, 6, 2, -2, -8, -9, -8,
					-- layer=2 filter=10 channel=33
					-2, -11, 0, -10, -4, -3, -1, -3, 6,
					-- layer=2 filter=10 channel=34
					0, -13, 1, 8, -5, -5, -8, 0, -8,
					-- layer=2 filter=10 channel=35
					0, -1, -4, -7, -2, 3, 7, -11, -11,
					-- layer=2 filter=10 channel=36
					-6, 0, -6, -11, 2, -4, -7, 2, -11,
					-- layer=2 filter=10 channel=37
					-7, 4, -16, -11, -10, -12, -19, -15, -12,
					-- layer=2 filter=10 channel=38
					-12, -11, 0, 1, -4, 5, -1, -6, 2,
					-- layer=2 filter=10 channel=39
					7, -5, 9, -8, -10, 0, -1, -1, 3,
					-- layer=2 filter=10 channel=40
					-6, -1, 0, -7, -1, -11, -6, 0, -8,
					-- layer=2 filter=10 channel=41
					12, -4, -11, 10, 0, -10, 3, -7, -1,
					-- layer=2 filter=10 channel=42
					0, 5, -7, 6, 10, 0, 3, -5, 0,
					-- layer=2 filter=10 channel=43
					4, -5, 3, 2, 8, -3, -9, -12, 7,
					-- layer=2 filter=10 channel=44
					-5, 9, 10, 0, -7, 3, 7, -9, 0,
					-- layer=2 filter=10 channel=45
					-10, -4, 7, -3, -7, -1, 5, -7, -7,
					-- layer=2 filter=10 channel=46
					0, -5, 5, 4, 6, -6, -7, 4, 5,
					-- layer=2 filter=10 channel=47
					-8, 3, 3, 1, -5, -1, -5, -5, -5,
					-- layer=2 filter=10 channel=48
					-9, 0, 2, -6, 11, -1, -8, 1, -2,
					-- layer=2 filter=10 channel=49
					-8, -7, -4, -12, -9, 0, -8, -11, 8,
					-- layer=2 filter=10 channel=50
					-9, 0, 2, -4, -8, 3, -8, 7, 0,
					-- layer=2 filter=10 channel=51
					-15, -4, -3, 4, -6, -6, -11, -1, -2,
					-- layer=2 filter=10 channel=52
					3, 0, -6, -14, -6, -16, -2, -14, -18,
					-- layer=2 filter=10 channel=53
					6, 9, 1, -4, 3, 6, -9, 3, 4,
					-- layer=2 filter=10 channel=54
					-8, -4, -8, -10, -9, -14, 0, -1, -7,
					-- layer=2 filter=10 channel=55
					0, 3, -5, -1, -6, -2, 2, -6, 6,
					-- layer=2 filter=10 channel=56
					5, -7, -13, 7, -7, -14, -13, 0, -10,
					-- layer=2 filter=10 channel=57
					-7, 6, 10, 3, 6, -1, -4, 7, 4,
					-- layer=2 filter=10 channel=58
					-5, -3, -1, -6, -6, -14, -12, 4, -3,
					-- layer=2 filter=10 channel=59
					-13, -4, 4, -11, -5, -1, 2, -17, -12,
					-- layer=2 filter=10 channel=60
					0, -9, 3, 0, -1, -5, -4, -8, -18,
					-- layer=2 filter=10 channel=61
					-13, 8, -12, -3, 0, 0, -15, -7, -4,
					-- layer=2 filter=10 channel=62
					-2, -7, -1, 0, -11, -2, -6, 0, -5,
					-- layer=2 filter=10 channel=63
					3, -3, -7, 0, 6, -4, 3, 5, -10,
					-- layer=2 filter=10 channel=64
					3, 4, -8, -9, -10, -1, 1, -4, -4,
					-- layer=2 filter=10 channel=65
					2, 4, -9, -15, -8, -9, 1, -4, 1,
					-- layer=2 filter=10 channel=66
					-10, -8, 6, 6, 5, -10, 7, 1, -3,
					-- layer=2 filter=10 channel=67
					-5, 3, -1, 2, -4, -4, 5, -5, -4,
					-- layer=2 filter=10 channel=68
					-9, 3, 1, -8, -7, 7, 3, -7, -9,
					-- layer=2 filter=10 channel=69
					8, -7, 5, -1, -9, -9, -1, -10, 1,
					-- layer=2 filter=10 channel=70
					0, -4, -6, -6, -14, -8, 3, 1, -9,
					-- layer=2 filter=10 channel=71
					6, -9, -6, -7, 0, -3, 5, 1, -7,
					-- layer=2 filter=10 channel=72
					-7, -10, 7, -6, -11, 3, -3, 1, -8,
					-- layer=2 filter=10 channel=73
					0, -5, 0, 2, -13, 6, 4, 1, -6,
					-- layer=2 filter=10 channel=74
					-11, -2, 0, 2, 5, -5, -9, 6, 4,
					-- layer=2 filter=10 channel=75
					-6, -4, 6, -2, -6, -1, 5, 4, 1,
					-- layer=2 filter=10 channel=76
					7, 2, -8, -8, 8, 2, 5, 2, -4,
					-- layer=2 filter=10 channel=77
					3, -10, 1, -6, -1, -1, -8, 7, 0,
					-- layer=2 filter=10 channel=78
					-10, -1, -7, -11, 1, -7, -14, -7, 1,
					-- layer=2 filter=10 channel=79
					2, -1, -6, 0, -5, -11, -9, -3, 0,
					-- layer=2 filter=10 channel=80
					-9, -11, 1, -3, -2, -5, -12, -10, 1,
					-- layer=2 filter=10 channel=81
					0, 6, -2, 1, -9, -8, 6, 4, -2,
					-- layer=2 filter=10 channel=82
					-10, -10, 8, 3, 3, 8, 3, -11, 8,
					-- layer=2 filter=10 channel=83
					0, -7, 0, -8, -8, 2, 1, 0, -4,
					-- layer=2 filter=10 channel=84
					-11, -11, 4, 1, 7, 5, 1, -9, 7,
					-- layer=2 filter=10 channel=85
					-10, -10, -7, -3, 6, -2, -8, -7, -3,
					-- layer=2 filter=10 channel=86
					0, -9, 2, 2, -6, -1, 9, 7, 3,
					-- layer=2 filter=10 channel=87
					-10, -8, 2, 9, 0, 8, -6, 2, -7,
					-- layer=2 filter=10 channel=88
					-8, -11, -3, 4, 1, -7, -3, 9, 8,
					-- layer=2 filter=10 channel=89
					4, 4, -12, 1, -3, -13, -7, 1, -5,
					-- layer=2 filter=10 channel=90
					3, 3, -11, 5, -8, -3, -2, -4, 6,
					-- layer=2 filter=10 channel=91
					3, -12, -10, -3, -10, -11, -11, -3, -9,
					-- layer=2 filter=10 channel=92
					-5, -7, -2, -2, 2, -4, -4, 2, -3,
					-- layer=2 filter=10 channel=93
					2, -10, -7, 1, 2, 7, -6, -5, 0,
					-- layer=2 filter=10 channel=94
					1, -9, -10, -2, -9, -11, -6, 9, -1,
					-- layer=2 filter=10 channel=95
					-11, 8, -1, 4, 0, 2, 3, -2, 2,
					-- layer=2 filter=10 channel=96
					0, -4, -12, 3, -1, -6, -4, 1, -7,
					-- layer=2 filter=10 channel=97
					7, -7, -6, -9, 0, 4, 5, -6, -10,
					-- layer=2 filter=10 channel=98
					-16, -17, -8, -4, -6, 3, -8, -1, -3,
					-- layer=2 filter=10 channel=99
					2, -5, -18, -1, -8, -14, -12, -9, 1,
					-- layer=2 filter=10 channel=100
					-8, 1, 0, -7, 7, 0, -3, -8, 0,
					-- layer=2 filter=10 channel=101
					1, -12, -12, 3, 9, -16, -4, 0, -5,
					-- layer=2 filter=10 channel=102
					-6, -13, 0, 5, -11, -9, -8, 6, 5,
					-- layer=2 filter=10 channel=103
					-6, 3, -9, 4, 5, -10, 7, 3, -6,
					-- layer=2 filter=10 channel=104
					0, 4, -4, 1, -1, -8, 0, -2, -1,
					-- layer=2 filter=10 channel=105
					8, 4, 4, -4, 0, -2, 0, -7, 5,
					-- layer=2 filter=10 channel=106
					-3, -3, -11, 0, -3, -2, 5, 7, 5,
					-- layer=2 filter=10 channel=107
					-5, 0, -6, 6, 4, -1, -4, -4, -5,
					-- layer=2 filter=10 channel=108
					2, -5, -2, 7, -14, -6, 8, -1, -4,
					-- layer=2 filter=10 channel=109
					0, -10, 0, -7, 1, -6, -1, -2, -12,
					-- layer=2 filter=10 channel=110
					-5, 3, -8, 0, -11, 6, -11, 6, 2,
					-- layer=2 filter=10 channel=111
					3, 8, -4, -12, 6, -2, 10, 1, 7,
					-- layer=2 filter=10 channel=112
					-14, 3, 3, 1, -3, -10, -1, -7, 2,
					-- layer=2 filter=10 channel=113
					-9, 4, 6, -7, -4, 8, -12, 0, 2,
					-- layer=2 filter=10 channel=114
					0, -5, 4, -7, -4, -8, -1, -1, 0,
					-- layer=2 filter=10 channel=115
					1, 2, -2, 0, 9, 2, 8, -10, 7,
					-- layer=2 filter=10 channel=116
					0, -16, -2, 3, -9, -9, -3, 0, 9,
					-- layer=2 filter=10 channel=117
					-4, -11, -19, 0, -5, -7, 5, 5, 0,
					-- layer=2 filter=10 channel=118
					8, 3, 4, 4, 1, -12, 7, -8, -6,
					-- layer=2 filter=10 channel=119
					-6, -7, -12, 3, 5, 5, -12, 3, -8,
					-- layer=2 filter=10 channel=120
					-8, 5, 9, -6, 2, -5, -7, 10, 1,
					-- layer=2 filter=10 channel=121
					2, 9, 7, 1, 3, -5, -9, -6, -7,
					-- layer=2 filter=10 channel=122
					-10, 0, 10, 7, 8, -6, -7, 1, -9,
					-- layer=2 filter=10 channel=123
					-3, -13, 1, -9, 2, 0, -4, -14, -5,
					-- layer=2 filter=10 channel=124
					-8, -6, 9, 7, 1, -12, 1, -1, -6,
					-- layer=2 filter=10 channel=125
					-8, 3, 2, 11, -5, -1, -4, -8, 3,
					-- layer=2 filter=10 channel=126
					8, 3, -8, 6, 5, -11, -10, 2, 5,
					-- layer=2 filter=10 channel=127
					-8, 0, 0, -2, -8, 0, 2, -6, 5,
					-- layer=2 filter=11 channel=0
					-1, 0, 0, -11, -15, 2, 2, 0, -12,
					-- layer=2 filter=11 channel=1
					-15, -12, -2, -15, -12, -8, -19, -25, -3,
					-- layer=2 filter=11 channel=2
					5, -9, 6, 7, -10, 3, 6, 10, -10,
					-- layer=2 filter=11 channel=3
					0, 10, -3, 0, 1, -15, 5, 0, 0,
					-- layer=2 filter=11 channel=4
					0, -6, -6, -3, 3, 9, -4, -2, 8,
					-- layer=2 filter=11 channel=5
					-8, -19, -5, -17, 0, 3, 4, -2, -3,
					-- layer=2 filter=11 channel=6
					-22, 8, -12, -19, -9, -15, 0, -10, -6,
					-- layer=2 filter=11 channel=7
					-1, -8, -10, 1, -12, -6, -5, -13, -12,
					-- layer=2 filter=11 channel=8
					-8, 2, 10, -10, 0, 2, -1, -8, 10,
					-- layer=2 filter=11 channel=9
					-12, -7, -17, 3, -9, -12, 0, -1, 2,
					-- layer=2 filter=11 channel=10
					2, -1, 4, 1, -8, -3, 5, -8, -5,
					-- layer=2 filter=11 channel=11
					-5, -21, -14, -9, -4, -8, -7, -5, -12,
					-- layer=2 filter=11 channel=12
					2, 0, -10, 3, -1, -13, -11, -20, -17,
					-- layer=2 filter=11 channel=13
					0, 3, -10, -2, 4, 6, 8, -1, -3,
					-- layer=2 filter=11 channel=14
					-11, 0, -8, -7, -2, -7, -12, -13, 3,
					-- layer=2 filter=11 channel=15
					0, 0, -9, 2, -3, -8, 0, -6, 7,
					-- layer=2 filter=11 channel=16
					-11, -3, -18, 0, -17, 1, -11, -14, -10,
					-- layer=2 filter=11 channel=17
					-7, 1, -6, -7, 1, -10, 0, 7, 8,
					-- layer=2 filter=11 channel=18
					-3, -15, 4, -7, 8, -8, -18, -8, -1,
					-- layer=2 filter=11 channel=19
					-10, -10, 1, -18, -10, -3, -6, -20, 1,
					-- layer=2 filter=11 channel=20
					-1, 0, -6, 4, 2, -7, 4, -8, -3,
					-- layer=2 filter=11 channel=21
					-2, 3, 1, 3, -3, 1, 0, -4, -1,
					-- layer=2 filter=11 channel=22
					10, -3, 0, 3, 1, -4, -8, 1, 3,
					-- layer=2 filter=11 channel=23
					-16, -11, 0, -9, 8, 2, -15, 2, 4,
					-- layer=2 filter=11 channel=24
					5, -4, -4, -3, 0, -13, -1, -1, -12,
					-- layer=2 filter=11 channel=25
					-14, -3, -11, -2, -5, -12, -9, -14, -15,
					-- layer=2 filter=11 channel=26
					0, 9, -2, -9, 1, -9, 0, 2, -2,
					-- layer=2 filter=11 channel=27
					6, 4, -1, -12, -17, -4, -11, -15, -6,
					-- layer=2 filter=11 channel=28
					0, 0, -1, 7, -5, 0, 1, 8, -1,
					-- layer=2 filter=11 channel=29
					7, 2, -7, 0, -10, -3, -8, 6, 3,
					-- layer=2 filter=11 channel=30
					-15, -18, -11, -17, -8, -2, -6, 4, -9,
					-- layer=2 filter=11 channel=31
					4, 4, -10, 0, 9, 1, -6, 3, 2,
					-- layer=2 filter=11 channel=32
					-1, 5, 2, -5, 1, -5, -7, -9, 6,
					-- layer=2 filter=11 channel=33
					-5, 19, 5, 14, -9, 2, 1, -4, 4,
					-- layer=2 filter=11 channel=34
					-5, 2, -15, -11, 0, -6, -10, -7, -5,
					-- layer=2 filter=11 channel=35
					5, -3, -8, -1, -19, 2, -11, -7, -5,
					-- layer=2 filter=11 channel=36
					2, -1, 7, -3, -8, 5, -2, -6, 3,
					-- layer=2 filter=11 channel=37
					-10, -12, -11, -5, -13, -11, 0, -10, 1,
					-- layer=2 filter=11 channel=38
					3, -7, -2, -14, -8, 7, -6, 0, 3,
					-- layer=2 filter=11 channel=39
					0, -4, -17, -7, -8, -9, -15, -17, 5,
					-- layer=2 filter=11 channel=40
					-9, -2, -13, -5, -2, -10, 10, -21, -1,
					-- layer=2 filter=11 channel=41
					5, 0, -5, -1, 8, -8, -8, 1, -1,
					-- layer=2 filter=11 channel=42
					4, -6, -3, -7, -15, -3, 2, -8, -12,
					-- layer=2 filter=11 channel=43
					12, -11, -2, -11, -9, 6, 0, -9, -2,
					-- layer=2 filter=11 channel=44
					-3, 5, 2, 6, 8, 8, -8, -3, -9,
					-- layer=2 filter=11 channel=45
					2, 0, 7, -8, 3, -2, 2, -6, -11,
					-- layer=2 filter=11 channel=46
					-7, 4, -10, -14, -13, 7, -6, -12, 3,
					-- layer=2 filter=11 channel=47
					-9, -2, 0, 1, -3, -1, -20, -8, -4,
					-- layer=2 filter=11 channel=48
					0, -3, -9, 1, -8, 8, -6, -9, 9,
					-- layer=2 filter=11 channel=49
					-4, -4, 7, -5, 2, -15, -1, 1, -5,
					-- layer=2 filter=11 channel=50
					2, -6, 4, 12, 9, -2, 5, 7, 11,
					-- layer=2 filter=11 channel=51
					-10, -14, -12, 0, -19, -20, -11, -6, -6,
					-- layer=2 filter=11 channel=52
					-19, -15, 5, -19, 0, 4, -12, -17, -7,
					-- layer=2 filter=11 channel=53
					11, 11, -2, -1, -11, 6, -8, -19, -6,
					-- layer=2 filter=11 channel=54
					-17, -18, -10, 0, -15, 0, -18, -3, 1,
					-- layer=2 filter=11 channel=55
					4, 10, 8, 7, 4, -11, -6, 9, 7,
					-- layer=2 filter=11 channel=56
					0, -1, -7, -7, -12, -17, -11, -3, 1,
					-- layer=2 filter=11 channel=57
					-4, 8, -3, 7, -6, -1, 0, 6, -5,
					-- layer=2 filter=11 channel=58
					-8, -14, -15, -11, -8, -1, -8, -11, -2,
					-- layer=2 filter=11 channel=59
					-8, 0, -9, 2, -21, -7, -20, -9, -9,
					-- layer=2 filter=11 channel=60
					-15, -17, -3, -10, -3, -9, -22, -10, 4,
					-- layer=2 filter=11 channel=61
					-5, -6, 8, -14, 2, -5, -7, -7, 0,
					-- layer=2 filter=11 channel=62
					-21, -15, -2, -9, -20, -22, -17, 6, -5,
					-- layer=2 filter=11 channel=63
					-13, -12, -9, -1, -1, -8, -11, -6, -2,
					-- layer=2 filter=11 channel=64
					-8, -3, -12, 3, -7, -4, -7, -4, -9,
					-- layer=2 filter=11 channel=65
					-10, 0, -11, -8, -10, -9, -16, -1, -7,
					-- layer=2 filter=11 channel=66
					0, 4, -10, 6, -4, 4, 5, 5, 10,
					-- layer=2 filter=11 channel=67
					-10, -12, -16, -16, -17, 2, -5, 2, -4,
					-- layer=2 filter=11 channel=68
					-6, -6, 4, 0, -6, -7, -11, -9, -2,
					-- layer=2 filter=11 channel=69
					-9, -12, -2, -14, 4, -6, 1, 1, -16,
					-- layer=2 filter=11 channel=70
					-1, -16, -1, -5, -12, 4, -11, -2, 6,
					-- layer=2 filter=11 channel=71
					-3, -6, 7, 0, -7, 5, -8, -7, -5,
					-- layer=2 filter=11 channel=72
					-3, -9, 6, -6, -4, 5, -7, -7, -17,
					-- layer=2 filter=11 channel=73
					-11, -15, -5, 8, -11, -8, -2, -1, 2,
					-- layer=2 filter=11 channel=74
					-9, -12, -19, 5, -13, 10, -10, -8, 8,
					-- layer=2 filter=11 channel=75
					-8, 6, 0, 0, -12, -10, -13, 12, -10,
					-- layer=2 filter=11 channel=76
					-7, -14, -20, 0, -13, 4, 1, 0, 5,
					-- layer=2 filter=11 channel=77
					-5, 5, 2, -8, -10, 0, -11, 6, 7,
					-- layer=2 filter=11 channel=78
					-14, 0, -10, -13, -13, -3, -19, -2, -13,
					-- layer=2 filter=11 channel=79
					-11, -3, 9, 1, -4, -8, -1, 5, 4,
					-- layer=2 filter=11 channel=80
					1, -12, -2, 0, -9, 8, -7, -8, 9,
					-- layer=2 filter=11 channel=81
					0, -9, 5, -10, -9, -6, 6, 4, 4,
					-- layer=2 filter=11 channel=82
					-11, -6, 8, 5, 6, -7, -8, -5, 0,
					-- layer=2 filter=11 channel=83
					-4, -6, -8, 2, 4, -1, -7, 6, -4,
					-- layer=2 filter=11 channel=84
					7, 4, 6, -3, 1, -3, -7, 1, -9,
					-- layer=2 filter=11 channel=85
					7, 9, 4, -8, -3, 3, 6, 0, -9,
					-- layer=2 filter=11 channel=86
					-5, 1, 5, -5, -9, 7, 4, 8, -3,
					-- layer=2 filter=11 channel=87
					-9, -6, 9, 1, -1, -12, -18, 4, 9,
					-- layer=2 filter=11 channel=88
					0, -4, -5, -9, 0, -3, -14, -8, -12,
					-- layer=2 filter=11 channel=89
					-7, -1, -7, 2, -14, -5, -6, 5, -8,
					-- layer=2 filter=11 channel=90
					8, -4, 0, -7, -7, 1, 3, -5, 7,
					-- layer=2 filter=11 channel=91
					5, -9, 4, 12, -3, -1, 1, -6, -9,
					-- layer=2 filter=11 channel=92
					-2, -2, 0, -7, -13, 6, -16, -17, -4,
					-- layer=2 filter=11 channel=93
					-16, 9, 3, -25, -9, -8, -7, 5, 5,
					-- layer=2 filter=11 channel=94
					-7, -13, 7, 0, -20, -2, -19, -10, -17,
					-- layer=2 filter=11 channel=95
					1, 2, 9, 4, -1, -3, 2, -4, 4,
					-- layer=2 filter=11 channel=96
					-7, -10, -16, -4, 8, 1, -17, -1, -15,
					-- layer=2 filter=11 channel=97
					3, 0, 4, -5, -19, -14, -7, 2, -4,
					-- layer=2 filter=11 channel=98
					-17, 3, 5, -9, -19, -19, -14, -18, 1,
					-- layer=2 filter=11 channel=99
					-3, -7, -19, -16, -13, 1, -13, -20, -2,
					-- layer=2 filter=11 channel=100
					4, -6, -2, 0, -6, -2, -1, -12, -5,
					-- layer=2 filter=11 channel=101
					-14, -8, -4, -3, -14, -7, -11, 3, 4,
					-- layer=2 filter=11 channel=102
					-17, -14, -7, 2, 0, -5, -2, 5, -11,
					-- layer=2 filter=11 channel=103
					-3, 5, 9, -10, -7, 0, 0, -8, -10,
					-- layer=2 filter=11 channel=104
					0, -15, 10, -3, 1, 6, 5, 1, 3,
					-- layer=2 filter=11 channel=105
					-8, 1, 0, -8, -5, 4, -10, -6, 10,
					-- layer=2 filter=11 channel=106
					8, -7, -12, 8, 5, -8, -8, -3, -7,
					-- layer=2 filter=11 channel=107
					-9, 0, -8, -2, 4, -6, -4, 3, 3,
					-- layer=2 filter=11 channel=108
					-1, -3, 2, 0, 0, 2, -5, -9, 0,
					-- layer=2 filter=11 channel=109
					2, -3, 8, -3, -3, -4, 1, -10, -4,
					-- layer=2 filter=11 channel=110
					-6, -13, -15, -7, -20, 4, -10, -1, 0,
					-- layer=2 filter=11 channel=111
					10, 2, -3, 4, 6, -6, -2, -3, -1,
					-- layer=2 filter=11 channel=112
					-7, -6, 8, -10, -4, -8, -12, -7, -4,
					-- layer=2 filter=11 channel=113
					-10, 8, -12, -7, -10, 0, -6, -9, -10,
					-- layer=2 filter=11 channel=114
					-2, -2, -4, 8, -6, 8, 5, -2, 0,
					-- layer=2 filter=11 channel=115
					7, 7, 5, -10, 1, -5, -3, 9, 2,
					-- layer=2 filter=11 channel=116
					-17, -11, 7, 9, 6, -9, 4, 3, -4,
					-- layer=2 filter=11 channel=117
					-3, -10, 2, -14, 2, -7, -7, -9, -7,
					-- layer=2 filter=11 channel=118
					2, 4, -8, -11, 0, 3, -11, -4, 1,
					-- layer=2 filter=11 channel=119
					-1, -6, -4, -16, -2, -6, -13, -8, 4,
					-- layer=2 filter=11 channel=120
					8, 5, 6, -6, -9, 0, 4, 3, 6,
					-- layer=2 filter=11 channel=121
					7, 0, 8, 8, 8, -10, -7, -2, 10,
					-- layer=2 filter=11 channel=122
					-2, 0, 2, -3, 6, 7, -3, -5, 1,
					-- layer=2 filter=11 channel=123
					-13, 17, -10, -8, -12, 4, -2, -13, -3,
					-- layer=2 filter=11 channel=124
					2, 2, 3, -14, -17, -4, -2, -2, -9,
					-- layer=2 filter=11 channel=125
					8, 5, 10, -1, 8, 8, 0, 5, -1,
					-- layer=2 filter=11 channel=126
					-4, 0, 0, -5, -3, -8, 1, -7, -3,
					-- layer=2 filter=11 channel=127
					-16, -5, -1, 0, 1, 0, -18, 3, -11,
					-- layer=2 filter=12 channel=0
					20, 18, 0, 19, 18, 8, 13, 22, 18,
					-- layer=2 filter=12 channel=1
					-51, 26, 14, -33, -23, 0, -16, -21, 0,
					-- layer=2 filter=12 channel=2
					3, -1, 4, -5, 0, 3, 6, 5, 5,
					-- layer=2 filter=12 channel=3
					32, 29, 11, 10, -2, -18, 1, -8, -15,
					-- layer=2 filter=12 channel=4
					-53, -55, 6, -34, -59, -37, -44, -61, -13,
					-- layer=2 filter=12 channel=5
					16, -7, -8, 39, 29, 15, 2, 7, 32,
					-- layer=2 filter=12 channel=6
					3, 39, 26, 30, 12, -1, 40, 18, 34,
					-- layer=2 filter=12 channel=7
					3, -35, 13, -45, -31, 38, -17, 0, 20,
					-- layer=2 filter=12 channel=8
					9, -7, -3, -4, -6, 0, -7, 6, 2,
					-- layer=2 filter=12 channel=9
					16, 6, -31, -16, 10, 3, -2, 29, -37,
					-- layer=2 filter=12 channel=10
					52, 12, 19, 32, 22, 17, 7, 24, 13,
					-- layer=2 filter=12 channel=11
					0, 9, 7, 20, 10, 1, 14, 14, 18,
					-- layer=2 filter=12 channel=12
					-13, 23, 8, -22, -3, -5, 18, -35, -8,
					-- layer=2 filter=12 channel=13
					4, 9, 0, 8, 7, 8, -8, -1, -5,
					-- layer=2 filter=12 channel=14
					-23, 0, 0, -27, -30, -18, 4, -22, -8,
					-- layer=2 filter=12 channel=15
					3, -9, -14, 0, -12, 44, -48, -16, -38,
					-- layer=2 filter=12 channel=16
					9, -59, -2, -6, 33, 49, 20, 58, 14,
					-- layer=2 filter=12 channel=17
					-7, -6, -5, 7, 9, -2, -9, -4, -10,
					-- layer=2 filter=12 channel=18
					-72, -41, 7, -27, -24, -21, -64, -57, -23,
					-- layer=2 filter=12 channel=19
					-18, 12, 55, -10, 19, 46, -16, -7, -16,
					-- layer=2 filter=12 channel=20
					5, 3, 0, 7, 0, -4, -2, -3, -5,
					-- layer=2 filter=12 channel=21
					14, -3, 16, 13, 6, 20, 19, 0, 18,
					-- layer=2 filter=12 channel=22
					13, 7, 0, -5, 9, 6, -4, -5, 4,
					-- layer=2 filter=12 channel=23
					-17, -22, -15, -37, -32, -51, -1, -38, -31,
					-- layer=2 filter=12 channel=24
					-8, 7, -11, 3, 9, -22, 25, 27, 9,
					-- layer=2 filter=12 channel=25
					1, 14, -12, 1, 3, -21, 8, 16, 18,
					-- layer=2 filter=12 channel=26
					5, 0, 7, -1, -8, 9, -6, 7, -5,
					-- layer=2 filter=12 channel=27
					21, -15, 20, 25, -1, 5, 6, 11, 23,
					-- layer=2 filter=12 channel=28
					-6, 27, -10, 12, 19, -4, 4, 11, 17,
					-- layer=2 filter=12 channel=29
					-5, 9, 0, -1, 0, -2, -5, 7, -5,
					-- layer=2 filter=12 channel=30
					-38, -71, -55, -6, -88, -11, -45, -49, -38,
					-- layer=2 filter=12 channel=31
					52, 24, -26, -7, 55, 19, 5, 2, -83,
					-- layer=2 filter=12 channel=32
					-9, 4, 5, -4, -5, 5, -5, -8, -3,
					-- layer=2 filter=12 channel=33
					27, 5, 19, -34, -30, 12, -31, -35, 21,
					-- layer=2 filter=12 channel=34
					-49, -3, 76, 9, 69, 39, -35, -26, 2,
					-- layer=2 filter=12 channel=35
					34, -8, 14, -26, -16, -30, -12, 0, -27,
					-- layer=2 filter=12 channel=36
					2, 9, 14, 8, 0, 8, -4, 0, 12,
					-- layer=2 filter=12 channel=37
					1, 12, 9, 28, 7, 17, 4, -3, 29,
					-- layer=2 filter=12 channel=38
					4, -12, 0, 12, 0, -8, 20, -6, 2,
					-- layer=2 filter=12 channel=39
					-25, -39, 34, -39, -9, 32, -39, -4, -19,
					-- layer=2 filter=12 channel=40
					7, -54, -22, -45, 35, 10, -38, -49, -2,
					-- layer=2 filter=12 channel=41
					11, -6, 6, 10, 3, -1, -1, 12, 3,
					-- layer=2 filter=12 channel=42
					-8, 11, 0, -59, -35, -50, 35, -44, -7,
					-- layer=2 filter=12 channel=43
					14, -1, 25, 36, 22, -12, -16, 21, -4,
					-- layer=2 filter=12 channel=44
					5, 6, 4, 5, -3, -2, -1, -7, 8,
					-- layer=2 filter=12 channel=45
					-9, -29, -40, -56, -65, -23, -54, -91, 13,
					-- layer=2 filter=12 channel=46
					-30, -21, -15, 9, -7, -19, -37, -3, -29,
					-- layer=2 filter=12 channel=47
					7, -23, -23, -25, -6, -14, -1, -44, 8,
					-- layer=2 filter=12 channel=48
					-2, 5, 0, -3, -10, -1, 10, 10, -9,
					-- layer=2 filter=12 channel=49
					-60, -27, 3, -22, -14, -18, -44, -65, -45,
					-- layer=2 filter=12 channel=50
					-10, -2, -1, -8, -5, -4, 9, 12, 15,
					-- layer=2 filter=12 channel=51
					6, 16, 11, 24, 5, 0, 10, 16, 15,
					-- layer=2 filter=12 channel=52
					-21, 16, 2, 5, 5, 33, 8, 26, 52,
					-- layer=2 filter=12 channel=53
					-96, 10, -1, -41, -17, -44, 6, -57, -12,
					-- layer=2 filter=12 channel=54
					-8, 19, 24, 2, 24, 28, 1, 25, 42,
					-- layer=2 filter=12 channel=55
					-1, 0, -3, 3, -7, -8, 1, 0, 4,
					-- layer=2 filter=12 channel=56
					9, -5, 13, 26, -3, 0, 12, -11, 8,
					-- layer=2 filter=12 channel=57
					-10, 0, -1, -13, -3, 0, 4, 11, 7,
					-- layer=2 filter=12 channel=58
					7, 40, 14, -20, 5, 20, 29, -10, 2,
					-- layer=2 filter=12 channel=59
					-38, 14, 28, -17, -10, 20, -19, 28, 4,
					-- layer=2 filter=12 channel=60
					-21, 24, 40, -24, 23, 38, 19, -12, 12,
					-- layer=2 filter=12 channel=61
					-33, 4, -24, -31, 9, -10, -7, 2, -14,
					-- layer=2 filter=12 channel=62
					-17, 22, 28, 6, 12, 22, -12, 30, 17,
					-- layer=2 filter=12 channel=63
					-22, 2, -32, -41, 36, -13, 0, -24, -17,
					-- layer=2 filter=12 channel=64
					1, -24, -10, 19, 0, -22, -1, 34, 5,
					-- layer=2 filter=12 channel=65
					0, 17, -2, 21, -23, 2, 19, 0, 12,
					-- layer=2 filter=12 channel=66
					7, -34, 3, 14, -21, 18, 54, -8, 73,
					-- layer=2 filter=12 channel=67
					-13, -33, 3, 27, 23, -14, -2, -8, -9,
					-- layer=2 filter=12 channel=68
					-2, 6, 9, 0, 0, -3, -8, 9, 2,
					-- layer=2 filter=12 channel=69
					-22, -13, 5, -5, -35, 4, -18, -20, -6,
					-- layer=2 filter=12 channel=70
					20, 12, 9, -6, 22, 10, -3, 0, 21,
					-- layer=2 filter=12 channel=71
					-1, -3, 15, -3, -41, -3, -1, -41, 16,
					-- layer=2 filter=12 channel=72
					7, 17, 58, -24, 0, -5, -3, -6, 37,
					-- layer=2 filter=12 channel=73
					0, -17, 15, 11, -6, 23, -26, -43, -1,
					-- layer=2 filter=12 channel=74
					-14, -54, -28, 9, 9, -54, -19, 7, -49,
					-- layer=2 filter=12 channel=75
					-18, 26, -19, -19, -6, 3, 15, 10, -35,
					-- layer=2 filter=12 channel=76
					-53, -20, -54, -14, -15, 21, -50, -70, -22,
					-- layer=2 filter=12 channel=77
					-2, 2, 12, -4, 0, 4, 9, -1, 12,
					-- layer=2 filter=12 channel=78
					-7, 4, 4, 13, 4, -11, 22, 14, -9,
					-- layer=2 filter=12 channel=79
					6, -7, 9, -2, -4, 11, -4, -8, 0,
					-- layer=2 filter=12 channel=80
					-37, -4, -17, -43, 20, -37, -19, -41, -30,
					-- layer=2 filter=12 channel=81
					-3, 5, -11, 9, -4, -5, 1, 5, 8,
					-- layer=2 filter=12 channel=82
					-4, 1, -1, 8, 8, -9, 4, -8, -2,
					-- layer=2 filter=12 channel=83
					-1, 1, 1, -26, -41, -34, 40, -31, -31,
					-- layer=2 filter=12 channel=84
					-1, 3, -5, 0, -4, -9, -9, 2, -10,
					-- layer=2 filter=12 channel=85
					-1, 9, 5, 5, 11, 6, 9, 6, 1,
					-- layer=2 filter=12 channel=86
					-2, 4, 14, 0, 7, 5, 2, 6, 5,
					-- layer=2 filter=12 channel=87
					23, -3, 46, -49, 42, -19, 0, -13, -28,
					-- layer=2 filter=12 channel=88
					-40, -63, -76, -34, -40, -57, -17, -28, -97,
					-- layer=2 filter=12 channel=89
					-37, 29, 20, -30, -18, -13, -20, 0, -16,
					-- layer=2 filter=12 channel=90
					3, 8, -6, 10, 3, 8, -1, 0, 9,
					-- layer=2 filter=12 channel=91
					-15, 32, 17, -20, 19, 12, 10, 5, 0,
					-- layer=2 filter=12 channel=92
					-16, 48, 12, -20, -25, -14, -1, -33, -42,
					-- layer=2 filter=12 channel=93
					8, -35, 12, 39, -20, -29, -6, -8, -2,
					-- layer=2 filter=12 channel=94
					-30, 18, 25, -16, 22, -10, 26, -12, -4,
					-- layer=2 filter=12 channel=95
					-12, -10, -4, -11, -11, 3, 2, -13, 3,
					-- layer=2 filter=12 channel=96
					-4, 25, 32, 0, 27, 5, 38, 30, 26,
					-- layer=2 filter=12 channel=97
					-1, -9, -1, -23, -30, -35, 6, 16, -23,
					-- layer=2 filter=12 channel=98
					11, 9, 27, 3, 24, 3, 16, 21, 22,
					-- layer=2 filter=12 channel=99
					-38, -7, 39, -5, 1, 46, -13, 32, 25,
					-- layer=2 filter=12 channel=100
					-4, 24, -12, 7, 16, 2, 15, 19, 51,
					-- layer=2 filter=12 channel=101
					15, -23, -6, -20, -38, -45, -25, -46, -47,
					-- layer=2 filter=12 channel=102
					-21, -11, -11, 14, -40, -15, 4, 0, -28,
					-- layer=2 filter=12 channel=103
					9, -38, -17, -13, 22, 15, -4, -22, -9,
					-- layer=2 filter=12 channel=104
					-52, -10, -2, 6, 16, -46, -40, -61, 0,
					-- layer=2 filter=12 channel=105
					-53, -16, 2, -70, 3, 35, 2, -5, -20,
					-- layer=2 filter=12 channel=106
					15, 12, 16, -6, 1, -14, -9, -4, 4,
					-- layer=2 filter=12 channel=107
					-21, -2, -39, -5, -35, 7, 3, 13, -44,
					-- layer=2 filter=12 channel=108
					-25, -4, 27, -18, -26, 0, -9, -9, -9,
					-- layer=2 filter=12 channel=109
					11, 10, -3, 5, 3, -12, 14, 1, 1,
					-- layer=2 filter=12 channel=110
					0, 8, 2, -3, 6, -25, -7, 30, 28,
					-- layer=2 filter=12 channel=111
					-5, -4, -6, 0, 8, -4, -10, 6, 4,
					-- layer=2 filter=12 channel=112
					8, 3, -16, 14, 2, -14, 9, -1, -4,
					-- layer=2 filter=12 channel=113
					-42, -38, -86, -30, -57, -17, -36, 8, -19,
					-- layer=2 filter=12 channel=114
					0, -2, 13, -10, -2, 2, 4, -11, 18,
					-- layer=2 filter=12 channel=115
					8, 1, 1, -3, -3, 7, -4, 4, -6,
					-- layer=2 filter=12 channel=116
					-10, 27, 47, -14, 11, -21, -12, -23, 18,
					-- layer=2 filter=12 channel=117
					5, -15, 12, -54, -27, 41, -41, -2, 7,
					-- layer=2 filter=12 channel=118
					28, 26, 32, 34, 29, -11, 5, 5, 10,
					-- layer=2 filter=12 channel=119
					-58, -62, -35, -11, -35, -15, -114, -106, -29,
					-- layer=2 filter=12 channel=120
					5, -4, 8, 0, 8, 0, 2, -9, 0,
					-- layer=2 filter=12 channel=121
					5, 4, 6, -1, 2, -7, -4, -5, -8,
					-- layer=2 filter=12 channel=122
					10, 0, 8, 6, -1, -6, 9, -1, 8,
					-- layer=2 filter=12 channel=123
					-23, 38, 33, -27, 14, 29, -7, -1, 44,
					-- layer=2 filter=12 channel=124
					-32, -20, -24, 0, -44, 49, -84, -8, -50,
					-- layer=2 filter=12 channel=125
					-7, -4, -8, 7, -11, 7, 1, -4, -5,
					-- layer=2 filter=12 channel=126
					-11, 12, -4, -34, -12, 11, -13, -1, -39,
					-- layer=2 filter=12 channel=127
					-44, 21, -7, -28, -46, -29, -8, -14, -11,
					-- layer=2 filter=13 channel=0
					1, 3, 9, 3, 14, 8, -3, -8, 14,
					-- layer=2 filter=13 channel=1
					9, 24, 40, -9, 24, 11, 8, -27, -15,
					-- layer=2 filter=13 channel=2
					1, 5, 7, -11, 2, -8, -6, -3, -10,
					-- layer=2 filter=13 channel=3
					-16, -21, -27, 28, 4, -14, 31, 55, 34,
					-- layer=2 filter=13 channel=4
					-15, 8, -3, 11, -22, -29, 27, -1, -31,
					-- layer=2 filter=13 channel=5
					9, -2, 20, -14, -3, 30, -20, -3, 14,
					-- layer=2 filter=13 channel=6
					21, 19, 12, 2, -22, -62, -50, -36, -42,
					-- layer=2 filter=13 channel=7
					-14, -4, 25, 0, -10, 18, -17, -16, -18,
					-- layer=2 filter=13 channel=8
					-5, -5, -6, 1, 1, -5, 8, 3, -3,
					-- layer=2 filter=13 channel=9
					-7, -10, 16, 12, 1, -23, 53, 61, 11,
					-- layer=2 filter=13 channel=10
					-12, -13, -22, 4, 11, -9, 29, 15, 30,
					-- layer=2 filter=13 channel=11
					-8, -12, -4, -13, -22, 17, -21, 12, 4,
					-- layer=2 filter=13 channel=12
					-7, 35, 48, -16, 8, 23, 2, -7, 6,
					-- layer=2 filter=13 channel=13
					-11, 5, 6, -3, 3, 2, -1, 0, 5,
					-- layer=2 filter=13 channel=14
					-8, 17, 26, -44, 0, -4, -12, -22, -15,
					-- layer=2 filter=13 channel=15
					-9, -1, 55, -53, 51, 34, -42, 8, 39,
					-- layer=2 filter=13 channel=16
					-8, 18, 24, -18, -6, -33, -24, -25, -54,
					-- layer=2 filter=13 channel=17
					0, 0, -4, 0, -2, -8, 0, 0, 0,
					-- layer=2 filter=13 channel=18
					37, 11, 20, 10, 35, 2, -1, 7, 16,
					-- layer=2 filter=13 channel=19
					38, 21, 27, -12, 24, 0, -41, -28, -24,
					-- layer=2 filter=13 channel=20
					-2, -8, 0, -3, 11, 4, 1, -8, 1,
					-- layer=2 filter=13 channel=21
					0, -6, -8, 11, 0, 0, 14, 6, -6,
					-- layer=2 filter=13 channel=22
					6, -5, 3, 10, 4, 5, -9, 7, -1,
					-- layer=2 filter=13 channel=23
					-28, 5, -4, 16, 12, 6, 24, 30, -31,
					-- layer=2 filter=13 channel=24
					1, -42, -11, 8, -29, -30, 28, 24, 6,
					-- layer=2 filter=13 channel=25
					-39, -71, -25, -17, -35, -42, -15, 2, -4,
					-- layer=2 filter=13 channel=26
					-8, 2, 5, 4, -10, 0, -2, -6, 8,
					-- layer=2 filter=13 channel=27
					18, 11, 11, -26, -14, -2, -32, -34, -18,
					-- layer=2 filter=13 channel=28
					-31, 11, -15, -29, 33, 7, -29, 7, -12,
					-- layer=2 filter=13 channel=29
					-7, 5, -3, 7, 6, -6, 2, -6, -7,
					-- layer=2 filter=13 channel=30
					-4, -16, -14, -3, 17, -13, 21, -13, 13,
					-- layer=2 filter=13 channel=31
					-3, -61, -32, 19, -52, -41, -29, 24, 33,
					-- layer=2 filter=13 channel=32
					9, 0, 3, 5, 5, -11, -2, -4, 1,
					-- layer=2 filter=13 channel=33
					-37, -5, -40, -54, -19, -13, 0, 22, 24,
					-- layer=2 filter=13 channel=34
					22, 23, -53, -49, 3, 12, -80, -9, 12,
					-- layer=2 filter=13 channel=35
					-6, -5, -3, -37, -12, -1, -21, -20, 29,
					-- layer=2 filter=13 channel=36
					1, -5, 2, -12, 1, -3, -5, 9, -7,
					-- layer=2 filter=13 channel=37
					7, -7, 18, -12, -13, 21, -13, 8, 7,
					-- layer=2 filter=13 channel=38
					2, -2, -5, -17, -14, -3, -54, -31, -2,
					-- layer=2 filter=13 channel=39
					-38, -32, -30, -3, -11, -25, 34, 34, -3,
					-- layer=2 filter=13 channel=40
					-1, -33, 15, -43, -16, 9, -38, 10, 0,
					-- layer=2 filter=13 channel=41
					-2, -9, -5, 8, -2, -2, -7, -6, 3,
					-- layer=2 filter=13 channel=42
					-12, -2, -12, -19, -22, -15, 38, 10, -4,
					-- layer=2 filter=13 channel=43
					-3, 15, 26, 15, 23, -13, 27, 0, 21,
					-- layer=2 filter=13 channel=44
					0, -6, 6, 2, -6, -4, 3, -7, 9,
					-- layer=2 filter=13 channel=45
					-18, 9, -15, -38, -23, 5, 11, -30, -22,
					-- layer=2 filter=13 channel=46
					15, -18, -3, -23, 14, -27, -8, 16, 19,
					-- layer=2 filter=13 channel=47
					-52, 0, 8, -61, -2, -5, -48, -24, -53,
					-- layer=2 filter=13 channel=48
					7, 5, -2, 6, 0, 8, -6, -6, -2,
					-- layer=2 filter=13 channel=49
					31, 43, 27, 4, 35, -18, 6, -22, -35,
					-- layer=2 filter=13 channel=50
					6, 17, 30, -10, -6, -10, 17, -16, 4,
					-- layer=2 filter=13 channel=51
					4, -2, -11, 6, -1, 3, -7, -9, -4,
					-- layer=2 filter=13 channel=52
					25, 10, 23, -44, 5, -13, -1, -15, 39,
					-- layer=2 filter=13 channel=53
					-3, -17, 52, -12, 1, 13, -38, 9, -25,
					-- layer=2 filter=13 channel=54
					2, -11, -6, -7, 15, 35, -31, -11, 21,
					-- layer=2 filter=13 channel=55
					11, 3, -1, -12, -5, -6, -7, 0, -4,
					-- layer=2 filter=13 channel=56
					0, 2, 1, 2, -5, 10, -11, 12, 23,
					-- layer=2 filter=13 channel=57
					-6, 0, 1, -6, -3, 11, -4, 11, 0,
					-- layer=2 filter=13 channel=58
					-17, 17, 37, 12, 4, 23, -23, 11, -8,
					-- layer=2 filter=13 channel=59
					19, 2, 19, 20, -3, 17, -44, -18, -45,
					-- layer=2 filter=13 channel=60
					38, 9, -3, 5, 34, 36, -10, -24, -8,
					-- layer=2 filter=13 channel=61
					24, 45, -5, 31, 30, 44, 20, -32, -17,
					-- layer=2 filter=13 channel=62
					3, -5, -4, -11, -25, -5, -53, -44, -31,
					-- layer=2 filter=13 channel=63
					-35, 14, -1, 0, 21, 1, 17, 26, -11,
					-- layer=2 filter=13 channel=64
					-29, -12, -16, -11, -11, -5, 47, 34, 6,
					-- layer=2 filter=13 channel=65
					44, 40, 19, 5, 8, 31, -18, -6, -34,
					-- layer=2 filter=13 channel=66
					-3, 82, 20, -46, 0, 16, 27, -3, 15,
					-- layer=2 filter=13 channel=67
					23, -4, -10, 12, 17, 0, 32, 36, 54,
					-- layer=2 filter=13 channel=68
					9, 0, -5, -11, -7, 2, 7, 6, 6,
					-- layer=2 filter=13 channel=69
					-37, 7, -8, -11, -11, -9, 33, 14, -20,
					-- layer=2 filter=13 channel=70
					-1, -2, -31, -12, 15, 22, -24, -5, 15,
					-- layer=2 filter=13 channel=71
					-6, -8, 7, -5, -10, -1, 1, -17, 28,
					-- layer=2 filter=13 channel=72
					-53, 1, -12, -17, 13, -12, -11, 34, 20,
					-- layer=2 filter=13 channel=73
					-19, 53, 29, -33, -1, 12, -16, 4, -23,
					-- layer=2 filter=13 channel=74
					-18, -25, 8, 2, 17, 0, 21, 38, 38,
					-- layer=2 filter=13 channel=75
					-31, 21, -28, -88, 18, -25, -56, -30, -19,
					-- layer=2 filter=13 channel=76
					-23, -2, 70, -62, -47, -5, -25, -28, -43,
					-- layer=2 filter=13 channel=77
					-5, -3, -3, 2, -7, 3, 2, 1, -7,
					-- layer=2 filter=13 channel=78
					38, -12, 8, -17, -20, -33, 0, -1, 5,
					-- layer=2 filter=13 channel=79
					1, -10, -1, 11, 1, 2, 2, -10, -11,
					-- layer=2 filter=13 channel=80
					3, -20, -19, 13, -2, -13, 38, 38, 6,
					-- layer=2 filter=13 channel=81
					7, -15, -7, -14, -7, 2, -10, -5, -14,
					-- layer=2 filter=13 channel=82
					-9, -7, 4, 6, 7, 8, -4, 7, 6,
					-- layer=2 filter=13 channel=83
					-45, 1, 6, 9, 7, -11, 3, 9, -45,
					-- layer=2 filter=13 channel=84
					1, 3, -7, 3, 5, 5, 0, -1, 0,
					-- layer=2 filter=13 channel=85
					0, -8, 6, -7, 4, -2, -1, 17, 0,
					-- layer=2 filter=13 channel=86
					-9, 10, 11, 4, 32, 0, -7, -10, -3,
					-- layer=2 filter=13 channel=87
					20, -1, 4, 34, -11, 18, -19, 0, 0,
					-- layer=2 filter=13 channel=88
					-1, -3, 33, -7, 20, -13, 22, 19, 14,
					-- layer=2 filter=13 channel=89
					-10, -3, 28, -42, -11, -3, -20, -16, -3,
					-- layer=2 filter=13 channel=90
					5, -9, 2, 3, -9, 8, -6, 8, 10,
					-- layer=2 filter=13 channel=91
					11, 21, 13, -28, -4, -38, -22, -1, -28,
					-- layer=2 filter=13 channel=92
					-5, -3, 41, -5, -13, -8, 2, 3, -1,
					-- layer=2 filter=13 channel=93
					47, 34, 38, 0, -7, -9, -23, -21, -19,
					-- layer=2 filter=13 channel=94
					-7, 33, 30, 47, 0, 11, -39, -22, -27,
					-- layer=2 filter=13 channel=95
					16, 20, -26, 0, 10, 10, 24, 18, 6,
					-- layer=2 filter=13 channel=96
					31, 29, -7, 13, -11, 11, -12, -36, -87,
					-- layer=2 filter=13 channel=97
					-1, 2, 18, 27, -24, -55, 38, 0, -20,
					-- layer=2 filter=13 channel=98
					-20, -1, -4, -33, 31, 30, 1, 2, 4,
					-- layer=2 filter=13 channel=99
					32, 33, 10, 3, 25, 30, -10, -32, -16,
					-- layer=2 filter=13 channel=100
					-17, -11, -7, -11, 5, -5, 17, 2, 33,
					-- layer=2 filter=13 channel=101
					9, -21, 30, -6, -28, -4, -1, 1, 22,
					-- layer=2 filter=13 channel=102
					42, 52, 17, -5, 23, 22, 2, -34, -27,
					-- layer=2 filter=13 channel=103
					33, 9, 3, -44, 12, 16, 0, -18, -9,
					-- layer=2 filter=13 channel=104
					15, 21, 57, 31, -1, 13, -27, -1, -13,
					-- layer=2 filter=13 channel=105
					-10, -20, 23, 50, -37, 14, 21, -51, -61,
					-- layer=2 filter=13 channel=106
					-10, 5, -15, -7, -48, 3, 19, 4, 20,
					-- layer=2 filter=13 channel=107
					13, -66, -13, 13, -29, 27, 33, -7, 35,
					-- layer=2 filter=13 channel=108
					-4, 16, 12, -39, 4, -11, -16, -68, -58,
					-- layer=2 filter=13 channel=109
					5, 0, 3, -17, 4, 0, 0, 5, -6,
					-- layer=2 filter=13 channel=110
					-10, -6, -8, -11, -10, -4, 36, 22, 34,
					-- layer=2 filter=13 channel=111
					8, 3, -8, -7, 10, 1, 4, 11, 0,
					-- layer=2 filter=13 channel=112
					38, 8, -20, -13, -13, 12, 35, -26, -7,
					-- layer=2 filter=13 channel=113
					-21, -6, -1, -6, 11, -5, -4, 6, -22,
					-- layer=2 filter=13 channel=114
					-2, 14, -13, 1, 0, 9, 2, 1, -4,
					-- layer=2 filter=13 channel=115
					1, 8, -7, -2, -9, -3, -6, 0, -8,
					-- layer=2 filter=13 channel=116
					30, 55, 28, 7, 37, 22, 0, -14, 9,
					-- layer=2 filter=13 channel=117
					19, 16, 32, -12, 19, 9, 32, 20, 44,
					-- layer=2 filter=13 channel=118
					14, 21, -7, 25, 15, -24, 20, 17, -2,
					-- layer=2 filter=13 channel=119
					-4, -2, 18, -13, -1, -12, 38, -21, -20,
					-- layer=2 filter=13 channel=120
					-3, 0, 6, 0, 0, 6, 6, -2, 5,
					-- layer=2 filter=13 channel=121
					-2, 10, -2, -3, 10, -5, 4, -5, 4,
					-- layer=2 filter=13 channel=122
					18, -2, 7, 1, 5, 18, -15, -4, 8,
					-- layer=2 filter=13 channel=123
					-17, 20, 0, 0, 22, 2, -22, 8, -29,
					-- layer=2 filter=13 channel=124
					6, 13, 2, -4, 44, 51, -21, 0, 31,
					-- layer=2 filter=13 channel=125
					-8, 0, 5, -6, 3, -2, 4, 0, -12,
					-- layer=2 filter=13 channel=126
					7, -57, -16, -63, -19, 9, -6, -51, -76,
					-- layer=2 filter=13 channel=127
					-7, 26, -7, -21, 3, -12, 42, 8, -22,
					-- layer=2 filter=14 channel=0
					-10, -7, -22, 18, -11, 1, 27, -22, 9,
					-- layer=2 filter=14 channel=1
					27, 13, 33, -10, 30, 6, 5, 19, 10,
					-- layer=2 filter=14 channel=2
					0, 0, 1, -6, 0, 7, -10, -2, -11,
					-- layer=2 filter=14 channel=3
					-35, -27, -25, 21, 13, 6, 56, -1, 19,
					-- layer=2 filter=14 channel=4
					-37, 28, -37, -1, -28, -62, -22, -22, -28,
					-- layer=2 filter=14 channel=5
					-18, -14, 49, -9, 2, 26, 17, -9, 10,
					-- layer=2 filter=14 channel=6
					36, 2, 20, 1, -8, -3, -23, 7, -83,
					-- layer=2 filter=14 channel=7
					-3, 30, -1, 8, 4, 4, -19, -9, -57,
					-- layer=2 filter=14 channel=8
					-8, -2, 0, -4, 2, 5, 7, -8, 0,
					-- layer=2 filter=14 channel=9
					-48, -54, -13, 20, -1, -16, 37, 43, 15,
					-- layer=2 filter=14 channel=10
					-21, -3, -37, 45, 7, 12, 55, -5, 35,
					-- layer=2 filter=14 channel=11
					-30, -10, 24, -33, -31, 21, -25, 10, 8,
					-- layer=2 filter=14 channel=12
					10, 1, 13, -15, 16, 24, 0, 14, -21,
					-- layer=2 filter=14 channel=13
					-7, -12, -4, -6, 9, -10, 4, -7, -6,
					-- layer=2 filter=14 channel=14
					-10, -22, 17, -11, 11, 7, -1, -1, -3,
					-- layer=2 filter=14 channel=15
					-81, 38, 18, -14, 42, 50, 45, -14, 53,
					-- layer=2 filter=14 channel=16
					23, 28, -41, 8, 18, -37, -12, -39, -22,
					-- layer=2 filter=14 channel=17
					-5, 3, 0, -6, -4, 3, -7, -1, -5,
					-- layer=2 filter=14 channel=18
					-3, 14, -1, -8, -11, 4, -36, 29, 41,
					-- layer=2 filter=14 channel=19
					38, 45, 63, -16, 5, 0, 2, 15, 9,
					-- layer=2 filter=14 channel=20
					3, 2, 3, 8, 7, 2, 7, 3, -11,
					-- layer=2 filter=14 channel=21
					19, -18, 0, 21, 19, -3, -14, 5, -16,
					-- layer=2 filter=14 channel=22
					11, 0, -7, 0, -1, -2, -10, -9, -8,
					-- layer=2 filter=14 channel=23
					11, 34, -7, 32, -20, -29, 23, -13, -14,
					-- layer=2 filter=14 channel=24
					32, 11, -37, 31, -9, -24, 67, 16, 8,
					-- layer=2 filter=14 channel=25
					-3, -22, -47, -59, -51, -39, -28, -34, -31,
					-- layer=2 filter=14 channel=26
					8, 2, -13, 1, -7, -10, -3, 3, 1,
					-- layer=2 filter=14 channel=27
					-26, 6, 47, -49, -11, 16, 4, -5, -19,
					-- layer=2 filter=14 channel=28
					-20, 9, -17, -4, 6, 5, -9, -11, -6,
					-- layer=2 filter=14 channel=29
					0, -1, -1, 6, -8, 5, -11, 2, 2,
					-- layer=2 filter=14 channel=30
					-12, -33, -8, -4, 5, -38, -10, -8, 5,
					-- layer=2 filter=14 channel=31
					-51, -63, -76, -8, -49, -1, 61, 26, 7,
					-- layer=2 filter=14 channel=32
					0, -11, 9, 3, -6, 9, -8, -5, 4,
					-- layer=2 filter=14 channel=33
					-61, -31, -30, -1, 3, -16, -2, -6, 18,
					-- layer=2 filter=14 channel=34
					-6, 33, 10, -18, 18, 8, -48, 38, 58,
					-- layer=2 filter=14 channel=35
					3, 21, 9, 11, 5, -7, -25, -5, -7,
					-- layer=2 filter=14 channel=36
					4, 12, -14, 2, 0, 9, 7, 6, -5,
					-- layer=2 filter=14 channel=37
					-18, -3, 39, -28, -13, 15, -7, -10, 8,
					-- layer=2 filter=14 channel=38
					-23, -23, 21, -20, 0, 17, -2, 1, -28,
					-- layer=2 filter=14 channel=39
					-9, 2, 9, 17, 4, -31, 37, -18, -19,
					-- layer=2 filter=14 channel=40
					41, 49, 12, -41, -38, -46, -18, 20, -1,
					-- layer=2 filter=14 channel=41
					-4, -1, 2, 9, -2, -3, 1, 5, -6,
					-- layer=2 filter=14 channel=42
					2, 2, -18, -3, 3, -20, 21, -18, -59,
					-- layer=2 filter=14 channel=43
					-39, 34, 91, -3, 14, 29, 32, 40, 46,
					-- layer=2 filter=14 channel=44
					-1, 0, 8, -8, 5, -3, -6, 9, 2,
					-- layer=2 filter=14 channel=45
					-18, -12, -38, -20, -7, -23, 18, -21, -45,
					-- layer=2 filter=14 channel=46
					-27, -20, -5, -37, -1, -11, 5, -14, -11,
					-- layer=2 filter=14 channel=47
					-24, 20, -39, 6, 13, -28, -21, -30, -13,
					-- layer=2 filter=14 channel=48
					-2, 3, -11, -3, 3, -3, -7, 5, -6,
					-- layer=2 filter=14 channel=49
					0, 6, -25, -94, -5, -9, -40, 10, -26,
					-- layer=2 filter=14 channel=50
					10, 19, 17, 29, 9, 1, 19, -1, -6,
					-- layer=2 filter=14 channel=51
					-4, -30, -4, -9, -23, 21, -10, -8, -28,
					-- layer=2 filter=14 channel=52
					46, -26, 17, 3, 10, 31, -23, 11, 0,
					-- layer=2 filter=14 channel=53
					-37, -33, -25, 4, -5, -4, 4, 27, -41,
					-- layer=2 filter=14 channel=54
					10, 7, -19, 0, 4, -2, -7, -5, -2,
					-- layer=2 filter=14 channel=55
					-9, 0, 4, -2, 13, 3, 3, 0, -7,
					-- layer=2 filter=14 channel=56
					-52, -17, 16, -26, -7, 37, 8, 4, 12,
					-- layer=2 filter=14 channel=57
					5, 1, 2, 12, 12, -11, -6, -1, 2,
					-- layer=2 filter=14 channel=58
					9, -13, -4, -12, 8, 5, -9, 40, 3,
					-- layer=2 filter=14 channel=59
					19, 5, 48, -15, 32, 6, -5, 44, 56,
					-- layer=2 filter=14 channel=60
					57, 4, 0, 19, 36, -9, 43, 23, -6,
					-- layer=2 filter=14 channel=61
					-1, -17, -8, 14, -4, 5, 20, -11, 5,
					-- layer=2 filter=14 channel=62
					23, 1, 7, -24, -15, -10, -57, 4, 20,
					-- layer=2 filter=14 channel=63
					-12, 7, 0, 23, -6, -12, 3, -12, -4,
					-- layer=2 filter=14 channel=64
					18, 32, -30, 16, 20, -54, 22, 12, -19,
					-- layer=2 filter=14 channel=65
					10, -46, 42, -19, 5, 22, -16, -21, -22,
					-- layer=2 filter=14 channel=66
					27, -53, -22, -7, -38, -6, 25, -16, -8,
					-- layer=2 filter=14 channel=67
					-33, -15, 20, -24, 16, 44, 29, 62, 80,
					-- layer=2 filter=14 channel=68
					-6, -2, -2, 7, -2, 3, 7, 1, -9,
					-- layer=2 filter=14 channel=69
					24, 31, 2, 35, 6, -47, 24, 2, -12,
					-- layer=2 filter=14 channel=70
					-15, -3, 10, 5, 20, -19, 3, -12, 1,
					-- layer=2 filter=14 channel=71
					-11, 35, 10, -50, 5, -4, -8, 1, 12,
					-- layer=2 filter=14 channel=72
					-17, 0, 5, 13, 16, 36, 0, -22, -2,
					-- layer=2 filter=14 channel=73
					-23, 23, 39, -37, -29, -23, 10, -8, -1,
					-- layer=2 filter=14 channel=74
					-32, -10, 17, -17, 16, 13, 1, -17, -11,
					-- layer=2 filter=14 channel=75
					-48, -1, -20, -28, -32, -39, -19, -18, -6,
					-- layer=2 filter=14 channel=76
					-42, -6, 21, 8, 9, -5, 16, -17, 4,
					-- layer=2 filter=14 channel=77
					-1, -5, -7, -11, -9, 7, -3, 0, 6,
					-- layer=2 filter=14 channel=78
					3, 13, 21, -46, -19, 16, -55, 2, 11,
					-- layer=2 filter=14 channel=79
					-7, -1, 1, -6, 3, -4, 3, -5, 7,
					-- layer=2 filter=14 channel=80
					-13, -5, -13, -4, -12, -44, 9, 26, -4,
					-- layer=2 filter=14 channel=81
					-2, 10, -1, -12, 7, -3, -2, 10, -9,
					-- layer=2 filter=14 channel=82
					-12, 1, -7, 0, 2, -5, -4, 6, -2,
					-- layer=2 filter=14 channel=83
					0, 8, 10, -1, -12, -13, 1, -8, -43,
					-- layer=2 filter=14 channel=84
					8, 1, 3, 7, 3, -9, 5, 0, 5,
					-- layer=2 filter=14 channel=85
					0, -8, 6, 0, 18, -4, 9, 0, -1,
					-- layer=2 filter=14 channel=86
					11, 4, -7, -5, 11, 0, 1, -14, 10,
					-- layer=2 filter=14 channel=87
					5, 20, -1, 43, 31, 49, -9, 28, 50,
					-- layer=2 filter=14 channel=88
					-12, 3, 39, 8, 8, 4, 20, -4, -31,
					-- layer=2 filter=14 channel=89
					-5, -1, 43, -33, 32, 34, -14, 18, 27,
					-- layer=2 filter=14 channel=90
					3, 7, -9, 0, -1, 4, 7, 8, 7,
					-- layer=2 filter=14 channel=91
					-10, 16, 5, -31, 1, 2, -19, -6, -18,
					-- layer=2 filter=14 channel=92
					11, 7, 45, -22, 30, 28, -22, 1, -13,
					-- layer=2 filter=14 channel=93
					39, -6, 17, -64, -25, -26, -27, -9, 9,
					-- layer=2 filter=14 channel=94
					-2, -21, -6, 36, -43, -16, 27, 20, -17,
					-- layer=2 filter=14 channel=95
					2, 14, 9, -10, 7, -4, 5, -2, 9,
					-- layer=2 filter=14 channel=96
					17, 15, 15, 1, -74, -28, -95, -41, -8,
					-- layer=2 filter=14 channel=97
					-22, -30, -44, -19, -38, -84, 15, -3, -51,
					-- layer=2 filter=14 channel=98
					0, 5, -6, 7, 10, 16, 8, -12, 3,
					-- layer=2 filter=14 channel=99
					35, 14, 13, 4, 8, -20, 33, 15, -13,
					-- layer=2 filter=14 channel=100
					-11, -28, 2, 2, 20, -11, 19, 5, 26,
					-- layer=2 filter=14 channel=101
					-38, -22, -6, -68, -33, -58, -18, -37, -8,
					-- layer=2 filter=14 channel=102
					26, 22, -20, -30, -51, -14, -30, 12, 29,
					-- layer=2 filter=14 channel=103
					7, 61, 17, -16, 22, 5, 24, -11, -6,
					-- layer=2 filter=14 channel=104
					-23, 8, -22, -32, -34, 5, -34, 33, -13,
					-- layer=2 filter=14 channel=105
					25, -22, -28, 23, 46, 14, -19, -46, 70,
					-- layer=2 filter=14 channel=106
					-50, -24, -59, -34, -36, -49, 0, -18, -35,
					-- layer=2 filter=14 channel=107
					7, 2, -14, -11, -47, 0, 36, 9, -11,
					-- layer=2 filter=14 channel=108
					21, 10, -8, -21, -7, -37, -9, -31, -45,
					-- layer=2 filter=14 channel=109
					-12, 4, -9, -6, 0, -6, -1, -5, 0,
					-- layer=2 filter=14 channel=110
					27, 28, -12, 13, 16, 4, -2, -29, -36,
					-- layer=2 filter=14 channel=111
					-7, -10, -9, 8, -7, 0, -8, 2, 0,
					-- layer=2 filter=14 channel=112
					0, 14, -4, -36, -26, -23, 26, -1, 26,
					-- layer=2 filter=14 channel=113
					7, -6, -27, -15, 7, -23, -31, -14, -3,
					-- layer=2 filter=14 channel=114
					3, 6, -7, -8, 4, -1, -3, -15, -25,
					-- layer=2 filter=14 channel=115
					7, 6, 6, 0, 1, -3, -3, -6, 1,
					-- layer=2 filter=14 channel=116
					-1, 42, 7, 41, 13, 47, -18, 39, 58,
					-- layer=2 filter=14 channel=117
					21, 10, 25, -1, -9, -14, 9, 0, -1,
					-- layer=2 filter=14 channel=118
					-8, 11, 5, 4, 36, 14, -10, 23, 29,
					-- layer=2 filter=14 channel=119
					-22, 31, 2, 1, -10, -41, -39, -20, 0,
					-- layer=2 filter=14 channel=120
					0, 3, -7, 3, -3, 0, -9, -2, 3,
					-- layer=2 filter=14 channel=121
					0, -1, 3, -6, -7, 9, -9, 8, -4,
					-- layer=2 filter=14 channel=122
					7, 1, -8, 14, 1, 0, 0, 12, -4,
					-- layer=2 filter=14 channel=123
					21, 11, -27, 30, 28, 29, 0, 9, 9,
					-- layer=2 filter=14 channel=124
					1, 40, 47, 48, 47, 36, 36, 16, 53,
					-- layer=2 filter=14 channel=125
					0, -3, -4, -9, 7, 6, 1, -7, 5,
					-- layer=2 filter=14 channel=126
					7, -39, 1, 1, -43, -26, -46, -16, 14,
					-- layer=2 filter=14 channel=127
					14, -8, 26, -11, 43, 1, -23, -2, -15,
					-- layer=2 filter=15 channel=0
					-26, -16, -17, -50, -55, -50, -35, -62, 12,
					-- layer=2 filter=15 channel=1
					-19, -16, -66, 19, -11, 7, 12, 27, 36,
					-- layer=2 filter=15 channel=2
					0, 5, -9, 3, -4, -5, -11, -8, 6,
					-- layer=2 filter=15 channel=3
					-25, -16, 0, 35, -8, -9, 28, 13, 2,
					-- layer=2 filter=15 channel=4
					-33, -6, -17, -26, 19, -50, 3, 9, -21,
					-- layer=2 filter=15 channel=5
					6, 6, 28, -37, -35, -15, -8, 5, -4,
					-- layer=2 filter=15 channel=6
					3, -3, -50, 23, 12, -5, 0, 7, 11,
					-- layer=2 filter=15 channel=7
					34, -19, 0, -55, -11, 12, -57, -57, 0,
					-- layer=2 filter=15 channel=8
					-4, 6, -7, -4, -1, -1, 6, 10, 7,
					-- layer=2 filter=15 channel=9
					-4, -21, -2, 50, -32, -24, 52, -17, -34,
					-- layer=2 filter=15 channel=10
					-29, -32, -2, -41, -37, -38, -3, 9, -10,
					-- layer=2 filter=15 channel=11
					18, 17, 11, -11, 6, -5, -13, -20, 18,
					-- layer=2 filter=15 channel=12
					-4, -1, -40, 3, -22, 14, -6, 7, -13,
					-- layer=2 filter=15 channel=13
					5, -8, 1, -8, -5, 6, -11, 0, 4,
					-- layer=2 filter=15 channel=14
					5, 6, -17, -7, -10, 12, -3, 9, 21,
					-- layer=2 filter=15 channel=15
					-28, -5, 15, -21, 7, -45, 39, 2, 21,
					-- layer=2 filter=15 channel=16
					-9, -5, -30, 32, 47, -9, 29, 37, -18,
					-- layer=2 filter=15 channel=17
					-2, -4, -9, 7, 7, 2, -2, -8, 9,
					-- layer=2 filter=15 channel=18
					9, -9, 16, -23, -4, 7, -1, 0, -36,
					-- layer=2 filter=15 channel=19
					-25, -41, -19, 41, -2, -12, 35, 7, 5,
					-- layer=2 filter=15 channel=20
					0, 8, -10, -5, -6, -5, 1, -4, 0,
					-- layer=2 filter=15 channel=21
					0, 9, 14, -3, -2, 14, 8, 12, -5,
					-- layer=2 filter=15 channel=22
					10, -3, -3, -2, 0, -3, -4, 7, 1,
					-- layer=2 filter=15 channel=23
					22, 8, -9, 30, 31, -17, 1, 17, 35,
					-- layer=2 filter=15 channel=24
					19, 19, 35, 15, 12, 14, -6, -23, -20,
					-- layer=2 filter=15 channel=25
					16, 43, 28, 8, 13, 16, -20, -20, -19,
					-- layer=2 filter=15 channel=26
					6, 7, 1, 0, 0, 9, -9, -9, 9,
					-- layer=2 filter=15 channel=27
					6, -23, -23, 7, -26, -37, 9, -43, -41,
					-- layer=2 filter=15 channel=28
					-10, -23, 1, -43, -16, -7, -25, -48, 5,
					-- layer=2 filter=15 channel=29
					-1, -6, 5, 0, -4, 2, -8, 6, 0,
					-- layer=2 filter=15 channel=30
					20, -26, -65, 22, 5, 0, -21, 70, -21,
					-- layer=2 filter=15 channel=31
					-29, -39, -36, -33, 37, 15, 9, 59, -19,
					-- layer=2 filter=15 channel=32
					-7, -9, 8, 4, 8, 0, 0, -1, -7,
					-- layer=2 filter=15 channel=33
					-16, -28, 9, -30, -65, -58, -3, -70, -29,
					-- layer=2 filter=15 channel=34
					-10, -9, -38, 21, 13, 39, -40, 29, -25,
					-- layer=2 filter=15 channel=35
					7, 2, 17, 5, 3, -16, -52, 12, 11,
					-- layer=2 filter=15 channel=36
					0, -13, -6, 15, -14, -16, -1, 0, -5,
					-- layer=2 filter=15 channel=37
					-8, 0, -1, 13, 9, 3, 14, -23, 22,
					-- layer=2 filter=15 channel=38
					12, -41, -66, -8, -50, -33, -15, -31, -33,
					-- layer=2 filter=15 channel=39
					-9, 3, -27, 19, 3, -23, -17, 30, -41,
					-- layer=2 filter=15 channel=40
					36, 33, 1, -5, -68, 24, -1, -15, -25,
					-- layer=2 filter=15 channel=41
					-6, 0, -8, -1, 0, 4, -1, 5, 0,
					-- layer=2 filter=15 channel=42
					-7, -2, -14, 38, 35, 16, 22, 26, 13,
					-- layer=2 filter=15 channel=43
					16, 6, -21, 39, -31, -49, 48, -54, -45,
					-- layer=2 filter=15 channel=44
					5, -8, -9, 8, 5, 0, 3, -6, -8,
					-- layer=2 filter=15 channel=45
					17, -60, -67, -6, -81, -51, -7, -24, -47,
					-- layer=2 filter=15 channel=46
					17, -102, -51, -23, -69, -47, -27, -23, -61,
					-- layer=2 filter=15 channel=47
					-31, -9, 0, -84, -57, -23, -2, -32, -24,
					-- layer=2 filter=15 channel=48
					-4, 7, -6, 5, 9, 0, -3, -2, -9,
					-- layer=2 filter=15 channel=49
					4, -46, 11, 62, -35, 19, 71, -10, 17,
					-- layer=2 filter=15 channel=50
					7, -10, -17, -13, 2, 13, 7, -4, 0,
					-- layer=2 filter=15 channel=51
					-8, 9, 0, -17, -18, -1, -33, -20, 8,
					-- layer=2 filter=15 channel=52
					21, -6, -39, -34, -2, -36, 15, -7, -19,
					-- layer=2 filter=15 channel=53
					-34, -52, -37, -10, -1, 12, -75, 7, 16,
					-- layer=2 filter=15 channel=54
					8, -7, 10, -26, -40, -6, -45, -43, 11,
					-- layer=2 filter=15 channel=55
					0, -1, 4, 3, -3, 3, -9, -5, -4,
					-- layer=2 filter=15 channel=56
					29, 16, 17, 5, -11, -11, 11, -1, 7,
					-- layer=2 filter=15 channel=57
					4, -5, 8, 3, 4, -11, -1, 8, -2,
					-- layer=2 filter=15 channel=58
					15, 18, -48, 14, -10, 7, -55, 6, -14,
					-- layer=2 filter=15 channel=59
					8, -57, -49, -12, -32, 7, -79, -48, 29,
					-- layer=2 filter=15 channel=60
					1, 18, -6, -40, -42, 29, -27, 4, -34,
					-- layer=2 filter=15 channel=61
					38, -5, 24, -64, 45, -8, -82, -39, 38,
					-- layer=2 filter=15 channel=62
					-16, -19, -40, 57, 7, 11, 43, -13, 40,
					-- layer=2 filter=15 channel=63
					18, -8, -11, -3, 10, -31, -6, 0, -8,
					-- layer=2 filter=15 channel=64
					-16, -18, 9, 23, 21, 0, 2, 5, 9,
					-- layer=2 filter=15 channel=65
					61, -27, 0, -5, 27, -13, 4, 6, 18,
					-- layer=2 filter=15 channel=66
					41, 18, 65, -18, 38, 34, 7, 18, 25,
					-- layer=2 filter=15 channel=67
					5, 2, -51, -3, -59, -77, -5, 3, -45,
					-- layer=2 filter=15 channel=68
					8, 7, 4, -3, -5, -7, 4, 6, 1,
					-- layer=2 filter=15 channel=69
					-19, 11, 8, 54, 31, 8, 18, 49, 5,
					-- layer=2 filter=15 channel=70
					19, 2, -1, -13, 4, -36, -38, 0, -22,
					-- layer=2 filter=15 channel=71
					44, 36, -6, 42, 18, -56, -10, -9, -52,
					-- layer=2 filter=15 channel=72
					3, -68, -9, -6, 11, 19, -2, -12, 34,
					-- layer=2 filter=15 channel=73
					30, 27, -4, 23, 61, 34, 39, 14, 14,
					-- layer=2 filter=15 channel=74
					-3, -32, -48, -11, -59, -73, -53, 2, -44,
					-- layer=2 filter=15 channel=75
					69, 40, 72, -10, -39, -13, 14, 12, -2,
					-- layer=2 filter=15 channel=76
					-27, 7, -29, -63, 15, 9, -66, -11, 39,
					-- layer=2 filter=15 channel=77
					-3, -7, -6, 4, -5, 5, 7, -4, 4,
					-- layer=2 filter=15 channel=78
					-7, -9, 15, -18, 2, -12, -25, -68, -8,
					-- layer=2 filter=15 channel=79
					6, -6, -10, 0, 0, 2, 7, -11, -1,
					-- layer=2 filter=15 channel=80
					-36, -37, -19, 17, 18, -30, 29, 36, -19,
					-- layer=2 filter=15 channel=81
					-8, -11, 3, -4, -9, 0, -9, -4, -5,
					-- layer=2 filter=15 channel=82
					10, 1, -3, 10, 1, -1, 7, -5, -4,
					-- layer=2 filter=15 channel=83
					1, -28, -9, 25, 39, -48, 6, 52, 37,
					-- layer=2 filter=15 channel=84
					-10, -7, -8, 8, -3, -9, 4, -9, -10,
					-- layer=2 filter=15 channel=85
					-13, -1, -5, -1, -3, 3, 14, -4, -6,
					-- layer=2 filter=15 channel=86
					-6, 0, 19, 8, 0, 17, 8, 6, 0,
					-- layer=2 filter=15 channel=87
					20, -5, -8, 26, -36, 37, 1, -28, 24,
					-- layer=2 filter=15 channel=88
					17, -11, -23, 26, -7, 7, -39, 30, 5,
					-- layer=2 filter=15 channel=89
					14, -27, -20, -11, -5, -3, -12, -14, 38,
					-- layer=2 filter=15 channel=90
					-8, -4, 10, 9, -1, 5, 0, -3, 5,
					-- layer=2 filter=15 channel=91
					-21, 11, -5, 29, -24, 2, -34, -18, -18,
					-- layer=2 filter=15 channel=92
					-1, -2, -80, 19, -29, -1, 2, 19, 1,
					-- layer=2 filter=15 channel=93
					40, -11, -17, 60, 37, -7, 68, 48, 35,
					-- layer=2 filter=15 channel=94
					36, 21, 18, 18, 11, 16, -44, -45, 68,
					-- layer=2 filter=15 channel=95
					-2, -17, 12, 0, 14, -20, 5, -5, -8,
					-- layer=2 filter=15 channel=96
					-7, 19, 22, -14, -28, -10, 18, -49, 65,
					-- layer=2 filter=15 channel=97
					-40, -42, 35, 20, -31, -48, 34, -45, -70,
					-- layer=2 filter=15 channel=98
					-17, -29, 33, -38, 0, -14, -39, -63, 8,
					-- layer=2 filter=15 channel=99
					-9, -7, 0, -12, -1, -12, -42, -64, -13,
					-- layer=2 filter=15 channel=100
					0, -2, -38, 17, -10, -65, 6, 18, -30,
					-- layer=2 filter=15 channel=101
					61, 53, 13, 20, 15, -25, -7, -3, -45,
					-- layer=2 filter=15 channel=102
					16, 43, 31, -21, 5, 2, 50, 3, 33,
					-- layer=2 filter=15 channel=103
					-17, -41, -37, -44, -13, 29, 4, 9, -14,
					-- layer=2 filter=15 channel=104
					13, -3, 13, 13, -5, 36, 19, -33, 47,
					-- layer=2 filter=15 channel=105
					-24, -29, 17, -69, 57, 0, -30, -91, 49,
					-- layer=2 filter=15 channel=106
					19, 38, 27, -14, 23, -9, -17, 5, 2,
					-- layer=2 filter=15 channel=107
					46, -16, -28, 6, 0, 45, 24, 27, 2,
					-- layer=2 filter=15 channel=108
					8, -10, -20, 4, 12, -3, 39, 15, 43,
					-- layer=2 filter=15 channel=109
					2, -3, 14, 10, -22, 0, -15, -14, 8,
					-- layer=2 filter=15 channel=110
					58, 1, 27, 52, 49, 42, 7, -2, 7,
					-- layer=2 filter=15 channel=111
					-7, 5, 0, 0, 6, 0, 7, -2, -10,
					-- layer=2 filter=15 channel=112
					11, -8, 25, -29, -19, -75, -51, -55, -46,
					-- layer=2 filter=15 channel=113
					25, -51, 1, 33, 37, -20, -44, 27, -9,
					-- layer=2 filter=15 channel=114
					-4, -8, -1, -9, -10, 12, 0, 0, 3,
					-- layer=2 filter=15 channel=115
					-5, 3, 1, -3, 7, -8, -7, 0, -3,
					-- layer=2 filter=15 channel=116
					-16, -13, -12, 0, -28, -20, -3, -27, 20,
					-- layer=2 filter=15 channel=117
					28, 8, -24, -19, -14, 10, -30, -40, 7,
					-- layer=2 filter=15 channel=118
					-59, -36, -6, 7, 4, -33, 66, -28, -17,
					-- layer=2 filter=15 channel=119
					-10, -6, 21, 7, 4, -16, 26, 18, -40,
					-- layer=2 filter=15 channel=120
					-3, -1, 10, 0, 0, 5, 1, 0, 5,
					-- layer=2 filter=15 channel=121
					-9, -3, -3, -1, -4, -6, 1, 6, 1,
					-- layer=2 filter=15 channel=122
					-6, -5, -9, 0, 5, 9, -8, 0, -6,
					-- layer=2 filter=15 channel=123
					22, -25, 28, -35, -1, -3, -27, -57, 36,
					-- layer=2 filter=15 channel=124
					-31, -11, -8, -28, -6, -31, 17, 0, 11,
					-- layer=2 filter=15 channel=125
					0, 4, 5, 0, -7, -10, 5, -1, -1,
					-- layer=2 filter=15 channel=126
					25, 13, -11, -6, -5, -23, -26, -49, 0,
					-- layer=2 filter=15 channel=127
					0, -20, -37, 12, 12, -13, -20, 9, -23,
					-- layer=2 filter=16 channel=0
					-24, 4, 5, -40, 15, 21, 11, -2, -10,
					-- layer=2 filter=16 channel=1
					-6, -10, -45, 19, 30, -34, 6, -1, 3,
					-- layer=2 filter=16 channel=2
					3, 5, 5, 2, 7, 0, -7, 1, -10,
					-- layer=2 filter=16 channel=3
					-37, 10, 65, -79, 15, 51, -7, -41, 19,
					-- layer=2 filter=16 channel=4
					-11, 0, -11, -7, 9, -23, -23, -29, -28,
					-- layer=2 filter=16 channel=5
					28, -27, -12, 6, 0, 19, 8, -4, -6,
					-- layer=2 filter=16 channel=6
					-33, -53, -23, 34, 3, -19, 5, 32, -5,
					-- layer=2 filter=16 channel=7
					5, 21, 36, 44, 36, -12, 8, -35, 18,
					-- layer=2 filter=16 channel=8
					-6, 10, -9, 3, -2, 2, -5, 4, 7,
					-- layer=2 filter=16 channel=9
					-18, 21, 47, -16, 0, 42, 0, 1, 6,
					-- layer=2 filter=16 channel=10
					-19, 11, 30, -32, -9, 4, 9, 6, 4,
					-- layer=2 filter=16 channel=11
					5, 0, -16, 9, 8, -2, -10, -7, -26,
					-- layer=2 filter=16 channel=12
					0, -17, -58, 16, 4, -22, 1, -2, -33,
					-- layer=2 filter=16 channel=13
					2, 11, -5, -4, -5, 8, 1, 7, 7,
					-- layer=2 filter=16 channel=14
					23, -10, -28, 16, 29, -9, -17, -7, -26,
					-- layer=2 filter=16 channel=15
					35, -34, -38, 24, 8, 33, 5, 12, -1,
					-- layer=2 filter=16 channel=16
					-14, 16, 20, -56, -50, 17, -2, -31, -9,
					-- layer=2 filter=16 channel=17
					8, -10, 9, 0, -2, 1, -6, 5, 0,
					-- layer=2 filter=16 channel=18
					27, -19, -9, 36, 18, 6, -13, 9, -47,
					-- layer=2 filter=16 channel=19
					28, 9, -6, 40, 38, -23, 5, 30, 6,
					-- layer=2 filter=16 channel=20
					-7, -3, 7, 9, 10, 9, 8, 1, 2,
					-- layer=2 filter=16 channel=21
					-1, 7, -4, -6, -7, -8, -3, -18, -13,
					-- layer=2 filter=16 channel=22
					3, -3, 10, 6, -2, 3, 0, 12, -10,
					-- layer=2 filter=16 channel=23
					-13, 17, 17, -8, -2, 1, 14, -5, -14,
					-- layer=2 filter=16 channel=24
					-43, 19, 62, -66, -12, 37, -44, -33, 54,
					-- layer=2 filter=16 channel=25
					-24, -4, 27, -33, -25, 2, -25, -22, 27,
					-- layer=2 filter=16 channel=26
					-5, -3, 5, -9, -8, -10, -8, -3, -8,
					-- layer=2 filter=16 channel=27
					28, 10, -26, 26, 7, -47, 5, 0, -29,
					-- layer=2 filter=16 channel=28
					-2, 12, -2, -5, -14, 17, 10, -7, -2,
					-- layer=2 filter=16 channel=29
					-8, -9, 7, 7, -5, -7, -1, 5, 4,
					-- layer=2 filter=16 channel=30
					1, -9, -5, 20, 14, 4, -19, -21, -14,
					-- layer=2 filter=16 channel=31
					40, -37, -4, 35, -13, -85, -35, -29, 5,
					-- layer=2 filter=16 channel=32
					1, 0, -6, 5, 7, 6, -9, 3, 8,
					-- layer=2 filter=16 channel=33
					-8, -13, 10, -2, 3, 4, 14, 2, 26,
					-- layer=2 filter=16 channel=34
					23, -4, -27, 19, 0, 3, 16, 25, -47,
					-- layer=2 filter=16 channel=35
					5, -3, 1, 21, 0, -9, 5, -12, -80,
					-- layer=2 filter=16 channel=36
					-5, 0, 2, -20, -3, -10, -7, 3, -7,
					-- layer=2 filter=16 channel=37
					36, -6, -10, 14, 1, 0, -8, 18, -15,
					-- layer=2 filter=16 channel=38
					31, -26, -50, 17, -14, -19, 4, -12, -15,
					-- layer=2 filter=16 channel=39
					-23, 23, 20, -29, -15, 14, 17, -28, -6,
					-- layer=2 filter=16 channel=40
					21, 4, -4, -2, -13, 65, -41, -8, 24,
					-- layer=2 filter=16 channel=41
					10, -3, -9, 11, -1, 10, 1, 11, 6,
					-- layer=2 filter=16 channel=42
					-18, 5, 20, -10, -11, 7, 4, -14, -16,
					-- layer=2 filter=16 channel=43
					-28, 1, 10, -19, -2, 13, -9, 21, -12,
					-- layer=2 filter=16 channel=44
					4, -6, -7, 8, 2, -7, 1, -1, 0,
					-- layer=2 filter=16 channel=45
					51, 16, -20, 3, -25, -81, 26, -15, -24,
					-- layer=2 filter=16 channel=46
					3, -8, 23, -42, -26, 7, -37, -5, 19,
					-- layer=2 filter=16 channel=47
					41, 21, -14, -11, 12, 7, -4, -33, 14,
					-- layer=2 filter=16 channel=48
					-5, 12, -8, -3, -4, 3, -4, -7, 3,
					-- layer=2 filter=16 channel=49
					10, -9, 8, 28, 24, -18, 2, 33, -58,
					-- layer=2 filter=16 channel=50
					10, 15, 10, -14, 11, 10, 27, -15, 0,
					-- layer=2 filter=16 channel=51
					-12, -7, -1, -6, 13, -13, -6, -3, -9,
					-- layer=2 filter=16 channel=52
					17, 12, -34, 9, 20, 0, 32, 12, -10,
					-- layer=2 filter=16 channel=53
					44, 20, 19, 14, 26, 12, 1, 0, 3,
					-- layer=2 filter=16 channel=54
					34, 5, -13, 35, 21, -22, 30, -13, -19,
					-- layer=2 filter=16 channel=55
					0, -5, 2, 4, -9, -10, -6, -1, 11,
					-- layer=2 filter=16 channel=56
					-18, -16, -5, 5, 11, -16, -22, -11, -3,
					-- layer=2 filter=16 channel=57
					-18, 9, -9, -10, 6, 0, 8, -12, 2,
					-- layer=2 filter=16 channel=58
					24, 10, -45, 8, 13, 6, 25, -4, -38,
					-- layer=2 filter=16 channel=59
					13, -18, -49, 40, 2, -43, -12, -27, -10,
					-- layer=2 filter=16 channel=60
					38, -42, -21, 9, -4, -31, 15, 34, -10,
					-- layer=2 filter=16 channel=61
					-21, 4, 22, 54, 0, 10, 16, 6, -6,
					-- layer=2 filter=16 channel=62
					12, -13, -27, 15, 12, -17, 5, 18, -19,
					-- layer=2 filter=16 channel=63
					-6, 21, 16, -1, 4, 18, -8, -4, -40,
					-- layer=2 filter=16 channel=64
					-46, 9, 26, -25, -29, 8, -7, 3, -10,
					-- layer=2 filter=16 channel=65
					-3, -34, 14, 32, -15, -13, 6, -9, 18,
					-- layer=2 filter=16 channel=66
					-38, 42, -38, 20, -12, -38, 33, -6, -9,
					-- layer=2 filter=16 channel=67
					-26, -8, 31, -39, -27, 67, -3, -28, 42,
					-- layer=2 filter=16 channel=68
					6, 8, 5, 10, 0, 2, 3, -2, 2,
					-- layer=2 filter=16 channel=69
					-34, 15, 18, -40, -7, 7, -26, -20, -15,
					-- layer=2 filter=16 channel=70
					24, -8, -42, 30, 14, -4, 16, -1, -82,
					-- layer=2 filter=16 channel=71
					30, 29, -13, 43, 1, -10, 20, 4, 21,
					-- layer=2 filter=16 channel=72
					0, -27, 10, 22, 6, -51, -18, -23, 36,
					-- layer=2 filter=16 channel=73
					14, 5, 23, 31, 28, -24, 30, -27, -30,
					-- layer=2 filter=16 channel=74
					-14, 13, 1, -50, -23, 21, -15, -10, -50,
					-- layer=2 filter=16 channel=75
					15, 4, -10, 40, 26, 30, -25, -79, -66,
					-- layer=2 filter=16 channel=76
					22, -23, -15, -18, 1, 19, 7, -20, -37,
					-- layer=2 filter=16 channel=77
					5, -1, -9, 8, 1, -5, 9, -3, -4,
					-- layer=2 filter=16 channel=78
					-1, -24, 2, -19, 19, 3, -11, 1, 5,
					-- layer=2 filter=16 channel=79
					6, -4, 0, -2, 6, 10, 5, -4, -6,
					-- layer=2 filter=16 channel=80
					-16, 16, 33, -65, -37, 11, -25, 16, -3,
					-- layer=2 filter=16 channel=81
					2, -6, -14, -6, -4, -3, 13, 10, -4,
					-- layer=2 filter=16 channel=82
					5, 5, -7, 1, -4, 1, 2, -4, 9,
					-- layer=2 filter=16 channel=83
					-6, 1, -5, 12, -29, -31, 13, -8, -46,
					-- layer=2 filter=16 channel=84
					4, 3, 3, 7, 7, 12, 7, -6, 4,
					-- layer=2 filter=16 channel=85
					1, 2, -4, -3, 6, 0, -8, -3, 2,
					-- layer=2 filter=16 channel=86
					10, 0, 13, 0, 27, -6, 9, 9, -4,
					-- layer=2 filter=16 channel=87
					0, -31, -22, -2, -9, -10, 26, -11, 1,
					-- layer=2 filter=16 channel=88
					-18, -13, 19, -7, -19, 19, 10, -16, -48,
					-- layer=2 filter=16 channel=89
					2, -30, -20, 29, 34, -25, 0, 4, -1,
					-- layer=2 filter=16 channel=90
					7, 7, -10, 9, 2, 6, 0, -4, 8,
					-- layer=2 filter=16 channel=91
					9, -26, -47, 11, -14, -1, 5, 0, 13,
					-- layer=2 filter=16 channel=92
					7, -25, -38, 53, 16, -27, 2, -14, 12,
					-- layer=2 filter=16 channel=93
					-34, -12, -29, -26, -31, -36, 50, -13, -40,
					-- layer=2 filter=16 channel=94
					-15, 19, -11, 48, 59, 38, 2, 30, 28,
					-- layer=2 filter=16 channel=95
					12, 14, 6, 6, -7, -7, 5, -2, 4,
					-- layer=2 filter=16 channel=96
					15, -2, -31, 29, 21, 10, 22, 24, 8,
					-- layer=2 filter=16 channel=97
					-25, 3, 49, -52, 6, 38, -75, -43, -1,
					-- layer=2 filter=16 channel=98
					17, 16, -1, -1, -27, -6, 8, -30, -11,
					-- layer=2 filter=16 channel=99
					37, -24, -29, 32, 17, -9, 28, 8, 0,
					-- layer=2 filter=16 channel=100
					-6, -10, -38, -4, -38, -21, 8, 24, -51,
					-- layer=2 filter=16 channel=101
					23, 24, 17, -9, -4, -2, 1, -5, 3,
					-- layer=2 filter=16 channel=102
					17, -8, 13, 6, 51, 20, 0, 0, 0,
					-- layer=2 filter=16 channel=103
					-4, -24, 8, 33, -12, 35, 36, 26, 11,
					-- layer=2 filter=16 channel=104
					2, -8, -6, 36, 29, 5, 6, -8, 4,
					-- layer=2 filter=16 channel=105
					54, 27, -1, 11, -49, 0, 15, -11, -38,
					-- layer=2 filter=16 channel=106
					-3, -6, 7, -37, -22, -4, -32, -33, 17,
					-- layer=2 filter=16 channel=107
					-15, -15, -15, -19, 0, -25, -25, 5, -18,
					-- layer=2 filter=16 channel=108
					9, 3, -15, 12, 13, -17, 2, 6, -22,
					-- layer=2 filter=16 channel=109
					-17, 3, -6, -10, -10, -1, -8, -9, 10,
					-- layer=2 filter=16 channel=110
					-25, -21, 35, 26, 2, 43, 15, 9, 28,
					-- layer=2 filter=16 channel=111
					11, 4, 0, 0, 1, 4, 9, -4, 3,
					-- layer=2 filter=16 channel=112
					-9, -5, 9, 0, -29, 4, -22, -10, 11,
					-- layer=2 filter=16 channel=113
					-10, 25, 1, -1, 18, -12, -12, -27, 4,
					-- layer=2 filter=16 channel=114
					5, 17, 11, 15, 5, 11, -6, 8, -1,
					-- layer=2 filter=16 channel=115
					4, -7, -5, 1, -2, 2, 0, 3, 4,
					-- layer=2 filter=16 channel=116
					35, 2, 0, 6, -12, 19, 27, 24, 2,
					-- layer=2 filter=16 channel=117
					-4, 35, -6, 15, 7, -47, 14, -69, -9,
					-- layer=2 filter=16 channel=118
					-5, 9, 48, -48, 3, 39, 10, 32, 5,
					-- layer=2 filter=16 channel=119
					-4, -3, -2, -2, 18, 22, 6, -33, -39,
					-- layer=2 filter=16 channel=120
					-7, -8, -7, 1, 0, 10, 4, 4, 1,
					-- layer=2 filter=16 channel=121
					7, 5, -10, -3, -6, -5, -2, 2, -6,
					-- layer=2 filter=16 channel=122
					-12, -2, 3, 9, 0, 5, 5, 5, 0,
					-- layer=2 filter=16 channel=123
					19, -6, 2, -1, 2, -49, -17, -29, 36,
					-- layer=2 filter=16 channel=124
					-25, -26, -7, -4, 19, -10, 22, 1, 2,
					-- layer=2 filter=16 channel=125
					2, -4, 6, -7, 3, -4, 12, -10, -5,
					-- layer=2 filter=16 channel=126
					10, -30, 21, 12, -23, 26, -2, -12, -7,
					-- layer=2 filter=16 channel=127
					5, 18, -1, 4, 15, -15, -9, -3, -41,
					-- layer=2 filter=17 channel=0
					-7, -13, -35, -21, -23, 0, 0, -14, -21,
					-- layer=2 filter=17 channel=1
					-3, -1, 6, 15, -4, 10, 3, 2, -12,
					-- layer=2 filter=17 channel=2
					-8, -3, 6, -9, -6, -9, 11, 5, -5,
					-- layer=2 filter=17 channel=3
					1, -15, -14, 8, 5, 11, 13, 0, 14,
					-- layer=2 filter=17 channel=4
					-5, -10, -17, -1, -14, -14, -21, -7, -3,
					-- layer=2 filter=17 channel=5
					-18, 0, -17, -10, -25, -17, -20, -1, -11,
					-- layer=2 filter=17 channel=6
					-11, -17, 1, 7, 0, 5, -9, -11, -2,
					-- layer=2 filter=17 channel=7
					-5, -13, -16, -4, -3, 2, 4, 9, -11,
					-- layer=2 filter=17 channel=8
					-8, 1, 7, -4, -6, -8, 8, 1, 0,
					-- layer=2 filter=17 channel=9
					-12, -15, -1, 19, 13, -10, 1, -4, 9,
					-- layer=2 filter=17 channel=10
					13, -16, -15, -6, 0, -21, -2, -17, -11,
					-- layer=2 filter=17 channel=11
					-19, -20, -22, -9, -16, -5, -12, -18, -18,
					-- layer=2 filter=17 channel=12
					-12, 2, 2, 0, -15, -15, 6, 12, -6,
					-- layer=2 filter=17 channel=13
					-2, 0, 4, 2, 1, -5, 8, -4, 9,
					-- layer=2 filter=17 channel=14
					-13, 0, -15, 0, -10, -12, 5, -5, 1,
					-- layer=2 filter=17 channel=15
					-6, -16, -24, 2, 2, -12, 0, -1, 14,
					-- layer=2 filter=17 channel=16
					-9, -17, -4, -22, -11, 7, -20, -6, 0,
					-- layer=2 filter=17 channel=17
					2, 0, -8, -9, -2, 6, 11, 3, 7,
					-- layer=2 filter=17 channel=18
					-12, -20, -33, -8, -11, -4, -9, 1, -14,
					-- layer=2 filter=17 channel=19
					-3, -5, -4, -1, -9, 3, -23, -11, 11,
					-- layer=2 filter=17 channel=20
					-8, 9, -6, 7, 8, 9, 10, -6, 7,
					-- layer=2 filter=17 channel=21
					-1, -8, 3, 1, 1, 5, -7, 7, -1,
					-- layer=2 filter=17 channel=22
					-6, -1, 3, 5, 0, 0, 7, -4, -4,
					-- layer=2 filter=17 channel=23
					-2, -5, -6, -6, -20, -10, -21, -12, -4,
					-- layer=2 filter=17 channel=24
					-13, -7, -5, -19, -2, -2, -15, 3, 0,
					-- layer=2 filter=17 channel=25
					-15, -9, -2, -13, -20, -14, 0, -3, 3,
					-- layer=2 filter=17 channel=26
					3, -2, -3, -6, 8, -9, -4, -3, 8,
					-- layer=2 filter=17 channel=27
					-15, -13, -5, -21, -18, -11, -9, -12, 1,
					-- layer=2 filter=17 channel=28
					15, 5, 0, 0, -14, -4, -13, -18, 10,
					-- layer=2 filter=17 channel=29
					4, -8, 1, 2, 7, -1, -5, 9, 0,
					-- layer=2 filter=17 channel=30
					-11, -1, -16, -14, 4, -35, -3, -12, -15,
					-- layer=2 filter=17 channel=31
					-19, -4, -17, -13, 7, -18, -13, -19, 0,
					-- layer=2 filter=17 channel=32
					4, -11, 8, 1, 2, 8, 0, -7, -10,
					-- layer=2 filter=17 channel=33
					-8, -18, 11, -9, 3, -11, 4, 19, -4,
					-- layer=2 filter=17 channel=34
					0, -5, -28, 2, -11, -28, -10, -23, -17,
					-- layer=2 filter=17 channel=35
					17, 28, -4, 0, -12, -11, -6, -16, -7,
					-- layer=2 filter=17 channel=36
					10, 8, 7, 1, 2, 3, -10, 0, -7,
					-- layer=2 filter=17 channel=37
					-15, -11, -14, -14, -28, -2, -10, -24, -10,
					-- layer=2 filter=17 channel=38
					-32, -10, -4, -9, -16, -2, -28, -17, -7,
					-- layer=2 filter=17 channel=39
					-17, -17, 1, 7, -8, -2, 12, -1, -13,
					-- layer=2 filter=17 channel=40
					-5, -17, 3, 4, -10, -4, -10, 10, -7,
					-- layer=2 filter=17 channel=41
					8, -7, 8, -6, -3, 0, -7, 11, -8,
					-- layer=2 filter=17 channel=42
					14, -1, 0, -2, -17, -2, 0, 1, 2,
					-- layer=2 filter=17 channel=43
					10, -8, -4, -7, -15, 4, -22, -13, 4,
					-- layer=2 filter=17 channel=44
					-10, 0, 0, 2, 0, -1, 1, -5, -2,
					-- layer=2 filter=17 channel=45
					-10, -23, 0, -8, 6, 9, -11, -4, -7,
					-- layer=2 filter=17 channel=46
					-13, -3, -10, -12, -2, -11, -12, -22, -22,
					-- layer=2 filter=17 channel=47
					-3, -26, -20, 8, -4, -1, -7, 6, 0,
					-- layer=2 filter=17 channel=48
					8, 3, 8, 4, 7, -5, 0, 4, 8,
					-- layer=2 filter=17 channel=49
					-20, -13, -12, -20, 3, -16, -25, -8, -4,
					-- layer=2 filter=17 channel=50
					0, 7, 4, 10, 0, -3, -8, -11, 12,
					-- layer=2 filter=17 channel=51
					-27, -26, -15, -15, -25, -6, -25, -7, -15,
					-- layer=2 filter=17 channel=52
					7, 2, -25, -21, -16, 0, 11, -4, -20,
					-- layer=2 filter=17 channel=53
					4, 5, -14, -19, -7, 4, -14, -16, -10,
					-- layer=2 filter=17 channel=54
					-7, -2, 0, 7, -12, -16, -23, -6, -19,
					-- layer=2 filter=17 channel=55
					2, 3, 6, -10, 1, -5, -4, -9, -5,
					-- layer=2 filter=17 channel=56
					-12, -19, -11, -15, -10, -11, -10, -17, -13,
					-- layer=2 filter=17 channel=57
					8, -5, 0, 7, 0, -2, 10, -2, -1,
					-- layer=2 filter=17 channel=58
					10, -2, -3, 3, -20, 0, -7, 1, -14,
					-- layer=2 filter=17 channel=59
					-8, -21, 0, -5, -13, 9, 4, -11, -10,
					-- layer=2 filter=17 channel=60
					-9, -18, -5, -8, -4, 0, -11, 5, -16,
					-- layer=2 filter=17 channel=61
					-1, -7, 3, -7, 3, -6, -4, 5, -14,
					-- layer=2 filter=17 channel=62
					-18, -6, -6, -10, -10, -7, -11, -7, -29,
					-- layer=2 filter=17 channel=63
					-12, -27, -18, -8, -6, 17, -4, -8, 0,
					-- layer=2 filter=17 channel=64
					-1, -18, -18, -4, -16, -19, 2, -5, -3,
					-- layer=2 filter=17 channel=65
					-5, -11, -10, -10, -6, -7, -4, -14, -7,
					-- layer=2 filter=17 channel=66
					-6, -10, -11, 1, 6, -6, 6, -5, 9,
					-- layer=2 filter=17 channel=67
					-9, -13, 0, -6, -7, -1, -15, -9, -22,
					-- layer=2 filter=17 channel=68
					-1, 2, -9, -2, 8, -11, 3, -2, -3,
					-- layer=2 filter=17 channel=69
					-6, -11, 9, 4, -2, -6, -7, -3, 7,
					-- layer=2 filter=17 channel=70
					22, 16, 5, 7, -2, -4, -7, -12, -10,
					-- layer=2 filter=17 channel=71
					-11, -5, -6, -16, -1, 0, -4, 0, -12,
					-- layer=2 filter=17 channel=72
					-19, -8, -3, -8, 7, -7, 1, 6, 18,
					-- layer=2 filter=17 channel=73
					-5, -7, -12, -11, -9, -13, -11, -6, -6,
					-- layer=2 filter=17 channel=74
					-1, -5, -1, 3, 7, 10, -2, -2, -20,
					-- layer=2 filter=17 channel=75
					-13, -14, -1, -8, 2, 0, 3, 7, 10,
					-- layer=2 filter=17 channel=76
					3, -6, -12, 3, -24, -9, -3, -23, -12,
					-- layer=2 filter=17 channel=77
					1, -5, 5, 9, -9, -8, 2, 2, -5,
					-- layer=2 filter=17 channel=78
					-20, -16, -38, -19, -18, -14, -23, -10, -7,
					-- layer=2 filter=17 channel=79
					2, 3, 0, 9, -6, 7, -8, 2, 5,
					-- layer=2 filter=17 channel=80
					-14, 0, -24, -9, -10, -5, -6, -9, -18,
					-- layer=2 filter=17 channel=81
					5, -8, -8, -6, 8, 4, -1, -9, 6,
					-- layer=2 filter=17 channel=82
					7, -1, 9, -7, 5, 8, -2, 9, 6,
					-- layer=2 filter=17 channel=83
					-3, -3, 0, -2, -11, -17, -2, -7, -8,
					-- layer=2 filter=17 channel=84
					-5, -10, -3, -10, -4, -11, 8, -8, -8,
					-- layer=2 filter=17 channel=85
					-3, 2, 2, 4, 8, 0, 0, 2, -9,
					-- layer=2 filter=17 channel=86
					5, 8, -3, -4, 4, -7, 1, 9, -6,
					-- layer=2 filter=17 channel=87
					-8, -26, -27, -10, 0, -1, -16, -15, -2,
					-- layer=2 filter=17 channel=88
					-14, -8, 3, 4, 19, 7, -4, -8, -28,
					-- layer=2 filter=17 channel=89
					-4, -14, -7, 4, 1, 8, 3, -2, 8,
					-- layer=2 filter=17 channel=90
					5, -8, 5, 10, -3, 4, -8, 9, -1,
					-- layer=2 filter=17 channel=91
					6, -13, 4, -8, -26, -6, -8, 4, 29,
					-- layer=2 filter=17 channel=92
					-13, -5, 11, 4, -5, -14, 0, 9, 2,
					-- layer=2 filter=17 channel=93
					-13, -6, -1, -9, -1, 3, 8, 0, -7,
					-- layer=2 filter=17 channel=94
					-11, 2, -9, 1, -8, 6, -5, -21, 17,
					-- layer=2 filter=17 channel=95
					2, -7, 3, -7, -6, -4, -3, 6, -8,
					-- layer=2 filter=17 channel=96
					12, -6, -15, -8, -3, -3, -1, -5, 5,
					-- layer=2 filter=17 channel=97
					-20, -34, -14, 23, -19, -6, -14, 12, 18,
					-- layer=2 filter=17 channel=98
					2, -20, -10, -10, -14, -5, -7, -9, 1,
					-- layer=2 filter=17 channel=99
					6, -5, -15, -17, -3, -6, 14, -2, -2,
					-- layer=2 filter=17 channel=100
					-11, -14, 15, -10, -13, -13, -21, -14, -21,
					-- layer=2 filter=17 channel=101
					-1, -16, -7, -8, -14, 0, 22, 8, -14,
					-- layer=2 filter=17 channel=102
					1, -3, -7, -18, 2, -1, 0, 2, 8,
					-- layer=2 filter=17 channel=103
					7, -4, 3, -6, -2, -17, 21, 7, -11,
					-- layer=2 filter=17 channel=104
					8, 0, -15, -21, -4, -14, -19, 1, 14,
					-- layer=2 filter=17 channel=105
					3, -22, -12, -12, 8, -7, -19, -28, -16,
					-- layer=2 filter=17 channel=106
					-12, -22, -13, -11, -5, -11, 7, -11, 4,
					-- layer=2 filter=17 channel=107
					-3, -13, 2, -1, -22, 8, 15, -5, 1,
					-- layer=2 filter=17 channel=108
					-25, -15, -1, -23, 9, 2, -10, 8, 4,
					-- layer=2 filter=17 channel=109
					-8, 2, 0, 5, -1, -10, -11, 5, -9,
					-- layer=2 filter=17 channel=110
					-7, -12, -8, -4, -9, -13, -14, 18, -1,
					-- layer=2 filter=17 channel=111
					0, 1, -7, 3, 8, -5, 11, 2, -4,
					-- layer=2 filter=17 channel=112
					-1, -17, -10, -8, -15, 1, -11, -4, -7,
					-- layer=2 filter=17 channel=113
					2, 8, 7, -10, -17, -17, -14, -1, -2,
					-- layer=2 filter=17 channel=114
					0, -6, 3, 1, 4, -2, 7, -11, 8,
					-- layer=2 filter=17 channel=115
					5, -8, 0, 4, -6, 6, -2, -5, 5,
					-- layer=2 filter=17 channel=116
					3, -18, -18, -18, -9, -4, -13, -8, -2,
					-- layer=2 filter=17 channel=117
					11, -17, -17, 7, 0, -6, -4, -8, -20,
					-- layer=2 filter=17 channel=118
					-14, -24, -18, -30, -18, -26, -30, -35, -32,
					-- layer=2 filter=17 channel=119
					0, 0, -20, -20, -1, -23, -23, -19, -7,
					-- layer=2 filter=17 channel=120
					-7, 1, 8, 4, 6, -8, 1, -3, -6,
					-- layer=2 filter=17 channel=121
					10, -7, 1, -8, 1, 0, 0, -8, -9,
					-- layer=2 filter=17 channel=122
					8, 1, -10, 2, 0, 4, -8, 4, -9,
					-- layer=2 filter=17 channel=123
					-12, -13, -12, -5, -7, -11, -7, -27, -16,
					-- layer=2 filter=17 channel=124
					-10, -4, -20, -4, -13, -13, -1, 1, -8,
					-- layer=2 filter=17 channel=125
					9, 1, 3, 7, 11, 8, 8, -1, -4,
					-- layer=2 filter=17 channel=126
					1, -3, -5, 7, 1, 19, -10, -18, 14,
					-- layer=2 filter=17 channel=127
					-24, 2, 1, -6, -12, 3, 0, 7, -1,
					-- layer=2 filter=18 channel=0
					-34, -11, 2, -14, 0, 18, -5, 25, 31,
					-- layer=2 filter=18 channel=1
					-12, -4, 1, -22, -39, -24, -7, -33, -21,
					-- layer=2 filter=18 channel=2
					6, 7, 4, -2, 5, 2, 7, -1, 1,
					-- layer=2 filter=18 channel=3
					7, -6, -8, -3, 10, -3, -29, 1, 16,
					-- layer=2 filter=18 channel=4
					-19, 12, 22, -25, 22, 11, -29, 44, -10,
					-- layer=2 filter=18 channel=5
					-25, 18, 7, -7, 13, 22, -12, 8, 12,
					-- layer=2 filter=18 channel=6
					23, -39, 3, -7, -70, -20, 4, 0, -1,
					-- layer=2 filter=18 channel=7
					10, 21, 3, 13, 19, 5, 29, 21, 6,
					-- layer=2 filter=18 channel=8
					-2, 7, 5, -1, 0, 0, 6, 10, -9,
					-- layer=2 filter=18 channel=9
					-29, -13, -5, -9, 10, 13, -33, -10, 7,
					-- layer=2 filter=18 channel=10
					-17, -3, -5, -4, 18, 15, -18, 17, 9,
					-- layer=2 filter=18 channel=11
					-2, 4, 8, -4, 7, 21, -14, 7, 13,
					-- layer=2 filter=18 channel=12
					-17, 4, 23, -19, -21, -9, 29, -9, -29,
					-- layer=2 filter=18 channel=13
					11, 0, 3, 5, -1, 3, -4, 7, 5,
					-- layer=2 filter=18 channel=14
					10, 10, 35, -3, 0, 17, 16, -3, 11,
					-- layer=2 filter=18 channel=15
					16, 0, -16, -16, -16, -24, 23, -4, -47,
					-- layer=2 filter=18 channel=16
					-36, -23, 5, 11, 20, 21, 6, 11, -8,
					-- layer=2 filter=18 channel=17
					1, -2, 8, 1, 5, -7, 7, -4, -7,
					-- layer=2 filter=18 channel=18
					77, 42, 22, 36, 32, 9, 46, 37, -5,
					-- layer=2 filter=18 channel=19
					5, -4, -7, -33, -29, -13, -12, -32, -37,
					-- layer=2 filter=18 channel=20
					1, 6, 9, 1, -4, -8, 4, -6, 7,
					-- layer=2 filter=18 channel=21
					4, 0, -5, -1, 3, 1, -3, 1, 2,
					-- layer=2 filter=18 channel=22
					-6, -12, 6, 8, -7, 7, -5, 4, 5,
					-- layer=2 filter=18 channel=23
					-34, -1, -18, 1, 9, 0, -26, 15, -29,
					-- layer=2 filter=18 channel=24
					-16, -33, -20, -12, -23, 12, -34, -26, 0,
					-- layer=2 filter=18 channel=25
					-17, -45, -7, -30, -44, -4, -29, -30, 12,
					-- layer=2 filter=18 channel=26
					6, -4, -3, 9, 0, 9, -3, 2, -6,
					-- layer=2 filter=18 channel=27
					19, 6, 13, 0, -13, 13, 5, -3, 6,
					-- layer=2 filter=18 channel=28
					21, 8, -9, 0, -14, -9, 20, 12, 38,
					-- layer=2 filter=18 channel=29
					-5, -7, -9, 6, -1, 5, -7, -1, 0,
					-- layer=2 filter=18 channel=30
					-13, 3, 29, -11, 6, 9, -1, 10, 34,
					-- layer=2 filter=18 channel=31
					-13, -3, -72, 17, 25, 37, 29, 1, -16,
					-- layer=2 filter=18 channel=32
					-6, 0, 4, 0, 7, -6, 2, -3, -8,
					-- layer=2 filter=18 channel=33
					36, 21, -10, 15, 1, 21, 48, 18, 5,
					-- layer=2 filter=18 channel=34
					31, 13, 3, -8, 21, -2, 40, 2, 13,
					-- layer=2 filter=18 channel=35
					16, 40, 17, 27, -9, -7, 34, 29, 36,
					-- layer=2 filter=18 channel=36
					1, 17, 8, 8, 10, 4, 7, 20, -12,
					-- layer=2 filter=18 channel=37
					4, 10, 2, -9, 9, 12, -16, 5, -2,
					-- layer=2 filter=18 channel=38
					-28, 6, 18, -24, 0, 28, -41, -14, 10,
					-- layer=2 filter=18 channel=39
					-7, -34, -24, 12, -7, 10, 36, 2, 6,
					-- layer=2 filter=18 channel=40
					-19, 5, -13, -3, 2, 27, -25, 38, -14,
					-- layer=2 filter=18 channel=41
					8, 9, 2, 10, 9, -1, 9, 10, 7,
					-- layer=2 filter=18 channel=42
					-16, 3, 10, -2, 2, -8, 15, -17, -49,
					-- layer=2 filter=18 channel=43
					16, 31, -18, -14, 2, -9, -30, 12, 21,
					-- layer=2 filter=18 channel=44
					-2, -7, 0, 6, 8, -6, 1, 0, 5,
					-- layer=2 filter=18 channel=45
					12, -1, 6, -25, 25, 33, 37, -3, 0,
					-- layer=2 filter=18 channel=46
					-37, -18, -4, -8, 0, 15, -2, 3, 13,
					-- layer=2 filter=18 channel=47
					-9, -4, -19, 13, -1, -21, 22, 4, 11,
					-- layer=2 filter=18 channel=48
					-7, -1, -2, 7, -2, 8, -1, 7, 8,
					-- layer=2 filter=18 channel=49
					50, 13, 12, 29, 21, 5, 30, -20, -21,
					-- layer=2 filter=18 channel=50
					-2, -2, 8, 27, 6, 6, 13, -7, -12,
					-- layer=2 filter=18 channel=51
					-23, -3, 17, -8, 17, 11, -28, 5, 12,
					-- layer=2 filter=18 channel=52
					28, 13, -6, 9, 7, -6, -40, -17, 15,
					-- layer=2 filter=18 channel=53
					32, 6, 55, 38, -33, -6, 7, -32, 8,
					-- layer=2 filter=18 channel=54
					12, -4, -20, 16, -6, -7, 23, 25, -14,
					-- layer=2 filter=18 channel=55
					11, -4, -5, 6, -10, -8, 1, 3, 12,
					-- layer=2 filter=18 channel=56
					-20, 7, -4, -14, -10, 9, -1, 4, 3,
					-- layer=2 filter=18 channel=57
					0, -2, 4, -11, 14, 2, -21, 5, 15,
					-- layer=2 filter=18 channel=58
					-47, -1, 29, -16, -45, -42, 47, -10, -20,
					-- layer=2 filter=18 channel=59
					1, -4, 5, 11, -44, -1, -11, -36, 2,
					-- layer=2 filter=18 channel=60
					-18, -65, -23, 24, -48, -19, -33, -86, -4,
					-- layer=2 filter=18 channel=61
					21, -18, 22, 40, 7, 7, -6, -17, 23,
					-- layer=2 filter=18 channel=62
					32, -34, -25, -12, -8, -2, 12, -6, -24,
					-- layer=2 filter=18 channel=63
					-4, -49, -9, 10, -21, 19, 0, -27, 3,
					-- layer=2 filter=18 channel=64
					-4, 0, 3, -5, 10, 16, 36, 17, 14,
					-- layer=2 filter=18 channel=65
					12, -21, 37, 19, -32, -5, 7, -9, 39,
					-- layer=2 filter=18 channel=66
					-21, -8, 3, -45, -15, -3, -16, -48, 2,
					-- layer=2 filter=18 channel=67
					-23, -7, -13, -17, 12, 17, -46, 6, 25,
					-- layer=2 filter=18 channel=68
					-3, -1, -3, -3, 1, -8, -8, -3, -5,
					-- layer=2 filter=18 channel=69
					-10, -11, -3, 2, -4, 10, 30, 17, 7,
					-- layer=2 filter=18 channel=70
					10, 0, 9, 4, 0, -25, 15, 13, 23,
					-- layer=2 filter=18 channel=71
					13, -19, 23, 5, -37, 12, -28, -38, 9,
					-- layer=2 filter=18 channel=72
					-15, 28, 8, -14, -2, 1, 12, -17, -18,
					-- layer=2 filter=18 channel=73
					9, -4, -14, 0, 48, 29, 35, -2, 18,
					-- layer=2 filter=18 channel=74
					-36, -6, -9, -17, -5, 8, -20, 11, 15,
					-- layer=2 filter=18 channel=75
					-50, -4, 3, 50, -69, -46, -5, 26, 12,
					-- layer=2 filter=18 channel=76
					33, -17, 11, 4, -5, -9, -9, 5, -4,
					-- layer=2 filter=18 channel=77
					3, 4, 2, 5, 6, 5, 7, 0, 0,
					-- layer=2 filter=18 channel=78
					9, 18, -13, 2, -5, 10, -17, 2, 33,
					-- layer=2 filter=18 channel=79
					7, 9, 5, -7, -10, -3, -6, 1, 7,
					-- layer=2 filter=18 channel=80
					-25, 18, 10, -8, 14, 5, -13, 9, -4,
					-- layer=2 filter=18 channel=81
					5, 5, -1, 11, -4, -1, -10, 10, 0,
					-- layer=2 filter=18 channel=82
					5, -10, 6, 5, 1, 10, -3, -3, 1,
					-- layer=2 filter=18 channel=83
					-30, -3, 15, -21, 13, -18, -19, 11, -20,
					-- layer=2 filter=18 channel=84
					3, 9, 2, 3, 1, 10, -10, 5, -7,
					-- layer=2 filter=18 channel=85
					9, 0, -8, 9, -4, -11, -2, 4, 4,
					-- layer=2 filter=18 channel=86
					2, -2, 11, 11, 16, -1, 10, 0, 0,
					-- layer=2 filter=18 channel=87
					49, 43, -21, 17, -34, -44, -17, 36, -12,
					-- layer=2 filter=18 channel=88
					-29, -9, 0, 4, -20, 33, 24, 6, 17,
					-- layer=2 filter=18 channel=89
					3, -3, 22, -20, -41, -27, 20, -16, -16,
					-- layer=2 filter=18 channel=90
					12, 9, 11, -1, 8, 3, -7, 7, -3,
					-- layer=2 filter=18 channel=91
					0, 11, 8, -44, -50, -77, -1, -37, -33,
					-- layer=2 filter=18 channel=92
					-8, -4, 6, -40, -19, -2, 23, -14, -9,
					-- layer=2 filter=18 channel=93
					51, 7, -31, 15, -82, -47, -31, -23, -36,
					-- layer=2 filter=18 channel=94
					5, -61, 2, 9, -34, 41, -21, -16, 17,
					-- layer=2 filter=18 channel=95
					-23, -31, -11, -42, -18, -12, -5, 1, -21,
					-- layer=2 filter=18 channel=96
					13, -22, 13, -2, -53, -4, 20, -11, -42,
					-- layer=2 filter=18 channel=97
					-14, -13, 0, 6, 24, 32, -10, 5, 18,
					-- layer=2 filter=18 channel=98
					6, 26, -32, 17, -8, -25, 24, 14, 4,
					-- layer=2 filter=18 channel=99
					15, -45, 0, 8, -41, 17, -20, -39, 27,
					-- layer=2 filter=18 channel=100
					-24, 0, 2, 20, -10, 5, -14, -30, -4,
					-- layer=2 filter=18 channel=101
					3, -10, 19, 3, -11, 14, 15, 24, 3,
					-- layer=2 filter=18 channel=102
					34, 18, 47, 31, 1, -10, 8, 17, -9,
					-- layer=2 filter=18 channel=103
					-2, -15, -2, -13, 26, 17, 18, 35, -2,
					-- layer=2 filter=18 channel=104
					72, 15, 2, 58, -5, 16, 39, 29, -29,
					-- layer=2 filter=18 channel=105
					0, -35, 27, -30, -33, -22, -36, 0, 9,
					-- layer=2 filter=18 channel=106
					-9, -20, 7, -4, -3, -16, -19, -1, 21,
					-- layer=2 filter=18 channel=107
					-24, 22, 18, 7, 62, 41, 9, 14, 8,
					-- layer=2 filter=18 channel=108
					0, -5, 2, -14, -28, -24, -34, -39, -12,
					-- layer=2 filter=18 channel=109
					-19, 15, 1, -21, 6, 0, 1, -15, -8,
					-- layer=2 filter=18 channel=110
					1, -26, 3, -9, -25, -21, 46, -6, -5,
					-- layer=2 filter=18 channel=111
					-5, 10, 6, -8, 11, -10, 0, 10, 6,
					-- layer=2 filter=18 channel=112
					-41, -6, -2, -32, 10, 15, -56, -17, 15,
					-- layer=2 filter=18 channel=113
					-26, -4, 35, 16, 9, 11, 14, -11, 36,
					-- layer=2 filter=18 channel=114
					-7, 13, 0, 3, 10, -8, 13, -4, -5,
					-- layer=2 filter=18 channel=115
					-5, 0, -6, 4, -5, 3, -4, -9, 0,
					-- layer=2 filter=18 channel=116
					49, 33, 0, -3, -47, -60, 11, 12, -32,
					-- layer=2 filter=18 channel=117
					-2, 3, 3, -5, 9, 18, 18, 21, -25,
					-- layer=2 filter=18 channel=118
					-3, 33, -6, 16, 12, 4, -23, 21, -9,
					-- layer=2 filter=18 channel=119
					-12, 8, 8, 19, 18, 18, 8, 27, 7,
					-- layer=2 filter=18 channel=120
					-1, -9, 9, -7, -4, 1, -5, -10, 0,
					-- layer=2 filter=18 channel=121
					-1, 1, 5, -5, -6, 7, 8, -3, 8,
					-- layer=2 filter=18 channel=122
					-1, 3, 0, 8, -6, 10, -2, 3, 4,
					-- layer=2 filter=18 channel=123
					-5, 7, -28, -7, -14, -18, 1, 10, -16,
					-- layer=2 filter=18 channel=124
					20, 4, -11, -3, -14, 6, -2, 15, -19,
					-- layer=2 filter=18 channel=125
					8, 2, 10, 2, -9, 2, -1, -10, 0,
					-- layer=2 filter=18 channel=126
					-13, -57, 15, 45, -50, 10, 24, -73, 0,
					-- layer=2 filter=18 channel=127
					-21, -43, 36, -3, -11, 16, -10, -37, 36,
					-- layer=2 filter=19 channel=0
					-26, -22, 0, -46, -20, 15, -37, -50, -6,
					-- layer=2 filter=19 channel=1
					-21, 32, 12, 0, -13, -38, -22, 15, 7,
					-- layer=2 filter=19 channel=2
					-4, -5, -7, 3, 5, -7, -7, 9, -8,
					-- layer=2 filter=19 channel=3
					-32, -25, 18, -40, -50, -42, -7, -25, 0,
					-- layer=2 filter=19 channel=4
					28, 13, 14, 13, 25, 1, 14, -13, -24,
					-- layer=2 filter=19 channel=5
					-28, -20, 31, -55, 7, 3, -13, 23, 2,
					-- layer=2 filter=19 channel=6
					2, 4, 5, 0, 18, 10, 4, 7, -21,
					-- layer=2 filter=19 channel=7
					-33, -35, 0, 51, 0, -19, -20, -75, 4,
					-- layer=2 filter=19 channel=8
					6, 6, 1, -2, 12, 5, -10, -3, -4,
					-- layer=2 filter=19 channel=9
					31, 17, 2, -42, -5, 19, -18, -26, -1,
					-- layer=2 filter=19 channel=10
					-31, -7, 3, -37, -26, 0, -6, -27, -23,
					-- layer=2 filter=19 channel=11
					-6, 17, 16, 24, 28, 11, 36, 7, 29,
					-- layer=2 filter=19 channel=12
					17, 13, -5, 7, -63, -16, 3, 13, 26,
					-- layer=2 filter=19 channel=13
					-5, -9, 6, -3, -7, 6, -1, 5, 8,
					-- layer=2 filter=19 channel=14
					30, 14, 4, 10, -4, 5, -5, 28, 44,
					-- layer=2 filter=19 channel=15
					-18, 22, -21, 35, 43, 5, 32, -8, -44,
					-- layer=2 filter=19 channel=16
					-17, 3, 3, 24, 22, 13, 18, 2, -23,
					-- layer=2 filter=19 channel=17
					-3, 6, -9, 2, 7, 6, 8, 1, 5,
					-- layer=2 filter=19 channel=18
					51, 12, 27, 6, 29, -37, 19, 14, -37,
					-- layer=2 filter=19 channel=19
					-81, -29, -47, -50, -4, -14, -39, 24, -44,
					-- layer=2 filter=19 channel=20
					-9, -5, 1, 6, 7, 6, -5, 5, -6,
					-- layer=2 filter=19 channel=21
					8, 9, 12, 8, 7, 4, -1, 19, 21,
					-- layer=2 filter=19 channel=22
					0, -6, 3, -5, -10, 7, 1, -8, -8,
					-- layer=2 filter=19 channel=23
					18, 20, -3, 20, 12, 6, 10, 1, -11,
					-- layer=2 filter=19 channel=24
					-24, -28, 14, -26, -59, -3, 6, -33, 13,
					-- layer=2 filter=19 channel=25
					12, -20, -13, 24, -19, 23, 40, 17, 52,
					-- layer=2 filter=19 channel=26
					0, 5, -6, 6, 3, -4, -4, 0, -5,
					-- layer=2 filter=19 channel=27
					-54, -48, 2, -70, -17, 25, -27, 12, 17,
					-- layer=2 filter=19 channel=28
					0, -8, -32, -9, -6, 6, 43, -63, -6,
					-- layer=2 filter=19 channel=29
					-1, -6, 8, -5, 6, -7, 8, 5, 6,
					-- layer=2 filter=19 channel=30
					-3, 26, 2, 9, 14, 7, -6, 35, -23,
					-- layer=2 filter=19 channel=31
					-65, -45, -64, -50, -20, 0, -9, 3, -4,
					-- layer=2 filter=19 channel=32
					5, -7, 7, 2, 0, -3, 8, -11, 0,
					-- layer=2 filter=19 channel=33
					-30, 22, 30, 45, 40, -39, -14, -23, -18,
					-- layer=2 filter=19 channel=34
					18, 16, 3, 18, 38, 12, 30, 18, -44,
					-- layer=2 filter=19 channel=35
					5, -8, -22, 17, 4, -6, 23, -64, -23,
					-- layer=2 filter=19 channel=36
					-4, -12, -6, 14, 5, 1, 12, -1, 1,
					-- layer=2 filter=19 channel=37
					-17, 15, -1, -26, 42, 18, 19, 34, 10,
					-- layer=2 filter=19 channel=38
					-52, 0, 13, -90, -31, 12, -31, 38, -3,
					-- layer=2 filter=19 channel=39
					-9, 28, 30, 30, -6, -3, 26, 6, 24,
					-- layer=2 filter=19 channel=40
					9, -59, 2, -9, 36, 37, 62, 31, 39,
					-- layer=2 filter=19 channel=41
					-5, -8, -7, 2, 0, -9, 0, -2, 0,
					-- layer=2 filter=19 channel=42
					18, 30, 0, 28, 10, -30, 15, 15, 3,
					-- layer=2 filter=19 channel=43
					-35, -12, 22, -40, -30, -40, 7, -61, -36,
					-- layer=2 filter=19 channel=44
					5, 3, 0, 6, -2, 1, -3, -7, -5,
					-- layer=2 filter=19 channel=45
					-129, -78, -41, -14, -38, -36, -33, 2, -23,
					-- layer=2 filter=19 channel=46
					-19, 2, 2, 10, -4, 7, 11, -37, 1,
					-- layer=2 filter=19 channel=47
					-18, -20, -11, 8, 25, 12, 5, -41, 1,
					-- layer=2 filter=19 channel=48
					9, 7, 4, 3, 5, 9, 1, 2, 6,
					-- layer=2 filter=19 channel=49
					46, 8, -4, 14, 8, -62, 36, 23, -4,
					-- layer=2 filter=19 channel=50
					21, 2, -18, -1, -8, -3, -4, -12, -9,
					-- layer=2 filter=19 channel=51
					-2, 16, -4, -9, 14, 14, 7, 11, 21,
					-- layer=2 filter=19 channel=52
					-31, 66, 14, 0, 20, -16, -4, 17, 30,
					-- layer=2 filter=19 channel=53
					11, 1, -50, 5, 6, -27, -2, 2, -56,
					-- layer=2 filter=19 channel=54
					22, 23, -9, -4, 5, 6, 2, -17, -11,
					-- layer=2 filter=19 channel=55
					-5, 8, 10, -5, -3, 11, 6, 12, 7,
					-- layer=2 filter=19 channel=56
					8, 4, 3, 4, 22, 20, 44, 22, 6,
					-- layer=2 filter=19 channel=57
					-6, 2, -13, 2, 2, 0, 11, 5, 13,
					-- layer=2 filter=19 channel=58
					-27, 4, -13, 13, -57, -1, 12, 20, 39,
					-- layer=2 filter=19 channel=59
					-76, -7, 8, -3, -19, -17, -38, 5, 21,
					-- layer=2 filter=19 channel=60
					-12, 22, 18, -67, 8, 50, -16, 16, 14,
					-- layer=2 filter=19 channel=61
					-14, -26, -10, -80, 3, 20, -86, 21, 22,
					-- layer=2 filter=19 channel=62
					13, 23, 22, 10, 7, -5, 15, 31, -24,
					-- layer=2 filter=19 channel=63
					-5, -3, -7, -11, 6, 2, -11, -30, -6,
					-- layer=2 filter=19 channel=64
					-13, -10, 3, -3, -7, 4, -22, -9, -27,
					-- layer=2 filter=19 channel=65
					-28, 3, -26, -36, 5, -10, -57, 30, 0,
					-- layer=2 filter=19 channel=66
					48, 56, 46, -52, -7, -38, -48, -22, 31,
					-- layer=2 filter=19 channel=67
					-22, 28, 26, -54, -22, 15, -44, -50, -21,
					-- layer=2 filter=19 channel=68
					-8, 8, -6, 11, 7, 11, -8, 4, -7,
					-- layer=2 filter=19 channel=69
					0, 17, 8, 12, 25, -17, 5, 12, -3,
					-- layer=2 filter=19 channel=70
					-22, -28, -39, -6, 15, 2, 17, -40, -12,
					-- layer=2 filter=19 channel=71
					-32, -34, -7, 0, 31, -2, 0, 47, 37,
					-- layer=2 filter=19 channel=72
					53, -7, 11, 0, 7, -23, 8, -1, 13,
					-- layer=2 filter=19 channel=73
					-37, -62, 0, 5, -51, 28, 8, 16, 20,
					-- layer=2 filter=19 channel=74
					-12, 36, 9, -17, -4, 29, 13, 25, -7,
					-- layer=2 filter=19 channel=75
					-56, -20, -76, -25, -21, 9, 26, 21, -53,
					-- layer=2 filter=19 channel=76
					19, 24, -80, -7, -12, -53, -3, 0, -91,
					-- layer=2 filter=19 channel=77
					-8, -2, -2, 0, 0, -4, 0, 9, -12,
					-- layer=2 filter=19 channel=78
					10, 11, 13, 12, 7, 0, 1, 7, -13,
					-- layer=2 filter=19 channel=79
					12, 4, 0, -8, -6, 2, 0, 1, -4,
					-- layer=2 filter=19 channel=80
					0, 18, 21, 45, 33, 37, 32, 4, 30,
					-- layer=2 filter=19 channel=81
					-4, 8, -8, 16, -4, -2, 1, 8, 11,
					-- layer=2 filter=19 channel=82
					6, 13, -6, -8, 13, 1, 11, 3, 8,
					-- layer=2 filter=19 channel=83
					15, -1, -1, 22, 25, 9, -10, 27, 7,
					-- layer=2 filter=19 channel=84
					-4, 10, -8, -1, -1, -4, -6, -1, -7,
					-- layer=2 filter=19 channel=85
					-1, -22, 5, -8, -3, 0, 0, 1, 13,
					-- layer=2 filter=19 channel=86
					4, -4, -10, 8, -17, 8, -8, -11, 1,
					-- layer=2 filter=19 channel=87
					24, 48, 28, 36, 36, -35, 6, 0, -55,
					-- layer=2 filter=19 channel=88
					3, 39, 8, -15, 3, 22, -13, 17, -5,
					-- layer=2 filter=19 channel=89
					32, 10, -20, 14, -16, -15, 24, 29, 54,
					-- layer=2 filter=19 channel=90
					8, 2, 7, -7, -4, -9, -4, 4, 1,
					-- layer=2 filter=19 channel=91
					-19, -4, -13, -18, -82, -9, 29, 31, 38,
					-- layer=2 filter=19 channel=92
					26, 0, 1, -5, -53, -16, -3, 36, 41,
					-- layer=2 filter=19 channel=93
					-16, 30, 22, 4, 48, 36, 17, 58, -5,
					-- layer=2 filter=19 channel=94
					22, 4, 1, -58, 33, 38, -61, -6, -8,
					-- layer=2 filter=19 channel=95
					-5, -9, -3, 5, 0, -3, 1, -17, -5,
					-- layer=2 filter=19 channel=96
					-43, -34, -34, -44, -4, 0, -45, 33, 37,
					-- layer=2 filter=19 channel=97
					-9, -27, 10, 0, -13, -22, -20, -4, -6,
					-- layer=2 filter=19 channel=98
					0, -48, -42, -8, 13, 25, -12, -77, -23,
					-- layer=2 filter=19 channel=99
					-61, 33, -48, -34, 20, 26, -15, 26, 36,
					-- layer=2 filter=19 channel=100
					5, 34, 43, -18, -18, 21, 22, 42, 27,
					-- layer=2 filter=19 channel=101
					-10, -40, -37, 24, -11, -8, 57, 15, 46,
					-- layer=2 filter=19 channel=102
					-9, 22, -55, 21, 58, -38, -7, 11, -21,
					-- layer=2 filter=19 channel=103
					-25, -23, 3, 42, -67, -29, 20, 28, 14,
					-- layer=2 filter=19 channel=104
					48, 21, 3, 21, 13, -27, 16, 19, -29,
					-- layer=2 filter=19 channel=105
					39, 30, -54, -35, 4, -42, -44, -31, -23,
					-- layer=2 filter=19 channel=106
					-39, 0, -23, -12, -35, -13, 36, 26, 22,
					-- layer=2 filter=19 channel=107
					12, 17, -23, 14, -26, -45, 0, 19, 38,
					-- layer=2 filter=19 channel=108
					-55, 4, -6, -33, 15, 1, -34, 0, -3,
					-- layer=2 filter=19 channel=109
					13, 6, 15, 10, 3, -1, 11, 15, 7,
					-- layer=2 filter=19 channel=110
					-1, -17, 1, -19, -3, 8, 4, 12, 35,
					-- layer=2 filter=19 channel=111
					-8, 0, -7, 2, 7, 2, 0, -11, -1,
					-- layer=2 filter=19 channel=112
					-18, -15, -38, -33, -35, 23, -25, -10, 1,
					-- layer=2 filter=19 channel=113
					12, 0, -28, 22, 0, -3, -23, -11, 14,
					-- layer=2 filter=19 channel=114
					-14, -23, -27, -20, -11, 1, -30, -8, -3,
					-- layer=2 filter=19 channel=115
					-8, 3, -10, -7, -11, 7, -2, -5, 3,
					-- layer=2 filter=19 channel=116
					-9, 23, 6, 29, 54, -3, 2, 18, -68,
					-- layer=2 filter=19 channel=117
					-7, -30, -20, 18, 18, 28, -17, -8, -35,
					-- layer=2 filter=19 channel=118
					-14, -1, 4, -7, -22, -35, -22, -31, -35,
					-- layer=2 filter=19 channel=119
					-4, 1, 14, 0, 7, -3, 1, -30, -35,
					-- layer=2 filter=19 channel=120
					1, 3, 9, 0, -1, 3, -5, 1, 7,
					-- layer=2 filter=19 channel=121
					-10, -2, 6, -9, -5, -7, -5, -10, -1,
					-- layer=2 filter=19 channel=122
					-6, -7, -9, 2, -2, 15, -5, 10, 4,
					-- layer=2 filter=19 channel=123
					-1, -10, 4, 18, 3, -4, -72, -36, -10,
					-- layer=2 filter=19 channel=124
					16, 53, -24, 32, -20, -88, 15, 0, -33,
					-- layer=2 filter=19 channel=125
					-3, 2, -1, 8, -2, 5, 4, 6, -5,
					-- layer=2 filter=19 channel=126
					20, -17, 53, -74, 0, 10, 5, -27, 8,
					-- layer=2 filter=19 channel=127
					-16, 49, -4, 19, 32, -20, -23, 18, 20,
					-- layer=2 filter=20 channel=0
					7, -14, 19, -1, -4, 24, -5, 5, -1,
					-- layer=2 filter=20 channel=1
					20, 31, -2, 36, 23, -17, -22, 34, -16,
					-- layer=2 filter=20 channel=2
					8, -8, -3, 1, -12, -3, -2, -2, 0,
					-- layer=2 filter=20 channel=3
					-9, -21, -11, 11, -5, -14, 58, 49, 23,
					-- layer=2 filter=20 channel=4
					-16, -25, 3, -6, 0, 21, -4, 1, -5,
					-- layer=2 filter=20 channel=5
					24, -3, -13, -7, -4, -2, 0, -4, -8,
					-- layer=2 filter=20 channel=6
					-10, 35, -30, -58, -99, -47, -86, -37, -120,
					-- layer=2 filter=20 channel=7
					37, 16, 52, 30, 48, 47, 4, 15, 1,
					-- layer=2 filter=20 channel=8
					-3, 7, -4, 0, -9, 5, 0, 0, -6,
					-- layer=2 filter=20 channel=9
					-12, -27, -43, 6, 0, -14, 56, 46, 0,
					-- layer=2 filter=20 channel=10
					-28, 2, 15, 14, 1, -1, 11, 45, 10,
					-- layer=2 filter=20 channel=11
					17, -19, -7, -2, -11, 6, -16, -1, 0,
					-- layer=2 filter=20 channel=12
					39, 31, 0, 25, 4, -6, 2, 29, -18,
					-- layer=2 filter=20 channel=13
					-4, 2, -5, -5, -5, 7, -3, -8, -5,
					-- layer=2 filter=20 channel=14
					26, 22, -7, 20, 23, 26, 5, 31, 14,
					-- layer=2 filter=20 channel=15
					5, -25, -17, -28, -12, -21, 0, -1, -25,
					-- layer=2 filter=20 channel=16
					-32, 8, 7, -49, 1, 8, -1, 29, 10,
					-- layer=2 filter=20 channel=17
					-5, 0, -2, 1, -5, -2, 0, 5, -1,
					-- layer=2 filter=20 channel=18
					-2, -11, -21, 0, 43, 19, -20, 38, 13,
					-- layer=2 filter=20 channel=19
					-24, 33, 13, -13, 6, -28, 5, 21, -18,
					-- layer=2 filter=20 channel=20
					10, -2, 8, -4, -8, -11, 9, -9, -7,
					-- layer=2 filter=20 channel=21
					10, -15, -11, -8, 4, -33, -19, -10, -2,
					-- layer=2 filter=20 channel=22
					-1, 13, -8, 11, -1, -3, -4, -10, 10,
					-- layer=2 filter=20 channel=23
					9, 26, -1, -15, 12, -9, -11, -7, -39,
					-- layer=2 filter=20 channel=24
					3, -31, -19, 27, 3, -5, 42, 38, 23,
					-- layer=2 filter=20 channel=25
					7, -41, -26, 5, -2, -5, 34, 37, 4,
					-- layer=2 filter=20 channel=26
					5, 9, 4, 0, 4, -9, 1, -6, 7,
					-- layer=2 filter=20 channel=27
					-20, -17, 14, 11, 17, -5, 9, 19, 36,
					-- layer=2 filter=20 channel=28
					5, 27, 14, 32, 17, 29, 27, 29, 32,
					-- layer=2 filter=20 channel=29
					-7, -1, 5, -7, -8, 2, 0, 3, 2,
					-- layer=2 filter=20 channel=30
					-24, -23, -4, -15, 22, -19, 17, -9, 44,
					-- layer=2 filter=20 channel=31
					-53, -59, -13, -34, 40, 44, 6, -10, -64,
					-- layer=2 filter=20 channel=32
					-9, 2, -4, 4, -4, 3, 3, -5, -10,
					-- layer=2 filter=20 channel=33
					1, 7, 22, 19, -6, 13, -18, 15, -3,
					-- layer=2 filter=20 channel=34
					17, -56, -22, -45, -15, -44, -22, -87, -1,
					-- layer=2 filter=20 channel=35
					27, 17, 12, -13, -5, -3, -4, 17, 26,
					-- layer=2 filter=20 channel=36
					12, 0, 5, 5, -15, 1, 8, -2, 18,
					-- layer=2 filter=20 channel=37
					8, 15, -3, -4, -16, -14, 19, 0, -9,
					-- layer=2 filter=20 channel=38
					20, 7, -9, 14, 19, -10, 0, 15, 11,
					-- layer=2 filter=20 channel=39
					-9, 11, 11, -14, 6, -13, -15, -9, -16,
					-- layer=2 filter=20 channel=40
					32, -18, -37, 17, -3, -62, 8, 42, 17,
					-- layer=2 filter=20 channel=41
					-3, 11, 0, -9, 8, 2, -2, -7, 10,
					-- layer=2 filter=20 channel=42
					5, 21, 0, -10, 7, 2, 11, -9, 0,
					-- layer=2 filter=20 channel=43
					-12, -62, -36, 0, -40, -24, 26, 15, 14,
					-- layer=2 filter=20 channel=44
					-9, -5, 5, -4, -2, 8, 0, 3, 3,
					-- layer=2 filter=20 channel=45
					-4, 29, 24, 22, 18, 2, 13, 32, 23,
					-- layer=2 filter=20 channel=46
					-26, -22, -12, -18, -5, -29, 21, 5, 4,
					-- layer=2 filter=20 channel=47
					6, 59, 55, 22, 5, 43, 13, 40, 41,
					-- layer=2 filter=20 channel=48
					-2, 5, -10, 5, -3, 2, 1, 5, 1,
					-- layer=2 filter=20 channel=49
					6, 48, -30, 12, 33, -9, -17, 69, 4,
					-- layer=2 filter=20 channel=50
					26, 14, 13, 4, 2, 16, 13, 5, 27,
					-- layer=2 filter=20 channel=51
					15, -4, -8, -10, -7, -8, -16, -2, 3,
					-- layer=2 filter=20 channel=52
					21, 7, 47, -15, -10, -24, -38, -22, 10,
					-- layer=2 filter=20 channel=53
					-10, -47, 14, -34, 15, -58, 37, -35, -51,
					-- layer=2 filter=20 channel=54
					0, 11, 42, -9, 0, 8, -42, -14, -11,
					-- layer=2 filter=20 channel=55
					11, 6, -7, 5, -2, 2, 8, -10, 0,
					-- layer=2 filter=20 channel=56
					41, -15, 3, 16, -14, -3, 0, 11, 2,
					-- layer=2 filter=20 channel=57
					-6, -13, 0, 0, -11, 0, 0, -3, -2,
					-- layer=2 filter=20 channel=58
					16, 46, 25, 15, -15, 19, -6, 18, -17,
					-- layer=2 filter=20 channel=59
					11, 25, 22, 42, -25, -12, -35, -12, -51,
					-- layer=2 filter=20 channel=60
					21, 0, -3, 4, 1, -33, -37, -17, -43,
					-- layer=2 filter=20 channel=61
					6, 32, -3, -12, -14, -20, -26, -42, -30,
					-- layer=2 filter=20 channel=62
					-7, 31, -7, -40, -18, -21, -37, -6, -11,
					-- layer=2 filter=20 channel=63
					24, 25, 9, 12, 7, 14, -32, -6, -12,
					-- layer=2 filter=20 channel=64
					-5, 30, 17, -25, 39, 5, 3, 28, 6,
					-- layer=2 filter=20 channel=65
					-10, 40, -24, -59, -45, -33, -86, -36, -85,
					-- layer=2 filter=20 channel=66
					-76, -19, 37, -23, -6, 17, 44, 27, 10,
					-- layer=2 filter=20 channel=67
					-36, -60, -41, -18, -23, -56, 17, 30, -1,
					-- layer=2 filter=20 channel=68
					-9, 0, -7, 4, -11, -8, -8, -2, 0,
					-- layer=2 filter=20 channel=69
					0, 43, -5, 5, 36, 14, -10, 2, 10,
					-- layer=2 filter=20 channel=70
					18, 18, 33, -5, 10, 21, -1, 1, 5,
					-- layer=2 filter=20 channel=71
					-16, -25, -18, 9, 22, 0, 8, 26, 31,
					-- layer=2 filter=20 channel=72
					11, 21, 25, 39, 5, 7, 15, 11, 45,
					-- layer=2 filter=20 channel=73
					-31, -3, 9, 12, 7, 16, 52, -2, -22,
					-- layer=2 filter=20 channel=74
					-10, -27, -15, -42, 6, 1, 17, 15, 11,
					-- layer=2 filter=20 channel=75
					0, 11, 43, -11, 0, 8, 0, 55, -15,
					-- layer=2 filter=20 channel=76
					46, -1, 19, 13, -19, -56, 35, -80, -88,
					-- layer=2 filter=20 channel=77
					-2, 0, -1, -4, -1, 4, -7, -4, -5,
					-- layer=2 filter=20 channel=78
					23, -7, 5, -36, -11, -8, 24, 20, -14,
					-- layer=2 filter=20 channel=79
					-7, 9, -6, -11, -1, -9, -9, -8, -9,
					-- layer=2 filter=20 channel=80
					-46, -12, 6, -22, 10, 16, 13, 28, 19,
					-- layer=2 filter=20 channel=81
					10, 10, 9, 3, 1, 0, -9, 2, 2,
					-- layer=2 filter=20 channel=82
					4, 6, -6, 0, 6, 0, -3, -9, -4,
					-- layer=2 filter=20 channel=83
					-29, 1, -14, -8, 5, -4, 8, 31, -19,
					-- layer=2 filter=20 channel=84
					-5, -3, 9, 5, 6, 10, -7, -10, 1,
					-- layer=2 filter=20 channel=85
					9, 8, 14, -18, 0, 13, -7, 0, 13,
					-- layer=2 filter=20 channel=86
					-8, -12, -9, 13, -26, 5, -5, 0, -5,
					-- layer=2 filter=20 channel=87
					-4, -21, -31, -24, -40, -21, -51, -55, -33,
					-- layer=2 filter=20 channel=88
					-4, -16, -6, -15, 24, 4, 5, 8, -14,
					-- layer=2 filter=20 channel=89
					-7, 24, 20, 43, 0, -5, 12, 28, -8,
					-- layer=2 filter=20 channel=90
					2, 7, 2, 2, -8, -4, 0, 0, 5,
					-- layer=2 filter=20 channel=91
					-11, 1, 4, 6, -38, -3, 2, 32, 5,
					-- layer=2 filter=20 channel=92
					31, 42, 1, 29, 12, 1, -21, 27, -14,
					-- layer=2 filter=20 channel=93
					0, 42, 36, -28, -14, -16, -44, 16, -5,
					-- layer=2 filter=20 channel=94
					18, 17, -31, 39, 10, -1, -10, 8, -45,
					-- layer=2 filter=20 channel=95
					0, 5, 15, 0, 2, -18, 20, -12, -3,
					-- layer=2 filter=20 channel=96
					-10, -37, -67, -61, -96, -111, -138, -146, -105,
					-- layer=2 filter=20 channel=97
					2, -10, -26, 15, 10, -8, 15, 30, -15,
					-- layer=2 filter=20 channel=98
					20, 44, 43, -3, 24, 36, 4, 7, 32,
					-- layer=2 filter=20 channel=99
					10, 8, -15, -44, -19, -23, -1, -69, -17,
					-- layer=2 filter=20 channel=100
					-21, -28, -13, 21, 0, -7, 27, 33, -28,
					-- layer=2 filter=20 channel=101
					0, -45, -40, 7, -28, 0, 38, 25, 10,
					-- layer=2 filter=20 channel=102
					-7, -42, -15, -62, -68, -74, -99, -60, -9,
					-- layer=2 filter=20 channel=103
					40, 16, -8, -20, 10, 0, 21, 18, 4,
					-- layer=2 filter=20 channel=104
					0, -2, -19, -10, -17, -7, -38, 34, -65,
					-- layer=2 filter=20 channel=105
					15, -50, -27, 39, 5, 24, -41, 36, -30,
					-- layer=2 filter=20 channel=106
					-4, -45, -45, 1, -16, -6, 13, 15, 21,
					-- layer=2 filter=20 channel=107
					16, -8, -22, 13, 17, 19, -9, -47, 41,
					-- layer=2 filter=20 channel=108
					15, 10, 13, 6, 29, -4, 7, -4, 19,
					-- layer=2 filter=20 channel=109
					18, 0, -2, 19, -4, 20, 20, -2, 9,
					-- layer=2 filter=20 channel=110
					-23, -7, 3, -20, 11, 11, 11, 18, 15,
					-- layer=2 filter=20 channel=111
					3, 1, -9, 4, 2, -1, 1, -4, -3,
					-- layer=2 filter=20 channel=112
					-13, 13, 0, -43, -11, -57, -36, 20, 17,
					-- layer=2 filter=20 channel=113
					-11, 26, 2, 0, 36, 1, -9, 11, 29,
					-- layer=2 filter=20 channel=114
					-7, 6, -13, 12, -4, 2, -6, -7, 0,
					-- layer=2 filter=20 channel=115
					-4, -1, 6, -11, -2, -3, -5, -7, -10,
					-- layer=2 filter=20 channel=116
					-13, -13, -36, -63, -29, -5, -28, -39, -45,
					-- layer=2 filter=20 channel=117
					17, 0, -12, 0, 27, 11, 7, 27, 50,
					-- layer=2 filter=20 channel=118
					-15, -4, 10, 0, -6, 0, 37, 20, 15,
					-- layer=2 filter=20 channel=119
					2, 24, 3, -1, 10, 27, -28, -11, 23,
					-- layer=2 filter=20 channel=120
					-9, 6, 2, 0, -6, 1, -5, -9, 7,
					-- layer=2 filter=20 channel=121
					9, -5, -5, -2, -9, 2, -2, -1, 4,
					-- layer=2 filter=20 channel=122
					0, -7, 8, -4, 2, 4, -10, -11, 0,
					-- layer=2 filter=20 channel=123
					28, 55, 17, 47, 20, 27, -4, 18, 17,
					-- layer=2 filter=20 channel=124
					26, 1, -22, 11, 2, 12, -14, 10, -41,
					-- layer=2 filter=20 channel=125
					0, 4, 8, 3, -6, 1, 9, 8, 8,
					-- layer=2 filter=20 channel=126
					32, -6, -56, 5, 37, -67, 3, 48, -41,
					-- layer=2 filter=20 channel=127
					23, 21, -4, 8, 0, 30, -28, -16, -14,
					-- layer=2 filter=21 channel=0
					-15, -18, -4, -8, -6, -10, -2, -1, 0,
					-- layer=2 filter=21 channel=1
					0, -3, -6, 0, -6, 0, -8, -3, -10,
					-- layer=2 filter=21 channel=2
					-7, 5, 7, 5, 5, 1, 0, -2, -5,
					-- layer=2 filter=21 channel=3
					-8, -14, -26, -22, -11, -9, -12, -13, -7,
					-- layer=2 filter=21 channel=4
					0, -11, -12, -11, -6, 0, 10, -4, -8,
					-- layer=2 filter=21 channel=5
					-7, -21, -16, 5, -28, -5, -6, -12, -19,
					-- layer=2 filter=21 channel=6
					-14, 1, -12, 6, -4, 0, -13, 0, -6,
					-- layer=2 filter=21 channel=7
					10, 13, -7, -15, -6, -2, -1, -15, -7,
					-- layer=2 filter=21 channel=8
					1, 1, -8, 3, -9, 2, -3, 0, 1,
					-- layer=2 filter=21 channel=9
					-22, -22, -1, -5, -19, -10, -3, -6, 0,
					-- layer=2 filter=21 channel=10
					0, -1, -3, -11, -13, -8, -8, -1, -3,
					-- layer=2 filter=21 channel=11
					-1, -4, -16, -17, -20, -14, -12, -4, -9,
					-- layer=2 filter=21 channel=12
					-9, -9, -1, 9, -5, 4, -3, -14, 0,
					-- layer=2 filter=21 channel=13
					10, 5, -5, 1, -8, 3, 2, 7, 5,
					-- layer=2 filter=21 channel=14
					-4, -3, -2, -3, -11, -3, -7, -25, -12,
					-- layer=2 filter=21 channel=15
					1, -26, -4, -16, -7, -26, 2, -22, 3,
					-- layer=2 filter=21 channel=16
					-11, 7, -11, -7, -3, -2, -8, -8, 2,
					-- layer=2 filter=21 channel=17
					-1, 0, -7, 6, -5, -10, 0, -5, -8,
					-- layer=2 filter=21 channel=18
					8, -4, 5, -11, -17, -2, -10, 6, -5,
					-- layer=2 filter=21 channel=19
					-5, -10, 6, 4, -11, -17, -12, -6, -12,
					-- layer=2 filter=21 channel=20
					9, -3, -5, 4, 8, -2, -6, 7, 9,
					-- layer=2 filter=21 channel=21
					0, -3, 0, -6, 5, 1, 10, -1, 7,
					-- layer=2 filter=21 channel=22
					-4, 4, 1, -7, -6, 6, -8, -1, -4,
					-- layer=2 filter=21 channel=23
					8, -5, 11, -3, -6, -1, 3, -2, -1,
					-- layer=2 filter=21 channel=24
					0, -6, -8, -5, -1, -15, -10, -21, -10,
					-- layer=2 filter=21 channel=25
					-10, -14, -9, -21, -5, -2, -2, -8, -13,
					-- layer=2 filter=21 channel=26
					3, -4, 9, -9, 4, -8, -10, 7, -2,
					-- layer=2 filter=21 channel=27
					-6, -4, -9, -21, -7, -2, -20, -10, -1,
					-- layer=2 filter=21 channel=28
					-8, -12, 0, -23, 0, 3, -4, -6, -10,
					-- layer=2 filter=21 channel=29
					-3, -5, -7, 7, -9, 8, -9, -1, 1,
					-- layer=2 filter=21 channel=30
					-12, -12, -11, -3, -7, -11, -10, 9, -6,
					-- layer=2 filter=21 channel=31
					-1, 6, 1, -11, 8, -1, 9, 3, -6,
					-- layer=2 filter=21 channel=32
					-5, -9, 1, 2, -6, -11, -1, -9, -8,
					-- layer=2 filter=21 channel=33
					1, 16, -6, 2, -10, 1, 0, -7, -7,
					-- layer=2 filter=21 channel=34
					7, -15, -6, -1, 2, -11, -6, 3, 4,
					-- layer=2 filter=21 channel=35
					-11, 0, 4, -16, 0, -7, -18, -7, -4,
					-- layer=2 filter=21 channel=36
					0, -9, 7, -1, -8, 1, -2, 6, -10,
					-- layer=2 filter=21 channel=37
					2, -11, 0, -10, -21, -21, -5, 0, -12,
					-- layer=2 filter=21 channel=38
					-15, -19, -18, -5, -12, -20, -10, -16, -2,
					-- layer=2 filter=21 channel=39
					-5, 1, 2, 2, 3, 1, -2, -2, -5,
					-- layer=2 filter=21 channel=40
					-3, 1, -12, -5, 3, 3, 0, -1, -13,
					-- layer=2 filter=21 channel=41
					-4, -7, -11, 0, 0, 0, 1, -5, -5,
					-- layer=2 filter=21 channel=42
					-10, -5, 2, 5, -10, -7, 4, -8, 10,
					-- layer=2 filter=21 channel=43
					-9, -22, -15, -1, 0, 7, -16, -4, 0,
					-- layer=2 filter=21 channel=44
					-2, -10, 9, -5, -7, -10, 6, 4, 2,
					-- layer=2 filter=21 channel=45
					15, 23, 2, 4, -13, 1, 11, -10, -5,
					-- layer=2 filter=21 channel=46
					1, 2, -20, -16, -11, 0, -3, 4, -7,
					-- layer=2 filter=21 channel=47
					6, -6, -6, -34, -6, -5, -10, -13, -10,
					-- layer=2 filter=21 channel=48
					-1, 4, -9, -6, -2, 0, -7, -6, -4,
					-- layer=2 filter=21 channel=49
					-5, -4, -10, -9, -7, 0, 7, -15, -6,
					-- layer=2 filter=21 channel=50
					-1, -2, -3, -4, -3, -3, -2, -12, 5,
					-- layer=2 filter=21 channel=51
					4, 0, 0, 2, -5, 0, 0, -6, -18,
					-- layer=2 filter=21 channel=52
					2, -11, -1, -6, 7, -7, 3, 0, -16,
					-- layer=2 filter=21 channel=53
					-4, -15, -8, 2, 0, -1, -4, -3, -20,
					-- layer=2 filter=21 channel=54
					-16, 3, -13, -5, -4, 0, -4, -8, 0,
					-- layer=2 filter=21 channel=55
					-8, -5, -10, 0, 8, 3, 9, 1, 5,
					-- layer=2 filter=21 channel=56
					1, -13, -12, -9, -5, -22, -11, -16, -18,
					-- layer=2 filter=21 channel=57
					-9, 5, -1, 4, 6, -3, -2, 0, -5,
					-- layer=2 filter=21 channel=58
					8, -13, -8, 2, 0, 2, 6, -10, -4,
					-- layer=2 filter=21 channel=59
					-16, -18, -12, -14, -14, -13, -9, -7, -3,
					-- layer=2 filter=21 channel=60
					-4, -19, -14, 3, -7, 0, -8, -4, 3,
					-- layer=2 filter=21 channel=61
					7, -7, 2, -8, 4, -16, -14, -1, -10,
					-- layer=2 filter=21 channel=62
					-3, 7, 5, 3, -16, -5, 8, 0, -12,
					-- layer=2 filter=21 channel=63
					-17, -19, -5, -1, -1, 2, 0, 4, 7,
					-- layer=2 filter=21 channel=64
					-4, -14, -1, -4, -5, -12, -10, -4, -15,
					-- layer=2 filter=21 channel=65
					0, 9, 6, 2, -6, -25, -5, -8, 6,
					-- layer=2 filter=21 channel=66
					0, 6, -5, 3, 5, -1, -3, -6, 1,
					-- layer=2 filter=21 channel=67
					-1, -14, -1, -13, -16, -5, -16, -15, -13,
					-- layer=2 filter=21 channel=68
					-8, -6, 1, -7, -7, -11, -10, -6, -9,
					-- layer=2 filter=21 channel=69
					-2, -7, -15, -7, -13, -9, 6, 3, -1,
					-- layer=2 filter=21 channel=70
					-14, -2, -5, 0, -6, -2, -14, -2, 3,
					-- layer=2 filter=21 channel=71
					-10, -12, -10, 3, -17, -4, -3, -13, -10,
					-- layer=2 filter=21 channel=72
					-5, 7, -1, -11, -3, -19, -19, 1, -8,
					-- layer=2 filter=21 channel=73
					-22, -17, -8, -24, 1, 2, 13, -17, 8,
					-- layer=2 filter=21 channel=74
					-18, -6, -13, -15, 0, -13, -4, -15, -1,
					-- layer=2 filter=21 channel=75
					-16, 0, -8, -19, 1, 4, -8, -16, -2,
					-- layer=2 filter=21 channel=76
					-18, 0, -12, -16, -3, 7, 7, -7, -10,
					-- layer=2 filter=21 channel=77
					7, 5, -5, -10, -6, -9, -7, 5, 0,
					-- layer=2 filter=21 channel=78
					7, -4, -11, -10, -11, -21, -6, -14, -11,
					-- layer=2 filter=21 channel=79
					8, -1, -4, 0, -1, -10, 0, 1, 1,
					-- layer=2 filter=21 channel=80
					-14, 3, 3, 0, 2, -9, -7, 1, -18,
					-- layer=2 filter=21 channel=81
					-5, -6, 8, -4, -4, 8, 1, -5, 4,
					-- layer=2 filter=21 channel=82
					8, 6, -7, 2, -2, 3, -5, 3, 2,
					-- layer=2 filter=21 channel=83
					-14, 1, -6, -4, -8, -9, -8, 7, -2,
					-- layer=2 filter=21 channel=84
					-3, 7, -5, 5, -6, -7, -1, -10, 0,
					-- layer=2 filter=21 channel=85
					-8, 7, 7, 9, 6, 4, -9, -10, 6,
					-- layer=2 filter=21 channel=86
					2, 2, 7, -10, 7, 9, -7, -9, -4,
					-- layer=2 filter=21 channel=87
					7, 2, 0, -23, 1, -2, 10, 1, -4,
					-- layer=2 filter=21 channel=88
					-17, -4, -7, 0, -3, -7, -8, -10, -10,
					-- layer=2 filter=21 channel=89
					-1, -1, -13, -8, -15, 0, -5, -10, -3,
					-- layer=2 filter=21 channel=90
					-7, 3, 0, 5, 7, 1, 0, -9, -5,
					-- layer=2 filter=21 channel=91
					-15, -2, 1, -13, -6, 0, 2, -21, -5,
					-- layer=2 filter=21 channel=92
					0, -4, -2, -1, -4, -6, 0, -9, 4,
					-- layer=2 filter=21 channel=93
					0, -7, 1, 4, 5, 2, -23, 0, 7,
					-- layer=2 filter=21 channel=94
					-2, 12, -11, -10, 1, 4, -14, -4, 0,
					-- layer=2 filter=21 channel=95
					-4, 1, -1, -10, -3, -8, 8, -5, 6,
					-- layer=2 filter=21 channel=96
					-1, -2, 4, 6, 8, -3, -8, 3, -13,
					-- layer=2 filter=21 channel=97
					-22, -18, -28, -18, -23, -19, -13, -2, -19,
					-- layer=2 filter=21 channel=98
					1, -2, -5, -14, -2, -5, -3, -7, -4,
					-- layer=2 filter=21 channel=99
					-10, -12, 8, 10, 0, -15, 4, -7, -6,
					-- layer=2 filter=21 channel=100
					-1, -2, -24, -10, -18, 5, -5, 5, -6,
					-- layer=2 filter=21 channel=101
					-14, -5, -8, -12, -11, -9, -13, -17, -12,
					-- layer=2 filter=21 channel=102
					5, -3, -9, 5, -1, -8, -4, 3, -9,
					-- layer=2 filter=21 channel=103
					-6, -8, -10, -1, -5, -12, -8, -5, -4,
					-- layer=2 filter=21 channel=104
					-5, 1, -25, -9, -13, -3, 2, -11, -16,
					-- layer=2 filter=21 channel=105
					9, 9, 15, -6, 3, -4, 5, -8, -5,
					-- layer=2 filter=21 channel=106
					-14, -14, -3, -13, -18, -11, -3, -13, -21,
					-- layer=2 filter=21 channel=107
					-2, -9, -9, 2, -10, 5, -6, 0, -5,
					-- layer=2 filter=21 channel=108
					-8, -21, -2, -8, -12, -13, -13, -21, -11,
					-- layer=2 filter=21 channel=109
					-12, -2, -7, -4, 6, -1, -9, -9, -1,
					-- layer=2 filter=21 channel=110
					-14, -10, -5, -4, -12, -3, -2, 3, -4,
					-- layer=2 filter=21 channel=111
					8, -5, -4, -6, 10, 0, -10, 1, -8,
					-- layer=2 filter=21 channel=112
					-5, -3, 0, 8, -13, -12, 0, -4, -19,
					-- layer=2 filter=21 channel=113
					0, 5, 10, 4, 0, -12, -5, 9, -12,
					-- layer=2 filter=21 channel=114
					-2, 10, -6, -1, 11, 8, 5, 8, 7,
					-- layer=2 filter=21 channel=115
					-4, 8, 8, 1, 7, 7, 10, 9, 10,
					-- layer=2 filter=21 channel=116
					11, 0, -18, -12, -6, -20, -2, -5, -18,
					-- layer=2 filter=21 channel=117
					0, 4, -1, -7, 0, -13, -5, 6, -7,
					-- layer=2 filter=21 channel=118
					-11, -22, -4, -9, -11, -3, -11, -13, -11,
					-- layer=2 filter=21 channel=119
					-9, 0, 7, 0, -16, 0, -1, -3, -13,
					-- layer=2 filter=21 channel=120
					0, -2, 6, 9, -6, 6, 4, 8, -8,
					-- layer=2 filter=21 channel=121
					-2, 4, 5, -9, 6, -2, 11, -3, 6,
					-- layer=2 filter=21 channel=122
					-8, -7, -4, 4, 11, 10, 9, 3, -4,
					-- layer=2 filter=21 channel=123
					7, -7, 0, -22, -11, -9, -2, -6, -9,
					-- layer=2 filter=21 channel=124
					4, -17, 4, -9, -4, -28, 21, -7, -9,
					-- layer=2 filter=21 channel=125
					1, 6, -8, 6, -6, 7, 1, -3, -7,
					-- layer=2 filter=21 channel=126
					-13, -16, 0, -6, -13, 9, -19, -4, -8,
					-- layer=2 filter=21 channel=127
					-16, -2, -9, -7, 6, 1, -15, -6, -6,
					-- layer=2 filter=22 channel=0
					5, 0, -15, 25, 9, 18, -8, -5, -2,
					-- layer=2 filter=22 channel=1
					-2, -8, 27, -13, -25, -22, 16, 26, 16,
					-- layer=2 filter=22 channel=2
					-2, -7, 0, -12, -10, 0, -8, -6, -9,
					-- layer=2 filter=22 channel=3
					11, 10, -18, -7, 7, 7, 10, -6, -4,
					-- layer=2 filter=22 channel=4
					1, 31, 0, -30, -7, 6, -42, -61, -16,
					-- layer=2 filter=22 channel=5
					-22, -36, -5, 21, 4, 15, -1, 9, 12,
					-- layer=2 filter=22 channel=6
					-13, 26, -1, -19, -113, -52, 15, 3, 10,
					-- layer=2 filter=22 channel=7
					53, 31, 31, 13, 36, 18, 6, -49, -22,
					-- layer=2 filter=22 channel=8
					0, 0, -2, 7, -5, 0, -9, 8, 0,
					-- layer=2 filter=22 channel=9
					-29, -8, 3, 36, 11, 29, 39, 17, 16,
					-- layer=2 filter=22 channel=10
					-2, -2, 7, 3, 11, 0, 7, 13, -9,
					-- layer=2 filter=22 channel=11
					-7, 1, -13, 12, 21, 15, 24, -13, 5,
					-- layer=2 filter=22 channel=12
					19, -11, 47, 6, 21, 11, 7, 17, 16,
					-- layer=2 filter=22 channel=13
					-1, -4, -5, 5, -6, -9, 8, 5, 5,
					-- layer=2 filter=22 channel=14
					0, -19, 0, 33, 12, 6, 5, 21, -9,
					-- layer=2 filter=22 channel=15
					-29, 17, -64, 59, 10, -26, -9, 22, 13,
					-- layer=2 filter=22 channel=16
					19, 16, -22, 20, 42, 0, -18, -25, 9,
					-- layer=2 filter=22 channel=17
					-5, -6, 9, 5, -8, -3, -10, -7, -9,
					-- layer=2 filter=22 channel=18
					-7, 9, 20, 12, -22, -27, 27, -15, -3,
					-- layer=2 filter=22 channel=19
					-24, 2, 12, 1, -17, -2, 21, 34, 11,
					-- layer=2 filter=22 channel=20
					-9, -3, 1, -4, 5, -4, -8, 1, -2,
					-- layer=2 filter=22 channel=21
					-13, -12, -7, 11, -1, 1, -2, -4, -4,
					-- layer=2 filter=22 channel=22
					-4, -6, 9, 4, -4, 4, 5, 3, 2,
					-- layer=2 filter=22 channel=23
					4, 38, 33, -11, 0, 26, -68, -30, 8,
					-- layer=2 filter=22 channel=24
					4, 4, -9, -8, -6, 11, -4, -16, 0,
					-- layer=2 filter=22 channel=25
					13, 3, -22, 1, 21, 8, 0, -2, -5,
					-- layer=2 filter=22 channel=26
					2, -8, -5, -9, 2, 9, 3, -2, -2,
					-- layer=2 filter=22 channel=27
					-35, -38, -26, 21, 25, 7, 10, -3, -23,
					-- layer=2 filter=22 channel=28
					14, 18, 18, 38, 59, 32, -65, -59, -56,
					-- layer=2 filter=22 channel=29
					-5, -8, 0, 0, -8, -7, 5, -3, -3,
					-- layer=2 filter=22 channel=30
					17, -13, 31, 2, 15, -1, 2, -4, -6,
					-- layer=2 filter=22 channel=31
					-3, 21, -4, -3, 30, 38, 26, -4, 16,
					-- layer=2 filter=22 channel=32
					-2, -2, 5, -6, 1, 9, 2, 8, 5,
					-- layer=2 filter=22 channel=33
					10, 16, -15, -8, 42, -9, -43, -50, -24,
					-- layer=2 filter=22 channel=34
					-15, -7, 20, 5, 4, -88, -8, 8, 3,
					-- layer=2 filter=22 channel=35
					21, 7, 18, 5, 13, -3, -14, -21, 2,
					-- layer=2 filter=22 channel=36
					6, 17, 11, 8, 7, -6, 8, 0, -5,
					-- layer=2 filter=22 channel=37
					-16, -36, -10, 4, 16, 7, 8, 2, -14,
					-- layer=2 filter=22 channel=38
					-36, -42, -23, 3, 1, 15, 18, 4, -6,
					-- layer=2 filter=22 channel=39
					26, 10, -6, -10, 21, 31, -7, -4, 6,
					-- layer=2 filter=22 channel=40
					-29, -7, -44, 21, -13, -39, 11, 13, -20,
					-- layer=2 filter=22 channel=41
					6, -10, 3, -4, -8, 5, 8, 8, -6,
					-- layer=2 filter=22 channel=42
					4, 37, 30, 0, 25, 42, -50, -9, 0,
					-- layer=2 filter=22 channel=43
					-18, 3, -7, 15, 0, 14, -2, -2, 14,
					-- layer=2 filter=22 channel=44
					0, 3, -2, -5, 3, -3, -10, 5, 0,
					-- layer=2 filter=22 channel=45
					12, 0, -27, 32, 34, -6, -2, -24, -53,
					-- layer=2 filter=22 channel=46
					0, -2, 6, 3, -5, -12, 1, -1, -31,
					-- layer=2 filter=22 channel=47
					15, 33, 19, 64, 96, 42, -46, -69, -90,
					-- layer=2 filter=22 channel=48
					2, -2, -10, -10, 1, -8, -1, 3, -4,
					-- layer=2 filter=22 channel=49
					-14, 17, 4, -6, -46, -46, 26, 6, 12,
					-- layer=2 filter=22 channel=50
					-2, -7, -2, -3, 8, 2, 9, 23, 0,
					-- layer=2 filter=22 channel=51
					-18, -36, -18, 25, 7, 12, 14, -6, -21,
					-- layer=2 filter=22 channel=52
					-30, -17, 14, 1, -13, 11, 14, -11, -3,
					-- layer=2 filter=22 channel=53
					39, -27, -14, 17, -64, 5, 45, 1, -22,
					-- layer=2 filter=22 channel=54
					36, 28, 48, -20, 16, 15, -56, -44, -14,
					-- layer=2 filter=22 channel=55
					0, -6, 1, -2, -13, 1, 5, 9, 5,
					-- layer=2 filter=22 channel=56
					-30, -23, -13, 20, 19, 28, 46, 10, 16,
					-- layer=2 filter=22 channel=57
					4, -5, 3, 14, 0, -14, -10, 16, -5,
					-- layer=2 filter=22 channel=58
					13, 1, 26, -5, 16, 50, -9, 32, 52,
					-- layer=2 filter=22 channel=59
					17, 5, -2, -19, -19, -50, 2, 4, 12,
					-- layer=2 filter=22 channel=60
					-35, -13, -10, -8, -11, 16, 6, 26, 44,
					-- layer=2 filter=22 channel=61
					-34, -24, -32, 19, -42, -47, 21, -31, -22,
					-- layer=2 filter=22 channel=62
					1, 20, -4, 20, -103, -24, 18, 15, 63,
					-- layer=2 filter=22 channel=63
					-7, 29, 15, 14, 0, -11, -35, 6, 12,
					-- layer=2 filter=22 channel=64
					7, 10, 11, -20, 8, 3, -59, -31, -5,
					-- layer=2 filter=22 channel=65
					-11, 0, -9, -37, -79, -45, 10, -47, 1,
					-- layer=2 filter=22 channel=66
					20, 37, 29, -30, -28, 46, 7, -53, 5,
					-- layer=2 filter=22 channel=67
					-35, -44, -54, -14, 6, -11, -32, 35, -3,
					-- layer=2 filter=22 channel=68
					0, -6, 7, -3, 6, 2, 8, -7, -1,
					-- layer=2 filter=22 channel=69
					16, 26, 5, 14, 10, 19, -33, -11, 26,
					-- layer=2 filter=22 channel=70
					-2, 15, 9, 34, 34, 0, -36, -18, -30,
					-- layer=2 filter=22 channel=71
					-29, -36, -47, 0, 27, 1, 16, 7, -6,
					-- layer=2 filter=22 channel=72
					-4, 8, 18, 19, 15, -12, 24, -4, -34,
					-- layer=2 filter=22 channel=73
					-21, -58, -26, -51, -91, -61, 69, 23, 36,
					-- layer=2 filter=22 channel=74
					-6, -13, -6, 3, 15, -17, -41, 6, -18,
					-- layer=2 filter=22 channel=75
					0, -45, -34, 8, 0, 8, 26, -9, 13,
					-- layer=2 filter=22 channel=76
					-38, -21, -7, 3, -88, -22, -30, -30, 13,
					-- layer=2 filter=22 channel=77
					-3, -7, -9, -9, -4, 6, 8, -4, -3,
					-- layer=2 filter=22 channel=78
					0, 10, -15, -19, -21, -9, 12, -28, 0,
					-- layer=2 filter=22 channel=79
					-5, -10, -5, -5, 2, -7, -2, -11, -9,
					-- layer=2 filter=22 channel=80
					-5, 0, -24, -10, -3, -10, -38, -9, -17,
					-- layer=2 filter=22 channel=81
					-4, -4, -5, 1, 2, 17, -3, 0, -4,
					-- layer=2 filter=22 channel=82
					1, 11, 10, -9, 6, 0, -8, -6, 7,
					-- layer=2 filter=22 channel=83
					-2, -5, 17, -11, 11, -5, -44, -10, -28,
					-- layer=2 filter=22 channel=84
					2, -1, -9, 1, 6, -12, -1, -3, -6,
					-- layer=2 filter=22 channel=85
					-14, -10, 7, -17, -3, 1, -5, 8, 5,
					-- layer=2 filter=22 channel=86
					-4, -1, 12, -2, 9, 3, 0, 15, 7,
					-- layer=2 filter=22 channel=87
					0, -19, -6, -61, -48, 24, -28, -68, 29,
					-- layer=2 filter=22 channel=88
					9, -1, 18, -8, -10, -3, -36, -8, -7,
					-- layer=2 filter=22 channel=89
					-12, 2, 17, 8, -9, 14, 6, 27, 31,
					-- layer=2 filter=22 channel=90
					10, 8, 8, -7, -9, -6, -5, 1, 7,
					-- layer=2 filter=22 channel=91
					-2, 8, -7, 19, 21, 31, 11, 36, 22,
					-- layer=2 filter=22 channel=92
					0, 3, 39, 14, 4, 13, 11, 37, 7,
					-- layer=2 filter=22 channel=93
					5, 42, 50, -13, -51, 21, 0, 60, 68,
					-- layer=2 filter=22 channel=94
					-11, 0, 7, -16, -63, -44, 31, 19, 47,
					-- layer=2 filter=22 channel=95
					-1, 5, -6, -8, 11, -5, 8, -1, 7,
					-- layer=2 filter=22 channel=96
					-37, -68, -23, -97, -105, -28, -73, -14, 8,
					-- layer=2 filter=22 channel=97
					-1, 3, -51, 9, 39, 5, -1, -15, 18,
					-- layer=2 filter=22 channel=98
					16, 5, 22, 46, 50, 22, -40, -66, -66,
					-- layer=2 filter=22 channel=99
					-16, -25, -19, -58, -51, -42, 51, 22, 31,
					-- layer=2 filter=22 channel=100
					-36, 11, 8, -12, 15, 28, -19, 21, 16,
					-- layer=2 filter=22 channel=101
					-14, 9, -5, 16, 33, 32, 13, -4, -16,
					-- layer=2 filter=22 channel=102
					-16, -27, 2, -32, -49, -19, 0, -19, 44,
					-- layer=2 filter=22 channel=103
					-53, -18, -17, -16, -18, 22, -27, -7, -10,
					-- layer=2 filter=22 channel=104
					-5, 10, -8, -53, -57, -29, -8, -10, -9,
					-- layer=2 filter=22 channel=105
					-24, 0, 59, -6, -31, -28, -51, -46, 6,
					-- layer=2 filter=22 channel=106
					-7, -13, -33, 23, 17, 26, 6, 3, 4,
					-- layer=2 filter=22 channel=107
					-26, -30, -6, 40, 65, 29, 81, 0, 13,
					-- layer=2 filter=22 channel=108
					-43, -35, -16, 31, 0, -27, 0, 32, -14,
					-- layer=2 filter=22 channel=109
					0, -7, 6, -8, -7, 9, 4, -4, 10,
					-- layer=2 filter=22 channel=110
					-31, 26, 20, -40, 3, 3, -54, -21, -3,
					-- layer=2 filter=22 channel=111
					0, 7, -6, -4, -6, 2, 7, -9, -5,
					-- layer=2 filter=22 channel=112
					-31, -23, 0, 26, 3, 6, 10, 10, -22,
					-- layer=2 filter=22 channel=113
					30, 3, -3, 6, -28, -13, -40, -24, 6,
					-- layer=2 filter=22 channel=114
					6, 11, 15, 3, -4, -5, -3, 7, 5,
					-- layer=2 filter=22 channel=115
					-8, 4, 6, -1, -13, 5, -4, 1, -13,
					-- layer=2 filter=22 channel=116
					11, -73, -16, -27, -38, 19, -41, -22, 19,
					-- layer=2 filter=22 channel=117
					-14, -5, 38, -11, 22, -4, 14, -16, -32,
					-- layer=2 filter=22 channel=118
					5, 10, -17, -24, -16, 31, -9, -24, 25,
					-- layer=2 filter=22 channel=119
					18, 45, 11, 24, 1, -23, -16, -35, -20,
					-- layer=2 filter=22 channel=120
					8, 0, -2, 8, 0, 4, 5, -9, -5,
					-- layer=2 filter=22 channel=121
					-7, 6, -9, 5, -6, -4, 8, 9, 2,
					-- layer=2 filter=22 channel=122
					-11, -9, -5, -7, -12, -12, -18, -1, -9,
					-- layer=2 filter=22 channel=123
					17, 22, 26, 6, 49, 28, -26, -49, -6,
					-- layer=2 filter=22 channel=124
					-38, 35, -9, 34, 17, 43, -48, -25, 10,
					-- layer=2 filter=22 channel=125
					8, 0, 9, 5, 8, 5, 5, 4, 6,
					-- layer=2 filter=22 channel=126
					-48, 26, -36, 18, 0, -5, 16, 43, 40,
					-- layer=2 filter=22 channel=127
					-1, 1, 7, -16, -14, -10, -16, -4, 19,
					-- layer=2 filter=23 channel=0
					27, 12, -6, 1, -17, -7, -2, -18, 12,
					-- layer=2 filter=23 channel=1
					-2, 29, -9, 7, -10, -21, 8, 21, 19,
					-- layer=2 filter=23 channel=2
					0, 4, 0, 0, -2, 12, -4, -2, 10,
					-- layer=2 filter=23 channel=3
					19, -7, -5, -30, -17, 5, 10, 3, 20,
					-- layer=2 filter=23 channel=4
					13, 10, 14, 11, -26, -14, 2, -5, -22,
					-- layer=2 filter=23 channel=5
					17, 32, 14, 19, 19, 12, 16, -20, 3,
					-- layer=2 filter=23 channel=6
					-23, -34, -14, -10, -59, -24, -9, -4, 13,
					-- layer=2 filter=23 channel=7
					32, -40, -5, 12, 40, -22, -2, 19, -19,
					-- layer=2 filter=23 channel=8
					-5, 7, 1, -7, 6, 9, 8, 4, 8,
					-- layer=2 filter=23 channel=9
					-4, -13, 14, -1, -1, 16, -3, -4, 12,
					-- layer=2 filter=23 channel=10
					25, 9, -1, 44, -8, -12, -12, -15, -1,
					-- layer=2 filter=23 channel=11
					-17, -17, 0, -3, 1, 27, -20, 3, 23,
					-- layer=2 filter=23 channel=12
					10, -9, -40, 9, 2, -13, 8, 1, 5,
					-- layer=2 filter=23 channel=13
					13, 0, 1, -7, 0, -6, -6, 3, 9,
					-- layer=2 filter=23 channel=14
					-27, -33, -58, 7, -15, -24, 4, -2, 27,
					-- layer=2 filter=23 channel=15
					-41, 13, 9, -8, 10, 55, -12, -20, -9,
					-- layer=2 filter=23 channel=16
					25, 12, -38, -27, -14, -44, -20, -29, -63,
					-- layer=2 filter=23 channel=17
					3, 1, -4, -10, -2, -6, 8, 2, 1,
					-- layer=2 filter=23 channel=18
					-10, -11, 12, -23, -23, 15, -11, -21, -27,
					-- layer=2 filter=23 channel=19
					13, 33, 0, 6, 17, -26, -2, -22, -11,
					-- layer=2 filter=23 channel=20
					-3, -7, 7, -7, 0, 5, 8, 7, -8,
					-- layer=2 filter=23 channel=21
					-12, 3, 5, -15, -20, -12, -1, -2, -4,
					-- layer=2 filter=23 channel=22
					-8, -5, -1, -8, 4, 6, 8, 7, -4,
					-- layer=2 filter=23 channel=23
					8, 4, -14, -17, -25, -1, -11, -7, 5,
					-- layer=2 filter=23 channel=24
					-6, 3, -17, -20, 0, 12, -8, 26, 41,
					-- layer=2 filter=23 channel=25
					-21, 3, -14, -32, 11, 34, -18, 27, 53,
					-- layer=2 filter=23 channel=26
					-6, -3, 5, 6, 7, -8, 3, 10, 0,
					-- layer=2 filter=23 channel=27
					-10, -24, 34, 16, -5, -5, 19, -6, -16,
					-- layer=2 filter=23 channel=28
					-2, 47, -2, 22, 24, 0, 47, 16, 10,
					-- layer=2 filter=23 channel=29
					-8, -4, 1, 10, 0, 4, -11, -1, -7,
					-- layer=2 filter=23 channel=30
					-7, 8, -15, -2, -14, 7, 11, -28, -21,
					-- layer=2 filter=23 channel=31
					14, -15, -30, -24, -38, 8, -12, -24, 14,
					-- layer=2 filter=23 channel=32
					-5, -7, 9, 2, 11, 4, -9, -6, 9,
					-- layer=2 filter=23 channel=33
					13, -26, -3, -23, -7, -23, -61, 31, 22,
					-- layer=2 filter=23 channel=34
					-2, 49, 14, -7, 48, 16, 0, 14, -11,
					-- layer=2 filter=23 channel=35
					-4, 12, -4, 8, 24, 4, -18, 39, -8,
					-- layer=2 filter=23 channel=36
					1, 2, 7, 8, 1, -7, -6, -6, -4,
					-- layer=2 filter=23 channel=37
					-13, 10, 13, -2, 20, 34, 16, -11, 10,
					-- layer=2 filter=23 channel=38
					13, 18, -13, 17, 11, 11, 36, 2, 1,
					-- layer=2 filter=23 channel=39
					24, 4, 22, 6, 35, 13, -41, -21, 9,
					-- layer=2 filter=23 channel=40
					14, 31, 37, -33, 3, 37, -9, -2, 17,
					-- layer=2 filter=23 channel=41
					-3, 3, -4, 7, 1, -5, -10, 0, 7,
					-- layer=2 filter=23 channel=42
					-16, -3, -20, -7, -8, -3, -23, -4, -11,
					-- layer=2 filter=23 channel=43
					14, 32, 62, -16, -3, 30, -25, -34, -4,
					-- layer=2 filter=23 channel=44
					-7, 1, 4, 7, 3, 11, 9, -11, -6,
					-- layer=2 filter=23 channel=45
					-21, -9, 0, -14, -6, 7, 19, -19, -12,
					-- layer=2 filter=23 channel=46
					0, 1, 40, 8, 14, 1, -6, -7, -23,
					-- layer=2 filter=23 channel=47
					-12, 28, -18, 20, -9, -9, 6, 16, 9,
					-- layer=2 filter=23 channel=48
					10, 3, 1, 5, -6, -8, 5, 0, 1,
					-- layer=2 filter=23 channel=49
					-53, -20, -11, -46, -31, -13, -1, -25, -28,
					-- layer=2 filter=23 channel=50
					-19, -22, 0, 27, 10, -2, 0, -2, 25,
					-- layer=2 filter=23 channel=51
					-4, -11, -14, -14, 5, 8, -17, -11, 14,
					-- layer=2 filter=23 channel=52
					1, 0, 43, 12, 8, 23, -7, 3, 3,
					-- layer=2 filter=23 channel=53
					-4, -56, -35, 0, -5, -46, -64, -35, -1,
					-- layer=2 filter=23 channel=54
					23, 19, -35, 16, 13, 22, -5, 22, 46,
					-- layer=2 filter=23 channel=55
					-8, -3, -3, 4, 9, 6, 8, -9, -9,
					-- layer=2 filter=23 channel=56
					-11, -3, 20, 14, -4, 15, -13, -16, 1,
					-- layer=2 filter=23 channel=57
					1, 12, 8, 1, -12, -19, -2, -12, -14,
					-- layer=2 filter=23 channel=58
					18, 13, -42, 62, 26, 10, 38, 3, 2,
					-- layer=2 filter=23 channel=59
					13, 28, 44, 61, 18, -10, 44, 25, 15,
					-- layer=2 filter=23 channel=60
					21, 29, -8, 44, 18, -27, 29, 10, -4,
					-- layer=2 filter=23 channel=61
					-36, -31, -68, 1, -30, -89, 3, -4, -21,
					-- layer=2 filter=23 channel=62
					-16, -8, -7, -5, 9, 16, 18, 7, 13,
					-- layer=2 filter=23 channel=63
					-12, 22, 5, -1, -11, -12, 20, -9, 18,
					-- layer=2 filter=23 channel=64
					-10, 9, 0, -18, 14, 4, -39, -1, -18,
					-- layer=2 filter=23 channel=65
					-6, -11, -24, -3, -19, -39, 5, -15, 20,
					-- layer=2 filter=23 channel=66
					31, 0, 10, 37, -10, -23, 31, 8, 25,
					-- layer=2 filter=23 channel=67
					-15, -9, 40, -3, -1, 27, -1, -2, 18,
					-- layer=2 filter=23 channel=68
					2, 0, 9, -4, -9, -3, 10, 8, -9,
					-- layer=2 filter=23 channel=69
					-29, 0, -1, -17, 3, -3, -14, 5, -11,
					-- layer=2 filter=23 channel=70
					15, 25, -12, 30, 2, 21, 24, -7, -15,
					-- layer=2 filter=23 channel=71
					-11, -16, 7, -1, -1, 7, -8, 13, 37,
					-- layer=2 filter=23 channel=72
					15, -22, -4, -29, -36, -29, -26, 34, 7,
					-- layer=2 filter=23 channel=73
					38, 19, 13, 11, 40, 34, 12, -10, 42,
					-- layer=2 filter=23 channel=74
					-1, 20, 20, -16, 10, 47, 8, 0, -8,
					-- layer=2 filter=23 channel=75
					-80, -92, -31, -56, 0, -62, -10, -58, -17,
					-- layer=2 filter=23 channel=76
					9, -28, -23, 28, -17, -23, -52, -55, 6,
					-- layer=2 filter=23 channel=77
					-6, -1, -1, 10, 0, 4, 8, 7, 3,
					-- layer=2 filter=23 channel=78
					-22, -21, -5, -26, 0, 7, -14, 4, 23,
					-- layer=2 filter=23 channel=79
					-1, 0, -1, -1, 8, -1, 0, -1, -10,
					-- layer=2 filter=23 channel=80
					48, -5, 2, 3, 16, -7, -10, -21, -16,
					-- layer=2 filter=23 channel=81
					3, -6, 6, -5, -3, 12, 5, -11, -9,
					-- layer=2 filter=23 channel=82
					-3, -9, 8, 2, -1, -9, 6, 1, -9,
					-- layer=2 filter=23 channel=83
					6, 31, -12, -12, -2, -33, 10, -17, -22,
					-- layer=2 filter=23 channel=84
					-5, 3, 6, 13, -2, 7, -2, -9, -8,
					-- layer=2 filter=23 channel=85
					8, 2, 0, -7, 11, 17, 1, -1, 0,
					-- layer=2 filter=23 channel=86
					7, 0, -5, 5, -8, -1, 6, 7, -10,
					-- layer=2 filter=23 channel=87
					44, 43, 23, 42, 49, 11, 39, 29, 7,
					-- layer=2 filter=23 channel=88
					-21, -6, 2, -3, -5, 2, 12, 27, -20,
					-- layer=2 filter=23 channel=89
					-9, -11, -20, 11, 0, -46, 5, -1, -4,
					-- layer=2 filter=23 channel=90
					7, 4, -6, -9, -7, -7, 0, -6, 8,
					-- layer=2 filter=23 channel=91
					10, -15, -16, 27, -13, -34, -2, -5, -30,
					-- layer=2 filter=23 channel=92
					0, -3, -9, 27, -39, -42, -4, 9, -13,
					-- layer=2 filter=23 channel=93
					15, 5, -31, -40, -18, -44, -13, 2, 14,
					-- layer=2 filter=23 channel=94
					-38, -21, -15, -12, -45, -35, 23, -4, 42,
					-- layer=2 filter=23 channel=95
					-7, -11, -2, -10, 9, -3, -1, -4, -5,
					-- layer=2 filter=23 channel=96
					-11, -27, -54, 8, -17, -35, 17, 24, -22,
					-- layer=2 filter=23 channel=97
					15, 1, -2, -2, 29, -7, -32, 21, 10,
					-- layer=2 filter=23 channel=98
					-10, 20, -3, 6, 11, -7, 20, 38, 9,
					-- layer=2 filter=23 channel=99
					-15, 12, 28, 36, 12, -3, 36, -13, 37,
					-- layer=2 filter=23 channel=100
					4, 20, 18, 29, 51, 23, 22, -9, -4,
					-- layer=2 filter=23 channel=101
					-28, -46, -6, -17, -9, 21, -16, 31, 63,
					-- layer=2 filter=23 channel=102
					-23, -9, -33, 2, -39, -35, 33, 0, -39,
					-- layer=2 filter=23 channel=103
					-66, -55, -83, -12, -46, -64, 14, -3, -1,
					-- layer=2 filter=23 channel=104
					-33, -33, -21, -37, -20, -45, -37, -4, -14,
					-- layer=2 filter=23 channel=105
					32, 0, -43, 38, -1, -18, 1, -25, -41,
					-- layer=2 filter=23 channel=106
					3, -10, -26, 9, -1, 9, -2, 4, 17,
					-- layer=2 filter=23 channel=107
					-56, -68, -7, -30, -17, -8, -15, -4, -32,
					-- layer=2 filter=23 channel=108
					-16, -30, -34, 10, -2, -19, 32, -3, 20,
					-- layer=2 filter=23 channel=109
					17, 13, -5, -1, 7, 6, -3, 4, 3,
					-- layer=2 filter=23 channel=110
					-31, 13, -5, -47, -7, 17, -23, 46, 9,
					-- layer=2 filter=23 channel=111
					-10, -3, -9, -2, 0, 9, 6, 3, -6,
					-- layer=2 filter=23 channel=112
					-35, -23, -27, -4, -21, -49, -15, -8, -17,
					-- layer=2 filter=23 channel=113
					-21, 2, -8, 3, -29, -40, -7, 13, -63,
					-- layer=2 filter=23 channel=114
					-6, 20, -4, 2, 15, 8, 12, 19, -3,
					-- layer=2 filter=23 channel=115
					3, 9, -4, -7, 3, -6, -3, 4, 2,
					-- layer=2 filter=23 channel=116
					1, 51, 18, 31, 29, 4, 51, 36, 28,
					-- layer=2 filter=23 channel=117
					18, -18, -13, 7, 42, -69, -16, 1, -13,
					-- layer=2 filter=23 channel=118
					46, -5, 45, -3, 0, 32, -24, 16, 11,
					-- layer=2 filter=23 channel=119
					-9, 0, -2, -22, 2, 2, -19, 25, -10,
					-- layer=2 filter=23 channel=120
					4, -8, 3, -6, 8, 5, -1, 6, 3,
					-- layer=2 filter=23 channel=121
					1, -6, 7, 8, 5, -4, 5, -7, -7,
					-- layer=2 filter=23 channel=122
					10, -1, 9, 22, 10, 8, -3, 0, 5,
					-- layer=2 filter=23 channel=123
					8, 8, 35, 25, 13, -26, 6, -11, 4,
					-- layer=2 filter=23 channel=124
					50, -2, 11, -4, -15, -7, -65, -29, -9,
					-- layer=2 filter=23 channel=125
					0, 2, 10, -7, -2, -2, 0, -7, 0,
					-- layer=2 filter=23 channel=126
					10, 37, 8, -9, -10, -7, -23, 11, 23,
					-- layer=2 filter=23 channel=127
					-10, 25, 0, 2, -5, -16, 4, 39, 16,
					-- layer=2 filter=24 channel=0
					-19, -8, -29, -16, 0, 11, 0, 22, 0,
					-- layer=2 filter=24 channel=1
					-9, -30, -11, 18, -66, -41, 2, -25, -31,
					-- layer=2 filter=24 channel=2
					-11, 8, -1, -1, 9, 0, -9, -1, -7,
					-- layer=2 filter=24 channel=3
					10, 16, 3, 26, 7, 24, 10, 17, 28,
					-- layer=2 filter=24 channel=4
					-21, -14, -20, -11, 8, -6, -1, 3, -13,
					-- layer=2 filter=24 channel=5
					-14, -17, 1, -18, 19, 28, -3, -2, 21,
					-- layer=2 filter=24 channel=6
					0, 28, -8, -1, -5, -12, -17, -20, 27,
					-- layer=2 filter=24 channel=7
					-9, 1, -31, -32, -71, -39, -16, -70, -18,
					-- layer=2 filter=24 channel=8
					-2, -6, 6, -9, 5, 7, 7, -4, -2,
					-- layer=2 filter=24 channel=9
					-1, -37, -14, -19, 5, -20, -10, -1, -40,
					-- layer=2 filter=24 channel=10
					-15, 3, -9, 10, 18, 18, 3, 34, 32,
					-- layer=2 filter=24 channel=11
					-10, -4, -4, -8, -5, 2, -8, -2, 12,
					-- layer=2 filter=24 channel=12
					14, -61, -37, -14, -24, -42, 16, 4, 0,
					-- layer=2 filter=24 channel=13
					0, -12, -2, -6, -11, -7, 8, 8, 2,
					-- layer=2 filter=24 channel=14
					-9, -27, 4, 0, -54, -12, -3, -33, -16,
					-- layer=2 filter=24 channel=15
					43, 14, 32, 8, 13, -2, 31, -50, -13,
					-- layer=2 filter=24 channel=16
					-48, -8, -44, -48, -4, -43, -28, -27, -47,
					-- layer=2 filter=24 channel=17
					1, -9, 0, 3, 6, 5, 7, 0, 2,
					-- layer=2 filter=24 channel=18
					0, 9, 18, 33, 11, 11, 17, -14, -52,
					-- layer=2 filter=24 channel=19
					10, 4, -55, 36, -33, -5, -14, -43, -1,
					-- layer=2 filter=24 channel=20
					8, 6, 7, -9, 6, 9, 11, -3, -1,
					-- layer=2 filter=24 channel=21
					-3, 15, 8, 19, 7, -2, 14, 7, 16,
					-- layer=2 filter=24 channel=22
					7, 8, 5, 0, 3, 0, 7, -5, 9,
					-- layer=2 filter=24 channel=23
					-4, 16, -28, 3, 52, -7, 27, 26, 13,
					-- layer=2 filter=24 channel=24
					-20, 0, 11, 5, -9, 19, -7, 3, 25,
					-- layer=2 filter=24 channel=25
					-21, 1, 26, -22, -18, 26, -33, 23, 47,
					-- layer=2 filter=24 channel=26
					2, 10, 5, -4, 6, -4, -1, 9, -3,
					-- layer=2 filter=24 channel=27
					-1, 0, -11, -2, 10, -9, -4, -12, 1,
					-- layer=2 filter=24 channel=28
					-26, 18, -3, -23, -31, -35, 17, 9, -13,
					-- layer=2 filter=24 channel=29
					1, 2, 3, 10, 8, 10, -7, 12, 4,
					-- layer=2 filter=24 channel=30
					-23, -48, 10, 14, -17, -13, 2, 13, -13,
					-- layer=2 filter=24 channel=31
					-65, -2, -19, -7, 22, -12, -10, -22, -7,
					-- layer=2 filter=24 channel=32
					-7, -10, -6, -6, 5, -7, 4, 10, -5,
					-- layer=2 filter=24 channel=33
					30, 23, -16, 9, 12, 21, -12, -16, -13,
					-- layer=2 filter=24 channel=34
					34, 8, 14, 39, 26, 29, 8, 24, -8,
					-- layer=2 filter=24 channel=35
					-13, 17, -21, -16, -28, -45, 32, -5, -27,
					-- layer=2 filter=24 channel=36
					3, -4, 2, -6, -6, -7, 3, -1, 15,
					-- layer=2 filter=24 channel=37
					-3, -9, 3, -4, 10, 0, 3, -13, 3,
					-- layer=2 filter=24 channel=38
					0, -54, 22, 15, -9, 0, -5, -14, 1,
					-- layer=2 filter=24 channel=39
					-43, -3, -36, -11, 47, 40, -19, -4, 31,
					-- layer=2 filter=24 channel=40
					17, -22, 12, 20, 26, 38, 1, 54, -38,
					-- layer=2 filter=24 channel=41
					1, -2, -9, 0, -1, 8, -9, -8, 1,
					-- layer=2 filter=24 channel=42
					1, 14, -7, 3, 7, 14, 36, 1, 31,
					-- layer=2 filter=24 channel=43
					6, 16, -6, 35, 29, -7, 26, 38, 1,
					-- layer=2 filter=24 channel=44
					4, 4, -11, 4, 8, 10, 0, -9, 5,
					-- layer=2 filter=24 channel=45
					-133, -45, -72, -86, -21, -7, -45, -27, -38,
					-- layer=2 filter=24 channel=46
					24, -24, -17, 16, 19, -3, -25, 7, -2,
					-- layer=2 filter=24 channel=47
					-54, -36, -27, -9, -25, -36, 5, 7, -16,
					-- layer=2 filter=24 channel=48
					7, 5, 4, 12, -10, 5, 7, -7, 0,
					-- layer=2 filter=24 channel=49
					-27, 19, 36, 18, -4, -32, -13, -45, -51,
					-- layer=2 filter=24 channel=50
					14, 22, 21, 0, -15, 2, 5, 9, 19,
					-- layer=2 filter=24 channel=51
					-26, 4, 24, -4, 11, 10, -21, 0, 12,
					-- layer=2 filter=24 channel=52
					-16, 14, 42, 7, -19, -17, 11, 21, -26,
					-- layer=2 filter=24 channel=53
					-14, 1, 19, -5, -10, -49, -75, -10, 30,
					-- layer=2 filter=24 channel=54
					-13, 12, -5, 9, 9, 13, 26, 9, 15,
					-- layer=2 filter=24 channel=55
					11, 6, -10, 2, 1, 8, -2, 4, 10,
					-- layer=2 filter=24 channel=56
					-11, -16, -19, -1, -15, 15, -5, -13, 16,
					-- layer=2 filter=24 channel=57
					-11, 6, -8, 6, -5, 6, -3, 7, 3,
					-- layer=2 filter=24 channel=58
					41, -78, -28, 3, -31, -40, 18, 9, 8,
					-- layer=2 filter=24 channel=59
					62, -15, -14, -8, -34, 22, -49, 33, 31,
					-- layer=2 filter=24 channel=60
					44, -32, 32, 13, -4, 25, -56, 3, 13,
					-- layer=2 filter=24 channel=61
					10, 21, 4, -12, -35, 13, -1, -18, -11,
					-- layer=2 filter=24 channel=62
					-4, 20, 2, 21, 27, -15, 0, -32, -3,
					-- layer=2 filter=24 channel=63
					-7, -19, -52, 14, 2, -1, 0, 22, -1,
					-- layer=2 filter=24 channel=64
					-9, -24, 6, 22, 24, -2, 46, 16, -1,
					-- layer=2 filter=24 channel=65
					14, 0, 8, 3, -26, 12, 23, 1, 10,
					-- layer=2 filter=24 channel=66
					19, 3, 43, 30, 36, 3, 16, 28, 10,
					-- layer=2 filter=24 channel=67
					24, 11, -5, -22, 23, 8, -26, 20, -9,
					-- layer=2 filter=24 channel=68
					-7, 2, -9, -1, 1, -7, 0, 0, 2,
					-- layer=2 filter=24 channel=69
					-28, -11, -13, 30, 9, 14, 26, 14, 11,
					-- layer=2 filter=24 channel=70
					-1, 12, 9, -10, 7, -24, 17, 10, 8,
					-- layer=2 filter=24 channel=71
					-9, 28, 31, -33, -7, 30, -9, -2, 20,
					-- layer=2 filter=24 channel=72
					-40, 3, -10, -8, -20, 21, -18, -26, -16,
					-- layer=2 filter=24 channel=73
					-41, 39, 47, 46, 38, 39, 16, 42, 51,
					-- layer=2 filter=24 channel=74
					-9, -11, -35, -9, 12, 0, -21, 28, 14,
					-- layer=2 filter=24 channel=75
					-44, -38, -4, -5, -29, 11, -41, -45, -10,
					-- layer=2 filter=24 channel=76
					-11, -23, 6, 13, 51, -4, 7, 12, 42,
					-- layer=2 filter=24 channel=77
					2, -3, -7, 2, 0, -1, 0, -7, -7,
					-- layer=2 filter=24 channel=78
					-12, 19, 10, 23, -28, 0, 2, -7, -7,
					-- layer=2 filter=24 channel=79
					-4, 10, 3, -1, -8, -3, 10, 11, 8,
					-- layer=2 filter=24 channel=80
					13, 3, -17, -9, 17, 0, 25, -14, -24,
					-- layer=2 filter=24 channel=81
					9, 4, 8, 0, -2, -1, 3, 8, 9,
					-- layer=2 filter=24 channel=82
					0, -8, -6, -1, -7, 2, -3, -2, 2,
					-- layer=2 filter=24 channel=83
					-8, -34, 18, -22, 12, -19, 22, -43, -26,
					-- layer=2 filter=24 channel=84
					-8, -11, 3, -4, -4, -3, 2, -6, -3,
					-- layer=2 filter=24 channel=85
					8, 9, -5, 6, -5, 0, -2, -6, 0,
					-- layer=2 filter=24 channel=86
					-10, 13, 11, -8, -10, 4, 7, -14, 10,
					-- layer=2 filter=24 channel=87
					36, 55, 18, 50, 40, 15, -1, 23, -8,
					-- layer=2 filter=24 channel=88
					-6, -12, -6, -3, -3, -1, -18, 25, 11,
					-- layer=2 filter=24 channel=89
					35, -24, -12, -13, -43, -36, -30, -3, 22,
					-- layer=2 filter=24 channel=90
					-1, 5, 8, -4, 4, 7, -5, 6, -4,
					-- layer=2 filter=24 channel=91
					16, -75, -35, -38, -67, -27, 5, 4, 41,
					-- layer=2 filter=24 channel=92
					12, -48, -47, -2, -39, -54, 3, -19, -28,
					-- layer=2 filter=24 channel=93
					-20, 11, -34, 10, 35, -34, -13, 3, 20,
					-- layer=2 filter=24 channel=94
					24, -6, -6, 20, -4, 0, -1, -52, -23,
					-- layer=2 filter=24 channel=95
					3, -3, -2, -11, -12, 2, -2, -13, 0,
					-- layer=2 filter=24 channel=96
					14, 44, 35, 24, 18, 18, -10, 10, 14,
					-- layer=2 filter=24 channel=97
					6, -28, -15, -2, -41, -8, 28, -5, -49,
					-- layer=2 filter=24 channel=98
					-26, 15, -34, -19, -23, -4, 25, 6, -46,
					-- layer=2 filter=24 channel=99
					21, -1, 18, 17, -20, -6, 10, 17, -2,
					-- layer=2 filter=24 channel=100
					6, -38, 25, 0, 4, 5, 0, 24, 45,
					-- layer=2 filter=24 channel=101
					-1, 23, -18, -13, -1, 10, -60, -6, 18,
					-- layer=2 filter=24 channel=102
					-3, 29, 14, 20, 19, 3, 30, 1, -37,
					-- layer=2 filter=24 channel=103
					-35, 20, 29, 69, 27, -24, 22, 45, -17,
					-- layer=2 filter=24 channel=104
					-13, 20, 14, 25, 14, -12, -13, -25, -23,
					-- layer=2 filter=24 channel=105
					23, 20, -15, -55, 0, -62, -23, -23, 10,
					-- layer=2 filter=24 channel=106
					9, -11, 6, -18, -13, 20, -37, 28, 47,
					-- layer=2 filter=24 channel=107
					-12, -4, 28, 52, 46, 7, 8, -15, 17,
					-- layer=2 filter=24 channel=108
					-31, 23, 13, -20, -19, 0, -29, -26, -48,
					-- layer=2 filter=24 channel=109
					-17, -3, 3, -3, 0, 12, 9, 10, 21,
					-- layer=2 filter=24 channel=110
					-15, -19, 9, -10, -8, 0, -2, -1, 5,
					-- layer=2 filter=24 channel=111
					-10, -5, 7, 8, -6, 8, 2, 10, 5,
					-- layer=2 filter=24 channel=112
					-5, -6, -14, -53, -13, 32, -34, -28, -2,
					-- layer=2 filter=24 channel=113
					11, -57, 22, -28, -12, -17, -8, 9, -29,
					-- layer=2 filter=24 channel=114
					0, 11, -3, 0, -7, -1, 5, 6, 0,
					-- layer=2 filter=24 channel=115
					-5, -1, -7, 4, 6, -2, -1, 3, -7,
					-- layer=2 filter=24 channel=116
					35, 25, 22, 64, 38, 9, 3, 7, 10,
					-- layer=2 filter=24 channel=117
					-25, 35, 7, 0, -67, -48, 40, -15, -22,
					-- layer=2 filter=24 channel=118
					10, 33, -11, 41, 33, 0, 17, 2, -15,
					-- layer=2 filter=24 channel=119
					-38, -30, 3, 13, -2, -35, 12, 6, -36,
					-- layer=2 filter=24 channel=120
					7, 1, -2, -5, -9, -4, 6, 8, -3,
					-- layer=2 filter=24 channel=121
					7, 7, 1, 2, 0, 4, 0, -2, 2,
					-- layer=2 filter=24 channel=122
					-2, 7, -6, -5, 0, 11, -1, 14, -6,
					-- layer=2 filter=24 channel=123
					-6, 3, -20, -12, -7, -4, 26, 16, -10,
					-- layer=2 filter=24 channel=124
					19, 12, -11, -29, 33, -45, 22, 5, 28,
					-- layer=2 filter=24 channel=125
					8, 4, 7, -5, -7, 3, -5, -1, -5,
					-- layer=2 filter=24 channel=126
					-15, 2, 41, 7, 30, 32, -44, 41, 14,
					-- layer=2 filter=24 channel=127
					-25, -32, -13, -18, -8, -11, -38, -27, 0,
					-- layer=2 filter=25 channel=0
					0, 12, 17, -18, -3, -15, -17, 10, -10,
					-- layer=2 filter=25 channel=1
					52, -7, -19, 15, 11, 12, 29, -22, -2,
					-- layer=2 filter=25 channel=2
					3, -11, 4, 3, 8, -3, 5, 3, 0,
					-- layer=2 filter=25 channel=3
					16, -3, 3, -2, 7, -9, -5, 27, 16,
					-- layer=2 filter=25 channel=4
					5, -20, 2, 18, -17, 16, 0, -31, -32,
					-- layer=2 filter=25 channel=5
					1, 13, 10, -20, 18, 3, 0, -1, -18,
					-- layer=2 filter=25 channel=6
					0, 14, 42, -30, -49, 8, -33, -50, -20,
					-- layer=2 filter=25 channel=7
					30, 39, 52, 28, 50, 49, 34, 58, 43,
					-- layer=2 filter=25 channel=8
					4, -7, -9, -4, -7, 5, 7, 2, 0,
					-- layer=2 filter=25 channel=9
					35, 14, 15, -4, -14, 0, 2, 38, 10,
					-- layer=2 filter=25 channel=10
					4, -2, -10, -8, -4, 1, 11, 15, 8,
					-- layer=2 filter=25 channel=11
					-4, 12, 0, -11, -10, -24, -31, -14, -24,
					-- layer=2 filter=25 channel=12
					56, 7, -8, 37, 21, 27, -7, -18, 14,
					-- layer=2 filter=25 channel=13
					-8, -1, 2, -2, 7, -10, 0, -4, 0,
					-- layer=2 filter=25 channel=14
					34, 24, 15, -5, 12, 28, -9, -13, -9,
					-- layer=2 filter=25 channel=15
					-16, -33, -10, -48, -26, -36, 4, -15, -59,
					-- layer=2 filter=25 channel=16
					-13, -31, -42, -47, -38, -14, 8, 25, -4,
					-- layer=2 filter=25 channel=17
					0, 0, 11, 2, -5, -7, 9, 0, 6,
					-- layer=2 filter=25 channel=18
					-34, -78, -29, -10, -29, -25, -18, -43, -44,
					-- layer=2 filter=25 channel=19
					17, 14, -4, -9, -29, -55, 24, 0, -24,
					-- layer=2 filter=25 channel=20
					-7, -10, 5, 4, 1, 6, 8, -5, 2,
					-- layer=2 filter=25 channel=21
					14, 0, 2, 19, 10, 6, -5, -2, 20,
					-- layer=2 filter=25 channel=22
					-8, 0, 0, 0, 11, -4, 0, 0, 0,
					-- layer=2 filter=25 channel=23
					8, -3, 8, 15, -25, -23, 14, 10, -7,
					-- layer=2 filter=25 channel=24
					19, 1, -6, 0, 12, 9, -1, 20, 27,
					-- layer=2 filter=25 channel=25
					-21, -30, -46, -47, -36, -38, -18, -1, -2,
					-- layer=2 filter=25 channel=26
					6, 6, -10, 0, 10, 0, -5, -10, 1,
					-- layer=2 filter=25 channel=27
					-15, -8, -14, 4, -20, 6, 14, 3, 21,
					-- layer=2 filter=25 channel=28
					-18, -8, 26, 17, 29, 23, 25, 3, -5,
					-- layer=2 filter=25 channel=29
					-4, 7, -2, 0, -2, 9, -1, 0, 6,
					-- layer=2 filter=25 channel=30
					0, 8, -13, -1, -17, -20, 1, -32, -21,
					-- layer=2 filter=25 channel=31
					56, 26, 52, 39, 10, 49, -3, 0, -40,
					-- layer=2 filter=25 channel=32
					-7, 7, -4, 8, 8, 6, -8, 7, -1,
					-- layer=2 filter=25 channel=33
					37, 33, 27, -15, 8, 79, 31, 48, 11,
					-- layer=2 filter=25 channel=34
					4, 8, -22, 18, 40, -52, 19, -26, -62,
					-- layer=2 filter=25 channel=35
					2, 42, 20, 9, 24, -12, 34, 8, 19,
					-- layer=2 filter=25 channel=36
					4, 15, 0, 2, 5, 11, -7, -8, -4,
					-- layer=2 filter=25 channel=37
					-7, 6, 2, 2, -18, -7, -21, 5, -14,
					-- layer=2 filter=25 channel=38
					13, 32, 10, 2, 10, 24, 12, -19, -6,
					-- layer=2 filter=25 channel=39
					-5, 7, -13, -6, 7, -4, -5, 0, 18,
					-- layer=2 filter=25 channel=40
					50, -9, -26, 10, -11, 27, 55, 32, 9,
					-- layer=2 filter=25 channel=41
					-9, 7, 0, 5, 5, 2, 10, 0, 7,
					-- layer=2 filter=25 channel=42
					36, 13, 10, 9, -3, -9, 15, 8, 0,
					-- layer=2 filter=25 channel=43
					2, 11, 7, -11, 7, 7, -10, 10, 5,
					-- layer=2 filter=25 channel=44
					5, -10, 8, -12, -3, 4, -9, 0, 0,
					-- layer=2 filter=25 channel=45
					-1, -18, -13, 16, -17, 22, 42, -2, 22,
					-- layer=2 filter=25 channel=46
					0, -24, -12, -15, -22, -23, -28, -36, -14,
					-- layer=2 filter=25 channel=47
					22, -22, 8, 1, 1, 26, 1, 36, 0,
					-- layer=2 filter=25 channel=48
					-3, 0, -7, -6, -1, -8, 2, -9, 4,
					-- layer=2 filter=25 channel=49
					-8, -33, -36, -34, -53, -27, -35, -64, -14,
					-- layer=2 filter=25 channel=50
					19, -5, -3, 4, 0, 19, 10, -7, -6,
					-- layer=2 filter=25 channel=51
					12, 12, 20, -12, -16, -10, -3, -3, -22,
					-- layer=2 filter=25 channel=52
					6, 3, 40, 46, -51, -15, -14, -16, -26,
					-- layer=2 filter=25 channel=53
					-48, -20, -20, -67, -19, -112, 10, -60, -65,
					-- layer=2 filter=25 channel=54
					17, 6, 7, 10, 7, 0, 2, 0, 10,
					-- layer=2 filter=25 channel=55
					0, 0, 13, -2, 7, -9, 0, 0, 0,
					-- layer=2 filter=25 channel=56
					1, 8, 9, 8, -6, 6, -22, -16, -19,
					-- layer=2 filter=25 channel=57
					5, 5, 3, -8, -2, 4, -5, 0, 1,
					-- layer=2 filter=25 channel=58
					46, 34, 20, 17, 28, 26, 9, 17, 21,
					-- layer=2 filter=25 channel=59
					-27, 24, -31, -5, 20, -4, 9, -3, -13,
					-- layer=2 filter=25 channel=60
					-3, -3, -14, -27, 0, -17, -25, -15, -31,
					-- layer=2 filter=25 channel=61
					-84, -7, 8, -48, -64, -37, -90, 1, -20,
					-- layer=2 filter=25 channel=62
					35, 25, 24, 28, -8, -12, 17, -23, -51,
					-- layer=2 filter=25 channel=63
					-2, 0, 0, -11, -17, -8, -29, 6, -18,
					-- layer=2 filter=25 channel=64
					7, 18, 17, 15, 9, 9, 19, 23, 16,
					-- layer=2 filter=25 channel=65
					-52, 13, 4, -14, -21, 4, -66, 10, -19,
					-- layer=2 filter=25 channel=66
					-46, 21, 40, 26, 31, 2, 11, 24, 5,
					-- layer=2 filter=25 channel=67
					4, -19, -14, 4, -26, 4, -17, 17, -18,
					-- layer=2 filter=25 channel=68
					12, -4, 2, 10, -8, 3, 8, 7, 1,
					-- layer=2 filter=25 channel=69
					4, 21, 3, -4, -18, 3, 12, 5, 0,
					-- layer=2 filter=25 channel=70
					-14, 17, 36, 24, 12, 1, 20, 0, 0,
					-- layer=2 filter=25 channel=71
					-15, 8, -7, 25, 22, 28, 11, 17, 28,
					-- layer=2 filter=25 channel=72
					12, 35, 33, 0, -1, 48, 43, 26, 14,
					-- layer=2 filter=25 channel=73
					-2, 1, 2, -12, 12, -1, 17, -18, 66,
					-- layer=2 filter=25 channel=74
					24, -2, -19, 1, -8, 4, -2, 13, 3,
					-- layer=2 filter=25 channel=75
					0, 14, 19, 42, 29, 19, 33, 60, -5,
					-- layer=2 filter=25 channel=76
					-30, 0, -5, 10, -18, -70, -12, -97, -45,
					-- layer=2 filter=25 channel=77
					-8, 3, -5, -5, 5, -8, 6, 9, 0,
					-- layer=2 filter=25 channel=78
					4, -15, -5, 0, -26, -27, 11, -3, -16,
					-- layer=2 filter=25 channel=79
					-6, -2, -4, 5, -2, -7, 0, -9, 10,
					-- layer=2 filter=25 channel=80
					-6, -22, 0, -13, 1, 19, -27, -11, -5,
					-- layer=2 filter=25 channel=81
					15, 4, 14, 10, 2, 0, 13, -5, 0,
					-- layer=2 filter=25 channel=82
					-11, 5, -8, 7, 8, -2, -3, -2, -7,
					-- layer=2 filter=25 channel=83
					-12, -30, -7, -9, -29, -16, 3, -19, 4,
					-- layer=2 filter=25 channel=84
					6, 4, -6, -6, -3, 1, 0, -4, -10,
					-- layer=2 filter=25 channel=85
					9, -7, 8, 7, 4, -3, 4, 1, 14,
					-- layer=2 filter=25 channel=86
					6, -6, -13, 1, -18, -11, 8, -15, -9,
					-- layer=2 filter=25 channel=87
					-1, -7, -8, -2, -41, -64, 6, -40, -83,
					-- layer=2 filter=25 channel=88
					38, 9, -10, 2, -18, 13, 23, -2, 11,
					-- layer=2 filter=25 channel=89
					10, 41, 11, 5, -8, 2, 11, -10, -27,
					-- layer=2 filter=25 channel=90
					-8, -3, -2, -11, 9, 1, 5, 8, 2,
					-- layer=2 filter=25 channel=91
					2, 25, -3, -13, -2, 5, 12, 11, 37,
					-- layer=2 filter=25 channel=92
					35, 29, 0, 13, 4, 12, -2, -20, -4,
					-- layer=2 filter=25 channel=93
					70, 26, 7, 59, 17, 47, 3, 86, 29,
					-- layer=2 filter=25 channel=94
					-53, 12, 11, -44, -69, -38, -13, -6, -47,
					-- layer=2 filter=25 channel=95
					-1, 6, 17, 19, -3, 3, -4, 5, 16,
					-- layer=2 filter=25 channel=96
					9, 1, 12, 17, -19, -76, 9, -41, -89,
					-- layer=2 filter=25 channel=97
					13, 23, 28, -5, -5, 12, -10, 22, 26,
					-- layer=2 filter=25 channel=98
					-13, 3, 18, 13, 9, 25, 5, 27, 4,
					-- layer=2 filter=25 channel=99
					-9, -11, 10, -14, -47, -29, -52, 10, -27,
					-- layer=2 filter=25 channel=100
					-7, -12, -46, -17, 17, -12, 4, 3, -28,
					-- layer=2 filter=25 channel=101
					17, -10, -21, -4, -19, -19, -19, 1, 0,
					-- layer=2 filter=25 channel=102
					11, -25, -47, 7, -22, -77, -20, -42, -68,
					-- layer=2 filter=25 channel=103
					26, -8, -4, -5, -2, 19, -56, -5, 3,
					-- layer=2 filter=25 channel=104
					-72, -39, -4, -24, -78, -48, -42, -114, -67,
					-- layer=2 filter=25 channel=105
					-7, -17, 11, 37, 27, -30, 14, -24, -41,
					-- layer=2 filter=25 channel=106
					2, 0, -15, -24, -15, -8, -25, -2, 0,
					-- layer=2 filter=25 channel=107
					-6, -12, -6, -2, 17, 21, -48, -45, -34,
					-- layer=2 filter=25 channel=108
					54, -2, 0, 10, -8, 11, 1, -12, -31,
					-- layer=2 filter=25 channel=109
					-4, -2, 12, -5, -4, 8, 6, 0, -3,
					-- layer=2 filter=25 channel=110
					-13, -4, 17, -17, 0, 13, 14, -6, 17,
					-- layer=2 filter=25 channel=111
					10, 5, 3, -5, -7, 8, -4, 0, 8,
					-- layer=2 filter=25 channel=112
					-37, 9, -1, -48, -36, -57, -36, 13, -18,
					-- layer=2 filter=25 channel=113
					-43, 11, -13, 1, 9, -4, -14, 0, 0,
					-- layer=2 filter=25 channel=114
					-6, 20, 6, -7, -11, 3, 0, 6, 14,
					-- layer=2 filter=25 channel=115
					1, 2, 8, 5, 2, 2, 0, -4, 6,
					-- layer=2 filter=25 channel=116
					-2, -4, -12, 4, -22, -50, 0, -21, -99,
					-- layer=2 filter=25 channel=117
					23, 15, 0, -6, -12, -9, 30, 3, 29,
					-- layer=2 filter=25 channel=118
					8, 1, 27, 20, 6, 18, 9, -1, 7,
					-- layer=2 filter=25 channel=119
					-7, -11, -13, 9, -21, -5, 12, -24, -30,
					-- layer=2 filter=25 channel=120
					3, 8, 7, -8, -2, 10, -8, 4, -8,
					-- layer=2 filter=25 channel=121
					7, -2, 0, 0, -5, -8, -6, 9, 2,
					-- layer=2 filter=25 channel=122
					12, 12, 8, 8, -10, 3, -9, -1, -13,
					-- layer=2 filter=25 channel=123
					-6, 27, 37, 24, 21, 50, 13, 19, 13,
					-- layer=2 filter=25 channel=124
					0, 13, -9, -9, -8, 17, 14, -47, -59,
					-- layer=2 filter=25 channel=125
					-6, -4, 0, 2, 6, -1, 0, -11, 10,
					-- layer=2 filter=25 channel=126
					-32, -70, 63, 9, -25, 8, -70, 34, 58,
					-- layer=2 filter=25 channel=127
					22, 15, 0, 3, 0, 20, -12, -21, -24,
					-- layer=2 filter=26 channel=0
					13, 12, 16, 24, 10, 21, 18, 11, 5,
					-- layer=2 filter=26 channel=1
					2, -9, 2, -11, -48, -39, -23, -19, 7,
					-- layer=2 filter=26 channel=2
					-5, 8, 0, 3, 9, -2, -3, 1, 10,
					-- layer=2 filter=26 channel=3
					10, 32, -14, 9, 16, 13, 51, 27, 38,
					-- layer=2 filter=26 channel=4
					-37, -35, -26, -13, -25, 3, -14, -14, 27,
					-- layer=2 filter=26 channel=5
					-10, -1, 21, 20, 16, -17, 14, 3, -6,
					-- layer=2 filter=26 channel=6
					61, 65, -25, 28, -34, -17, -58, -14, -67,
					-- layer=2 filter=26 channel=7
					-94, -28, 20, -45, 7, 13, -34, -36, 24,
					-- layer=2 filter=26 channel=8
					-6, 6, -7, 5, 5, 6, 0, -5, 5,
					-- layer=2 filter=26 channel=9
					-11, 6, -13, -1, 50, 2, 13, 25, 44,
					-- layer=2 filter=26 channel=10
					1, 4, 10, -2, 12, 24, 27, 1, 47,
					-- layer=2 filter=26 channel=11
					19, 12, 0, 25, 7, -14, 0, 22, 1,
					-- layer=2 filter=26 channel=12
					23, -3, 1, -31, -64, -31, -66, -29, -20,
					-- layer=2 filter=26 channel=13
					2, -2, 5, -3, -3, 2, -6, -1, 8,
					-- layer=2 filter=26 channel=14
					0, 0, -1, -29, -27, -80, -41, -16, -3,
					-- layer=2 filter=26 channel=15
					38, 0, -85, 58, -4, -38, 29, 51, 4,
					-- layer=2 filter=26 channel=16
					-24, -46, -44, -10, -41, -25, 21, 4, -1,
					-- layer=2 filter=26 channel=17
					0, 9, -8, -7, 0, -2, -5, -3, 5,
					-- layer=2 filter=26 channel=18
					-75, -51, -98, -77, -37, -72, -65, -17, -55,
					-- layer=2 filter=26 channel=19
					-20, -3, 0, 11, -45, -59, 38, -2, 8,
					-- layer=2 filter=26 channel=20
					3, -8, -9, 0, 7, 3, -9, -8, -1,
					-- layer=2 filter=26 channel=21
					7, 3, 14, 7, -1, 20, 0, 0, 9,
					-- layer=2 filter=26 channel=22
					9, 7, -7, 7, 6, 0, 0, 8, -8,
					-- layer=2 filter=26 channel=23
					13, 19, 12, 9, -2, 17, 11, -2, 25,
					-- layer=2 filter=26 channel=24
					6, 11, -6, 26, 39, -3, 39, 47, 37,
					-- layer=2 filter=26 channel=25
					-2, 16, -25, 8, 3, -26, 31, 52, 17,
					-- layer=2 filter=26 channel=26
					-5, 8, 1, 0, 6, -7, -3, 4, 9,
					-- layer=2 filter=26 channel=27
					27, 6, 6, 22, 6, 9, 29, 14, 35,
					-- layer=2 filter=26 channel=28
					-1, -5, -1, -23, -21, -21, 36, -51, -65,
					-- layer=2 filter=26 channel=29
					2, 2, 2, 2, 2, -8, 2, -1, -1,
					-- layer=2 filter=26 channel=30
					-27, -6, -16, -16, 19, -6, -26, -18, 18,
					-- layer=2 filter=26 channel=31
					1, 31, 5, 46, 7, -23, 29, -19, -44,
					-- layer=2 filter=26 channel=32
					10, 10, 3, -9, 7, 9, 6, 0, 9,
					-- layer=2 filter=26 channel=33
					-28, 10, -5, -61, -46, -48, 10, -20, 31,
					-- layer=2 filter=26 channel=34
					-60, -66, -2, -37, 6, -7, -32, -56, 9,
					-- layer=2 filter=26 channel=35
					-12, -25, -10, -27, 12, 2, 30, -25, -32,
					-- layer=2 filter=26 channel=36
					-4, 14, -6, 6, 0, -8, -1, 7, -8,
					-- layer=2 filter=26 channel=37
					20, 9, 12, 30, -1, -3, 14, -5, 21,
					-- layer=2 filter=26 channel=38
					14, -18, 14, 1, 3, -5, 13, -13, -5,
					-- layer=2 filter=26 channel=39
					-4, 8, -1, 14, -13, 16, 10, -8, 23,
					-- layer=2 filter=26 channel=40
					-11, -72, -52, -9, -14, -30, 52, 36, 4,
					-- layer=2 filter=26 channel=41
					-1, -3, 4, 2, -10, -1, 2, -3, 3,
					-- layer=2 filter=26 channel=42
					14, 4, -15, -11, -5, 15, 1, 24, 17,
					-- layer=2 filter=26 channel=43
					7, 19, 14, 14, 48, 33, 19, 34, 30,
					-- layer=2 filter=26 channel=44
					2, 0, -10, -4, 8, 7, 0, 7, -8,
					-- layer=2 filter=26 channel=45
					20, -4, 6, 8, -11, 20, 7, 4, 22,
					-- layer=2 filter=26 channel=46
					-16, -23, -17, -23, 15, 19, -11, 18, 28,
					-- layer=2 filter=26 channel=47
					-15, 25, -15, 20, -44, -18, 4, -17, 6,
					-- layer=2 filter=26 channel=48
					-9, 3, -1, -5, 2, -5, -1, 2, 8,
					-- layer=2 filter=26 channel=49
					-18, -29, -78, 7, 0, -58, -46, 34, 4,
					-- layer=2 filter=26 channel=50
					5, 6, -15, 18, -5, -7, 2, -10, -7,
					-- layer=2 filter=26 channel=51
					17, 17, 3, 3, 7, -4, 14, 6, 19,
					-- layer=2 filter=26 channel=52
					5, 9, 44, -28, -26, 0, -20, 4, 7,
					-- layer=2 filter=26 channel=53
					18, -1, -53, -6, -6, -67, -11, 26, 51,
					-- layer=2 filter=26 channel=54
					-36, 15, -16, -23, 7, -51, -8, 13, 39,
					-- layer=2 filter=26 channel=55
					1, -8, 7, -9, 5, 0, 1, 6, -1,
					-- layer=2 filter=26 channel=56
					36, 19, 0, 32, 14, 0, 0, 1, -11,
					-- layer=2 filter=26 channel=57
					0, -8, -8, 6, 3, 1, 9, -2, -16,
					-- layer=2 filter=26 channel=58
					30, 19, -18, -29, -21, -1, -50, -29, -20,
					-- layer=2 filter=26 channel=59
					18, -44, -32, -15, -45, 2, -28, 19, -6,
					-- layer=2 filter=26 channel=60
					0, -54, -17, -2, -55, -18, -10, -11, -47,
					-- layer=2 filter=26 channel=61
					-7, -22, -39, 12, -90, -9, -16, -69, -75,
					-- layer=2 filter=26 channel=62
					-13, 7, -3, -45, -15, 0, -96, -23, 2,
					-- layer=2 filter=26 channel=63
					19, -1, -17, 20, -23, 2, 6, -3, -3,
					-- layer=2 filter=26 channel=64
					4, 13, -6, -14, 8, 16, 0, 21, 22,
					-- layer=2 filter=26 channel=65
					-1, 4, -33, 6, -70, 1, 0, -28, -59,
					-- layer=2 filter=26 channel=66
					-49, -35, -7, -6, -15, -3, -6, 23, 33,
					-- layer=2 filter=26 channel=67
					6, -8, -20, 14, 35, 22, 10, 25, 5,
					-- layer=2 filter=26 channel=68
					1, -6, -11, 7, 3, -7, -2, 6, 5,
					-- layer=2 filter=26 channel=69
					-5, -7, -10, 12, -9, 10, -4, 6, 29,
					-- layer=2 filter=26 channel=70
					3, -10, 2, -7, 2, -18, 39, 0, -15,
					-- layer=2 filter=26 channel=71
					54, 17, 28, 43, 13, 12, 34, 13, 26,
					-- layer=2 filter=26 channel=72
					-19, 37, 19, -50, -51, -23, 27, -20, -18,
					-- layer=2 filter=26 channel=73
					-17, -57, -17, 4, -15, -36, 4, -32, 0,
					-- layer=2 filter=26 channel=74
					0, -12, -8, 6, 8, 4, 24, 11, 10,
					-- layer=2 filter=26 channel=75
					-7, 19, -47, 17, -8, -5, 27, -32, 16,
					-- layer=2 filter=26 channel=76
					-19, -15, -38, -16, -42, -3, -48, 0, 53,
					-- layer=2 filter=26 channel=77
					2, -9, -4, 9, -5, 7, 5, 8, -6,
					-- layer=2 filter=26 channel=78
					-31, 21, -1, 7, -3, -10, -10, 48, -9,
					-- layer=2 filter=26 channel=79
					8, -7, 11, -3, 6, -3, -7, 6, 0,
					-- layer=2 filter=26 channel=80
					-3, 0, -7, -6, 5, 4, 17, -8, 32,
					-- layer=2 filter=26 channel=81
					-3, -8, 3, 9, 3, 1, 7, 7, 8,
					-- layer=2 filter=26 channel=82
					-5, 4, 7, 3, 9, -8, -2, -10, 2,
					-- layer=2 filter=26 channel=83
					-6, -9, -29, -1, -19, -18, 28, 5, 17,
					-- layer=2 filter=26 channel=84
					7, 0, 2, 0, -4, 2, -4, -5, -2,
					-- layer=2 filter=26 channel=85
					-11, -6, -17, 7, 0, 11, 6, 1, 3,
					-- layer=2 filter=26 channel=86
					0, 26, 4, 2, 13, 6, -15, 16, 3,
					-- layer=2 filter=26 channel=87
					-46, -56, -51, -27, -76, -50, -4, 13, -6,
					-- layer=2 filter=26 channel=88
					0, -21, -26, 6, 2, -18, 13, 5, -5,
					-- layer=2 filter=26 channel=89
					0, 21, 11, -38, -39, -16, -28, -3, -22,
					-- layer=2 filter=26 channel=90
					-8, -3, 7, 2, 0, 9, -1, 3, -2,
					-- layer=2 filter=26 channel=91
					13, -3, 15, -13, -15, 7, -11, -16, -26,
					-- layer=2 filter=26 channel=92
					16, -6, 0, -49, -56, -40, -49, -22, -23,
					-- layer=2 filter=26 channel=93
					1, 31, 41, 29, 40, 24, 96, 20, 12,
					-- layer=2 filter=26 channel=94
					34, 38, -20, 48, -59, -22, -41, -45, -7,
					-- layer=2 filter=26 channel=95
					-4, -8, -5, -17, -4, 0, 2, -4, 0,
					-- layer=2 filter=26 channel=96
					10, 9, -46, 48, -53, -39, 20, -6, -22,
					-- layer=2 filter=26 channel=97
					-6, 1, -23, 4, 8, -4, 34, 27, 32,
					-- layer=2 filter=26 channel=98
					-19, 6, -31, 25, -51, -23, 28, -26, -4,
					-- layer=2 filter=26 channel=99
					5, -27, -32, 27, -30, -47, 15, 4, -35,
					-- layer=2 filter=26 channel=100
					-5, -7, 9, -36, 12, 14, 6, 24, 1,
					-- layer=2 filter=26 channel=101
					53, 24, 36, 21, 17, -3, 27, 13, 10,
					-- layer=2 filter=26 channel=102
					-58, -13, -30, -34, 8, -25, -36, -54, 9,
					-- layer=2 filter=26 channel=103
					15, 39, 9, 2, -16, -5, -13, 22, -50,
					-- layer=2 filter=26 channel=104
					-27, -28, -91, 20, -28, -85, -71, -7, -31,
					-- layer=2 filter=26 channel=105
					-37, -35, -13, -49, -4, 7, -12, 55, 70,
					-- layer=2 filter=26 channel=106
					22, 5, -25, 13, -1, -34, 36, 36, 7,
					-- layer=2 filter=26 channel=107
					-6, 51, 11, 9, -39, -2, 0, -34, -51,
					-- layer=2 filter=26 channel=108
					19, 19, -14, 8, -1, -21, 23, -25, -4,
					-- layer=2 filter=26 channel=109
					0, -10, 8, 0, 6, -3, 0, 7, 9,
					-- layer=2 filter=26 channel=110
					-5, -8, 4, -18, 8, 7, 15, 29, -2,
					-- layer=2 filter=26 channel=111
					-11, -7, -6, 0, -7, -7, 2, 10, 4,
					-- layer=2 filter=26 channel=112
					25, -22, -15, 26, -1, 14, 9, -9, -4,
					-- layer=2 filter=26 channel=113
					-22, -6, -26, 16, -10, 30, -6, -3, 35,
					-- layer=2 filter=26 channel=114
					-1, -15, -17, 3, 3, -3, -3, -2, -4,
					-- layer=2 filter=26 channel=115
					-7, 7, -9, 6, 4, 7, -2, -3, -2,
					-- layer=2 filter=26 channel=116
					-33, -52, -83, -45, -60, -55, -59, -4, 6,
					-- layer=2 filter=26 channel=117
					-12, 2, -12, -10, -61, -32, -9, -44, -43,
					-- layer=2 filter=26 channel=118
					8, 14, 15, 20, 33, 17, 22, 13, 17,
					-- layer=2 filter=26 channel=119
					-27, -33, -43, -36, -26, 0, -22, -27, 26,
					-- layer=2 filter=26 channel=120
					10, -9, 6, 0, -6, -7, 9, 8, -9,
					-- layer=2 filter=26 channel=121
					-1, -1, -1, 3, -5, 0, -5, -4, 5,
					-- layer=2 filter=26 channel=122
					-9, 1, 8, -3, 5, 10, -7, 1, 6,
					-- layer=2 filter=26 channel=123
					-69, 6, -3, -19, -64, 0, 0, -2, 37,
					-- layer=2 filter=26 channel=124
					-17, -16, -71, -36, -6, -29, -8, 19, 41,
					-- layer=2 filter=26 channel=125
					-3, -3, -3, 0, 6, -4, -8, 2, 0,
					-- layer=2 filter=26 channel=126
					33, 5, 7, 18, 25, 38, 0, 43, 9,
					-- layer=2 filter=26 channel=127
					1, -20, -8, 1, -30, -17, -9, -15, 16,
					-- layer=2 filter=27 channel=0
					6, -2, 19, -27, -8, 9, 29, -9, -17,
					-- layer=2 filter=27 channel=1
					5, 9, -6, 24, 28, -16, -71, -12, 31,
					-- layer=2 filter=27 channel=2
					-6, -8, 1, -5, 0, -4, 0, 10, 4,
					-- layer=2 filter=27 channel=3
					-6, 22, 30, -8, 8, 4, 13, 21, 6,
					-- layer=2 filter=27 channel=4
					11, 21, 8, -5, -14, 15, -25, -22, 18,
					-- layer=2 filter=27 channel=5
					-8, 20, 26, -40, 6, 17, -18, -25, -16,
					-- layer=2 filter=27 channel=6
					-55, -12, -8, -19, -50, -7, -44, -8, -21,
					-- layer=2 filter=27 channel=7
					-3, 21, 10, -1, -4, 3, 8, 6, -43,
					-- layer=2 filter=27 channel=8
					2, 0, -5, -2, -1, 0, -5, 5, -5,
					-- layer=2 filter=27 channel=9
					-24, -12, 10, -24, 9, 21, -1, 21, 30,
					-- layer=2 filter=27 channel=10
					0, 6, 19, -10, -1, 4, 25, 24, -4,
					-- layer=2 filter=27 channel=11
					3, 11, 0, -14, 11, 19, -26, -28, -37,
					-- layer=2 filter=27 channel=12
					27, 33, 14, 40, 30, 12, -61, 10, 54,
					-- layer=2 filter=27 channel=13
					-9, -4, 5, 7, -9, 9, -7, 1, 1,
					-- layer=2 filter=27 channel=14
					20, 32, 3, 34, 40, -1, -37, 14, 14,
					-- layer=2 filter=27 channel=15
					31, 17, 26, -31, 34, 23, -73, -29, -45,
					-- layer=2 filter=27 channel=16
					-18, -4, -23, -12, -11, -11, -1, -15, 9,
					-- layer=2 filter=27 channel=17
					-1, 0, -2, 4, 2, 5, 0, 1, 9,
					-- layer=2 filter=27 channel=18
					23, 31, -10, 56, 30, 33, -9, 26, 9,
					-- layer=2 filter=27 channel=19
					-8, -34, 0, -21, 26, 1, -53, -61, -27,
					-- layer=2 filter=27 channel=20
					9, -4, -6, 5, 4, 12, -2, 8, 4,
					-- layer=2 filter=27 channel=21
					4, -4, 0, 9, 15, -11, 2, 1, 3,
					-- layer=2 filter=27 channel=22
					-2, 6, 7, -7, 4, 1, -6, 0, -1,
					-- layer=2 filter=27 channel=23
					-17, -11, -4, -30, -5, 30, 8, -7, 28,
					-- layer=2 filter=27 channel=24
					-28, 1, -12, 4, 26, 12, 35, -4, 6,
					-- layer=2 filter=27 channel=25
					-55, -6, -14, -33, -13, -25, -50, -39, -37,
					-- layer=2 filter=27 channel=26
					-3, -1, 3, 2, 0, 5, 0, -3, 2,
					-- layer=2 filter=27 channel=27
					-20, 16, 29, -45, 15, 17, -28, -7, -11,
					-- layer=2 filter=27 channel=28
					4, 14, 12, 17, -8, -15, -31, 1, -11,
					-- layer=2 filter=27 channel=29
					2, 0, 10, -1, -1, 7, 6, 9, 3,
					-- layer=2 filter=27 channel=30
					-25, 15, -2, -12, -1, 0, -12, -9, 34,
					-- layer=2 filter=27 channel=31
					-21, -27, 5, -40, -9, 57, -17, -66, -9,
					-- layer=2 filter=27 channel=32
					7, 0, -3, -4, 2, -3, -8, -3, -7,
					-- layer=2 filter=27 channel=33
					40, 61, 23, -17, -9, 4, -49, -7, -49,
					-- layer=2 filter=27 channel=34
					-3, 27, 12, -20, -37, 31, -18, -53, 21,
					-- layer=2 filter=27 channel=35
					30, 36, 21, 4, 2, 30, -34, 13, -8,
					-- layer=2 filter=27 channel=36
					3, 14, 11, 12, -2, 0, 12, -5, 10,
					-- layer=2 filter=27 channel=37
					-13, 7, 4, -6, 19, 9, -22, -16, -2,
					-- layer=2 filter=27 channel=38
					13, 16, 9, -23, 15, 31, -28, -40, -6,
					-- layer=2 filter=27 channel=39
					-36, -11, -15, 3, -13, 7, 19, -2, -2,
					-- layer=2 filter=27 channel=40
					40, 8, -36, 9, 19, 51, -30, 1, -61,
					-- layer=2 filter=27 channel=41
					4, -6, -6, 3, 0, 2, 7, -4, -10,
					-- layer=2 filter=27 channel=42
					6, -9, 9, -21, 10, 26, -16, -7, 49,
					-- layer=2 filter=27 channel=43
					-22, 65, 40, -45, 42, 68, -23, -25, -10,
					-- layer=2 filter=27 channel=44
					10, -4, 5, -1, 4, 0, 10, -4, 8,
					-- layer=2 filter=27 channel=45
					1, 12, 15, 3, 12, 33, -42, -4, -23,
					-- layer=2 filter=27 channel=46
					0, -19, 4, -50, -6, 27, -23, -33, 0,
					-- layer=2 filter=27 channel=47
					-8, 13, 0, 19, -14, 20, 14, -4, -57,
					-- layer=2 filter=27 channel=48
					2, 7, 0, 2, 2, -7, -7, -9, 9,
					-- layer=2 filter=27 channel=49
					4, -30, 11, 27, 16, 48, -3, 56, 28,
					-- layer=2 filter=27 channel=50
					25, -5, 16, -13, 2, 15, 13, 3, 2,
					-- layer=2 filter=27 channel=51
					2, 2, 7, -9, 6, 8, 3, -9, -28,
					-- layer=2 filter=27 channel=52
					-10, -6, -10, 19, -21, 11, -33, -48, -51,
					-- layer=2 filter=27 channel=53
					0, -59, -7, 2, 36, 2, -7, -23, -44,
					-- layer=2 filter=27 channel=54
					-20, -5, 0, -22, -31, -24, -37, -4, -27,
					-- layer=2 filter=27 channel=55
					9, -5, 6, -9, 13, -5, 12, 3, 12,
					-- layer=2 filter=27 channel=56
					-15, 7, 3, -19, 8, 8, -10, -5, -2,
					-- layer=2 filter=27 channel=57
					10, 13, -8, 1, 9, 2, 2, 2, -2,
					-- layer=2 filter=27 channel=58
					30, 16, 0, 25, 22, 11, -75, -29, 33,
					-- layer=2 filter=27 channel=59
					56, 20, 24, 10, 5, 1, -27, -59, -1,
					-- layer=2 filter=27 channel=60
					39, -9, -6, 46, -2, 0, 51, -12, 26,
					-- layer=2 filter=27 channel=61
					-3, -42, -41, 37, 5, -41, 86, 17, 4,
					-- layer=2 filter=27 channel=62
					25, -4, 9, -2, -22, 27, -49, -12, -24,
					-- layer=2 filter=27 channel=63
					14, -9, -2, -1, -4, -11, 10, -18, -13,
					-- layer=2 filter=27 channel=64
					-41, -42, -27, -1, -8, 2, 12, 21, 37,
					-- layer=2 filter=27 channel=65
					-23, -6, -31, 11, -60, -49, 20, -54, -25,
					-- layer=2 filter=27 channel=66
					-10, -1, -7, 11, -27, 15, 13, 7, 51,
					-- layer=2 filter=27 channel=67
					-17, -13, -18, -45, 1, 1, -6, -8, 0,
					-- layer=2 filter=27 channel=68
					-3, 1, -4, -1, 11, 5, -9, 3, 1,
					-- layer=2 filter=27 channel=69
					-43, -52, -4, -6, 3, 4, 11, 5, 30,
					-- layer=2 filter=27 channel=70
					0, 23, 17, -14, -13, 0, -21, -22, -11,
					-- layer=2 filter=27 channel=71
					-6, -5, 5, -79, 3, 17, -54, 2, 4,
					-- layer=2 filter=27 channel=72
					47, 54, 10, 18, 8, 21, 28, 57, 3,
					-- layer=2 filter=27 channel=73
					8, 29, 27, 11, 62, 41, -7, -17, 5,
					-- layer=2 filter=27 channel=74
					18, -16, 2, -16, -1, 14, -46, -19, -10,
					-- layer=2 filter=27 channel=75
					-9, 14, -12, -12, 18, -38, -2, 2, 20,
					-- layer=2 filter=27 channel=76
					15, -56, 45, -22, 96, 41, 13, -15, -14,
					-- layer=2 filter=27 channel=77
					-6, -3, 5, -3, -3, 8, -1, -9, -9,
					-- layer=2 filter=27 channel=78
					0, -2, 11, -4, 1, 20, -37, -26, -20,
					-- layer=2 filter=27 channel=79
					6, 3, 0, 3, 0, -5, -6, -6, 4,
					-- layer=2 filter=27 channel=80
					5, -1, -1, -13, -12, 19, 4, -8, 24,
					-- layer=2 filter=27 channel=81
					0, 7, 0, 8, 16, 20, 8, 13, 3,
					-- layer=2 filter=27 channel=82
					-5, 0, 0, -6, 11, 5, -4, 4, 9,
					-- layer=2 filter=27 channel=83
					9, 0, 0, -22, 7, 5, -28, -34, 6,
					-- layer=2 filter=27 channel=84
					0, 1, -3, -6, 7, -6, 6, 12, 9,
					-- layer=2 filter=27 channel=85
					-10, -7, -3, 4, -8, 5, -5, 0, 8,
					-- layer=2 filter=27 channel=86
					1, 0, -1, 3, -3, 11, 6, 1, 12,
					-- layer=2 filter=27 channel=87
					21, -14, 19, -22, -18, 48, -16, 7, -23,
					-- layer=2 filter=27 channel=88
					-1, 18, 1, 2, 13, -14, -13, -14, 6,
					-- layer=2 filter=27 channel=89
					17, 27, 12, 24, 12, -11, -50, -16, 18,
					-- layer=2 filter=27 channel=90
					6, -4, -2, 2, 6, 2, 1, -6, 4,
					-- layer=2 filter=27 channel=91
					21, 4, 19, 4, -6, 14, -13, -7, 52,
					-- layer=2 filter=27 channel=92
					24, 4, 10, 14, 27, 5, -29, 4, 44,
					-- layer=2 filter=27 channel=93
					-45, 8, -51, -50, -48, -19, -39, -24, -8,
					-- layer=2 filter=27 channel=94
					-20, -82, -69, 0, -25, -60, 33, -34, 5,
					-- layer=2 filter=27 channel=95
					7, 16, 15, 9, 3, 1, -2, 10, 0,
					-- layer=2 filter=27 channel=96
					-33, -63, 13, 11, -98, -26, 16, -3, 35,
					-- layer=2 filter=27 channel=97
					-29, 3, 24, 0, 58, 43, -26, -18, -16,
					-- layer=2 filter=27 channel=98
					28, 19, 10, 26, 5, 30, 10, -1, -30,
					-- layer=2 filter=27 channel=99
					-55, -60, 6, 37, -20, -43, -1, -51, -44,
					-- layer=2 filter=27 channel=100
					9, 30, 12, -4, 34, 4, -41, -33, 0,
					-- layer=2 filter=27 channel=101
					0, 29, -11, -43, 19, 10, -61, 0, -4,
					-- layer=2 filter=27 channel=102
					-67, -68, 9, 6, -69, 2, -21, 18, 12,
					-- layer=2 filter=27 channel=103
					15, -4, 19, -12, -6, -10, -20, 23, 19,
					-- layer=2 filter=27 channel=104
					6, -59, 2, 16, -11, -9, 2, 38, 0,
					-- layer=2 filter=27 channel=105
					0, 16, -56, -31, 52, 73, -19, -2, -39,
					-- layer=2 filter=27 channel=106
					-26, 19, 35, -39, -7, 29, -45, -61, -4,
					-- layer=2 filter=27 channel=107
					-18, 5, 13, 35, -77, 0, -1, -11, 8,
					-- layer=2 filter=27 channel=108
					-25, -20, 8, -22, -17, -26, -85, -29, -46,
					-- layer=2 filter=27 channel=109
					-14, 9, 13, -9, 1, -2, 18, 6, 0,
					-- layer=2 filter=27 channel=110
					-12, -27, -46, 3, 16, -20, 42, 12, -4,
					-- layer=2 filter=27 channel=111
					6, -5, 0, -3, -8, 6, 5, -8, 3,
					-- layer=2 filter=27 channel=112
					-10, -32, -5, 8, -46, -27, 25, -11, -38,
					-- layer=2 filter=27 channel=113
					0, -3, -1, 10, -6, 21, -14, -17, -4,
					-- layer=2 filter=27 channel=114
					-1, 19, 5, 6, 13, -9, -3, -11, -10,
					-- layer=2 filter=27 channel=115
					4, -7, 4, -3, -1, 9, 12, -3, 0,
					-- layer=2 filter=27 channel=116
					24, -4, 17, -8, -27, 42, -10, 3, -12,
					-- layer=2 filter=27 channel=117
					-19, -3, -18, 18, 38, 13, -3, 29, -13,
					-- layer=2 filter=27 channel=118
					0, 2, 35, -8, 8, 46, 20, 23, 28,
					-- layer=2 filter=27 channel=119
					-4, 27, 19, -20, 13, 8, -61, -18, 14,
					-- layer=2 filter=27 channel=120
					2, 4, 5, -3, 0, -8, -6, 3, 2,
					-- layer=2 filter=27 channel=121
					2, -7, 5, 3, -4, 5, 4, 4, 0,
					-- layer=2 filter=27 channel=122
					-4, -17, -1, -1, 11, 3, 3, 0, -12,
					-- layer=2 filter=27 channel=123
					-1, 0, -6, 20, 21, -2, 16, 6, -43,
					-- layer=2 filter=27 channel=124
					-1, -36, 10, -56, -16, 22, -51, -23, -46,
					-- layer=2 filter=27 channel=125
					9, 12, -8, 4, 5, 0, 6, -8, 2,
					-- layer=2 filter=27 channel=126
					-23, -83, 3, -25, -21, -12, -19, -28, 20,
					-- layer=2 filter=27 channel=127
					-16, 34, -6, 3, -27, 9, -15, -45, 1,
					-- layer=2 filter=28 channel=0
					-10, -12, 6, -2, 0, 4, -6, -6, -11,
					-- layer=2 filter=28 channel=1
					7, 2, -5, -7, -3, 0, 0, 1, -1,
					-- layer=2 filter=28 channel=2
					1, 3, -12, -7, 4, -11, -3, -7, -4,
					-- layer=2 filter=28 channel=3
					1, 1, 0, 2, 8, 3, -11, 5, -3,
					-- layer=2 filter=28 channel=4
					-3, -5, -1, -20, -16, -7, -7, 0, -8,
					-- layer=2 filter=28 channel=5
					-10, -3, -2, -6, -6, -6, 1, 0, -5,
					-- layer=2 filter=28 channel=6
					4, -1, 5, -1, -4, 4, -12, 3, -3,
					-- layer=2 filter=28 channel=7
					-5, 4, -6, 8, 7, -3, -19, -7, -4,
					-- layer=2 filter=28 channel=8
					7, -3, 8, -3, -6, 3, 7, -11, 2,
					-- layer=2 filter=28 channel=9
					5, 5, -10, -7, 7, -8, -5, -7, -2,
					-- layer=2 filter=28 channel=10
					-2, -6, -8, -14, -12, 3, -11, -8, -16,
					-- layer=2 filter=28 channel=11
					-8, -16, -13, 0, -10, -17, 0, 3, -15,
					-- layer=2 filter=28 channel=12
					14, 8, -2, 13, 12, -11, -1, -1, -1,
					-- layer=2 filter=28 channel=13
					6, 4, -10, 8, 3, -6, -3, 1, -4,
					-- layer=2 filter=28 channel=14
					-11, -11, -5, -5, 4, 1, -9, -11, 0,
					-- layer=2 filter=28 channel=15
					0, -7, 1, -3, -3, 0, 9, -6, 7,
					-- layer=2 filter=28 channel=16
					-6, 0, 2, 6, -11, 0, -1, -1, -2,
					-- layer=2 filter=28 channel=17
					-8, 0, -6, -1, -3, 2, 5, -6, 6,
					-- layer=2 filter=28 channel=18
					-2, -6, 2, -18, 1, -2, -4, -1, -5,
					-- layer=2 filter=28 channel=19
					-8, -6, -11, -11, 0, 0, -2, -3, -18,
					-- layer=2 filter=28 channel=20
					-4, 2, 7, -2, -11, -7, -9, 5, -8,
					-- layer=2 filter=28 channel=21
					3, -7, 2, 0, 5, 0, -7, -5, -2,
					-- layer=2 filter=28 channel=22
					9, -9, -3, 1, 6, -5, 5, 8, -1,
					-- layer=2 filter=28 channel=23
					0, -2, -9, 4, 1, -14, 0, -9, -7,
					-- layer=2 filter=28 channel=24
					-11, 0, 4, -4, 2, -5, -8, -7, 1,
					-- layer=2 filter=28 channel=25
					-1, -5, -5, 0, 10, 4, 0, 5, -1,
					-- layer=2 filter=28 channel=26
					-10, 7, 6, 2, -4, 4, -5, 9, -6,
					-- layer=2 filter=28 channel=27
					-14, -13, -16, -2, -7, -5, -12, 1, -3,
					-- layer=2 filter=28 channel=28
					-1, 1, 3, 2, 15, -4, 0, -15, -5,
					-- layer=2 filter=28 channel=29
					7, -6, 3, -1, 4, 8, 5, -8, -10,
					-- layer=2 filter=28 channel=30
					-14, -10, 0, -11, 5, -2, 3, -6, 0,
					-- layer=2 filter=28 channel=31
					4, -1, -10, -1, -6, -9, -1, 8, 2,
					-- layer=2 filter=28 channel=32
					9, -3, 0, -9, -10, 9, -3, 7, 1,
					-- layer=2 filter=28 channel=33
					-3, -1, 8, 0, 0, -4, -6, -6, 6,
					-- layer=2 filter=28 channel=34
					11, -7, -2, 1, 3, -11, 4, -10, 7,
					-- layer=2 filter=28 channel=35
					0, -8, 1, -20, 6, -1, 5, 0, 8,
					-- layer=2 filter=28 channel=36
					-12, -8, 2, -7, -2, -10, 2, 1, -10,
					-- layer=2 filter=28 channel=37
					-13, -2, -12, -10, -17, -15, -14, -6, 0,
					-- layer=2 filter=28 channel=38
					0, -4, -7, -8, -1, -17, -14, 0, -3,
					-- layer=2 filter=28 channel=39
					-10, 6, 0, -10, 3, 0, -6, 6, 1,
					-- layer=2 filter=28 channel=40
					-8, -2, 4, -3, -11, -7, -1, -12, 7,
					-- layer=2 filter=28 channel=41
					7, -6, -12, 7, 3, -6, -10, 5, -2,
					-- layer=2 filter=28 channel=42
					14, -12, -12, -4, 0, -3, -8, -9, -9,
					-- layer=2 filter=28 channel=43
					3, -3, 8, -1, 5, -10, -2, 5, 7,
					-- layer=2 filter=28 channel=44
					6, 7, 1, 7, 9, 1, 0, 5, 8,
					-- layer=2 filter=28 channel=45
					-2, 0, 6, -2, 9, 0, -5, -4, -5,
					-- layer=2 filter=28 channel=46
					1, -8, -6, -6, -6, -1, -8, 3, 0,
					-- layer=2 filter=28 channel=47
					-14, -7, -7, -4, 0, -11, -2, -4, -5,
					-- layer=2 filter=28 channel=48
					7, -9, -2, 9, -3, -4, 3, 8, -2,
					-- layer=2 filter=28 channel=49
					-13, -2, -5, -3, 4, 5, 0, 1, 12,
					-- layer=2 filter=28 channel=50
					-8, 3, -10, -3, 0, 4, 2, 3, -4,
					-- layer=2 filter=28 channel=51
					-12, -13, 3, -15, -13, -12, -8, -11, -17,
					-- layer=2 filter=28 channel=52
					-9, -4, -3, -13, 2, -15, -14, -17, -13,
					-- layer=2 filter=28 channel=53
					5, -13, 2, 2, -7, -7, -4, -5, 5,
					-- layer=2 filter=28 channel=54
					10, -18, -22, -3, -5, -4, -12, -14, -2,
					-- layer=2 filter=28 channel=55
					-2, -10, -6, -4, 0, -5, -3, -6, 9,
					-- layer=2 filter=28 channel=56
					-15, -4, 7, -12, -13, -3, -10, -10, -8,
					-- layer=2 filter=28 channel=57
					-4, 6, 10, -5, -2, 6, -7, -8, 10,
					-- layer=2 filter=28 channel=58
					5, 0, -16, -3, -7, 5, -15, -11, -15,
					-- layer=2 filter=28 channel=59
					-15, -2, -9, -13, -10, 0, -14, 0, -4,
					-- layer=2 filter=28 channel=60
					-9, -11, 2, -8, 8, -5, -5, -3, -6,
					-- layer=2 filter=28 channel=61
					-10, 0, -5, 2, -6, -11, -14, -7, -2,
					-- layer=2 filter=28 channel=62
					5, 0, -4, 6, 3, 3, 4, 2, -2,
					-- layer=2 filter=28 channel=63
					8, 3, -11, -5, 0, -6, 5, -11, -5,
					-- layer=2 filter=28 channel=64
					-6, 4, -4, -1, -1, 4, 6, 5, 4,
					-- layer=2 filter=28 channel=65
					-2, -12, -12, 9, -4, -11, -4, 7, 1,
					-- layer=2 filter=28 channel=66
					1, 0, -4, -7, -6, 1, -5, -9, -7,
					-- layer=2 filter=28 channel=67
					0, -6, -1, 3, -8, -4, -4, -7, -2,
					-- layer=2 filter=28 channel=68
					-7, 6, -10, 3, -4, -10, -8, 0, 0,
					-- layer=2 filter=28 channel=69
					5, -2, -7, -9, -12, 2, -3, 0, -11,
					-- layer=2 filter=28 channel=70
					-1, -2, -5, -16, 0, -11, -12, -16, -15,
					-- layer=2 filter=28 channel=71
					-16, -11, -1, -2, -7, -5, -13, 3, 2,
					-- layer=2 filter=28 channel=72
					3, -4, -13, 2, 6, 6, -19, 0, -8,
					-- layer=2 filter=28 channel=73
					-7, 5, 11, 2, 18, 13, 5, 7, 14,
					-- layer=2 filter=28 channel=74
					-6, 4, 0, -12, 3, -7, 6, 2, 7,
					-- layer=2 filter=28 channel=75
					-1, -11, 3, -13, -1, -15, 10, -6, -2,
					-- layer=2 filter=28 channel=76
					-12, 1, 2, 5, -8, -3, 4, -8, 1,
					-- layer=2 filter=28 channel=77
					-6, -1, 6, 0, 8, -10, 0, 5, 0,
					-- layer=2 filter=28 channel=78
					-7, -9, 5, 3, -13, -1, -4, -12, 0,
					-- layer=2 filter=28 channel=79
					0, 6, 2, -11, -9, 4, 5, -3, 5,
					-- layer=2 filter=28 channel=80
					-2, 4, 1, 2, 3, -5, -6, 7, -4,
					-- layer=2 filter=28 channel=81
					6, -5, 6, -11, 8, 4, 8, -4, -9,
					-- layer=2 filter=28 channel=82
					-10, 0, 0, -2, 5, -5, 3, -2, 0,
					-- layer=2 filter=28 channel=83
					-3, 4, -2, -2, 3, 1, 2, -13, -5,
					-- layer=2 filter=28 channel=84
					-8, 1, 2, -8, 8, -12, 4, 0, 1,
					-- layer=2 filter=28 channel=85
					3, 10, -2, 2, -1, 2, 0, 0, 9,
					-- layer=2 filter=28 channel=86
					-8, 8, 0, -4, -1, 1, -2, -1, -5,
					-- layer=2 filter=28 channel=87
					-3, -9, -5, -5, -17, -3, -7, -11, -1,
					-- layer=2 filter=28 channel=88
					-13, -1, -10, -5, 1, -19, -9, -10, 0,
					-- layer=2 filter=28 channel=89
					9, 6, -11, 5, 1, -9, -1, -15, -18,
					-- layer=2 filter=28 channel=90
					9, 6, -7, -1, 0, -4, -2, 6, -8,
					-- layer=2 filter=28 channel=91
					4, -6, -7, -1, -2, -11, -2, 0, 5,
					-- layer=2 filter=28 channel=92
					14, -2, 6, 0, 4, -3, 0, -12, -7,
					-- layer=2 filter=28 channel=93
					9, -1, 2, 18, -5, -3, 2, -10, 8,
					-- layer=2 filter=28 channel=94
					13, -5, 2, 2, -3, -9, -10, 3, 6,
					-- layer=2 filter=28 channel=95
					-6, 5, 0, -11, -2, -4, -6, 1, 3,
					-- layer=2 filter=28 channel=96
					-17, -19, -9, -19, 0, -10, -1, 3, -1,
					-- layer=2 filter=28 channel=97
					-12, -11, -9, -7, 3, 4, -6, 0, -1,
					-- layer=2 filter=28 channel=98
					-12, -5, -12, 12, 13, 0, -3, -11, -13,
					-- layer=2 filter=28 channel=99
					-2, -6, -13, -13, -5, -1, -9, -9, -7,
					-- layer=2 filter=28 channel=100
					-8, 0, -3, -13, 0, -3, -1, -12, 0,
					-- layer=2 filter=28 channel=101
					0, -3, -6, -9, 0, 0, 0, 1, -7,
					-- layer=2 filter=28 channel=102
					-11, -7, 0, -13, 0, 10, -19, -14, 3,
					-- layer=2 filter=28 channel=103
					-10, 1, 2, -6, 5, 7, 0, 7, -11,
					-- layer=2 filter=28 channel=104
					-15, -2, -5, 0, -9, 3, -3, -8, 2,
					-- layer=2 filter=28 channel=105
					-5, -9, 0, -1, -4, 8, 0, -6, 6,
					-- layer=2 filter=28 channel=106
					-13, -6, -9, -4, 2, 5, -6, -8, -4,
					-- layer=2 filter=28 channel=107
					-3, 10, 6, -6, 1, 4, 0, -4, -8,
					-- layer=2 filter=28 channel=108
					-16, -13, -1, -8, -8, 2, -5, -13, -7,
					-- layer=2 filter=28 channel=109
					-2, -6, 0, 0, -4, 4, 7, -4, 0,
					-- layer=2 filter=28 channel=110
					-9, 2, -9, -10, -11, -14, -1, -13, -8,
					-- layer=2 filter=28 channel=111
					-5, -3, 4, 0, 5, -6, -4, -4, 0,
					-- layer=2 filter=28 channel=112
					0, 6, -2, 0, 6, 4, 0, 10, -8,
					-- layer=2 filter=28 channel=113
					-4, 0, -4, -9, -8, -10, 0, -10, -13,
					-- layer=2 filter=28 channel=114
					3, 0, 3, 8, 2, 5, -6, -7, 0,
					-- layer=2 filter=28 channel=115
					-2, 1, -2, 0, -3, -7, 10, -4, -3,
					-- layer=2 filter=28 channel=116
					-6, 2, -9, -6, -6, 2, 1, -8, 15,
					-- layer=2 filter=28 channel=117
					-12, 0, -4, 5, 23, 0, 5, -17, -15,
					-- layer=2 filter=28 channel=118
					-11, 2, 1, 2, 0, -5, -3, 3, -4,
					-- layer=2 filter=28 channel=119
					1, 1, -9, -1, -6, -8, 2, -5, 2,
					-- layer=2 filter=28 channel=120
					7, 8, -3, 4, -3, -1, 1, 5, 6,
					-- layer=2 filter=28 channel=121
					-1, 10, -4, 4, -11, -3, 7, -10, 8,
					-- layer=2 filter=28 channel=122
					-6, 8, 6, 1, 5, 6, 3, 0, 4,
					-- layer=2 filter=28 channel=123
					-13, -14, -5, -2, 16, -4, -5, -19, -16,
					-- layer=2 filter=28 channel=124
					0, -10, 2, 4, -8, 5, -3, -3, 7,
					-- layer=2 filter=28 channel=125
					9, -9, 3, -5, 11, 6, 3, -11, 5,
					-- layer=2 filter=28 channel=126
					2, -7, -1, 3, -3, 0, 2, -5, 0,
					-- layer=2 filter=28 channel=127
					9, 2, -5, -6, 1, -9, -10, -12, 0,
					-- layer=2 filter=29 channel=0
					0, -22, -15, 17, -2, -11, -2, 22, 7,
					-- layer=2 filter=29 channel=1
					-4, 15, -5, -17, -7, 9, -14, 0, 4,
					-- layer=2 filter=29 channel=2
					6, 0, 3, -3, -9, 2, 4, -4, 4,
					-- layer=2 filter=29 channel=3
					-14, -12, 37, 0, -25, 3, -11, 0, 28,
					-- layer=2 filter=29 channel=4
					-26, -14, -9, 0, -26, 7, 18, -9, 19,
					-- layer=2 filter=29 channel=5
					19, 4, -17, -8, -10, -21, 33, -15, -3,
					-- layer=2 filter=29 channel=6
					31, -25, -32, 10, -6, -30, 15, 0, -7,
					-- layer=2 filter=29 channel=7
					-21, -78, -66, -36, -52, -31, -23, -43, 4,
					-- layer=2 filter=29 channel=8
					7, -2, -6, 5, -5, -6, 0, 3, -9,
					-- layer=2 filter=29 channel=9
					-9, 10, 25, 16, 9, 11, 9, -12, 19,
					-- layer=2 filter=29 channel=10
					-20, -14, 0, 1, 8, 8, -10, 4, 5,
					-- layer=2 filter=29 channel=11
					20, 3, -8, 14, -11, -11, 27, 26, 1,
					-- layer=2 filter=29 channel=12
					5, 24, -7, -33, -30, -23, -30, -47, -31,
					-- layer=2 filter=29 channel=13
					-8, -5, 7, -3, 5, 5, -1, 10, -11,
					-- layer=2 filter=29 channel=14
					24, 5, -10, -6, -30, -28, 23, -19, -20,
					-- layer=2 filter=29 channel=15
					-23, -6, -49, 0, -45, 26, -52, 31, 51,
					-- layer=2 filter=29 channel=16
					-16, -14, -21, 9, -10, -5, 24, 7, 10,
					-- layer=2 filter=29 channel=17
					-8, 1, -4, -8, -2, -9, 1, -2, -4,
					-- layer=2 filter=29 channel=18
					-39, -12, -26, -20, -40, -11, -19, -9, -12,
					-- layer=2 filter=29 channel=19
					0, 0, 13, 0, -19, -6, -1, -19, 27,
					-- layer=2 filter=29 channel=20
					8, 8, 1, 7, 4, -1, -7, -4, -1,
					-- layer=2 filter=29 channel=21
					-7, -5, -15, 2, 5, -2, 2, -13, 12,
					-- layer=2 filter=29 channel=22
					0, 3, 1, -4, 1, 3, -5, 0, 9,
					-- layer=2 filter=29 channel=23
					0, -9, -3, -17, 6, -16, -13, 6, 32,
					-- layer=2 filter=29 channel=24
					25, -4, 35, 0, 18, 23, -3, 26, 54,
					-- layer=2 filter=29 channel=25
					-3, 7, 29, 16, 27, 13, 5, 51, 44,
					-- layer=2 filter=29 channel=26
					-2, 4, 0, 4, 3, 2, 4, 0, 0,
					-- layer=2 filter=29 channel=27
					56, 34, 1, 60, 43, 12, 55, 28, 0,
					-- layer=2 filter=29 channel=28
					-66, -34, -55, -47, -43, -53, -23, -44, -31,
					-- layer=2 filter=29 channel=29
					2, -9, -1, 12, -3, 1, 5, 9, -2,
					-- layer=2 filter=29 channel=30
					-34, -1, -2, 16, -3, 11, 14, 12, -11,
					-- layer=2 filter=29 channel=31
					7, 3, -43, 37, -15, -32, -50, 9, 30,
					-- layer=2 filter=29 channel=32
					0, -3, -5, 7, -6, 11, -6, 13, -5,
					-- layer=2 filter=29 channel=33
					-46, -13, -57, -46, -80, -39, -49, -74, -2,
					-- layer=2 filter=29 channel=34
					-5, -13, -37, 0, -3, 20, 27, 13, 40,
					-- layer=2 filter=29 channel=35
					-40, -45, -40, -40, -12, -27, -39, -66, -2,
					-- layer=2 filter=29 channel=36
					4, 15, 7, 3, 1, 2, -3, -1, -7,
					-- layer=2 filter=29 channel=37
					13, -1, -8, 19, -5, -26, 21, 14, -19,
					-- layer=2 filter=29 channel=38
					25, 9, -18, 17, 16, -26, 26, 6, -20,
					-- layer=2 filter=29 channel=39
					-22, -12, -10, -3, 1, -1, -5, -9, 20,
					-- layer=2 filter=29 channel=40
					-35, 10, -9, -32, -24, 33, 7, 12, 77,
					-- layer=2 filter=29 channel=41
					11, -1, -10, -9, -6, -2, -5, -9, -10,
					-- layer=2 filter=29 channel=42
					-20, -10, 10, 0, -23, 13, 5, -16, 19,
					-- layer=2 filter=29 channel=43
					16, -10, -26, -10, -19, -49, 18, -20, 26,
					-- layer=2 filter=29 channel=44
					-3, -5, 8, 9, 5, -3, 0, 11, -3,
					-- layer=2 filter=29 channel=45
					-20, -4, -2, 11, -8, 20, -3, -17, -4,
					-- layer=2 filter=29 channel=46
					-2, -7, -19, -12, 13, -15, 17, 27, -13,
					-- layer=2 filter=29 channel=47
					-2, -19, -67, -22, -40, -32, -2, -14, 5,
					-- layer=2 filter=29 channel=48
					-2, -6, 1, 2, 1, -9, -7, 8, 9,
					-- layer=2 filter=29 channel=49
					28, 7, 29, 40, 26, -18, 24, 25, 16,
					-- layer=2 filter=29 channel=50
					2, 16, 12, 18, -7, -12, -3, -3, 10,
					-- layer=2 filter=29 channel=51
					24, -4, 0, 26, 4, -29, 31, 23, -3,
					-- layer=2 filter=29 channel=52
					16, 0, -18, -11, -66, -35, 13, 8, -21,
					-- layer=2 filter=29 channel=53
					-11, -21, 5, -5, -12, -15, -14, 54, 2,
					-- layer=2 filter=29 channel=54
					-6, -57, -68, -31, -28, -43, 3, 8, 50,
					-- layer=2 filter=29 channel=55
					-13, -3, -3, 0, -8, 6, 4, -6, -9,
					-- layer=2 filter=29 channel=56
					15, -5, -3, 23, -10, -21, 33, 14, -19,
					-- layer=2 filter=29 channel=57
					-2, -11, 4, 5, 4, -9, -4, 3, 1,
					-- layer=2 filter=29 channel=58
					-9, -15, -8, -45, -39, -4, -55, -21, -42,
					-- layer=2 filter=29 channel=59
					-7, -13, -7, -20, 0, 0, -8, 13, 18,
					-- layer=2 filter=29 channel=60
					-6, -11, -1, 6, 11, 47, -10, 9, 30,
					-- layer=2 filter=29 channel=61
					45, -5, 21, 35, 17, 46, 32, 34, 23,
					-- layer=2 filter=29 channel=62
					16, -14, 0, 0, -5, -16, 28, 7, 27,
					-- layer=2 filter=29 channel=63
					2, -25, -23, 2, -17, 0, 6, 21, 13,
					-- layer=2 filter=29 channel=64
					2, 1, -14, -19, -14, 2, 9, 16, 9,
					-- layer=2 filter=29 channel=65
					22, 11, 2, 32, 25, 25, 29, 26, -8,
					-- layer=2 filter=29 channel=66
					1, 27, 1, -4, 0, 2, -20, 25, 37,
					-- layer=2 filter=29 channel=67
					-9, -13, -5, 6, 9, -23, 45, -7, -9,
					-- layer=2 filter=29 channel=68
					6, 8, -9, 9, -5, -10, 3, 4, -3,
					-- layer=2 filter=29 channel=69
					-1, 2, -6, 0, -3, -1, 14, 4, 27,
					-- layer=2 filter=29 channel=70
					-12, -13, -51, -10, -16, -6, -8, -23, -6,
					-- layer=2 filter=29 channel=71
					51, 17, -14, 36, 1, -27, 39, -7, -14,
					-- layer=2 filter=29 channel=72
					-62, -16, -22, -7, -16, -36, -19, -63, 0,
					-- layer=2 filter=29 channel=73
					-29, 16, 38, -1, 0, 6, 52, 11, 42,
					-- layer=2 filter=29 channel=74
					-40, -13, -10, -7, -6, -4, 0, 10, -2,
					-- layer=2 filter=29 channel=75
					0, -25, -11, -4, -29, 24, -30, -57, -76,
					-- layer=2 filter=29 channel=76
					20, 24, -16, -2, -38, -50, 28, -1, -22,
					-- layer=2 filter=29 channel=77
					2, -10, -11, 5, -4, -7, -3, -1, 6,
					-- layer=2 filter=29 channel=78
					-6, -27, 3, 26, -26, -20, -8, 4, 14,
					-- layer=2 filter=29 channel=79
					4, -4, 0, 0, 0, 0, 11, 7, -7,
					-- layer=2 filter=29 channel=80
					-18, -8, 13, 1, 7, 20, 17, 0, 4,
					-- layer=2 filter=29 channel=81
					8, 17, 2, 9, 7, 0, 5, 18, -2,
					-- layer=2 filter=29 channel=82
					-8, 1, 6, 10, -11, -6, -10, 6, -9,
					-- layer=2 filter=29 channel=83
					9, -7, 0, 19, 17, 15, 11, 19, 15,
					-- layer=2 filter=29 channel=84
					-1, -2, -9, -4, -2, 9, -5, 4, -7,
					-- layer=2 filter=29 channel=85
					-7, -7, -14, 0, -6, -1, 4, 0, 7,
					-- layer=2 filter=29 channel=86
					-8, 5, -10, 15, -3, 0, 15, 14, 0,
					-- layer=2 filter=29 channel=87
					-27, -89, -19, -19, -80, -22, -8, -38, 23,
					-- layer=2 filter=29 channel=88
					-31, -16, -11, -16, 5, -1, -9, 27, 21,
					-- layer=2 filter=29 channel=89
					3, -9, 1, -13, -47, -25, -20, -29, -19,
					-- layer=2 filter=29 channel=90
					-7, 4, -1, -7, -5, 4, -6, 0, -8,
					-- layer=2 filter=29 channel=91
					3, 2, -5, -35, -35, 7, -43, -73, -4,
					-- layer=2 filter=29 channel=92
					-9, 17, -13, -19, -11, -12, -29, -41, 20,
					-- layer=2 filter=29 channel=93
					16, 30, 2, -42, 8, 17, -4, 11, -33,
					-- layer=2 filter=29 channel=94
					57, -37, 34, 26, 2, -4, -7, 28, 65,
					-- layer=2 filter=29 channel=95
					-4, 5, 10, -3, -5, 4, 7, 3, 12,
					-- layer=2 filter=29 channel=96
					-19, 5, -41, -5, -36, -21, 31, 24, -3,
					-- layer=2 filter=29 channel=97
					-14, -12, 30, -16, -18, -14, -32, -19, 9,
					-- layer=2 filter=29 channel=98
					2, 3, -20, 23, -22, 5, 7, 13, 1,
					-- layer=2 filter=29 channel=99
					17, 13, -33, -9, -60, -12, 0, 32, -23,
					-- layer=2 filter=29 channel=100
					-2, -15, -12, 8, 4, 7, 5, 0, 2,
					-- layer=2 filter=29 channel=101
					30, 10, 30, 22, 32, -15, 44, 30, -23,
					-- layer=2 filter=29 channel=102
					-39, -5, -50, 10, -54, -1, 31, -11, 9,
					-- layer=2 filter=29 channel=103
					13, 46, -17, -24, 7, -15, 15, -54, 26,
					-- layer=2 filter=29 channel=104
					-15, -13, 18, 3, -2, -40, -30, -15, -3,
					-- layer=2 filter=29 channel=105
					-57, 0, 28, -50, -17, 28, 34, 34, 17,
					-- layer=2 filter=29 channel=106
					29, -1, 24, -12, 4, 8, 4, 26, 15,
					-- layer=2 filter=29 channel=107
					51, -14, -36, 19, 62, 15, -20, -14, 23,
					-- layer=2 filter=29 channel=108
					24, -2, -2, 36, -10, 3, 48, -5, -33,
					-- layer=2 filter=29 channel=109
					13, -12, 2, 27, 3, -12, -4, -1, -2,
					-- layer=2 filter=29 channel=110
					-1, -5, -13, -15, 6, -20, 0, 17, 15,
					-- layer=2 filter=29 channel=111
					6, 1, 1, 6, 0, -12, 10, 4, 6,
					-- layer=2 filter=29 channel=112
					13, -4, 2, 35, 3, -31, 38, 19, -3,
					-- layer=2 filter=29 channel=113
					-16, -14, -6, 17, 7, 14, 10, 19, 4,
					-- layer=2 filter=29 channel=114
					-11, 9, -3, 4, -8, -4, 7, -15, 1,
					-- layer=2 filter=29 channel=115
					-5, 10, -5, -8, -1, 7, 9, -4, -6,
					-- layer=2 filter=29 channel=116
					-39, -26, -34, -15, -66, 4, -15, -12, 27,
					-- layer=2 filter=29 channel=117
					25, -36, -17, -20, -35, -32, 47, -9, 51,
					-- layer=2 filter=29 channel=118
					9, 1, 26, 15, -16, 2, 7, -12, 29,
					-- layer=2 filter=29 channel=119
					-26, -6, -3, 18, 2, 13, 12, 2, 23,
					-- layer=2 filter=29 channel=120
					-5, 0, -4, 10, -5, -5, 9, 6, 8,
					-- layer=2 filter=29 channel=121
					-1, -5, 4, 1, 8, 9, 0, -7, -1,
					-- layer=2 filter=29 channel=122
					-8, 9, 11, -6, -5, -5, -5, -1, 0,
					-- layer=2 filter=29 channel=123
					-35, -66, -60, -18, -8, -15, -15, -30, 1,
					-- layer=2 filter=29 channel=124
					-65, -97, -88, -65, -69, -34, -43, -39, 20,
					-- layer=2 filter=29 channel=125
					0, 1, -10, -5, -7, 4, 8, -6, -3,
					-- layer=2 filter=29 channel=126
					0, 1, 5, -28, 13, -24, -1, 28, 22,
					-- layer=2 filter=29 channel=127
					-8, -5, -7, 6, -16, -3, -28, 4, 19,
					-- layer=2 filter=30 channel=0
					3, 18, -3, -7, 11, -5, 16, -4, -9,
					-- layer=2 filter=30 channel=1
					17, 4, -13, -20, 0, 3, -4, -20, -28,
					-- layer=2 filter=30 channel=2
					1, 6, 1, -6, 7, -9, -2, -5, -8,
					-- layer=2 filter=30 channel=3
					-19, -10, 6, 42, -1, 5, -16, -22, -14,
					-- layer=2 filter=30 channel=4
					-14, -43, -4, -7, -28, -4, 13, -21, 16,
					-- layer=2 filter=30 channel=5
					9, 27, 29, -2, 25, 16, -22, 18, -7,
					-- layer=2 filter=30 channel=6
					-5, -57, -22, -13, -15, -16, 28, 4, 39,
					-- layer=2 filter=30 channel=7
					-28, 6, -2, 9, -5, 6, 6, 8, 33,
					-- layer=2 filter=30 channel=8
					-6, -7, -2, 2, 5, 7, 3, -9, -6,
					-- layer=2 filter=30 channel=9
					-14, -22, -8, 11, -43, -32, -23, -28, -10,
					-- layer=2 filter=30 channel=10
					14, 6, 12, 21, 24, 9, 14, 8, -25,
					-- layer=2 filter=30 channel=11
					0, 26, 16, -5, 11, 17, -12, -1, 22,
					-- layer=2 filter=30 channel=12
					20, 26, 6, -10, -22, 24, -15, -7, 18,
					-- layer=2 filter=30 channel=13
					0, 8, 9, 4, 2, -8, 2, -5, 11,
					-- layer=2 filter=30 channel=14
					20, 11, 16, -27, -14, 12, -30, -38, -20,
					-- layer=2 filter=30 channel=15
					-7, 27, 11, 27, -7, -20, -31, -13, -24,
					-- layer=2 filter=30 channel=16
					-17, -35, 6, 6, -23, 0, 23, -20, -36,
					-- layer=2 filter=30 channel=17
					1, 2, -1, -2, 0, -7, 4, -2, -6,
					-- layer=2 filter=30 channel=18
					16, 6, 32, -2, 13, 43, -39, -21, 9,
					-- layer=2 filter=30 channel=19
					-8, -38, -26, -4, -31, 2, 0, 10, -19,
					-- layer=2 filter=30 channel=20
					6, 2, 0, 10, 0, 1, -6, 4, 2,
					-- layer=2 filter=30 channel=21
					19, 13, 11, -3, -16, -2, 5, 2, 6,
					-- layer=2 filter=30 channel=22
					8, 0, -2, 1, 0, -2, 4, 0, 5,
					-- layer=2 filter=30 channel=23
					0, -53, -33, 39, -8, -19, 0, -5, 5,
					-- layer=2 filter=30 channel=24
					4, 18, 14, 15, 2, 36, 3, -8, 13,
					-- layer=2 filter=30 channel=25
					-11, 29, 0, -1, 15, 25, 17, 22, 25,
					-- layer=2 filter=30 channel=26
					0, -1, 11, 2, 6, 5, 9, 8, 9,
					-- layer=2 filter=30 channel=27
					-8, -3, 0, 8, 1, 10, 10, 1, 18,
					-- layer=2 filter=30 channel=28
					-16, 11, -38, 3, 8, 34, -7, -48, -8,
					-- layer=2 filter=30 channel=29
					8, 2, -4, 4, -8, 8, 6, -1, -7,
					-- layer=2 filter=30 channel=30
					-4, -10, -36, 26, -23, 4, 1, -14, -40,
					-- layer=2 filter=30 channel=31
					6, -15, -46, -41, 13, -74, -34, 21, -20,
					-- layer=2 filter=30 channel=32
					-7, 1, -4, -6, -7, 7, 10, 10, -4,
					-- layer=2 filter=30 channel=33
					-29, 3, 12, 4, 6, -29, -18, -59, 4,
					-- layer=2 filter=30 channel=34
					5, 3, 1, -20, 16, 4, 37, 18, 27,
					-- layer=2 filter=30 channel=35
					-12, -1, -24, 26, 20, 29, -2, -18, 17,
					-- layer=2 filter=30 channel=36
					11, 6, 6, -10, 9, -2, 0, -3, 12,
					-- layer=2 filter=30 channel=37
					0, 19, 4, -10, 10, 10, 6, 29, 8,
					-- layer=2 filter=30 channel=38
					-21, -14, 3, 0, -3, -8, 12, 4, 5,
					-- layer=2 filter=30 channel=39
					-13, -42, -29, 31, -28, 11, -5, -5, -12,
					-- layer=2 filter=30 channel=40
					14, 23, -6, -34, 4, -9, -39, -29, 20,
					-- layer=2 filter=30 channel=41
					10, 2, 7, 6, 6, -12, 0, -2, -2,
					-- layer=2 filter=30 channel=42
					-7, -36, 4, 33, -17, 4, -19, -33, -2,
					-- layer=2 filter=30 channel=43
					-14, -18, -7, -2, 3, -43, -30, -32, -37,
					-- layer=2 filter=30 channel=44
					4, -10, -6, -6, -2, -9, -2, 6, -10,
					-- layer=2 filter=30 channel=45
					-48, -69, -62, -53, -87, -58, -24, -38, -65,
					-- layer=2 filter=30 channel=46
					-33, -58, -27, 1, -45, -47, -1, -36, -18,
					-- layer=2 filter=30 channel=47
					-52, -34, -41, -39, -14, -17, -4, -19, 14,
					-- layer=2 filter=30 channel=48
					5, -1, 11, 0, 5, 6, 4, 2, -9,
					-- layer=2 filter=30 channel=49
					21, -1, 37, 5, -19, 23, -11, -9, -2,
					-- layer=2 filter=30 channel=50
					-21, -12, -10, -10, -20, -4, 0, -10, 1,
					-- layer=2 filter=30 channel=51
					11, 11, 14, -8, 18, 10, 7, 7, 12,
					-- layer=2 filter=30 channel=52
					2, 23, -2, 40, 0, 0, 11, -5, 15,
					-- layer=2 filter=30 channel=53
					-71, -5, -51, -30, -38, 15, -24, -51, 24,
					-- layer=2 filter=30 channel=54
					39, 13, 3, 10, 20, 8, 31, 32, 42,
					-- layer=2 filter=30 channel=55
					8, 2, 0, 5, 2, -4, 5, 12, 10,
					-- layer=2 filter=30 channel=56
					-6, -1, 8, -19, 11, 21, -36, 4, 1,
					-- layer=2 filter=30 channel=57
					-1, 4, -12, -6, -7, -11, 0, 14, -4,
					-- layer=2 filter=30 channel=58
					11, 13, -12, 14, -9, 12, 35, 8, 7,
					-- layer=2 filter=30 channel=59
					-18, 8, -33, -14, 6, 39, 11, 16, 9,
					-- layer=2 filter=30 channel=60
					2, 23, 12, -13, 27, 22, 6, 6, 6,
					-- layer=2 filter=30 channel=61
					13, 12, -3, -32, 11, -16, 2, 0, 13,
					-- layer=2 filter=30 channel=62
					-11, 13, -7, -58, -17, 11, 7, 0, 34,
					-- layer=2 filter=30 channel=63
					-2, -48, -39, 18, -31, -60, 4, -21, -4,
					-- layer=2 filter=30 channel=64
					18, -43, -4, 24, -15, 5, 27, -18, -14,
					-- layer=2 filter=30 channel=65
					26, -19, 30, 8, 16, -1, 28, 7, 49,
					-- layer=2 filter=30 channel=66
					74, 26, 21, -10, -10, -40, -9, 41, -8,
					-- layer=2 filter=30 channel=67
					-26, -52, -36, -27, -72, -73, -23, -49, -14,
					-- layer=2 filter=30 channel=68
					1, 5, 2, 4, 9, -1, 0, -7, -5,
					-- layer=2 filter=30 channel=69
					-8, -33, 8, 27, -21, -8, 11, -18, -13,
					-- layer=2 filter=30 channel=70
					19, 7, 4, 26, 9, 0, 10, 9, 37,
					-- layer=2 filter=30 channel=71
					-35, -56, -60, -34, -51, 0, -26, -38, -40,
					-- layer=2 filter=30 channel=72
					6, -8, 32, 7, 47, 23, 0, -24, 20,
					-- layer=2 filter=30 channel=73
					-17, 30, 35, 25, -46, 18, 12, 9, -13,
					-- layer=2 filter=30 channel=74
					0, -19, -13, 12, -36, -71, 13, -30, -16,
					-- layer=2 filter=30 channel=75
					-24, 16, -50, -26, -20, -16, -9, -29, -24,
					-- layer=2 filter=30 channel=76
					-79, -24, -21, -13, 1, -30, 19, 17, -8,
					-- layer=2 filter=30 channel=77
					9, 5, 0, 12, 4, 0, 11, 12, -7,
					-- layer=2 filter=30 channel=78
					9, 14, 21, -7, 25, -4, 14, 11, 7,
					-- layer=2 filter=30 channel=79
					7, 5, -2, -7, -2, -11, -5, -8, 6,
					-- layer=2 filter=30 channel=80
					19, -19, 3, 38, -28, -60, 22, -20, -33,
					-- layer=2 filter=30 channel=81
					-3, 4, -5, -11, 0, -16, 6, 5, 5,
					-- layer=2 filter=30 channel=82
					0, 5, -6, -3, -5, 5, -8, 4, 12,
					-- layer=2 filter=30 channel=83
					18, -46, -8, 42, -22, -19, 2, 20, 9,
					-- layer=2 filter=30 channel=84
					-10, -3, 2, -5, -3, -11, -5, -5, -3,
					-- layer=2 filter=30 channel=85
					-2, -4, -9, -1, -7, 9, -1, 2, -14,
					-- layer=2 filter=30 channel=86
					14, -3, 2, -5, 3, -16, 9, -11, -9,
					-- layer=2 filter=30 channel=87
					31, 19, 14, 11, 15, 0, 13, 12, 7,
					-- layer=2 filter=30 channel=88
					-3, -25, -27, 28, -18, -64, 19, -36, -31,
					-- layer=2 filter=30 channel=89
					-14, 5, -3, 4, 4, 18, -15, -19, -23,
					-- layer=2 filter=30 channel=90
					2, 3, 5, 1, -5, 3, -2, 0, -11,
					-- layer=2 filter=30 channel=91
					-26, -5, -15, -11, -6, -17, 0, -6, -13,
					-- layer=2 filter=30 channel=92
					4, 2, 16, 7, 2, 24, -13, -5, 11,
					-- layer=2 filter=30 channel=93
					37, -31, 8, -80, -54, -45, -40, -18, -32,
					-- layer=2 filter=30 channel=94
					-45, 12, -23, -26, -20, 9, -3, -3, 23,
					-- layer=2 filter=30 channel=95
					-3, -1, 0, -2, -6, -1, 0, 6, -11,
					-- layer=2 filter=30 channel=96
					-6, -3, -58, 1, -31, 22, 47, 34, 22,
					-- layer=2 filter=30 channel=97
					-17, -14, 32, 27, -8, -1, 16, 13, 4,
					-- layer=2 filter=30 channel=98
					11, 12, -3, -7, 26, 32, 22, -4, 47,
					-- layer=2 filter=30 channel=99
					3, 6, 7, -27, 6, 3, -7, 3, 38,
					-- layer=2 filter=30 channel=100
					-8, 18, 19, 41, 11, -11, 2, 27, 9,
					-- layer=2 filter=30 channel=101
					-44, -39, -28, -18, -43, -22, -12, -20, -6,
					-- layer=2 filter=30 channel=102
					-32, -30, 11, 10, -33, 25, -18, -18, 18,
					-- layer=2 filter=30 channel=103
					4, -31, -21, -52, -3, -53, -12, 29, 7,
					-- layer=2 filter=30 channel=104
					-33, -11, 10, 2, -5, 50, -30, 11, 12,
					-- layer=2 filter=30 channel=105
					-29, -18, -18, -38, 17, -52, -41, 4, 16,
					-- layer=2 filter=30 channel=106
					0, 3, -13, -41, 7, 3, -8, 2, 19,
					-- layer=2 filter=30 channel=107
					-20, -38, 21, -15, 25, 20, -25, 36, 19,
					-- layer=2 filter=30 channel=108
					-15, -16, -14, -12, -32, 24, -25, -26, -11,
					-- layer=2 filter=30 channel=109
					-4, -11, 5, -1, -5, -12, -1, -3, 4,
					-- layer=2 filter=30 channel=110
					38, -31, -10, 48, 23, -2, 23, 2, 8,
					-- layer=2 filter=30 channel=111
					8, 6, 5, 3, 0, 6, 7, 9, 0,
					-- layer=2 filter=30 channel=112
					23, 14, -20, -40, 7, -10, -16, -33, -7,
					-- layer=2 filter=30 channel=113
					17, -19, -9, 8, -5, 4, -17, -5, 15,
					-- layer=2 filter=30 channel=114
					1, -1, 6, 8, 4, -1, 11, 2, 2,
					-- layer=2 filter=30 channel=115
					-1, 11, -7, -10, -6, -1, 0, 8, 7,
					-- layer=2 filter=30 channel=116
					21, -4, -16, 18, -10, -38, 22, 15, 1,
					-- layer=2 filter=30 channel=117
					-16, -12, 32, -15, -31, -13, -29, -12, 30,
					-- layer=2 filter=30 channel=118
					0, -5, 24, 26, 30, 10, 17, 29, 1,
					-- layer=2 filter=30 channel=119
					-33, -17, -2, -12, -10, 18, -33, -29, 3,
					-- layer=2 filter=30 channel=120
					7, 6, 8, -2, 6, 2, -9, -6, -1,
					-- layer=2 filter=30 channel=121
					-8, -7, 2, 2, -3, -10, -4, 0, 5,
					-- layer=2 filter=30 channel=122
					10, 6, -12, -6, 6, 8, 6, -3, 3,
					-- layer=2 filter=30 channel=123
					-2, -2, 11, -9, 12, 15, -6, 25, 34,
					-- layer=2 filter=30 channel=124
					36, 24, -8, 9, -25, -28, -9, -10, -15,
					-- layer=2 filter=30 channel=125
					-5, -3, 6, -9, 8, -10, 6, 13, 0,
					-- layer=2 filter=30 channel=126
					-45, -31, -53, -18, -129, -69, -11, -61, -114,
					-- layer=2 filter=30 channel=127
					7, -13, -28, 21, -30, 0, -20, -44, 0,
					-- layer=2 filter=31 channel=0
					-27, -12, -13, -8, 13, -6, 7, 42, 7,
					-- layer=2 filter=31 channel=1
					-20, -81, -16, -25, -6, -5, -17, -7, -4,
					-- layer=2 filter=31 channel=2
					1, 4, -6, 6, 5, 3, -5, -9, 0,
					-- layer=2 filter=31 channel=3
					10, 22, 15, -18, -1, 48, 26, -10, -40,
					-- layer=2 filter=31 channel=4
					-17, -34, -50, -1, -17, -19, 23, 26, -2,
					-- layer=2 filter=31 channel=5
					-21, -5, -7, -6, 6, -11, 10, 38, 0,
					-- layer=2 filter=31 channel=6
					42, 31, 11, 26, 6, 14, 57, 7, 30,
					-- layer=2 filter=31 channel=7
					27, 48, 41, 22, 26, 36, -17, -10, 7,
					-- layer=2 filter=31 channel=8
					11, 3, -3, 2, 0, -3, 4, -5, 4,
					-- layer=2 filter=31 channel=9
					4, 12, 11, -70, -24, -42, 26, 37, 20,
					-- layer=2 filter=31 channel=10
					-22, -16, -3, -31, 3, -4, 9, 1, -14,
					-- layer=2 filter=31 channel=11
					16, -9, -20, 8, -9, -21, -15, 21, 1,
					-- layer=2 filter=31 channel=12
					-22, -67, 8, -2, -13, -25, 16, 26, 38,
					-- layer=2 filter=31 channel=13
					10, -9, 3, 10, 4, 2, 4, -1, 8,
					-- layer=2 filter=31 channel=14
					-13, -77, -27, -22, -25, -39, -18, 8, 5,
					-- layer=2 filter=31 channel=15
					-35, -17, -51, 21, -4, -30, -41, 10, 21,
					-- layer=2 filter=31 channel=16
					-26, -3, 17, -28, 0, -15, -39, -29, -31,
					-- layer=2 filter=31 channel=17
					7, 5, 8, 4, -7, 1, -7, 0, -1,
					-- layer=2 filter=31 channel=18
					22, -29, -34, 17, 5, -16, 7, 17, 23,
					-- layer=2 filter=31 channel=19
					0, -43, -31, 6, 9, 13, -15, 0, -23,
					-- layer=2 filter=31 channel=20
					-2, -1, 0, 1, -7, 6, 4, -3, 7,
					-- layer=2 filter=31 channel=21
					-5, 0, 3, 6, -15, -11, 10, -4, -10,
					-- layer=2 filter=31 channel=22
					-4, -8, 1, 4, 4, 5, 4, -1, 7,
					-- layer=2 filter=31 channel=23
					20, -24, 24, -1, -29, 14, 37, 30, 51,
					-- layer=2 filter=31 channel=24
					11, 12, 11, -6, -24, 0, 2, -14, -51,
					-- layer=2 filter=31 channel=25
					-35, -10, -5, -8, -7, -14, -8, -19, -51,
					-- layer=2 filter=31 channel=26
					-10, -2, 7, 5, -4, 3, 10, 1, 5,
					-- layer=2 filter=31 channel=27
					-25, -28, -65, -55, -44, -45, -20, 2, 3,
					-- layer=2 filter=31 channel=28
					26, 4, 23, 30, 26, 42, 34, 4, 3,
					-- layer=2 filter=31 channel=29
					-6, -11, 4, 3, 3, -8, 0, -4, 7,
					-- layer=2 filter=31 channel=30
					-69, -39, -71, -6, 2, 13, 22, 8, 23,
					-- layer=2 filter=31 channel=31
					-18, 56, -15, -4, -5, -35, -14, 42, 79,
					-- layer=2 filter=31 channel=32
					-4, -9, -4, -9, 10, 4, 8, -4, 5,
					-- layer=2 filter=31 channel=33
					15, 1, -18, 17, 7, 4, 21, 4, -32,
					-- layer=2 filter=31 channel=34
					48, 22, 5, -6, 36, 11, -37, 0, 0,
					-- layer=2 filter=31 channel=35
					62, 10, 29, 13, 27, 22, 17, -9, 15,
					-- layer=2 filter=31 channel=36
					1, 9, -7, -2, 0, 8, 21, 10, -7,
					-- layer=2 filter=31 channel=37
					2, -11, -13, 7, -19, -25, 3, 3, -17,
					-- layer=2 filter=31 channel=38
					-10, -21, -30, -19, 11, -18, -15, 30, 33,
					-- layer=2 filter=31 channel=39
					-27, -13, -3, 12, -30, -3, -21, -5, 19,
					-- layer=2 filter=31 channel=40
					17, 9, -12, 49, 17, 54, 23, 36, -20,
					-- layer=2 filter=31 channel=41
					3, -4, -11, 8, -3, 5, -8, -2, -4,
					-- layer=2 filter=31 channel=42
					-4, 5, 2, 3, -25, 10, 21, -25, 3,
					-- layer=2 filter=31 channel=43
					-50, -46, -66, -10, -8, -15, 2, -33, -13,
					-- layer=2 filter=31 channel=44
					2, 3, -1, -8, -9, 9, -4, 10, 5,
					-- layer=2 filter=31 channel=45
					-71, -16, 9, -7, -7, -8, -29, -17, -18,
					-- layer=2 filter=31 channel=46
					-36, -30, -69, -16, 1, -23, -7, 8, -6,
					-- layer=2 filter=31 channel=47
					21, 1, 60, 12, 22, 25, 39, 17, 25,
					-- layer=2 filter=31 channel=48
					-8, -5, 8, 9, -2, 9, 4, 6, 0,
					-- layer=2 filter=31 channel=49
					2, -4, -35, 23, -31, -12, -24, -23, 0,
					-- layer=2 filter=31 channel=50
					-17, 2, -16, 1, -1, 21, -4, 3, -11,
					-- layer=2 filter=31 channel=51
					-16, -13, -3, 4, -7, -5, 7, 8, 4,
					-- layer=2 filter=31 channel=52
					3, -40, -12, -15, 8, -18, -1, -12, 10,
					-- layer=2 filter=31 channel=53
					-7, 16, -52, -16, 50, 10, -14, 52, -22,
					-- layer=2 filter=31 channel=54
					11, 24, 29, 38, 19, 32, 17, 10, 20,
					-- layer=2 filter=31 channel=55
					0, -8, 14, -1, 16, 17, 8, 16, -2,
					-- layer=2 filter=31 channel=56
					10, -17, -15, 18, -16, -35, -11, 24, 15,
					-- layer=2 filter=31 channel=57
					9, -5, -3, 3, -5, 7, -1, -7, 0,
					-- layer=2 filter=31 channel=58
					-11, -74, 1, 12, -12, -14, 8, 16, 54,
					-- layer=2 filter=31 channel=59
					-2, -27, -44, -23, 13, 1, -27, 32, 23,
					-- layer=2 filter=31 channel=60
					-26, -10, -3, 29, 29, 11, 13, 14, 7,
					-- layer=2 filter=31 channel=61
					-13, -7, 20, 8, 0, 28, -8, 5, 6,
					-- layer=2 filter=31 channel=62
					25, -17, -40, -7, 5, 13, -3, 15, -1,
					-- layer=2 filter=31 channel=63
					-28, -30, -13, 1, -20, 6, -12, 3, 49,
					-- layer=2 filter=31 channel=64
					-8, -7, 13, 2, -6, 10, 16, 8, 0,
					-- layer=2 filter=31 channel=65
					18, -10, 13, 12, 0, -5, 0, 0, 15,
					-- layer=2 filter=31 channel=66
					29, 40, 72, 0, 24, 33, 12, 24, -46,
					-- layer=2 filter=31 channel=67
					-57, -4, -73, -79, -55, -81, -16, -2, 0,
					-- layer=2 filter=31 channel=68
					-9, 5, 0, 4, 2, 2, -4, 5, -11,
					-- layer=2 filter=31 channel=69
					4, -21, 7, 7, -18, 21, 13, -10, -10,
					-- layer=2 filter=31 channel=70
					39, 8, 33, 31, 28, 31, -2, 3, 26,
					-- layer=2 filter=31 channel=71
					0, -3, -25, -69, -87, -64, -32, -1, 0,
					-- layer=2 filter=31 channel=72
					18, -41, -11, 31, -2, -11, 0, 12, -28,
					-- layer=2 filter=31 channel=73
					28, 73, 19, -14, -9, 13, -15, 3, 2,
					-- layer=2 filter=31 channel=74
					-55, -37, -76, -42, -20, -12, -7, -13, 40,
					-- layer=2 filter=31 channel=75
					-34, -45, -51, 10, 36, -23, -12, -33, -57,
					-- layer=2 filter=31 channel=76
					-3, 10, 21, 57, 13, 69, 5, 37, 36,
					-- layer=2 filter=31 channel=77
					-3, -5, -7, -4, 6, 5, -5, -6, 2,
					-- layer=2 filter=31 channel=78
					1, 1, -10, -7, -9, 5, -10, -17, -18,
					-- layer=2 filter=31 channel=79
					-2, 0, -2, 2, -10, -3, 6, -7, 8,
					-- layer=2 filter=31 channel=80
					1, 4, 13, 0, -5, 18, 22, -3, -13,
					-- layer=2 filter=31 channel=81
					-6, -6, 2, -18, -5, 3, -3, -12, 0,
					-- layer=2 filter=31 channel=82
					0, 7, 4, -7, 9, 12, -6, -2, 0,
					-- layer=2 filter=31 channel=83
					-12, -6, -19, 29, -23, -17, 17, -21, 6,
					-- layer=2 filter=31 channel=84
					-11, 5, 6, 5, 4, -6, 8, 3, 5,
					-- layer=2 filter=31 channel=85
					1, -14, -19, -16, -9, -3, -6, -18, -2,
					-- layer=2 filter=31 channel=86
					-2, 0, 19, 16, 2, 4, 0, 7, 5,
					-- layer=2 filter=31 channel=87
					26, 4, -9, 58, 39, 25, 18, 37, 23,
					-- layer=2 filter=31 channel=88
					-37, -59, -68, -8, -14, -22, 18, -17, 17,
					-- layer=2 filter=31 channel=89
					-26, -66, -21, 4, -3, -32, -30, -6, 3,
					-- layer=2 filter=31 channel=90
					-3, 8, 4, 3, -5, -4, -2, 3, -11,
					-- layer=2 filter=31 channel=91
					-55, -94, -21, 5, -13, -30, 12, -30, -37,
					-- layer=2 filter=31 channel=92
					-20, -42, 0, -42, -25, -50, -16, -10, 9,
					-- layer=2 filter=31 channel=93
					52, -46, -11, -35, -46, -15, -24, -55, -25,
					-- layer=2 filter=31 channel=94
					12, 24, 17, 40, 13, 47, 36, 39, 24,
					-- layer=2 filter=31 channel=95
					3, -9, -8, 6, 14, -1, 6, -3, -2,
					-- layer=2 filter=31 channel=96
					23, -59, 9, 33, 15, 12, 12, 20, 27,
					-- layer=2 filter=31 channel=97
					18, -5, -17, -18, -16, -4, 41, 1, -13,
					-- layer=2 filter=31 channel=98
					26, 9, 55, 20, 44, 49, 10, 1, 13,
					-- layer=2 filter=31 channel=99
					13, -12, 21, 8, 20, 3, -8, -27, -21,
					-- layer=2 filter=31 channel=100
					-41, -42, -28, 15, -18, -30, -6, 9, 40,
					-- layer=2 filter=31 channel=101
					-43, -42, -9, -42, -31, -44, -8, -19, -28,
					-- layer=2 filter=31 channel=102
					-2, -62, 13, 3, -11, -20, -13, -17, 36,
					-- layer=2 filter=31 channel=103
					-13, -23, 26, -11, 23, -62, 29, 15, -17,
					-- layer=2 filter=31 channel=104
					-4, -16, -50, 40, 2, -12, 19, 28, 40,
					-- layer=2 filter=31 channel=105
					-63, -78, 29, 57, 12, 40, -44, 3, 18,
					-- layer=2 filter=31 channel=106
					-16, -77, -27, -20, -24, -44, -1, 2, -18,
					-- layer=2 filter=31 channel=107
					-2, 45, 35, 6, -10, -43, 25, 0, 83,
					-- layer=2 filter=31 channel=108
					-34, -40, -4, -29, -30, -27, -37, -34, -1,
					-- layer=2 filter=31 channel=109
					-1, -7, -15, 6, 8, 4, -5, 0, -15,
					-- layer=2 filter=31 channel=110
					-11, 8, 35, -12, -4, -22, 0, -53, -35,
					-- layer=2 filter=31 channel=111
					4, 5, 7, 3, 1, 9, 4, 0, 2,
					-- layer=2 filter=31 channel=112
					-22, -40, -4, -9, -14, -32, -14, -11, -12,
					-- layer=2 filter=31 channel=113
					-44, -22, 0, 4, -2, 5, 30, -13, 27,
					-- layer=2 filter=31 channel=114
					-3, 2, -14, 4, -11, 7, 9, -5, 0,
					-- layer=2 filter=31 channel=115
					-7, -3, 0, -3, 2, -10, 11, 5, 6,
					-- layer=2 filter=31 channel=116
					23, 0, -11, 46, 15, 12, 21, -14, 48,
					-- layer=2 filter=31 channel=117
					7, 0, -9, 3, 0, -17, -20, -27, -24,
					-- layer=2 filter=31 channel=118
					21, 23, -6, 6, -2, -10, 15, -9, -33,
					-- layer=2 filter=31 channel=119
					20, -32, -24, 18, 3, -29, -4, 21, -2,
					-- layer=2 filter=31 channel=120
					2, -5, -2, -7, -9, -7, -6, -10, -3,
					-- layer=2 filter=31 channel=121
					-10, 2, 1, -10, -8, 2, -1, -3, 3,
					-- layer=2 filter=31 channel=122
					-7, 9, 14, 1, 0, 3, 10, 16, 9,
					-- layer=2 filter=31 channel=123
					46, 0, 37, 34, 26, 41, -6, 20, 22,
					-- layer=2 filter=31 channel=124
					-16, -1, -26, 8, 31, -11, -7, 5, 3,
					-- layer=2 filter=31 channel=125
					4, 7, 9, 6, -3, -11, 6, 0, -9,
					-- layer=2 filter=31 channel=126
					-27, -36, -34, -29, 13, 3, -58, -4, -62,
					-- layer=2 filter=31 channel=127
					-18, -59, -33, -9, -27, 28, 38, 8, 36,
					-- layer=2 filter=32 channel=0
					-12, 3, -5, -2, -6, 7, 3, -9, -6,
					-- layer=2 filter=32 channel=1
					-10, 0, 0, -10, 8, -7, -8, -3, -8,
					-- layer=2 filter=32 channel=2
					7, -1, 5, -10, 0, 0, 2, 7, -8,
					-- layer=2 filter=32 channel=3
					-11, -5, -9, -7, -6, -2, 5, -9, 7,
					-- layer=2 filter=32 channel=4
					-12, 0, 0, -13, -2, 0, -8, 6, -8,
					-- layer=2 filter=32 channel=5
					-9, 0, -7, -3, 2, 6, -11, -7, -5,
					-- layer=2 filter=32 channel=6
					2, -6, -3, 6, -11, 2, -8, -3, 4,
					-- layer=2 filter=32 channel=7
					7, 0, -8, 6, 0, -6, 0, -7, -1,
					-- layer=2 filter=32 channel=8
					4, -8, -9, 7, 0, -1, 5, 3, 0,
					-- layer=2 filter=32 channel=9
					1, 5, -1, 0, 1, -9, 4, -6, -4,
					-- layer=2 filter=32 channel=10
					-12, -2, 0, -2, 5, 0, 5, -3, -4,
					-- layer=2 filter=32 channel=11
					3, 1, 4, -2, -11, 4, -7, -16, -7,
					-- layer=2 filter=32 channel=12
					6, 4, -11, -12, -10, 1, -1, 5, -3,
					-- layer=2 filter=32 channel=13
					-6, 4, -8, -1, -6, -11, -7, -4, 10,
					-- layer=2 filter=32 channel=14
					-12, -3, 7, -6, -12, 6, 1, -1, -5,
					-- layer=2 filter=32 channel=15
					3, -8, -10, 6, -3, -3, -8, -9, -12,
					-- layer=2 filter=32 channel=16
					-4, -9, -8, -5, -8, 4, -3, 2, 2,
					-- layer=2 filter=32 channel=17
					-10, -5, 0, -1, -1, 8, -4, -9, -6,
					-- layer=2 filter=32 channel=18
					-7, 0, -3, -5, 2, -4, 3, -6, 4,
					-- layer=2 filter=32 channel=19
					-12, 5, 0, -14, 2, -12, -2, 0, -16,
					-- layer=2 filter=32 channel=20
					5, 4, 2, -6, -5, 4, 0, -10, 4,
					-- layer=2 filter=32 channel=21
					1, -7, 2, -11, -4, 9, 6, -2, 8,
					-- layer=2 filter=32 channel=22
					-1, 8, 6, 6, 1, -10, 0, 7, -7,
					-- layer=2 filter=32 channel=23
					7, 7, -7, 0, 0, 0, 0, -2, 4,
					-- layer=2 filter=32 channel=24
					7, -10, -8, -9, -12, 6, 4, -10, -10,
					-- layer=2 filter=32 channel=25
					3, -1, -1, 8, -9, 2, -1, 7, -10,
					-- layer=2 filter=32 channel=26
					-8, 0, 0, -1, -2, 4, 7, 8, 4,
					-- layer=2 filter=32 channel=27
					-1, -11, -14, -7, 2, -11, -4, 0, -2,
					-- layer=2 filter=32 channel=28
					-5, 3, -5, 0, -14, -11, 3, 0, 6,
					-- layer=2 filter=32 channel=29
					4, -2, 6, 4, -8, -4, -3, -8, 3,
					-- layer=2 filter=32 channel=30
					-11, -12, 1, 7, 4, -10, 3, 0, 0,
					-- layer=2 filter=32 channel=31
					-7, -7, 8, 4, 5, -1, 4, -9, 5,
					-- layer=2 filter=32 channel=32
					-4, 2, 7, -12, 7, -3, -7, 7, 0,
					-- layer=2 filter=32 channel=33
					7, 5, 2, -14, -4, 5, 4, 4, 4,
					-- layer=2 filter=32 channel=34
					7, 5, -6, -1, -15, -8, -1, -10, 1,
					-- layer=2 filter=32 channel=35
					-9, 7, 3, 1, 6, 0, 0, 2, 2,
					-- layer=2 filter=32 channel=36
					-8, 0, -3, -11, 0, 4, 7, 0, -5,
					-- layer=2 filter=32 channel=37
					0, -13, -8, -10, -10, 5, -3, -2, -9,
					-- layer=2 filter=32 channel=38
					-1, 0, -10, -1, -10, -12, -8, -12, 6,
					-- layer=2 filter=32 channel=39
					-1, -4, -9, 7, -12, 5, -4, -1, -10,
					-- layer=2 filter=32 channel=40
					-5, -7, 0, -7, 1, 9, -4, -7, 7,
					-- layer=2 filter=32 channel=41
					5, 6, 3, -5, 6, -2, -11, 3, 0,
					-- layer=2 filter=32 channel=42
					-1, 6, -5, -10, 7, 8, -9, 0, 2,
					-- layer=2 filter=32 channel=43
					-8, -10, 6, -3, -6, -3, 0, 0, -6,
					-- layer=2 filter=32 channel=44
					-3, 2, 3, 10, 9, 3, 7, -8, 6,
					-- layer=2 filter=32 channel=45
					1, -10, 8, -8, -1, 0, 3, -4, -8,
					-- layer=2 filter=32 channel=46
					-6, -6, 6, 4, -9, 0, 0, -1, -11,
					-- layer=2 filter=32 channel=47
					2, -10, -9, -3, -4, -8, -5, -1, -8,
					-- layer=2 filter=32 channel=48
					-10, 7, 5, 7, -1, 2, -8, 7, -1,
					-- layer=2 filter=32 channel=49
					-6, 1, 2, -6, 1, 9, -3, -6, 6,
					-- layer=2 filter=32 channel=50
					0, -7, -4, 8, 3, -4, -8, 0, -8,
					-- layer=2 filter=32 channel=51
					2, 0, -5, -11, -15, -12, -3, -11, -8,
					-- layer=2 filter=32 channel=52
					-12, -2, 5, -8, -16, 3, -12, -6, -7,
					-- layer=2 filter=32 channel=53
					-6, 2, -7, 5, -1, -15, 2, 5, -1,
					-- layer=2 filter=32 channel=54
					-6, -2, -5, -5, 0, -8, -9, 4, 1,
					-- layer=2 filter=32 channel=55
					-6, 5, -9, -7, -4, -2, 2, 8, -8,
					-- layer=2 filter=32 channel=56
					6, -7, 5, -14, -6, 4, -11, -8, 2,
					-- layer=2 filter=32 channel=57
					4, 5, 7, 6, -2, 0, 4, 1, 6,
					-- layer=2 filter=32 channel=58
					-2, 8, -11, 2, 0, 8, -9, 3, 3,
					-- layer=2 filter=32 channel=59
					-5, 8, 3, -1, 2, 7, 2, 1, -11,
					-- layer=2 filter=32 channel=60
					-6, 6, -12, -5, -6, -6, -2, 4, 2,
					-- layer=2 filter=32 channel=61
					-4, -11, -7, 5, -2, -8, 0, -11, -3,
					-- layer=2 filter=32 channel=62
					-10, -12, 1, -6, -4, 8, 9, -3, 8,
					-- layer=2 filter=32 channel=63
					-1, -7, -5, -4, 0, 0, -1, -7, -5,
					-- layer=2 filter=32 channel=64
					-6, 6, 0, -10, -5, -8, -3, 2, -12,
					-- layer=2 filter=32 channel=65
					3, 5, 1, 2, -5, -12, -9, -10, -7,
					-- layer=2 filter=32 channel=66
					4, 9, -3, -3, 4, 3, -4, -7, -10,
					-- layer=2 filter=32 channel=67
					-6, -5, 4, 2, 1, 6, 0, -9, 2,
					-- layer=2 filter=32 channel=68
					-6, -10, -6, -1, -8, 1, 0, -8, -3,
					-- layer=2 filter=32 channel=69
					-5, 8, 11, 9, -3, 5, 0, 7, 5,
					-- layer=2 filter=32 channel=70
					3, -13, -6, -4, -14, -7, -14, 1, -4,
					-- layer=2 filter=32 channel=71
					-2, -3, 0, 1, -12, 4, -2, -5, 3,
					-- layer=2 filter=32 channel=72
					-5, -1, 5, -1, -1, -11, 1, -11, -6,
					-- layer=2 filter=32 channel=73
					-5, -1, 0, -7, -10, 2, 0, 0, -3,
					-- layer=2 filter=32 channel=74
					6, -2, -4, 2, 0, -4, 2, -12, -8,
					-- layer=2 filter=32 channel=75
					-13, 0, 7, -7, 7, 7, -2, -6, 0,
					-- layer=2 filter=32 channel=76
					-4, -14, -11, -2, -6, 2, -2, -6, 1,
					-- layer=2 filter=32 channel=77
					7, 1, 3, -7, 7, -3, -9, -8, 7,
					-- layer=2 filter=32 channel=78
					-10, -6, -6, -2, -13, -12, -1, 0, 0,
					-- layer=2 filter=32 channel=79
					0, -9, -5, 5, -1, -10, 5, 3, -7,
					-- layer=2 filter=32 channel=80
					3, -2, -8, -1, 4, -2, -9, 4, -6,
					-- layer=2 filter=32 channel=81
					-6, -6, -2, 0, -4, -6, 2, -9, -5,
					-- layer=2 filter=32 channel=82
					2, -8, 0, 5, -1, -7, 7, 9, -9,
					-- layer=2 filter=32 channel=83
					-9, 2, -9, -9, -4, 4, -9, -5, -12,
					-- layer=2 filter=32 channel=84
					-6, 5, 5, -6, 8, 8, -1, -10, 1,
					-- layer=2 filter=32 channel=85
					-4, -7, 0, -2, 9, -9, 5, 0, 5,
					-- layer=2 filter=32 channel=86
					9, -2, 6, -10, 5, -1, -6, 0, -3,
					-- layer=2 filter=32 channel=87
					-8, 4, 8, 7, 1, 6, -5, -9, 6,
					-- layer=2 filter=32 channel=88
					-3, 5, -8, -13, -12, -9, -2, 1, -9,
					-- layer=2 filter=32 channel=89
					-8, -11, -1, 5, 2, -2, -9, -10, -8,
					-- layer=2 filter=32 channel=90
					-2, 0, -10, 2, 0, 3, -9, -2, -9,
					-- layer=2 filter=32 channel=91
					-13, -10, -2, -9, 9, -2, -9, -4, 3,
					-- layer=2 filter=32 channel=92
					-17, -4, -1, 3, 1, 5, 4, -10, 1,
					-- layer=2 filter=32 channel=93
					-1, -8, -3, 1, 0, 9, 4, -2, 4,
					-- layer=2 filter=32 channel=94
					-1, -14, 3, -2, 7, -10, 1, 2, -1,
					-- layer=2 filter=32 channel=95
					-1, 6, 0, -8, 3, -3, -2, 5, -10,
					-- layer=2 filter=32 channel=96
					4, -9, 4, 0, -1, -5, 4, 5, -12,
					-- layer=2 filter=32 channel=97
					0, -9, -12, 4, -5, -1, 2, 1, -1,
					-- layer=2 filter=32 channel=98
					0, -12, -6, -6, -4, 0, -6, 0, -2,
					-- layer=2 filter=32 channel=99
					-7, -12, -14, -14, -9, -6, -12, -11, -9,
					-- layer=2 filter=32 channel=100
					-5, 5, 3, -11, -8, -10, 4, -3, 7,
					-- layer=2 filter=32 channel=101
					-9, -5, 0, 2, 0, -9, 0, 4, 8,
					-- layer=2 filter=32 channel=102
					-4, -16, 0, -1, -7, -4, -5, 0, -11,
					-- layer=2 filter=32 channel=103
					6, 2, 2, 4, 0, 1, 3, 4, -10,
					-- layer=2 filter=32 channel=104
					-2, -11, -7, 0, 0, 0, 2, -2, 4,
					-- layer=2 filter=32 channel=105
					-4, -4, 0, -5, 0, 3, 2, 0, -4,
					-- layer=2 filter=32 channel=106
					1, -9, -3, 6, -3, 1, -3, -6, 4,
					-- layer=2 filter=32 channel=107
					0, 1, 7, 0, -6, -7, -8, -8, -8,
					-- layer=2 filter=32 channel=108
					-6, 6, 0, -2, -11, -6, -3, -2, -10,
					-- layer=2 filter=32 channel=109
					-2, -3, 8, -9, 2, -5, -5, 2, 7,
					-- layer=2 filter=32 channel=110
					-4, 7, -5, 5, 0, -10, -9, -11, 4,
					-- layer=2 filter=32 channel=111
					0, -1, -2, 7, 8, -9, -11, 4, -9,
					-- layer=2 filter=32 channel=112
					-7, -2, 6, -7, -8, 0, 8, -3, -7,
					-- layer=2 filter=32 channel=113
					6, -6, -13, 5, 0, -8, -2, -1, 7,
					-- layer=2 filter=32 channel=114
					-8, -5, 4, -3, 6, -8, 0, 8, 1,
					-- layer=2 filter=32 channel=115
					2, 5, -7, 5, 6, 8, 8, 5, -10,
					-- layer=2 filter=32 channel=116
					3, -3, 6, -3, -11, 6, 0, -2, -1,
					-- layer=2 filter=32 channel=117
					6, 1, -4, -8, -5, -7, -7, -10, -12,
					-- layer=2 filter=32 channel=118
					-2, -7, -12, -5, 2, -11, 5, -8, -3,
					-- layer=2 filter=32 channel=119
					-5, 5, 6, -11, 6, -6, 0, -10, 0,
					-- layer=2 filter=32 channel=120
					-9, 6, -3, 1, 0, 3, 4, 3, 1,
					-- layer=2 filter=32 channel=121
					9, 0, 1, -2, -2, 3, 11, -9, -5,
					-- layer=2 filter=32 channel=122
					5, 6, 3, -9, 7, 2, -4, -6, -4,
					-- layer=2 filter=32 channel=123
					0, -4, -10, -6, -11, -3, 0, -7, -14,
					-- layer=2 filter=32 channel=124
					-6, 0, -7, 5, 2, -11, 5, -9, -11,
					-- layer=2 filter=32 channel=125
					-2, -4, 10, -3, -7, -2, -7, -2, -4,
					-- layer=2 filter=32 channel=126
					2, -3, -7, -3, 0, -5, -8, -9, -7,
					-- layer=2 filter=32 channel=127
					-14, -6, 0, -12, 7, 7, 1, 6, 1,
					-- layer=2 filter=33 channel=0
					4, -11, -2, 8, -2, 1, -4, 1, 0,
					-- layer=2 filter=33 channel=1
					5, 2, -5, -5, 0, -9, 5, -3, -8,
					-- layer=2 filter=33 channel=2
					0, 8, 5, 0, 8, -9, 3, 6, -3,
					-- layer=2 filter=33 channel=3
					5, 9, -4, 3, -9, 8, -10, 8, -2,
					-- layer=2 filter=33 channel=4
					-3, 8, 6, -7, -9, -7, 6, 7, 5,
					-- layer=2 filter=33 channel=5
					5, -11, -10, 1, -10, -4, -10, 0, 1,
					-- layer=2 filter=33 channel=6
					-9, 0, -6, -7, -5, -2, 6, 3, -11,
					-- layer=2 filter=33 channel=7
					9, 4, -11, -7, -7, 0, -10, -5, -10,
					-- layer=2 filter=33 channel=8
					2, -3, -1, -8, -6, 0, 2, -9, 0,
					-- layer=2 filter=33 channel=9
					-2, 3, 0, 2, 2, 6, -3, -5, 1,
					-- layer=2 filter=33 channel=10
					3, -2, -9, -6, -1, -7, -3, 5, 1,
					-- layer=2 filter=33 channel=11
					5, -1, -5, 8, 1, 1, 7, 10, 3,
					-- layer=2 filter=33 channel=12
					-5, 2, -13, 9, 0, -7, 7, 0, -8,
					-- layer=2 filter=33 channel=13
					-1, -8, 0, -2, -11, -4, -7, -1, -12,
					-- layer=2 filter=33 channel=14
					4, 0, -12, 0, 0, -6, 5, 2, -4,
					-- layer=2 filter=33 channel=15
					4, -10, -11, -7, 0, 6, -7, 0, 1,
					-- layer=2 filter=33 channel=16
					5, -9, 3, -2, 8, -5, 6, 0, 4,
					-- layer=2 filter=33 channel=17
					-9, 4, 3, -7, 9, -3, -9, -2, 6,
					-- layer=2 filter=33 channel=18
					-13, 4, -8, 1, -8, 10, 5, 0, -12,
					-- layer=2 filter=33 channel=19
					0, -11, 4, -12, -1, 5, 2, -3, 3,
					-- layer=2 filter=33 channel=20
					-5, -6, 2, 8, -6, 0, 1, -8, 0,
					-- layer=2 filter=33 channel=21
					-5, 2, 0, 7, -9, 1, 8, 5, -5,
					-- layer=2 filter=33 channel=22
					7, -3, 7, -5, -4, -3, 5, -10, -10,
					-- layer=2 filter=33 channel=23
					-5, -7, 6, -2, -11, 7, -1, -10, -8,
					-- layer=2 filter=33 channel=24
					3, -8, -2, -4, 4, 0, 0, -9, 0,
					-- layer=2 filter=33 channel=25
					-10, 5, 0, 9, -12, 2, 2, 0, -2,
					-- layer=2 filter=33 channel=26
					-5, -1, 5, -4, 2, 6, -8, 5, 4,
					-- layer=2 filter=33 channel=27
					-9, -10, 1, 8, 7, 1, -4, 5, -7,
					-- layer=2 filter=33 channel=28
					3, -4, -2, -7, -8, 7, 6, 2, -8,
					-- layer=2 filter=33 channel=29
					3, 6, 4, 6, -3, -7, 0, 3, -12,
					-- layer=2 filter=33 channel=30
					-9, 0, -9, -5, 8, 4, 2, -8, -7,
					-- layer=2 filter=33 channel=31
					-5, -2, -4, -5, 5, -4, -6, 0, 5,
					-- layer=2 filter=33 channel=32
					6, 2, 7, 4, 0, 8, 7, 6, -10,
					-- layer=2 filter=33 channel=33
					3, 1, -6, -7, 7, -5, -4, -4, 2,
					-- layer=2 filter=33 channel=34
					-6, -3, 0, 6, -12, -10, 0, -7, 7,
					-- layer=2 filter=33 channel=35
					1, 0, 4, -3, -6, -2, 5, -10, 4,
					-- layer=2 filter=33 channel=36
					6, 3, 3, 8, -10, -11, 4, 2, -2,
					-- layer=2 filter=33 channel=37
					-3, 2, 2, -8, -9, -6, 7, 3, -1,
					-- layer=2 filter=33 channel=38
					0, -10, 5, 7, 0, 7, -5, 0, 3,
					-- layer=2 filter=33 channel=39
					4, -8, 8, -9, 4, 0, -2, -6, -5,
					-- layer=2 filter=33 channel=40
					-2, 3, 0, -6, -5, -7, 7, -5, 1,
					-- layer=2 filter=33 channel=41
					-6, -5, -8, 0, 8, -8, 7, 1, 9,
					-- layer=2 filter=33 channel=42
					0, -4, 2, 0, 3, -7, -7, 7, -6,
					-- layer=2 filter=33 channel=43
					7, 6, 5, 4, -10, 3, 5, -8, 2,
					-- layer=2 filter=33 channel=44
					-6, 3, 10, -2, 1, -5, 5, 4, -7,
					-- layer=2 filter=33 channel=45
					-3, -10, -1, 1, -6, 7, 3, 4, -11,
					-- layer=2 filter=33 channel=46
					-6, -4, -8, 0, 0, -8, -5, 7, 6,
					-- layer=2 filter=33 channel=47
					-6, 1, 0, -11, -7, 1, -4, 0, -9,
					-- layer=2 filter=33 channel=48
					-6, 8, -4, -2, -5, -5, 4, -6, -7,
					-- layer=2 filter=33 channel=49
					-11, 8, -2, -11, 2, -8, -4, -1, -1,
					-- layer=2 filter=33 channel=50
					1, 6, -6, 8, 7, -2, -6, 8, -6,
					-- layer=2 filter=33 channel=51
					-5, 6, 0, -7, -3, 3, -5, -3, -8,
					-- layer=2 filter=33 channel=52
					0, -7, 3, -12, -2, -7, 1, 0, -9,
					-- layer=2 filter=33 channel=53
					0, 6, 8, -11, -2, 4, 1, -6, -8,
					-- layer=2 filter=33 channel=54
					-12, 8, -10, -10, -6, -9, -12, 1, -8,
					-- layer=2 filter=33 channel=55
					4, 9, -1, 4, 7, 6, 0, -6, -1,
					-- layer=2 filter=33 channel=56
					-11, 0, -9, -4, 8, -3, 1, 8, 0,
					-- layer=2 filter=33 channel=57
					-7, 4, 5, 0, 5, -8, 4, -9, 1,
					-- layer=2 filter=33 channel=58
					1, -2, 4, -5, -11, 5, -4, 0, -2,
					-- layer=2 filter=33 channel=59
					-2, -5, 5, -12, -5, 0, -10, -7, 8,
					-- layer=2 filter=33 channel=60
					1, 1, 2, 1, 0, -3, 6, -2, 0,
					-- layer=2 filter=33 channel=61
					-2, -9, -3, -1, -1, 7, -7, -6, -8,
					-- layer=2 filter=33 channel=62
					0, 9, 7, 5, 6, 2, 4, 8, -2,
					-- layer=2 filter=33 channel=63
					4, -8, -3, -2, -9, -11, 7, 0, 0,
					-- layer=2 filter=33 channel=64
					-6, 5, -10, 2, -8, -3, -6, -1, -6,
					-- layer=2 filter=33 channel=65
					2, 6, -10, 0, 0, -6, -4, -9, -6,
					-- layer=2 filter=33 channel=66
					-10, 8, 1, -10, 8, 4, -5, 5, 1,
					-- layer=2 filter=33 channel=67
					-10, 0, 5, 0, -8, -3, 2, 0, 0,
					-- layer=2 filter=33 channel=68
					3, -4, 0, 6, -2, -5, -10, -1, 5,
					-- layer=2 filter=33 channel=69
					-6, -6, 2, 6, 6, -4, -9, -4, -8,
					-- layer=2 filter=33 channel=70
					-3, -5, -9, 6, -7, 1, 0, -5, 0,
					-- layer=2 filter=33 channel=71
					0, -7, -5, 3, -6, -10, -4, -4, 0,
					-- layer=2 filter=33 channel=72
					-6, 7, -4, -11, -9, -2, -3, -11, -2,
					-- layer=2 filter=33 channel=73
					-5, 8, 3, -5, 9, 0, 1, -2, 4,
					-- layer=2 filter=33 channel=74
					0, 8, -4, -5, -10, 2, -8, -1, 2,
					-- layer=2 filter=33 channel=75
					8, 5, 6, 5, 8, -8, -2, -4, 1,
					-- layer=2 filter=33 channel=76
					-3, -3, 4, -11, 7, 1, 5, -11, -13,
					-- layer=2 filter=33 channel=77
					-1, -5, 0, 7, -5, -3, -4, 6, 4,
					-- layer=2 filter=33 channel=78
					4, -2, -1, 6, -7, -5, 6, 7, -11,
					-- layer=2 filter=33 channel=79
					5, 8, -1, 3, 7, -1, -2, 6, -3,
					-- layer=2 filter=33 channel=80
					-5, 3, -5, 0, -12, -1, -8, -7, -11,
					-- layer=2 filter=33 channel=81
					0, 4, 4, 1, -11, 6, -7, -1, -4,
					-- layer=2 filter=33 channel=82
					3, -6, 3, 7, -5, 7, -9, -9, 0,
					-- layer=2 filter=33 channel=83
					6, -6, 3, 2, 0, -9, 0, 6, -6,
					-- layer=2 filter=33 channel=84
					3, 0, 0, 11, 4, 5, 7, -3, 6,
					-- layer=2 filter=33 channel=85
					1, -7, -1, -7, 0, 0, 1, 4, 6,
					-- layer=2 filter=33 channel=86
					-11, 9, 9, 9, -5, 0, 4, 6, 8,
					-- layer=2 filter=33 channel=87
					6, -7, 8, 3, -6, 3, 8, -10, -4,
					-- layer=2 filter=33 channel=88
					-2, -8, 6, -10, -4, -11, -8, -1, -3,
					-- layer=2 filter=33 channel=89
					-8, 9, -5, -4, 9, 7, -4, 9, 3,
					-- layer=2 filter=33 channel=90
					-7, 8, -5, 1, 6, 0, -5, 0, 8,
					-- layer=2 filter=33 channel=91
					-13, -16, -9, -8, -7, 1, -5, 4, 1,
					-- layer=2 filter=33 channel=92
					0, -2, -7, -8, -11, 4, -6, -7, -8,
					-- layer=2 filter=33 channel=93
					-3, -8, 8, 7, -8, 7, 2, 1, -8,
					-- layer=2 filter=33 channel=94
					-16, -3, -6, -7, 2, -6, 4, 1, -10,
					-- layer=2 filter=33 channel=95
					-6, 4, -6, 5, 3, -3, 5, -2, -5,
					-- layer=2 filter=33 channel=96
					3, -5, -1, -6, -1, 0, 0, 1, 0,
					-- layer=2 filter=33 channel=97
					0, 1, 7, -10, -6, -4, 7, -3, -8,
					-- layer=2 filter=33 channel=98
					-2, -8, -4, 3, -2, -7, -3, 0, -8,
					-- layer=2 filter=33 channel=99
					7, 6, 7, -15, -2, -7, -11, -11, 3,
					-- layer=2 filter=33 channel=100
					-6, 4, 4, 8, -1, 8, 0, 0, -4,
					-- layer=2 filter=33 channel=101
					-9, 0, -2, -2, -13, 10, -5, 0, 7,
					-- layer=2 filter=33 channel=102
					-8, -10, -4, 2, 7, -8, 7, 6, 5,
					-- layer=2 filter=33 channel=103
					-8, -1, -10, -9, 0, 6, -4, 3, -5,
					-- layer=2 filter=33 channel=104
					0, -1, -7, 0, 2, -7, 7, 0, -11,
					-- layer=2 filter=33 channel=105
					-5, -2, -8, -5, 4, 6, 2, 8, 5,
					-- layer=2 filter=33 channel=106
					-3, -8, 3, 8, 1, -4, 2, 2, 3,
					-- layer=2 filter=33 channel=107
					-3, 0, -8, 2, 3, 6, 11, -5, 7,
					-- layer=2 filter=33 channel=108
					-2, -4, -4, -5, 7, -1, -10, 0, -7,
					-- layer=2 filter=33 channel=109
					-2, 6, -1, 2, 7, 5, 1, 7, -4,
					-- layer=2 filter=33 channel=110
					2, -4, -5, -8, 6, 0, -2, -10, -11,
					-- layer=2 filter=33 channel=111
					-6, 1, 6, -8, 9, 6, 1, 6, -9,
					-- layer=2 filter=33 channel=112
					8, -9, 0, -5, 0, -5, 0, -11, -9,
					-- layer=2 filter=33 channel=113
					4, 1, -4, 8, 1, 2, -3, -11, -5,
					-- layer=2 filter=33 channel=114
					4, 8, -7, 1, -3, 0, 0, -3, -2,
					-- layer=2 filter=33 channel=115
					9, 5, -8, -2, 5, 3, -6, -9, -10,
					-- layer=2 filter=33 channel=116
					-7, 4, -5, -4, -7, -7, 5, -4, -1,
					-- layer=2 filter=33 channel=117
					-5, -2, 2, 0, 4, -11, 6, 6, 4,
					-- layer=2 filter=33 channel=118
					-12, 2, -10, 0, 0, 3, 2, -10, 3,
					-- layer=2 filter=33 channel=119
					0, -1, 6, 1, -4, -5, 4, 0, 4,
					-- layer=2 filter=33 channel=120
					4, 1, 0, 3, 0, 6, 1, 0, 0,
					-- layer=2 filter=33 channel=121
					-1, 4, 5, 3, -5, 4, 4, 3, -2,
					-- layer=2 filter=33 channel=122
					9, -4, -8, 7, 3, -11, 7, 0, 2,
					-- layer=2 filter=33 channel=123
					5, -4, 0, -12, -15, -6, 10, -8, -1,
					-- layer=2 filter=33 channel=124
					0, -9, 2, -7, 8, 5, -5, -1, -2,
					-- layer=2 filter=33 channel=125
					7, -4, -6, 6, 1, -9, -2, 7, -10,
					-- layer=2 filter=33 channel=126
					4, 1, 2, -1, -12, -9, 0, -5, 0,
					-- layer=2 filter=33 channel=127
					2, 5, -10, -10, -7, -6, -1, 0, 2,
					-- layer=2 filter=34 channel=0
					-5, -8, 4, -2, -3, -4, -3, -1, -2,
					-- layer=2 filter=34 channel=1
					-21, -2, -20, -16, -12, 1, 7, -10, 0,
					-- layer=2 filter=34 channel=2
					4, -2, 4, 7, 5, 7, -2, -10, 4,
					-- layer=2 filter=34 channel=3
					-10, 1, 15, -12, -8, -1, 6, 2, 6,
					-- layer=2 filter=34 channel=4
					-25, -10, 15, -13, 4, 10, -1, -6, -3,
					-- layer=2 filter=34 channel=5
					-18, -10, -11, -10, -17, 7, -17, -21, -3,
					-- layer=2 filter=34 channel=6
					17, -28, -16, -23, -19, 2, -26, -34, 0,
					-- layer=2 filter=34 channel=7
					9, 6, -11, 15, 0, -11, -22, -1, -9,
					-- layer=2 filter=34 channel=8
					0, 5, 4, 8, -9, 2, -6, 9, 5,
					-- layer=2 filter=34 channel=9
					-12, -7, 0, -6, -17, -3, 0, -5, -2,
					-- layer=2 filter=34 channel=10
					-13, -11, 4, -18, 4, -10, -8, -3, -15,
					-- layer=2 filter=34 channel=11
					-3, -16, 0, -1, -4, -11, -6, -5, -7,
					-- layer=2 filter=34 channel=12
					-4, -20, -19, -8, -17, -9, -25, -14, -4,
					-- layer=2 filter=34 channel=13
					-7, 7, 4, 4, -3, -9, 2, 6, 4,
					-- layer=2 filter=34 channel=14
					1, -18, -4, -9, -15, -1, -2, -10, -7,
					-- layer=2 filter=34 channel=15
					-4, 9, -6, 22, -4, -13, 0, -7, 6,
					-- layer=2 filter=34 channel=16
					-20, -18, -3, -19, -32, -12, -16, -12, -3,
					-- layer=2 filter=34 channel=17
					0, -7, 8, -5, -7, 4, -11, 9, -5,
					-- layer=2 filter=34 channel=18
					3, -21, 7, 5, -4, -21, 17, -23, 2,
					-- layer=2 filter=34 channel=19
					-35, -24, -9, -12, -1, -3, -12, -13, -22,
					-- layer=2 filter=34 channel=20
					4, 5, 5, 0, 2, -5, 3, -5, -4,
					-- layer=2 filter=34 channel=21
					8, 11, 3, -4, -4, 4, -7, -2, -3,
					-- layer=2 filter=34 channel=22
					-1, -4, 9, 8, 0, -1, 9, 1, -7,
					-- layer=2 filter=34 channel=23
					-8, -7, 11, -28, -7, -12, -5, -5, -12,
					-- layer=2 filter=34 channel=24
					-22, -11, 8, -26, -11, -17, 4, 0, -7,
					-- layer=2 filter=34 channel=25
					-39, -23, -8, -13, -15, -7, -5, -19, -36,
					-- layer=2 filter=34 channel=26
					8, 2, 0, 1, -2, 2, 6, -4, -3,
					-- layer=2 filter=34 channel=27
					5, 0, -1, -3, -17, -26, -22, -7, -7,
					-- layer=2 filter=34 channel=28
					-19, -9, 17, 5, -6, 21, 0, -20, -5,
					-- layer=2 filter=34 channel=29
					7, 2, -5, 7, -7, -4, 9, 2, -3,
					-- layer=2 filter=34 channel=30
					-5, -6, -2, -11, -6, -9, 2, -11, -16,
					-- layer=2 filter=34 channel=31
					0, 0, 6, 10, -4, -2, 3, 5, 1,
					-- layer=2 filter=34 channel=32
					-4, -7, 9, 3, 1, 3, 7, 4, -2,
					-- layer=2 filter=34 channel=33
					0, 0, -18, 9, -18, -13, -14, -12, 0,
					-- layer=2 filter=34 channel=34
					11, -6, -2, 29, 6, 19, 16, -15, 9,
					-- layer=2 filter=34 channel=35
					-6, -9, 34, -4, -6, 25, 14, -6, -15,
					-- layer=2 filter=34 channel=36
					8, 3, -5, 5, 10, 1, 0, 7, -1,
					-- layer=2 filter=34 channel=37
					0, -9, -16, -2, -8, -20, -15, -3, -18,
					-- layer=2 filter=34 channel=38
					-8, 8, -39, -22, -21, -19, -23, -13, -7,
					-- layer=2 filter=34 channel=39
					-4, -10, -6, -23, -11, -8, -15, -14, -5,
					-- layer=2 filter=34 channel=40
					-22, -6, 10, -7, -2, -6, 7, -15, 0,
					-- layer=2 filter=34 channel=41
					-7, -9, -3, 1, 3, 0, 0, -4, -1,
					-- layer=2 filter=34 channel=42
					-16, -1, -13, -15, -5, 3, -1, 8, -9,
					-- layer=2 filter=34 channel=43
					-11, -10, 3, 20, 8, 12, 12, -29, -19,
					-- layer=2 filter=34 channel=44
					-3, -2, -6, -3, 0, 5, -8, 4, 10,
					-- layer=2 filter=34 channel=45
					19, 16, -22, 5, -7, -8, -4, -6, 2,
					-- layer=2 filter=34 channel=46
					11, -3, 1, 2, -5, -1, -8, 12, -13,
					-- layer=2 filter=34 channel=47
					-20, -30, -15, 1, -5, 7, -30, -29, 0,
					-- layer=2 filter=34 channel=48
					5, 6, 11, -4, 2, 8, 9, -2, 7,
					-- layer=2 filter=34 channel=49
					13, -32, -7, 8, -30, -7, 6, -25, -15,
					-- layer=2 filter=34 channel=50
					0, 9, 1, 7, -3, 5, 3, 5, -10,
					-- layer=2 filter=34 channel=51
					-14, -10, -19, -6, -28, -14, -10, -9, -20,
					-- layer=2 filter=34 channel=52
					-8, -18, 13, -14, -13, -4, -8, 8, -19,
					-- layer=2 filter=34 channel=53
					3, 17, 12, 0, 2, -6, 2, -13, -3,
					-- layer=2 filter=34 channel=54
					-10, -13, 13, -31, -18, -8, -27, -17, -26,
					-- layer=2 filter=34 channel=55
					7, 8, 2, 7, 1, 0, -2, 5, -7,
					-- layer=2 filter=34 channel=56
					4, -11, 6, -10, -9, 0, -16, -13, -18,
					-- layer=2 filter=34 channel=57
					6, 3, -3, -8, -4, -9, -9, 8, -1,
					-- layer=2 filter=34 channel=58
					-19, -12, -1, 0, 0, -21, -13, -8, -17,
					-- layer=2 filter=34 channel=59
					0, -4, -8, -20, -11, -35, -17, -26, -6,
					-- layer=2 filter=34 channel=60
					1, 10, -15, -19, -13, -6, -16, -13, -26,
					-- layer=2 filter=34 channel=61
					4, 1, 2, -13, -12, -5, -2, -39, -8,
					-- layer=2 filter=34 channel=62
					25, -20, -1, 15, -13, 10, 3, -25, -6,
					-- layer=2 filter=34 channel=63
					11, -4, 0, -1, 4, 0, -11, 1, -15,
					-- layer=2 filter=34 channel=64
					-15, -5, -6, -11, -23, -11, 8, -19, 0,
					-- layer=2 filter=34 channel=65
					8, 7, -11, -21, -6, -16, -5, -19, 7,
					-- layer=2 filter=34 channel=66
					0, -11, -15, 5, 1, -2, 4, -3, -6,
					-- layer=2 filter=34 channel=67
					-8, -8, -17, -1, -11, -6, -16, 2, -4,
					-- layer=2 filter=34 channel=68
					-6, -9, -8, -3, 4, 9, 0, 5, 0,
					-- layer=2 filter=34 channel=69
					-15, -2, -7, -4, -15, -8, -12, -1, 0,
					-- layer=2 filter=34 channel=70
					-29, -2, 36, -5, -1, 28, -8, -1, -10,
					-- layer=2 filter=34 channel=71
					8, 13, -22, 0, 0, -5, 3, 12, 3,
					-- layer=2 filter=34 channel=72
					-19, -29, -22, -11, 12, 23, -9, -12, -6,
					-- layer=2 filter=34 channel=73
					8, 1, -11, -4, 2, -10, -6, 2, -1,
					-- layer=2 filter=34 channel=74
					-11, -3, -20, -14, 1, -10, -4, 17, 5,
					-- layer=2 filter=34 channel=75
					-6, -18, 3, 1, -5, -12, 0, 3, -6,
					-- layer=2 filter=34 channel=76
					-2, 13, 29, -1, -11, -21, -8, -14, -25,
					-- layer=2 filter=34 channel=77
					-4, 8, -8, 1, 2, -9, 6, 2, 3,
					-- layer=2 filter=34 channel=78
					5, 2, -2, -4, -18, 4, -4, -9, -6,
					-- layer=2 filter=34 channel=79
					-10, 0, -4, 7, -3, 8, 3, -7, -4,
					-- layer=2 filter=34 channel=80
					-1, -12, -8, -21, -18, -1, 0, -6, 7,
					-- layer=2 filter=34 channel=81
					9, -6, -3, -1, 4, -2, 9, -3, 11,
					-- layer=2 filter=34 channel=82
					-8, 1, -2, 5, 0, 0, -9, -5, -4,
					-- layer=2 filter=34 channel=83
					-2, 10, 14, -19, -3, -1, -17, -12, 0,
					-- layer=2 filter=34 channel=84
					-5, 9, 10, 6, -4, -8, 11, 0, -6,
					-- layer=2 filter=34 channel=85
					-2, -10, 4, 1, 5, -8, -3, 0, -4,
					-- layer=2 filter=34 channel=86
					-11, -6, 4, -3, 3, 0, 3, -6, -9,
					-- layer=2 filter=34 channel=87
					-46, -15, 33, -29, 0, -20, -10, -19, 1,
					-- layer=2 filter=34 channel=88
					-21, -13, -19, 0, -10, -7, -19, -19, -6,
					-- layer=2 filter=34 channel=89
					-16, -31, -8, -21, -7, -5, -16, -12, -25,
					-- layer=2 filter=34 channel=90
					0, -2, -4, 0, -5, -4, 3, -6, 9,
					-- layer=2 filter=34 channel=91
					-5, -11, -6, -5, -12, 2, -5, -4, -30,
					-- layer=2 filter=34 channel=92
					-36, -8, -40, -7, -12, -15, 9, -20, -24,
					-- layer=2 filter=34 channel=93
					-6, -5, -20, -1, -10, -28, 11, -9, -5,
					-- layer=2 filter=34 channel=94
					11, -7, 20, -9, -32, 11, -14, -22, -12,
					-- layer=2 filter=34 channel=95
					4, -4, -10, 5, 9, -1, 3, -5, -2,
					-- layer=2 filter=34 channel=96
					-39, 5, 37, -25, -4, 0, -27, -18, 3,
					-- layer=2 filter=34 channel=97
					-16, -7, -10, -24, -8, -15, -16, -10, 10,
					-- layer=2 filter=34 channel=98
					1, -33, 22, -4, -30, -4, -26, -29, -17,
					-- layer=2 filter=34 channel=99
					12, -20, -12, -1, 5, -3, -3, 4, -32,
					-- layer=2 filter=34 channel=100
					-15, 0, -1, -8, -6, 7, -13, 2, 8,
					-- layer=2 filter=34 channel=101
					11, 9, 4, 0, -17, -4, 11, 0, -6,
					-- layer=2 filter=34 channel=102
					-30, -11, 31, -17, -34, -17, -3, -29, -17,
					-- layer=2 filter=34 channel=103
					-13, 1, 7, -10, 7, 3, 4, -2, -5,
					-- layer=2 filter=34 channel=104
					-21, 9, 9, -20, -18, 8, -3, -26, -9,
					-- layer=2 filter=34 channel=105
					3, -2, -7, -2, -2, -13, 5, 3, -3,
					-- layer=2 filter=34 channel=106
					-16, -9, -17, -12, -22, -26, -18, -16, -6,
					-- layer=2 filter=34 channel=107
					0, 0, -7, -16, -1, 9, 6, -1, 2,
					-- layer=2 filter=34 channel=108
					24, 13, -5, -1, -32, -18, 14, -5, -8,
					-- layer=2 filter=34 channel=109
					-8, 2, 8, -2, 4, 10, -6, 6, -4,
					-- layer=2 filter=34 channel=110
					-17, -24, -15, -15, -20, -19, -3, -17, -18,
					-- layer=2 filter=34 channel=111
					11, 1, -4, -1, -6, -8, 9, -6, 0,
					-- layer=2 filter=34 channel=112
					0, -7, -15, -21, -24, -24, -11, -26, -40,
					-- layer=2 filter=34 channel=113
					0, -6, -8, -1, -10, -5, -3, 1, -21,
					-- layer=2 filter=34 channel=114
					7, 0, 11, 10, -1, -9, -8, 8, -5,
					-- layer=2 filter=34 channel=115
					-8, 3, 7, -1, 0, -3, 4, 9, 4,
					-- layer=2 filter=34 channel=116
					-15, -9, 25, -18, -8, -13, -2, -8, -10,
					-- layer=2 filter=34 channel=117
					-14, -45, -19, -12, -15, -11, -17, -15, -7,
					-- layer=2 filter=34 channel=118
					-2, -14, -18, -12, -4, -3, 1, 2, 18,
					-- layer=2 filter=34 channel=119
					2, -19, 8, 6, -10, 14, -1, -22, -5,
					-- layer=2 filter=34 channel=120
					3, 0, -3, -2, 6, 7, -9, 5, -7,
					-- layer=2 filter=34 channel=121
					2, -12, 1, 0, -1, 9, 7, 6, 4,
					-- layer=2 filter=34 channel=122
					0, -3, -3, 10, 2, 1, 0, 0, 10,
					-- layer=2 filter=34 channel=123
					-34, -37, -4, -8, -3, -1, -18, -9, -17,
					-- layer=2 filter=34 channel=124
					-24, 5, -26, -11, -8, -18, -12, 1, -18,
					-- layer=2 filter=34 channel=125
					4, -11, 0, 4, -10, 0, 0, 2, -1,
					-- layer=2 filter=34 channel=126
					0, 4, 18, -12, -11, -21, 0, -13, -17,
					-- layer=2 filter=34 channel=127
					-2, 4, 6, -10, -7, -8, -11, -4, 9,
					-- layer=2 filter=35 channel=0
					-12, -6, -9, -17, -4, -7, -9, 4, -1,
					-- layer=2 filter=35 channel=1
					-8, 4, -3, -12, 0, -20, -17, -6, -9,
					-- layer=2 filter=35 channel=2
					-8, 2, 8, -11, 7, -9, 4, 2, 1,
					-- layer=2 filter=35 channel=3
					-1, -28, -16, -9, -14, -9, -6, 9, 13,
					-- layer=2 filter=35 channel=4
					6, -31, -11, -18, -22, -18, -10, -14, -16,
					-- layer=2 filter=35 channel=5
					-18, -3, -3, -3, -4, -4, -18, -4, -8,
					-- layer=2 filter=35 channel=6
					-14, -8, 19, -18, 2, 1, -7, 5, -11,
					-- layer=2 filter=35 channel=7
					7, -21, -8, -3, -10, 5, 11, 8, 11,
					-- layer=2 filter=35 channel=8
					-8, -8, 2, 0, 11, 9, -3, -8, -2,
					-- layer=2 filter=35 channel=9
					6, -20, -34, -11, -24, -23, -9, -22, -31,
					-- layer=2 filter=35 channel=10
					15, -2, -16, -23, -12, 0, 4, 2, 11,
					-- layer=2 filter=35 channel=11
					-13, -10, -8, 0, 0, -4, 11, -13, 0,
					-- layer=2 filter=35 channel=12
					1, -3, -7, 8, -14, -6, -7, -14, -7,
					-- layer=2 filter=35 channel=13
					-2, -7, -1, -9, 9, 9, 6, -5, 0,
					-- layer=2 filter=35 channel=14
					-12, -11, -22, -15, -15, -12, -5, -17, -24,
					-- layer=2 filter=35 channel=15
					-15, -17, 1, -10, 7, -2, -19, -11, -19,
					-- layer=2 filter=35 channel=16
					-14, -14, -25, -10, -11, -5, 3, 6, 8,
					-- layer=2 filter=35 channel=17
					2, 8, -9, 10, 4, -6, -6, 10, -7,
					-- layer=2 filter=35 channel=18
					3, -22, 1, -22, -38, -12, 6, -18, -21,
					-- layer=2 filter=35 channel=19
					4, 15, 7, 3, 10, 10, -14, 0, -15,
					-- layer=2 filter=35 channel=20
					6, 3, -10, -10, -1, -2, 0, -5, -3,
					-- layer=2 filter=35 channel=21
					2, -5, 8, -11, 3, -3, 7, 9, -4,
					-- layer=2 filter=35 channel=22
					-7, 3, 3, -2, 1, 3, -6, -3, 8,
					-- layer=2 filter=35 channel=23
					-28, -5, -23, -16, -10, -11, -5, -8, 4,
					-- layer=2 filter=35 channel=24
					-12, -12, -4, -5, -25, -22, -2, 0, -5,
					-- layer=2 filter=35 channel=25
					-20, -27, -29, -16, -28, -20, 9, -8, -6,
					-- layer=2 filter=35 channel=26
					6, 4, -2, 2, -2, 1, 10, 0, -10,
					-- layer=2 filter=35 channel=27
					3, 1, -3, -11, -11, -15, -10, -12, -3,
					-- layer=2 filter=35 channel=28
					-3, -12, -12, -14, -6, -11, 10, 0, 12,
					-- layer=2 filter=35 channel=29
					-11, -12, -6, 0, -9, 1, -12, -7, -4,
					-- layer=2 filter=35 channel=30
					6, -19, -33, 0, -18, -12, 1, -17, -28,
					-- layer=2 filter=35 channel=31
					3, -5, 7, -5, -10, -13, -23, -2, -14,
					-- layer=2 filter=35 channel=32
					0, -8, -4, -3, 0, 1, 4, 0, 2,
					-- layer=2 filter=35 channel=33
					-13, -8, -20, -21, -23, -17, 11, -3, 8,
					-- layer=2 filter=35 channel=34
					-2, -7, -16, -25, -20, -10, 0, -2, -8,
					-- layer=2 filter=35 channel=35
					27, -5, -5, 6, 0, 11, -1, -2, 12,
					-- layer=2 filter=35 channel=36
					-8, 0, 1, -7, -10, -11, 5, -2, -5,
					-- layer=2 filter=35 channel=37
					-11, -19, -21, -22, -10, -4, -16, -18, -16,
					-- layer=2 filter=35 channel=38
					-20, -6, -13, -20, -20, -25, -26, -3, -10,
					-- layer=2 filter=35 channel=39
					-33, -10, -11, -7, -18, -20, -7, -1, 9,
					-- layer=2 filter=35 channel=40
					-7, -12, 0, -5, -16, 12, 15, -11, 11,
					-- layer=2 filter=35 channel=41
					4, -10, -9, 4, -9, 0, -2, -2, -1,
					-- layer=2 filter=35 channel=42
					-23, -23, 0, -12, -18, -13, -15, -6, 7,
					-- layer=2 filter=35 channel=43
					3, -26, -25, -18, -31, -15, -8, -7, -7,
					-- layer=2 filter=35 channel=44
					-9, 1, -5, 10, -10, -6, 3, -9, 4,
					-- layer=2 filter=35 channel=45
					-9, -7, -7, -8, -20, -19, -20, -3, 0,
					-- layer=2 filter=35 channel=46
					-2, -7, -8, -14, -16, -33, -35, -15, -26,
					-- layer=2 filter=35 channel=47
					-18, 0, -33, 0, -2, -8, 5, -11, 12,
					-- layer=2 filter=35 channel=48
					-3, -4, 9, 2, 0, 7, -5, -9, 1,
					-- layer=2 filter=35 channel=49
					0, -19, -7, -17, -20, -19, -14, -17, -32,
					-- layer=2 filter=35 channel=50
					6, 3, 2, -9, -9, -12, 0, 3, 9,
					-- layer=2 filter=35 channel=51
					-1, -3, -10, 3, -11, -14, -12, 0, -12,
					-- layer=2 filter=35 channel=52
					-15, -8, -15, -14, -13, 21, 20, -5, 1,
					-- layer=2 filter=35 channel=53
					0, -2, -7, -6, 4, 2, -1, -10, -14,
					-- layer=2 filter=35 channel=54
					0, -17, -23, -4, -21, -11, 4, 10, -5,
					-- layer=2 filter=35 channel=55
					0, -8, -8, -6, -7, 4, 6, 1, 2,
					-- layer=2 filter=35 channel=56
					-3, -2, -9, -10, 2, -10, -9, -11, -10,
					-- layer=2 filter=35 channel=57
					-6, 5, 7, -2, -7, -2, -5, -3, -8,
					-- layer=2 filter=35 channel=58
					-16, 2, -21, 0, -3, -6, -21, -21, -28,
					-- layer=2 filter=35 channel=59
					-20, 22, -15, -26, -2, -5, -25, -1, -11,
					-- layer=2 filter=35 channel=60
					-28, 13, -15, -1, 9, -5, -2, 4, -29,
					-- layer=2 filter=35 channel=61
					-23, 0, -19, -20, 19, 1, -7, 23, -13,
					-- layer=2 filter=35 channel=62
					-18, -8, 19, -16, 15, -4, 5, 9, -11,
					-- layer=2 filter=35 channel=63
					-42, 6, -19, -14, 9, 5, -15, 15, -9,
					-- layer=2 filter=35 channel=64
					-12, -12, -31, 0, -15, -10, -12, -14, -6,
					-- layer=2 filter=35 channel=65
					-20, 4, 2, -14, 1, -7, 7, 4, -10,
					-- layer=2 filter=35 channel=66
					5, 3, -4, -4, 0, 3, 1, 0, -10,
					-- layer=2 filter=35 channel=67
					-16, -14, -7, -28, -24, -8, -15, -19, -15,
					-- layer=2 filter=35 channel=68
					-6, 4, 7, 2, -9, 0, 4, -5, -3,
					-- layer=2 filter=35 channel=69
					-41, -26, -22, -5, -9, -16, -15, -31, -10,
					-- layer=2 filter=35 channel=70
					12, -10, -18, -7, -1, 0, 15, 9, 4,
					-- layer=2 filter=35 channel=71
					3, 7, -2, 5, -11, -3, -22, -6, -14,
					-- layer=2 filter=35 channel=72
					-10, -4, -1, -6, -22, -14, 5, -1, -8,
					-- layer=2 filter=35 channel=73
					-9, 1, 0, -13, 0, 3, -34, 8, -22,
					-- layer=2 filter=35 channel=74
					-19, 7, -18, -4, -19, -11, -13, -31, -25,
					-- layer=2 filter=35 channel=75
					2, 0, -16, 4, -13, -1, -2, -1, -14,
					-- layer=2 filter=35 channel=76
					9, 3, -17, -4, 3, 11, -20, 11, -19,
					-- layer=2 filter=35 channel=77
					-5, 5, -2, -5, 0, -8, -1, -10, -6,
					-- layer=2 filter=35 channel=78
					0, -22, -10, -20, -11, -4, 12, 13, -3,
					-- layer=2 filter=35 channel=79
					-11, -3, -5, -11, -10, 7, -10, -10, -12,
					-- layer=2 filter=35 channel=80
					-5, -21, -37, -36, -27, -18, -19, -17, -4,
					-- layer=2 filter=35 channel=81
					-8, -4, -7, 5, 0, 5, 0, -12, -11,
					-- layer=2 filter=35 channel=82
					-3, -7, 0, 1, -11, 4, 5, -10, -6,
					-- layer=2 filter=35 channel=83
					4, -6, -9, -4, -10, -14, -10, -6, -6,
					-- layer=2 filter=35 channel=84
					-5, 5, 10, 11, 5, 4, -6, -5, 7,
					-- layer=2 filter=35 channel=85
					2, -5, 2, -1, 8, 9, -3, 1, 6,
					-- layer=2 filter=35 channel=86
					10, 4, 0, 4, -8, -4, 0, -6, 10,
					-- layer=2 filter=35 channel=87
					-2, -21, -8, -17, 4, 0, 18, -20, 6,
					-- layer=2 filter=35 channel=88
					-18, 9, -31, 4, -3, 11, -28, -10, -24,
					-- layer=2 filter=35 channel=89
					-9, -1, -4, 20, 5, -12, -4, -6, -25,
					-- layer=2 filter=35 channel=90
					3, 3, -1, 3, -4, -9, 0, -5, -5,
					-- layer=2 filter=35 channel=91
					-10, 3, -1, 13, 8, 15, -6, -12, -28,
					-- layer=2 filter=35 channel=92
					2, 24, 2, 9, -16, -13, -26, -16, -20,
					-- layer=2 filter=35 channel=93
					-9, -1, 7, -15, -4, -8, -8, -18, -11,
					-- layer=2 filter=35 channel=94
					-14, -9, 5, -16, 4, 22, -7, 25, 0,
					-- layer=2 filter=35 channel=95
					-9, -2, -10, 2, -7, -4, 3, -2, 6,
					-- layer=2 filter=35 channel=96
					0, 13, -18, -4, 17, -10, -21, -3, -6,
					-- layer=2 filter=35 channel=97
					-12, -28, -24, -30, -12, -23, -23, -15, -8,
					-- layer=2 filter=35 channel=98
					-16, -28, -22, -9, -16, -2, 16, 0, -3,
					-- layer=2 filter=35 channel=99
					-17, -18, -20, 1, 17, 0, -15, 12, -18,
					-- layer=2 filter=35 channel=100
					9, 6, -10, -8, -8, -20, -30, 6, -13,
					-- layer=2 filter=35 channel=101
					11, 1, -20, 0, -7, -10, -1, -13, -11,
					-- layer=2 filter=35 channel=102
					-3, 1, -16, -11, 13, -28, 0, -13, -6,
					-- layer=2 filter=35 channel=103
					9, -2, 7, -7, -4, 7, 3, -12, -7,
					-- layer=2 filter=35 channel=104
					-20, -11, 4, 5, -7, -7, -5, -4, -17,
					-- layer=2 filter=35 channel=105
					14, 12, 0, -4, 21, 11, 6, -16, -17,
					-- layer=2 filter=35 channel=106
					-15, -29, -30, -17, 0, -11, -8, -22, -3,
					-- layer=2 filter=35 channel=107
					-1, 4, 18, 16, 15, 11, -8, 7, 7,
					-- layer=2 filter=35 channel=108
					-8, 4, -1, -15, -4, -10, -1, -13, -20,
					-- layer=2 filter=35 channel=109
					4, 7, -12, 0, -6, -3, -7, -1, -3,
					-- layer=2 filter=35 channel=110
					-16, -1, -15, 18, -7, -9, -1, -13, -23,
					-- layer=2 filter=35 channel=111
					5, 7, -7, 4, 7, 2, 4, 9, -6,
					-- layer=2 filter=35 channel=112
					-16, -10, -21, -15, -11, -5, -5, 3, 0,
					-- layer=2 filter=35 channel=113
					-6, 3, -35, 7, -10, -14, 10, -11, -28,
					-- layer=2 filter=35 channel=114
					-8, -3, 3, -5, -6, 5, -6, 5, 6,
					-- layer=2 filter=35 channel=115
					7, 4, 8, 7, 4, -10, -10, -4, 3,
					-- layer=2 filter=35 channel=116
					-3, -17, -12, -20, -1, -3, 21, -23, 12,
					-- layer=2 filter=35 channel=117
					17, -4, -2, 0, 0, -2, 3, 4, 0,
					-- layer=2 filter=35 channel=118
					-8, -22, -17, -22, -8, 5, -4, -6, 0,
					-- layer=2 filter=35 channel=119
					-8, -26, 1, -30, -29, -2, -9, -25, -18,
					-- layer=2 filter=35 channel=120
					4, 6, 1, 9, 2, 3, -4, 0, 7,
					-- layer=2 filter=35 channel=121
					-7, -7, -8, -7, -3, 6, -8, -5, 3,
					-- layer=2 filter=35 channel=122
					1, 5, -1, 9, -6, 0, -5, 2, -3,
					-- layer=2 filter=35 channel=123
					-27, -19, -27, -9, -10, 11, 36, 16, -2,
					-- layer=2 filter=35 channel=124
					-17, -15, -7, -10, -3, -11, -17, -13, -7,
					-- layer=2 filter=35 channel=125
					2, -2, -2, -3, 2, -7, -1, 9, 7,
					-- layer=2 filter=35 channel=126
					-20, -3, 11, -2, 8, 14, -22, -11, -7,
					-- layer=2 filter=35 channel=127
					-22, 10, -9, -6, -5, -27, -6, -6, -6,
					-- layer=2 filter=36 channel=0
					7, 4, 6, -10, -4, -8, -9, -9, -4,
					-- layer=2 filter=36 channel=1
					1, -12, -1, 10, 0, -8, 0, -9, 0,
					-- layer=2 filter=36 channel=2
					-5, 5, -1, -8, -4, 3, 3, -1, 10,
					-- layer=2 filter=36 channel=3
					-3, -11, 2, 9, 8, -6, 10, 1, 0,
					-- layer=2 filter=36 channel=4
					0, 2, -8, -9, 5, 0, -3, 8, 1,
					-- layer=2 filter=36 channel=5
					-12, -2, -9, -10, -6, -8, -9, -2, 7,
					-- layer=2 filter=36 channel=6
					7, 0, -12, -9, -5, -10, 7, -2, -3,
					-- layer=2 filter=36 channel=7
					6, -11, -12, 1, -7, 3, 6, -3, 7,
					-- layer=2 filter=36 channel=8
					-3, 4, -2, -4, 8, 2, -4, -10, 9,
					-- layer=2 filter=36 channel=9
					5, -3, 4, 0, 0, 3, -5, 2, 6,
					-- layer=2 filter=36 channel=10
					-2, 8, -10, 4, -6, 2, -7, 2, -9,
					-- layer=2 filter=36 channel=11
					0, -3, -7, 9, -13, -3, 0, -9, -7,
					-- layer=2 filter=36 channel=12
					0, -3, 1, -1, -3, -5, 0, 0, -14,
					-- layer=2 filter=36 channel=13
					9, -6, -4, 8, 1, 7, 4, -6, -4,
					-- layer=2 filter=36 channel=14
					5, -6, 0, -9, -3, -4, -9, -13, 4,
					-- layer=2 filter=36 channel=15
					-4, 2, 4, -3, 0, -8, -4, 3, -8,
					-- layer=2 filter=36 channel=16
					-12, -8, -10, -1, 0, 2, -11, 1, 2,
					-- layer=2 filter=36 channel=17
					9, 4, 0, 1, 1, 6, -7, 5, 10,
					-- layer=2 filter=36 channel=18
					-3, 0, 3, 8, -3, 2, 2, -8, -3,
					-- layer=2 filter=36 channel=19
					-6, 11, 0, 1, 0, -6, 3, -6, 1,
					-- layer=2 filter=36 channel=20
					8, -4, 3, -2, 0, 1, -6, -1, 5,
					-- layer=2 filter=36 channel=21
					5, -2, 7, 5, 1, -1, -6, -4, 4,
					-- layer=2 filter=36 channel=22
					-9, 0, 5, -7, 5, -3, 4, 0, 0,
					-- layer=2 filter=36 channel=23
					-8, 3, -8, 7, -7, -1, -7, -7, 0,
					-- layer=2 filter=36 channel=24
					5, -15, -1, -9, 3, -13, -10, -7, 5,
					-- layer=2 filter=36 channel=25
					11, -6, -5, 2, -6, -10, 4, -8, 2,
					-- layer=2 filter=36 channel=26
					-8, -4, -1, 10, 8, -4, 0, 0, 3,
					-- layer=2 filter=36 channel=27
					-11, -2, -4, 2, 3, 2, 6, 6, -8,
					-- layer=2 filter=36 channel=28
					2, 8, -2, 3, -8, -6, -15, -7, -15,
					-- layer=2 filter=36 channel=29
					5, -5, -11, -8, 2, 2, 7, -10, -8,
					-- layer=2 filter=36 channel=30
					0, -10, -1, 9, -10, -6, -12, -1, -6,
					-- layer=2 filter=36 channel=31
					7, -10, -10, -8, 2, 0, -11, -6, 2,
					-- layer=2 filter=36 channel=32
					-3, -7, -1, 2, -2, 4, 0, 6, 6,
					-- layer=2 filter=36 channel=33
					-4, -10, -9, 6, 0, -14, -5, -6, 3,
					-- layer=2 filter=36 channel=34
					0, -7, 4, -11, -5, 1, -6, -10, -3,
					-- layer=2 filter=36 channel=35
					1, 6, 8, -6, -4, 4, -19, 0, -1,
					-- layer=2 filter=36 channel=36
					-5, -1, 2, -4, -10, -7, -8, -12, -3,
					-- layer=2 filter=36 channel=37
					2, 0, -6, 2, -4, -1, -6, -10, 0,
					-- layer=2 filter=36 channel=38
					-1, -5, -2, 0, 6, -6, -4, -9, 7,
					-- layer=2 filter=36 channel=39
					5, -10, -7, -11, -9, -10, 7, -2, -7,
					-- layer=2 filter=36 channel=40
					-4, -5, -1, -2, 0, 0, 5, -12, -13,
					-- layer=2 filter=36 channel=41
					5, -6, 4, -5, -9, -2, 2, 1, 7,
					-- layer=2 filter=36 channel=42
					6, 2, -10, 4, 3, 0, -16, 0, -4,
					-- layer=2 filter=36 channel=43
					0, -4, 4, -13, -5, -6, -8, 0, -1,
					-- layer=2 filter=36 channel=44
					-5, 0, 9, -3, 6, 6, -8, 0, -10,
					-- layer=2 filter=36 channel=45
					-8, 2, -8, -3, -6, 8, -6, -1, 7,
					-- layer=2 filter=36 channel=46
					0, -2, -10, 5, -4, -2, -5, 6, 0,
					-- layer=2 filter=36 channel=47
					-4, -7, 8, 3, 3, -12, 1, -2, -6,
					-- layer=2 filter=36 channel=48
					-1, -9, 8, -3, -7, 0, -1, 1, -3,
					-- layer=2 filter=36 channel=49
					-8, -1, -8, 1, -5, -5, -1, 6, -8,
					-- layer=2 filter=36 channel=50
					0, 0, -3, 0, -10, -10, 7, -1, 4,
					-- layer=2 filter=36 channel=51
					-11, -11, -16, 6, -9, -1, -10, -1, -8,
					-- layer=2 filter=36 channel=52
					0, 4, 9, 0, 3, -2, -7, -4, -5,
					-- layer=2 filter=36 channel=53
					-7, 11, 8, -4, -5, 2, 8, -8, -2,
					-- layer=2 filter=36 channel=54
					-3, 1, -7, -11, -5, -8, -5, 1, 4,
					-- layer=2 filter=36 channel=55
					-8, -5, 1, 2, 6, 10, 0, -9, 4,
					-- layer=2 filter=36 channel=56
					6, 9, 0, -5, 6, -11, 8, 1, 3,
					-- layer=2 filter=36 channel=57
					2, -5, -7, 4, -7, 3, 4, 8, 0,
					-- layer=2 filter=36 channel=58
					-6, -6, 0, 6, 4, -5, -6, 0, -1,
					-- layer=2 filter=36 channel=59
					5, -6, 12, 9, -5, -2, -4, 2, -4,
					-- layer=2 filter=36 channel=60
					2, 1, 0, -1, -6, 1, -6, -11, -9,
					-- layer=2 filter=36 channel=61
					3, -3, 3, -14, -15, 2, -11, -6, 0,
					-- layer=2 filter=36 channel=62
					-4, -4, 2, 4, 9, -2, 5, 1, -8,
					-- layer=2 filter=36 channel=63
					-10, -5, -11, -3, -5, -13, -2, 0, 2,
					-- layer=2 filter=36 channel=64
					0, -10, -1, 5, -1, -6, 1, -4, -9,
					-- layer=2 filter=36 channel=65
					-1, -7, 0, -3, -2, -3, -1, -9, -6,
					-- layer=2 filter=36 channel=66
					3, -10, 0, 8, -9, 5, -5, -3, -11,
					-- layer=2 filter=36 channel=67
					-8, -7, -5, -6, 0, 1, -6, -3, -7,
					-- layer=2 filter=36 channel=68
					4, -2, 1, -2, 3, 8, 2, 3, 1,
					-- layer=2 filter=36 channel=69
					0, -7, 6, -2, -6, 1, -1, 3, 1,
					-- layer=2 filter=36 channel=70
					-6, -7, -4, 1, 4, 2, -2, 0, 2,
					-- layer=2 filter=36 channel=71
					-2, 4, -10, -10, 4, -6, -1, -4, -9,
					-- layer=2 filter=36 channel=72
					-10, 1, -9, -12, 2, -15, -2, -11, -12,
					-- layer=2 filter=36 channel=73
					-2, 5, -6, -8, -6, -2, -6, -6, 6,
					-- layer=2 filter=36 channel=74
					0, -14, -3, 1, -7, 1, -7, 3, -3,
					-- layer=2 filter=36 channel=75
					2, -1, -2, 11, 6, -8, -14, -6, -2,
					-- layer=2 filter=36 channel=76
					-3, -2, -7, 0, -8, 7, -5, -11, 8,
					-- layer=2 filter=36 channel=77
					-3, 5, -3, -3, 6, -10, -5, 9, 7,
					-- layer=2 filter=36 channel=78
					-2, -11, 4, 3, 1, -5, 3, -2, -6,
					-- layer=2 filter=36 channel=79
					-5, 8, -5, -8, -2, -5, -9, 6, 7,
					-- layer=2 filter=36 channel=80
					6, -11, -9, 6, -3, -4, -3, -1, -4,
					-- layer=2 filter=36 channel=81
					-6, -3, 3, -3, -10, -1, 8, 4, -8,
					-- layer=2 filter=36 channel=82
					5, -10, -3, -10, -8, 3, -9, 4, -5,
					-- layer=2 filter=36 channel=83
					0, -5, 2, -12, 4, 0, -11, 0, -14,
					-- layer=2 filter=36 channel=84
					-7, 1, 6, 8, -4, 0, 2, -6, 11,
					-- layer=2 filter=36 channel=85
					6, 4, -6, 10, -3, 0, 0, -3, 0,
					-- layer=2 filter=36 channel=86
					-1, 7, 10, -4, -9, 6, 0, 8, -3,
					-- layer=2 filter=36 channel=87
					-12, -5, -8, -2, 1, -3, -6, 1, 0,
					-- layer=2 filter=36 channel=88
					-14, -6, -10, -3, -5, 2, -11, -1, 0,
					-- layer=2 filter=36 channel=89
					-8, -6, 1, -8, 6, 2, -12, 0, -2,
					-- layer=2 filter=36 channel=90
					6, 8, 0, -9, 0, 2, -3, 0, 9,
					-- layer=2 filter=36 channel=91
					-9, -2, -6, 3, -3, -5, -8, 0, -1,
					-- layer=2 filter=36 channel=92
					4, -5, -9, 3, -5, -2, -2, -7, 3,
					-- layer=2 filter=36 channel=93
					0, -5, -2, -10, -9, 8, -3, 3, -6,
					-- layer=2 filter=36 channel=94
					-9, -6, -2, 2, -10, 2, 0, -9, 1,
					-- layer=2 filter=36 channel=95
					-12, 6, 5, -3, 0, -3, -7, -8, 7,
					-- layer=2 filter=36 channel=96
					0, -3, -11, -2, -15, 6, 8, 5, 9,
					-- layer=2 filter=36 channel=97
					3, 1, -2, 6, 0, -8, 0, -8, -1,
					-- layer=2 filter=36 channel=98
					-7, -9, -14, -11, -14, -10, 0, -9, -4,
					-- layer=2 filter=36 channel=99
					0, -3, 4, 2, 7, 2, -5, -11, 2,
					-- layer=2 filter=36 channel=100
					-11, 0, -13, -3, -10, -4, -1, 3, -17,
					-- layer=2 filter=36 channel=101
					0, -13, -10, -11, -2, 2, -9, -4, 1,
					-- layer=2 filter=36 channel=102
					8, 7, -8, -2, -6, 2, -3, 6, -7,
					-- layer=2 filter=36 channel=103
					-5, 6, -3, 6, -11, -2, -1, -3, 2,
					-- layer=2 filter=36 channel=104
					2, 0, -4, 4, -2, 3, -6, 5, 5,
					-- layer=2 filter=36 channel=105
					0, 5, -9, 4, -1, 9, 9, -8, -3,
					-- layer=2 filter=36 channel=106
					-8, -8, -9, 0, 3, -9, -12, 0, -2,
					-- layer=2 filter=36 channel=107
					5, -8, -6, 10, 0, -2, -4, -7, -11,
					-- layer=2 filter=36 channel=108
					1, -2, 0, -13, -3, 2, -11, -8, -10,
					-- layer=2 filter=36 channel=109
					2, -1, 1, 0, 3, 4, 9, 0, 0,
					-- layer=2 filter=36 channel=110
					1, 1, -13, -7, 0, -8, -16, -1, -4,
					-- layer=2 filter=36 channel=111
					6, 7, -3, -2, -3, 9, 5, -5, 2,
					-- layer=2 filter=36 channel=112
					-3, -5, -10, 5, 1, -5, -8, 1, 2,
					-- layer=2 filter=36 channel=113
					0, 0, 3, 4, -5, 6, -9, -12, -6,
					-- layer=2 filter=36 channel=114
					8, 1, 1, 2, 0, -7, -8, -2, 4,
					-- layer=2 filter=36 channel=115
					7, -1, 4, 0, 8, -6, 7, 1, 1,
					-- layer=2 filter=36 channel=116
					-10, -13, -2, -6, -8, -8, 13, 0, -11,
					-- layer=2 filter=36 channel=117
					-11, 8, -10, 6, -11, 2, 7, -10, -1,
					-- layer=2 filter=36 channel=118
					-11, -1, -2, 0, 6, -12, -11, 0, 0,
					-- layer=2 filter=36 channel=119
					-11, -4, 8, -5, -11, -9, -6, 0, 0,
					-- layer=2 filter=36 channel=120
					8, 9, -3, 9, 3, 0, -9, 2, -8,
					-- layer=2 filter=36 channel=121
					0, 10, 1, -2, 11, 9, -1, 0, 0,
					-- layer=2 filter=36 channel=122
					2, 6, -8, 1, -10, 0, -4, 7, 6,
					-- layer=2 filter=36 channel=123
					0, -2, 5, -12, -8, 5, 10, -6, -5,
					-- layer=2 filter=36 channel=124
					3, 4, 0, 2, -4, -7, 0, -3, -9,
					-- layer=2 filter=36 channel=125
					-1, -2, 6, -3, 2, -8, -5, -1, 2,
					-- layer=2 filter=36 channel=126
					-3, 3, -6, 4, 0, 4, 5, 5, -1,
					-- layer=2 filter=36 channel=127
					0, -4, 0, -2, -9, -11, 1, -12, 2,
					-- layer=2 filter=37 channel=0
					-6, -13, -9, -7, -9, -5, -7, -15, -5,
					-- layer=2 filter=37 channel=1
					-9, -7, -1, 5, 0, 7, -8, -11, 6,
					-- layer=2 filter=37 channel=2
					6, 6, 2, -8, -2, 0, 3, -11, -9,
					-- layer=2 filter=37 channel=3
					-10, -6, -11, -9, 6, -1, 2, 4, -9,
					-- layer=2 filter=37 channel=4
					8, 3, -13, -2, 1, -10, 1, -1, -2,
					-- layer=2 filter=37 channel=5
					4, 1, -5, 0, -2, -9, 3, -3, 1,
					-- layer=2 filter=37 channel=6
					9, -6, -8, -12, 8, 5, -7, 0, -3,
					-- layer=2 filter=37 channel=7
					3, -3, -5, 3, -6, -3, 11, -4, 5,
					-- layer=2 filter=37 channel=8
					-3, -9, -3, 5, 2, -9, 8, 6, 0,
					-- layer=2 filter=37 channel=9
					-14, -12, -7, -12, 0, -9, -6, 1, -5,
					-- layer=2 filter=37 channel=10
					-10, 5, -12, -8, 0, -7, -9, -12, -11,
					-- layer=2 filter=37 channel=11
					0, 4, -2, 3, -2, -8, 0, -7, -1,
					-- layer=2 filter=37 channel=12
					-8, 4, -15, 5, 2, 9, -4, 0, -3,
					-- layer=2 filter=37 channel=13
					-10, 1, 10, 5, 7, -9, -7, 0, -5,
					-- layer=2 filter=37 channel=14
					5, -7, -2, -6, -7, 4, 4, -11, 4,
					-- layer=2 filter=37 channel=15
					-9, 5, 6, 0, -3, -1, 1, 3, 1,
					-- layer=2 filter=37 channel=16
					7, 6, 0, -15, -1, -5, -1, -3, -2,
					-- layer=2 filter=37 channel=17
					6, 4, -6, -3, 0, -7, 0, 9, 0,
					-- layer=2 filter=37 channel=18
					-1, 0, 6, -3, 0, -5, 4, -3, -1,
					-- layer=2 filter=37 channel=19
					0, -10, -7, -9, -12, -10, -7, -12, -3,
					-- layer=2 filter=37 channel=20
					-10, -1, 2, -9, -7, 2, 3, 9, 3,
					-- layer=2 filter=37 channel=21
					2, -3, -4, 3, -7, 2, 3, 3, 4,
					-- layer=2 filter=37 channel=22
					8, 7, 5, -1, 0, 7, 6, -7, 6,
					-- layer=2 filter=37 channel=23
					-9, 5, 0, 0, 2, -5, 1, 5, 5,
					-- layer=2 filter=37 channel=24
					-10, -4, 0, 5, -13, 4, 4, -2, -10,
					-- layer=2 filter=37 channel=25
					1, -4, 1, -1, -13, -12, -8, 5, -2,
					-- layer=2 filter=37 channel=26
					-8, 6, 5, 0, 4, -4, 7, 10, 5,
					-- layer=2 filter=37 channel=27
					1, -8, -11, -1, -8, -6, 2, -7, -18,
					-- layer=2 filter=37 channel=28
					5, -14, -1, -3, 0, -11, -10, 0, 0,
					-- layer=2 filter=37 channel=29
					-10, -7, 7, -2, 1, 5, 6, 5, -8,
					-- layer=2 filter=37 channel=30
					-13, -7, -6, -10, -11, -5, -12, 1, -12,
					-- layer=2 filter=37 channel=31
					-3, -2, -1, 0, 8, -2, 1, 1, -6,
					-- layer=2 filter=37 channel=32
					1, 7, -10, -3, -2, 0, -2, -2, 4,
					-- layer=2 filter=37 channel=33
					-8, 5, -8, 4, -5, -11, 3, -2, -12,
					-- layer=2 filter=37 channel=34
					9, -1, 9, 10, 4, 8, 1, -6, -1,
					-- layer=2 filter=37 channel=35
					10, -9, 8, -5, -8, -5, -1, -13, -2,
					-- layer=2 filter=37 channel=36
					2, -4, -1, 7, 2, 0, 5, -1, -3,
					-- layer=2 filter=37 channel=37
					-8, -4, 2, 4, -9, -7, 0, 2, -10,
					-- layer=2 filter=37 channel=38
					0, -10, 2, -15, -4, -1, -10, 0, 3,
					-- layer=2 filter=37 channel=39
					-6, -13, -12, 0, -11, -5, 3, -4, -9,
					-- layer=2 filter=37 channel=40
					8, 3, -6, 1, 2, -8, 9, -4, -10,
					-- layer=2 filter=37 channel=41
					0, 8, -5, 5, 4, -4, -8, -4, -5,
					-- layer=2 filter=37 channel=42
					1, -1, -5, -1, -13, 1, -14, 0, 0,
					-- layer=2 filter=37 channel=43
					-14, -1, 0, 5, 5, 0, 1, -5, 0,
					-- layer=2 filter=37 channel=44
					6, 8, 7, -8, -8, 1, 0, 2, -7,
					-- layer=2 filter=37 channel=45
					-9, -12, -2, 5, -14, 2, -1, 1, 0,
					-- layer=2 filter=37 channel=46
					3, 0, -15, -8, 2, -7, 4, -8, 4,
					-- layer=2 filter=37 channel=47
					-9, -4, -8, -4, 4, 2, 0, -9, -3,
					-- layer=2 filter=37 channel=48
					7, 8, -8, -2, 2, 5, -5, 5, 7,
					-- layer=2 filter=37 channel=49
					-6, 6, 5, 7, 1, -4, 7, -2, 5,
					-- layer=2 filter=37 channel=50
					-1, -15, -6, 6, -8, 6, -10, -8, 11,
					-- layer=2 filter=37 channel=51
					-4, 1, 5, 2, 4, -10, -5, -14, -10,
					-- layer=2 filter=37 channel=52
					-12, -14, 1, 4, 4, -10, 1, -7, 6,
					-- layer=2 filter=37 channel=53
					-6, -5, -4, 2, -11, -11, 6, 4, 7,
					-- layer=2 filter=37 channel=54
					13, -7, -10, 3, -1, -6, 10, -3, -13,
					-- layer=2 filter=37 channel=55
					4, 6, 2, 6, 4, 7, 7, 1, 0,
					-- layer=2 filter=37 channel=56
					6, 1, -13, -9, 4, -7, -5, -1, 3,
					-- layer=2 filter=37 channel=57
					7, -9, 11, 8, 7, 6, 7, 4, 1,
					-- layer=2 filter=37 channel=58
					2, -12, -1, -6, 0, 0, -10, 5, -5,
					-- layer=2 filter=37 channel=59
					-1, -15, -14, 3, 2, -9, 3, 8, -12,
					-- layer=2 filter=37 channel=60
					2, -5, -6, -2, 3, 11, -7, 4, 5,
					-- layer=2 filter=37 channel=61
					0, 2, -9, -16, 1, -9, -12, 2, -1,
					-- layer=2 filter=37 channel=62
					4, -12, 2, 0, 2, 5, 0, -6, -4,
					-- layer=2 filter=37 channel=63
					0, 8, 4, -9, 11, -2, -12, -6, 0,
					-- layer=2 filter=37 channel=64
					-6, -9, -3, -9, -13, -4, -12, -3, -5,
					-- layer=2 filter=37 channel=65
					-1, -10, -3, -17, -15, 7, -14, -5, 9,
					-- layer=2 filter=37 channel=66
					9, -2, 4, 0, -2, 6, 4, -3, -11,
					-- layer=2 filter=37 channel=67
					-2, -14, -8, 0, -7, -6, -3, -4, 0,
					-- layer=2 filter=37 channel=68
					8, 4, 1, -12, -8, -10, -2, 7, 0,
					-- layer=2 filter=37 channel=69
					4, 1, 1, -9, 2, -12, 3, -5, 8,
					-- layer=2 filter=37 channel=70
					-12, -4, 1, -9, 11, -4, -4, -3, -3,
					-- layer=2 filter=37 channel=71
					-12, -2, -12, 2, -9, -3, 0, -2, -8,
					-- layer=2 filter=37 channel=72
					-6, -4, -7, -10, -4, -6, 5, 7, -2,
					-- layer=2 filter=37 channel=73
					1, 3, 11, 3, 0, 2, -10, -7, -7,
					-- layer=2 filter=37 channel=74
					0, -2, -14, -14, -4, 2, -9, -11, 4,
					-- layer=2 filter=37 channel=75
					9, -8, -3, 5, 4, 6, -8, 4, -5,
					-- layer=2 filter=37 channel=76
					7, 10, -2, -10, 1, -7, 6, -7, 1,
					-- layer=2 filter=37 channel=77
					-6, -8, 0, 8, 2, 0, 2, 5, -12,
					-- layer=2 filter=37 channel=78
					-9, -2, -11, -5, -5, -4, -6, 4, -14,
					-- layer=2 filter=37 channel=79
					-9, -3, 0, -1, -4, 7, 6, -8, 6,
					-- layer=2 filter=37 channel=80
					-10, -12, -8, -16, 3, -2, -11, -6, 0,
					-- layer=2 filter=37 channel=81
					-9, 8, 6, 2, -9, 0, 4, -11, 4,
					-- layer=2 filter=37 channel=82
					2, -5, -7, 10, -9, -5, 6, 8, 10,
					-- layer=2 filter=37 channel=83
					-10, 2, -11, 6, -2, 4, -10, 2, -14,
					-- layer=2 filter=37 channel=84
					-1, 6, -7, 0, 0, 2, 7, -1, 3,
					-- layer=2 filter=37 channel=85
					5, 8, -6, -8, 2, 7, 3, -8, 9,
					-- layer=2 filter=37 channel=86
					-11, -1, 0, -2, -10, -9, -2, -4, 2,
					-- layer=2 filter=37 channel=87
					7, 0, 2, 8, -5, -4, -4, -14, -7,
					-- layer=2 filter=37 channel=88
					-1, -11, -11, 5, -4, 6, -7, -10, -10,
					-- layer=2 filter=37 channel=89
					3, -3, -13, 2, -6, -4, 4, -3, 3,
					-- layer=2 filter=37 channel=90
					6, 4, 5, 6, 0, -3, -8, -1, 2,
					-- layer=2 filter=37 channel=91
					0, -12, 4, 3, -2, 7, -4, 1, 5,
					-- layer=2 filter=37 channel=92
					0, 2, 0, -6, -9, 6, -3, -10, 7,
					-- layer=2 filter=37 channel=93
					7, -11, 2, -10, -4, 5, -2, -7, -5,
					-- layer=2 filter=37 channel=94
					7, 4, 6, -8, 3, 5, -1, -9, 5,
					-- layer=2 filter=37 channel=95
					0, -1, -12, 8, 6, 0, -1, 7, 3,
					-- layer=2 filter=37 channel=96
					-9, 11, 0, 2, -8, -14, -2, -3, -12,
					-- layer=2 filter=37 channel=97
					0, -8, -2, 3, 2, -13, 0, -11, 2,
					-- layer=2 filter=37 channel=98
					0, -4, 0, 9, 8, -4, -4, -6, -1,
					-- layer=2 filter=37 channel=99
					3, 0, -6, -12, 0, -10, -14, -8, -6,
					-- layer=2 filter=37 channel=100
					-1, -8, -12, 6, -17, 1, 3, -14, 0,
					-- layer=2 filter=37 channel=101
					-11, -6, -4, 6, 2, 9, -9, 5, 0,
					-- layer=2 filter=37 channel=102
					7, 5, 2, -7, 4, 2, -8, 7, -8,
					-- layer=2 filter=37 channel=103
					-7, -7, 7, -6, -6, -11, 3, 2, 3,
					-- layer=2 filter=37 channel=104
					-7, -14, -2, -9, -4, 5, -1, -7, -3,
					-- layer=2 filter=37 channel=105
					0, -2, -11, 5, 5, 1, -4, -11, -5,
					-- layer=2 filter=37 channel=106
					-8, 2, 3, -12, 4, -3, 3, 0, -2,
					-- layer=2 filter=37 channel=107
					6, -5, -5, -6, -5, -7, 4, 0, -1,
					-- layer=2 filter=37 channel=108
					-13, 4, -8, -1, 4, -1, -1, 0, -14,
					-- layer=2 filter=37 channel=109
					-4, 7, -8, 6, -1, 1, -2, -12, 0,
					-- layer=2 filter=37 channel=110
					-3, 1, -4, -15, -11, -2, -4, 3, 7,
					-- layer=2 filter=37 channel=111
					9, 3, 10, -5, 4, -2, 1, 0, -7,
					-- layer=2 filter=37 channel=112
					-10, -10, -10, -5, -5, -11, -10, -11, -4,
					-- layer=2 filter=37 channel=113
					-12, 2, 0, 6, 0, -11, -1, 4, -12,
					-- layer=2 filter=37 channel=114
					-3, -6, 1, -2, -2, -2, 1, 3, 2,
					-- layer=2 filter=37 channel=115
					9, 8, 1, 5, 8, -4, 7, 4, 2,
					-- layer=2 filter=37 channel=116
					5, 1, 11, -2, -1, 0, 8, -5, -6,
					-- layer=2 filter=37 channel=117
					-12, -4, -3, -1, 9, 3, 0, -2, 7,
					-- layer=2 filter=37 channel=118
					-11, 4, -4, -4, -8, 1, -4, 2, -15,
					-- layer=2 filter=37 channel=119
					5, 0, -14, -7, -10, -2, 4, -2, 0,
					-- layer=2 filter=37 channel=120
					0, -2, -2, 8, 10, 7, 4, 1, 0,
					-- layer=2 filter=37 channel=121
					8, -8, 2, 0, -8, -6, 3, 0, 8,
					-- layer=2 filter=37 channel=122
					0, 5, 1, -7, 1, -9, 6, 4, -10,
					-- layer=2 filter=37 channel=123
					-3, 8, -7, -4, -2, -10, 6, 6, -10,
					-- layer=2 filter=37 channel=124
					-3, -13, 2, 2, -1, 5, -2, -8, -10,
					-- layer=2 filter=37 channel=125
					0, 3, -1, -6, -10, 7, -1, 7, 6,
					-- layer=2 filter=37 channel=126
					-10, -8, 3, -4, -5, 0, 2, -6, 4,
					-- layer=2 filter=37 channel=127
					-1, -10, -3, -3, 6, 2, 0, -9, 5,
					-- layer=2 filter=38 channel=0
					10, 22, -9, 16, 10, -47, 9, 24, 38,
					-- layer=2 filter=38 channel=1
					0, 7, -6, 6, -11, 21, -22, -27, -45,
					-- layer=2 filter=38 channel=2
					7, 3, 1, -2, 1, -11, -9, -9, -10,
					-- layer=2 filter=38 channel=3
					-5, -22, -33, 11, -19, -21, -27, -29, -25,
					-- layer=2 filter=38 channel=4
					0, -26, 0, -4, -65, 2, -1, -4, -15,
					-- layer=2 filter=38 channel=5
					-2, -6, -12, 12, -5, -13, -1, 1, 29,
					-- layer=2 filter=38 channel=6
					34, 15, 8, 14, 20, 8, -2, 32, 9,
					-- layer=2 filter=38 channel=7
					42, 0, -15, -45, 7, 21, -25, -25, -21,
					-- layer=2 filter=38 channel=8
					2, 2, -2, -3, 7, 5, 2, 2, 4,
					-- layer=2 filter=38 channel=9
					13, 34, 0, 43, 16, 29, -30, -83, -48,
					-- layer=2 filter=38 channel=10
					11, -5, 1, 16, -14, -28, 7, 4, 27,
					-- layer=2 filter=38 channel=11
					16, 0, 17, 6, 19, 12, 23, 9, 15,
					-- layer=2 filter=38 channel=12
					11, 24, 3, 15, 33, 47, -4, -29, -32,
					-- layer=2 filter=38 channel=13
					12, -7, 2, 10, 5, 3, 7, 5, -4,
					-- layer=2 filter=38 channel=14
					4, 0, 17, 12, 23, 13, -26, -21, -10,
					-- layer=2 filter=38 channel=15
					-17, -6, 22, 7, -31, 10, 39, 10, 26,
					-- layer=2 filter=38 channel=16
					9, 20, 18, 35, -32, 4, -18, -18, 1,
					-- layer=2 filter=38 channel=17
					-2, -9, 3, -10, -3, -3, 5, 2, -9,
					-- layer=2 filter=38 channel=18
					-1, -7, 30, -24, -35, 1, -12, 1, 10,
					-- layer=2 filter=38 channel=19
					33, 36, 56, -2, -9, 24, -19, -16, 6,
					-- layer=2 filter=38 channel=20
					-5, -8, 4, -6, 5, 1, -4, 1, 6,
					-- layer=2 filter=38 channel=21
					8, 16, -10, 9, -4, -4, -17, -5, 2,
					-- layer=2 filter=38 channel=22
					7, 5, -5, 0, 7, 4, 1, 2, -4,
					-- layer=2 filter=38 channel=23
					8, 3, -27, 7, -6, 12, -16, -20, -53,
					-- layer=2 filter=38 channel=24
					-28, -22, -28, -44, -39, -57, -57, -51, -46,
					-- layer=2 filter=38 channel=25
					-6, -9, -35, -23, -8, -23, -20, -10, 13,
					-- layer=2 filter=38 channel=26
					8, -7, -9, 0, -7, 8, 4, 10, 7,
					-- layer=2 filter=38 channel=27
					-12, 0, 29, 15, 0, -1, -26, -36, 0,
					-- layer=2 filter=38 channel=28
					18, 0, -17, -22, -35, -34, -5, 34, 21,
					-- layer=2 filter=38 channel=29
					1, 1, 1, 5, 6, -6, -10, -4, 2,
					-- layer=2 filter=38 channel=30
					-9, 17, -1, 32, -34, -35, -24, -10, 21,
					-- layer=2 filter=38 channel=31
					33, 20, -10, 26, 24, -54, -22, 56, 51,
					-- layer=2 filter=38 channel=32
					-7, -3, -1, 1, -5, -8, 4, 2, -2,
					-- layer=2 filter=38 channel=33
					0, -36, 21, 1, 37, 61, 12, 12, -27,
					-- layer=2 filter=38 channel=34
					-8, 33, 51, -25, 16, 17, -11, -10, 16,
					-- layer=2 filter=38 channel=35
					23, 15, 9, 2, -39, -9, 8, -5, 1,
					-- layer=2 filter=38 channel=36
					5, -9, -4, -4, 0, -15, -4, 2, 6,
					-- layer=2 filter=38 channel=37
					-16, -7, 0, 20, -13, 3, 7, -12, 18,
					-- layer=2 filter=38 channel=38
					-8, 12, 1, 17, 3, 24, -7, -55, -6,
					-- layer=2 filter=38 channel=39
					-9, 0, -11, -3, -7, -16, -7, -34, -39,
					-- layer=2 filter=38 channel=40
					-9, -8, 39, -2, 9, -5, -2, 4, 38,
					-- layer=2 filter=38 channel=41
					-7, -6, -6, -6, -3, 11, -11, -3, 11,
					-- layer=2 filter=38 channel=42
					-5, -24, -21, 16, -30, -10, -27, -11, -73,
					-- layer=2 filter=38 channel=43
					18, 2, 17, 2, -38, -6, 8, 2, 12,
					-- layer=2 filter=38 channel=44
					-6, 1, 5, -7, -8, 2, -6, -3, 5,
					-- layer=2 filter=38 channel=45
					-2, -15, -15, -17, -53, -11, -63, -53, -27,
					-- layer=2 filter=38 channel=46
					0, -17, 23, 22, -3, -33, -28, 8, 22,
					-- layer=2 filter=38 channel=47
					-5, -38, -34, -22, 8, -16, -7, 3, 38,
					-- layer=2 filter=38 channel=48
					3, 2, -5, -6, 7, 4, 0, -5, 8,
					-- layer=2 filter=38 channel=49
					31, 16, -7, 9, -39, -11, -9, -18, 10,
					-- layer=2 filter=38 channel=50
					-2, -6, -9, 7, 4, -3, 10, 20, 11,
					-- layer=2 filter=38 channel=51
					23, 0, -9, 18, -3, 0, 19, 16, 17,
					-- layer=2 filter=38 channel=52
					-17, 16, 7, 18, -4, 6, -4, -13, 14,
					-- layer=2 filter=38 channel=53
					4, 62, 9, 41, 19, -18, 17, 32, 17,
					-- layer=2 filter=38 channel=54
					12, 20, 5, 6, 2, 52, -5, 17, 28,
					-- layer=2 filter=38 channel=55
					-11, -6, 7, 8, -15, -14, 0, -7, -15,
					-- layer=2 filter=38 channel=56
					16, 11, 14, 9, 8, 3, 18, -6, 6,
					-- layer=2 filter=38 channel=57
					-4, -9, 4, 0, 3, 10, -10, -7, 3,
					-- layer=2 filter=38 channel=58
					-8, -4, 0, 31, 54, 38, 1, -40, -40,
					-- layer=2 filter=38 channel=59
					-11, 9, 4, 13, 25, -2, -10, -20, -36,
					-- layer=2 filter=38 channel=60
					-12, 9, 24, 16, 11, -12, 28, -10, -16,
					-- layer=2 filter=38 channel=61
					9, 22, -18, 2, -11, -60, -20, -31, -31,
					-- layer=2 filter=38 channel=62
					2, 30, 21, -11, -16, 4, -12, 2, 27,
					-- layer=2 filter=38 channel=63
					25, 0, 1, 12, -14, -17, 11, -22, -12,
					-- layer=2 filter=38 channel=64
					-26, -19, -16, -26, -22, -47, -23, -47, -19,
					-- layer=2 filter=38 channel=65
					26, 17, -3, 21, -7, 3, 4, -10, 3,
					-- layer=2 filter=38 channel=66
					33, -32, 35, -21, 23, 6, -23, 1, -38,
					-- layer=2 filter=38 channel=67
					-2, -12, 18, 61, -12, -32, 14, -25, -30,
					-- layer=2 filter=38 channel=68
					-8, -6, -8, 8, -6, -5, -10, 0, -7,
					-- layer=2 filter=38 channel=69
					-19, -2, -38, 9, -21, -1, 17, -25, -7,
					-- layer=2 filter=38 channel=70
					5, 9, -5, -10, -13, 13, 9, 18, 24,
					-- layer=2 filter=38 channel=71
					3, 24, 17, 9, 7, -3, 6, -18, 26,
					-- layer=2 filter=38 channel=72
					5, -28, -4, -52, 18, 21, 7, 7, -19,
					-- layer=2 filter=38 channel=73
					32, 33, 15, -27, 7, -31, -35, 31, -14,
					-- layer=2 filter=38 channel=74
					-33, 4, 29, 24, -9, -32, 37, 3, -30,
					-- layer=2 filter=38 channel=75
					21, 4, 19, 7, 52, -12, -13, -20, 15,
					-- layer=2 filter=38 channel=76
					24, 16, 0, 35, 19, -12, -47, -5, 1,
					-- layer=2 filter=38 channel=77
					3, 4, -7, 0, 11, -7, -1, 1, -6,
					-- layer=2 filter=38 channel=78
					-8, 2, -28, -20, -34, -19, -12, -27, 21,
					-- layer=2 filter=38 channel=79
					-9, -10, -1, 11, 6, -8, -6, -1, -2,
					-- layer=2 filter=38 channel=80
					-14, -22, 5, 22, -35, -63, -33, -3, -11,
					-- layer=2 filter=38 channel=81
					0, 0, -1, -7, 12, -8, 3, -10, 0,
					-- layer=2 filter=38 channel=82
					-4, 7, -1, -9, -4, 6, 8, -7, -8,
					-- layer=2 filter=38 channel=83
					-18, -23, 11, -11, -83, -3, 21, -41, 16,
					-- layer=2 filter=38 channel=84
					-6, -6, 0, -6, -8, 3, -4, 4, -7,
					-- layer=2 filter=38 channel=85
					-2, 0, 10, 8, -6, 3, 7, -3, -8,
					-- layer=2 filter=38 channel=86
					2, 1, 6, -3, -8, -9, 1, -5, 9,
					-- layer=2 filter=38 channel=87
					-40, -15, 18, 15, -20, -22, 12, 2, -27,
					-- layer=2 filter=38 channel=88
					-19, 12, -9, 25, -16, 20, 11, -28, -45,
					-- layer=2 filter=38 channel=89
					-8, 6, 14, 0, 26, 14, -11, -13, -16,
					-- layer=2 filter=38 channel=90
					4, -1, -3, 7, -1, -10, -3, -10, 6,
					-- layer=2 filter=38 channel=91
					-12, 3, -8, -35, 25, -4, -17, -3, -57,
					-- layer=2 filter=38 channel=92
					6, -1, -19, -11, 13, 28, -19, -37, -59,
					-- layer=2 filter=38 channel=93
					32, 28, 20, -26, -11, -31, -27, -24, 11,
					-- layer=2 filter=38 channel=94
					-9, -1, 14, 23, 35, -34, -16, 0, -46,
					-- layer=2 filter=38 channel=95
					4, -10, -13, -12, 5, 0, -11, -5, -3,
					-- layer=2 filter=38 channel=96
					-14, 16, 1, 14, 38, 8, 26, 52, 57,
					-- layer=2 filter=38 channel=97
					22, 19, 42, -9, -1, 2, -24, -50, -35,
					-- layer=2 filter=38 channel=98
					10, -6, 6, -28, -11, -19, -2, 9, 27,
					-- layer=2 filter=38 channel=99
					-14, 2, 2, 20, 0, 17, 18, 4, -2,
					-- layer=2 filter=38 channel=100
					-40, -5, 1, -25, 1, -1, -1, -20, -22,
					-- layer=2 filter=38 channel=101
					10, 7, 24, 18, -3, -2, 24, -9, 31,
					-- layer=2 filter=38 channel=102
					-15, 5, 15, -7, -50, 10, 4, -2, 0,
					-- layer=2 filter=38 channel=103
					25, -27, -29, -11, -13, 18, -14, -29, -8,
					-- layer=2 filter=38 channel=104
					1, 10, 6, 14, -30, -16, -17, -23, -25,
					-- layer=2 filter=38 channel=105
					9, 32, 76, -13, 16, -3, 20, -6, 11,
					-- layer=2 filter=38 channel=106
					0, 1, 2, 13, 14, 20, 15, -24, 5,
					-- layer=2 filter=38 channel=107
					11, 24, 11, -11, 12, -21, 10, 4, -4,
					-- layer=2 filter=38 channel=108
					-23, 0, 16, 25, -13, 23, -23, -38, 19,
					-- layer=2 filter=38 channel=109
					13, 12, 8, -10, 11, -3, -15, 9, 15,
					-- layer=2 filter=38 channel=110
					10, 17, -18, -43, -20, -13, -55, -66, -50,
					-- layer=2 filter=38 channel=111
					9, -5, -6, 8, 4, 5, 3, 3, -1,
					-- layer=2 filter=38 channel=112
					22, -16, -2, 30, -12, -1, 26, 15, 29,
					-- layer=2 filter=38 channel=113
					16, 17, -31, 34, -42, -43, 18, 10, -15,
					-- layer=2 filter=38 channel=114
					15, -1, 9, 12, 8, 13, 12, 20, 20,
					-- layer=2 filter=38 channel=115
					-7, -5, 8, -6, 4, 6, 11, -3, -3,
					-- layer=2 filter=38 channel=116
					-58, 0, 48, 10, -29, 18, 22, -8, 23,
					-- layer=2 filter=38 channel=117
					26, 23, 19, -15, -11, 21, -17, -31, -3,
					-- layer=2 filter=38 channel=118
					-14, -11, 10, 7, -37, 0, -9, -17, -16,
					-- layer=2 filter=38 channel=119
					4, -28, 2, -6, -65, 8, 15, -28, -35,
					-- layer=2 filter=38 channel=120
					0, 0, 0, -5, -6, -5, 3, -3, -3,
					-- layer=2 filter=38 channel=121
					3, -1, 7, -8, -3, 6, -2, 10, 9,
					-- layer=2 filter=38 channel=122
					13, 10, 10, -5, 5, -3, 7, 12, 1,
					-- layer=2 filter=38 channel=123
					-3, 14, 0, -45, 5, 33, 12, -1, 11,
					-- layer=2 filter=38 channel=124
					31, -28, 29, -24, -47, 28, 10, 19, -19,
					-- layer=2 filter=38 channel=125
					-11, 2, 8, 5, -1, -1, 0, 1, 1,
					-- layer=2 filter=38 channel=126
					-11, 12, -41, 41, 5, -37, 20, 16, -43,
					-- layer=2 filter=38 channel=127
					-31, -6, -38, -9, -44, 3, -3, -17, -27,
					-- layer=2 filter=39 channel=0
					23, 15, 32, 5, -3, -1, -19, -41, -23,
					-- layer=2 filter=39 channel=1
					-14, 8, 1, 0, 42, -13, 12, 17, 21,
					-- layer=2 filter=39 channel=2
					6, 1, -8, -8, -1, 1, -1, 10, -7,
					-- layer=2 filter=39 channel=3
					26, 16, -9, 11, -1, -14, -20, -22, -44,
					-- layer=2 filter=39 channel=4
					19, -8, 12, 23, 48, -8, 1, -4, -5,
					-- layer=2 filter=39 channel=5
					8, 10, 28, -33, -3, -21, -10, -1, -2,
					-- layer=2 filter=39 channel=6
					-11, -16, -42, -6, -29, -43, 27, 46, 31,
					-- layer=2 filter=39 channel=7
					-3, 13, 48, -46, 10, -15, -6, 5, 5,
					-- layer=2 filter=39 channel=8
					2, -1, -4, 4, 2, 4, 1, 7, 0,
					-- layer=2 filter=39 channel=9
					-19, -8, -10, -14, 19, -6, -11, -1, -7,
					-- layer=2 filter=39 channel=10
					43, 24, 0, 8, 11, 0, -31, -15, -36,
					-- layer=2 filter=39 channel=11
					16, -2, 12, -8, -26, -13, -27, -13, -18,
					-- layer=2 filter=39 channel=12
					13, 15, 31, 35, 21, -9, 16, 11, 24,
					-- layer=2 filter=39 channel=13
					-4, -6, -5, -6, 2, -3, 3, -7, 0,
					-- layer=2 filter=39 channel=14
					-5, 1, 0, 3, 42, 0, 29, 21, 16,
					-- layer=2 filter=39 channel=15
					-21, -6, -7, -56, -9, 42, -63, -53, 6,
					-- layer=2 filter=39 channel=16
					-19, 12, 12, 19, 16, 19, 14, 10, 11,
					-- layer=2 filter=39 channel=17
					-10, 4, -10, 9, 4, -1, 0, 7, -4,
					-- layer=2 filter=39 channel=18
					0, -15, 36, -16, -19, -12, -7, 0, 14,
					-- layer=2 filter=39 channel=19
					-19, -1, 13, -23, 36, 3, 12, 5, 7,
					-- layer=2 filter=39 channel=20
					-3, 0, 5, 9, -6, -6, 4, 1, 2,
					-- layer=2 filter=39 channel=21
					-26, -16, -27, -15, 6, 4, -16, -27, -15,
					-- layer=2 filter=39 channel=22
					-5, 2, 8, 3, 8, -3, -5, 0, 7,
					-- layer=2 filter=39 channel=23
					-7, -19, -7, -4, -11, -6, 29, 10, 24,
					-- layer=2 filter=39 channel=24
					34, 31, -1, 39, 36, 12, 4, -5, -9,
					-- layer=2 filter=39 channel=25
					60, 41, 7, 39, -1, 6, -14, -31, -20,
					-- layer=2 filter=39 channel=26
					-2, -5, -3, -2, 1, 0, 0, -8, -11,
					-- layer=2 filter=39 channel=27
					5, 3, -12, 2, 45, -13, -37, -7, -15,
					-- layer=2 filter=39 channel=28
					8, 35, 3, 0, 33, 20, -2, -27, -20,
					-- layer=2 filter=39 channel=29
					-8, 0, -4, 8, -1, 0, -5, 0, -9,
					-- layer=2 filter=39 channel=30
					-14, -15, 19, 27, -8, 23, 33, -18, 20,
					-- layer=2 filter=39 channel=31
					-5, 17, -53, -143, -54, -56, -68, -107, -54,
					-- layer=2 filter=39 channel=32
					6, 6, 2, -4, 4, -7, -6, -4, 0,
					-- layer=2 filter=39 channel=33
					-16, -15, -26, -48, -18, -27, -28, -13, -2,
					-- layer=2 filter=39 channel=34
					-45, -11, 8, -6, -8, 37, 5, -5, -24,
					-- layer=2 filter=39 channel=35
					46, 45, 18, -13, 7, 30, -30, 2, -45,
					-- layer=2 filter=39 channel=36
					10, 0, 10, 11, -10, 5, -6, -1, -4,
					-- layer=2 filter=39 channel=37
					1, -12, 7, -24, -10, -17, -20, 8, 2,
					-- layer=2 filter=39 channel=38
					-24, 0, -7, -5, 19, -16, -27, 3, -9,
					-- layer=2 filter=39 channel=39
					-21, -5, -10, -1, 4, 5, 12, 30, 18,
					-- layer=2 filter=39 channel=40
					21, -39, 16, -35, -62, -37, -55, 2, 50,
					-- layer=2 filter=39 channel=41
					-3, -8, 6, 0, 1, 1, 5, -12, -8,
					-- layer=2 filter=39 channel=42
					15, -15, -6, 25, 14, 14, 7, 3, 23,
					-- layer=2 filter=39 channel=43
					62, 13, -47, -34, -22, -17, -37, -18, -17,
					-- layer=2 filter=39 channel=44
					-3, 8, 10, -4, 5, 5, -1, -7, 9,
					-- layer=2 filter=39 channel=45
					7, 21, -34, 31, 69, 12, -13, -7, -10,
					-- layer=2 filter=39 channel=46
					26, -13, -18, 10, -20, -2, -20, -68, 11,
					-- layer=2 filter=39 channel=47
					-3, 36, 14, 34, 20, 13, -35, -5, -19,
					-- layer=2 filter=39 channel=48
					-1, 4, -7, 10, -9, 3, -8, -2, -6,
					-- layer=2 filter=39 channel=49
					-3, 15, -24, -15, 10, -21, 18, 23, 18,
					-- layer=2 filter=39 channel=50
					-24, -19, 5, -9, 4, 24, -5, -6, 11,
					-- layer=2 filter=39 channel=51
					10, 15, 27, -19, -9, -5, -16, -23, -9,
					-- layer=2 filter=39 channel=52
					-52, -26, -4, -16, -19, -26, -14, -1, 15,
					-- layer=2 filter=39 channel=53
					-11, 18, -44, -53, 46, 10, -50, -28, 20,
					-- layer=2 filter=39 channel=54
					3, 32, 8, -40, -15, -21, -26, -7, 25,
					-- layer=2 filter=39 channel=55
					1, 9, -10, -11, -7, -11, 14, -4, -11,
					-- layer=2 filter=39 channel=56
					19, 11, 0, -6, -28, -7, -23, 0, 1,
					-- layer=2 filter=39 channel=57
					-5, 12, 2, 13, 9, 6, 3, 2, 3,
					-- layer=2 filter=39 channel=58
					6, 23, 27, 31, 31, 14, 1, 16, 5,
					-- layer=2 filter=39 channel=59
					-21, 15, -2, 62, 43, -16, -6, -8, 4,
					-- layer=2 filter=39 channel=60
					12, 3, 33, 9, 11, -12, 13, 27, 30,
					-- layer=2 filter=39 channel=61
					-35, -3, -17, -14, -71, -21, -2, 2, 5,
					-- layer=2 filter=39 channel=62
					-21, -1, -1, -25, -26, 1, 10, 34, 18,
					-- layer=2 filter=39 channel=63
					-8, 1, -6, 29, 7, 15, 3, 7, 35,
					-- layer=2 filter=39 channel=64
					-27, 0, -17, 22, 15, 27, 19, 15, 14,
					-- layer=2 filter=39 channel=65
					-7, -16, -5, -31, -50, -34, 13, 23, 38,
					-- layer=2 filter=39 channel=66
					19, -6, -42, 0, 6, -36, -34, -20, -62,
					-- layer=2 filter=39 channel=67
					-13, -54, -43, 19, 11, 8, -23, -56, -43,
					-- layer=2 filter=39 channel=68
					-12, 5, 3, -2, 10, -4, 5, -11, 1,
					-- layer=2 filter=39 channel=69
					-28, -22, -15, 20, 15, 7, 31, 25, 31,
					-- layer=2 filter=39 channel=70
					23, 29, 16, -25, 32, 22, -33, -30, -20,
					-- layer=2 filter=39 channel=71
					-1, -24, -39, 17, 37, -24, -6, 22, -6,
					-- layer=2 filter=39 channel=72
					2, -21, 15, -39, 0, 29, 20, 15, 27,
					-- layer=2 filter=39 channel=73
					17, 52, -50, 48, 6, -29, -2, 0, -19,
					-- layer=2 filter=39 channel=74
					5, -15, -33, 41, -15, 4, -13, -21, -4,
					-- layer=2 filter=39 channel=75
					-26, 1, 34, -31, 32, -43, 21, 22, 1,
					-- layer=2 filter=39 channel=76
					-65, 29, -44, -15, -73, -20, 0, 29, -14,
					-- layer=2 filter=39 channel=77
					-1, 10, 6, 7, 0, -3, 2, -11, 9,
					-- layer=2 filter=39 channel=78
					37, 36, 9, -10, -35, -24, -31, -14, -20,
					-- layer=2 filter=39 channel=79
					-3, -9, 5, 6, 6, 1, -9, -1, 6,
					-- layer=2 filter=39 channel=80
					5, -28, -12, 32, 23, -1, 3, -18, -8,
					-- layer=2 filter=39 channel=81
					-4, -12, 8, 9, -5, 4, 2, -4, 0,
					-- layer=2 filter=39 channel=82
					-10, 10, -4, 4, -2, -6, 0, -6, 4,
					-- layer=2 filter=39 channel=83
					16, -4, -25, 28, 38, -5, 9, -5, 10,
					-- layer=2 filter=39 channel=84
					4, -11, -1, 6, 4, -2, -9, 5, -8,
					-- layer=2 filter=39 channel=85
					2, 0, 0, -18, 12, 13, 8, -2, 3,
					-- layer=2 filter=39 channel=86
					5, -13, 4, 2, 0, 32, 6, -1, 6,
					-- layer=2 filter=39 channel=87
					10, 36, -13, 28, -55, -29, 33, -6, -1,
					-- layer=2 filter=39 channel=88
					-6, -18, -9, 54, -4, 14, 26, 6, 4,
					-- layer=2 filter=39 channel=89
					-11, -1, 17, 19, 19, -4, 28, 12, 11,
					-- layer=2 filter=39 channel=90
					4, 9, 5, -2, 6, -3, -4, -9, 9,
					-- layer=2 filter=39 channel=91
					14, 11, 43, 9, 12, 13, -15, 34, 11,
					-- layer=2 filter=39 channel=92
					18, 1, 32, 20, 40, 1, 12, 11, 49,
					-- layer=2 filter=39 channel=93
					-38, 14, -6, -52, -34, -55, 0, 1, -34,
					-- layer=2 filter=39 channel=94
					-93, -41, -25, -45, -11, -52, 39, -28, 24,
					-- layer=2 filter=39 channel=95
					5, 8, 9, 1, 0, -8, 3, 0, 14,
					-- layer=2 filter=39 channel=96
					-52, -10, -34, -3, -71, -23, 14, 37, 13,
					-- layer=2 filter=39 channel=97
					0, 12, 0, 15, 9, -6, 1, 19, -2,
					-- layer=2 filter=39 channel=98
					5, 21, 0, -2, 2, 22, -12, 26, 14,
					-- layer=2 filter=39 channel=99
					-33, 1, -19, 6, 6, -32, 1, 41, 12,
					-- layer=2 filter=39 channel=100
					6, -5, 15, 6, 13, 6, -21, 19, -38,
					-- layer=2 filter=39 channel=101
					9, 6, 5, 14, 27, 8, -11, 14, 7,
					-- layer=2 filter=39 channel=102
					-41, -44, 16, -37, -67, -28, 23, 34, 19,
					-- layer=2 filter=39 channel=103
					-7, -7, 54, -32, -39, -44, -69, -44, 28,
					-- layer=2 filter=39 channel=104
					-3, -20, -19, -77, -35, -5, 28, -35, 1,
					-- layer=2 filter=39 channel=105
					-24, -8, 72, 39, 13, 19, 16, 19, -25,
					-- layer=2 filter=39 channel=106
					29, 18, 40, 25, 20, 29, -22, -9, -11,
					-- layer=2 filter=39 channel=107
					-7, -53, -6, -1, -10, -32, 17, -49, -6,
					-- layer=2 filter=39 channel=108
					-33, -17, -41, -8, 36, -1, -29, 6, 9,
					-- layer=2 filter=39 channel=109
					-1, 3, 14, -3, 8, 6, 9, -15, -3,
					-- layer=2 filter=39 channel=110
					9, -16, -16, 11, 3, 14, 58, 7, 0,
					-- layer=2 filter=39 channel=111
					-8, -5, -1, 11, -6, 1, 8, -8, 0,
					-- layer=2 filter=39 channel=112
					29, 21, 25, -6, -7, 0, -5, -49, 12,
					-- layer=2 filter=39 channel=113
					-31, -2, -15, 21, -9, 33, 8, 3, 2,
					-- layer=2 filter=39 channel=114
					7, 28, 7, 3, -5, -14, -26, 2, 6,
					-- layer=2 filter=39 channel=115
					0, 1, -3, 10, 4, 6, -4, -12, -9,
					-- layer=2 filter=39 channel=116
					-13, 2, -2, -5, -43, -16, 27, 9, -14,
					-- layer=2 filter=39 channel=117
					-33, 9, 6, -51, -5, -21, -29, -19, -3,
					-- layer=2 filter=39 channel=118
					41, 11, 3, 2, 5, -20, 4, -26, -24,
					-- layer=2 filter=39 channel=119
					-13, 30, 23, -4, 29, 10, -14, 11, -27,
					-- layer=2 filter=39 channel=120
					0, 6, -3, -9, 7, 7, 1, 3, 5,
					-- layer=2 filter=39 channel=121
					-5, -5, 6, -8, 2, 0, 0, -3, 9,
					-- layer=2 filter=39 channel=122
					-5, -8, -2, 6, 0, -4, -9, -9, -2,
					-- layer=2 filter=39 channel=123
					-36, 18, 27, -34, 25, 3, 3, 11, 11,
					-- layer=2 filter=39 channel=124
					19, 1, -33, 5, -26, 14, -37, -68, -3,
					-- layer=2 filter=39 channel=125
					3, 7, 5, -10, -3, 3, 2, 9, 13,
					-- layer=2 filter=39 channel=126
					-22, 22, -113, 31, 2, -26, -19, 33, -1,
					-- layer=2 filter=39 channel=127
					-31, -3, -6, 18, 14, 15, 8, 9, 23,
					-- layer=2 filter=40 channel=0
					-11, -11, -7, 0, 4, 22, 0, 13, -3,
					-- layer=2 filter=40 channel=1
					11, 2, -3, -39, -84, -28, -39, -30, -16,
					-- layer=2 filter=40 channel=2
					-3, 7, 6, 7, -9, 10, -11, 8, -9,
					-- layer=2 filter=40 channel=3
					14, 17, 5, 38, 32, 26, -12, 7, 23,
					-- layer=2 filter=40 channel=4
					-2, -20, -32, -4, -9, -52, -3, 6, -15,
					-- layer=2 filter=40 channel=5
					-8, -12, -2, 5, 0, 13, 32, 27, 3,
					-- layer=2 filter=40 channel=6
					4, -12, -29, -13, -18, 25, -9, -11, 20,
					-- layer=2 filter=40 channel=7
					1, 28, 50, 59, 23, 41, 9, 43, 65,
					-- layer=2 filter=40 channel=8
					-2, -4, -9, 8, 2, 4, -7, 9, 6,
					-- layer=2 filter=40 channel=9
					10, 12, -8, 13, 17, 13, 8, 11, -9,
					-- layer=2 filter=40 channel=10
					-6, 4, 2, 18, 19, 26, -6, 21, 17,
					-- layer=2 filter=40 channel=11
					9, -12, -4, 18, 0, -4, 3, 19, 14,
					-- layer=2 filter=40 channel=12
					21, 17, -4, 14, -5, 5, -2, -3, 34,
					-- layer=2 filter=40 channel=13
					9, -7, 3, -3, 8, -9, -2, -10, 2,
					-- layer=2 filter=40 channel=14
					20, 9, -8, -25, -33, -21, -21, -18, -17,
					-- layer=2 filter=40 channel=15
					16, 28, -57, 32, -43, -26, 5, 43, 17,
					-- layer=2 filter=40 channel=16
					-26, -35, -30, -63, -31, -51, -77, -13, -25,
					-- layer=2 filter=40 channel=17
					-1, -4, 4, -6, 4, 6, 6, 7, 10,
					-- layer=2 filter=40 channel=18
					-25, -47, -66, -39, -24, -50, 0, -27, -38,
					-- layer=2 filter=40 channel=19
					-30, -23, -33, -21, -77, -53, 3, -10, -12,
					-- layer=2 filter=40 channel=20
					3, 5, 7, -2, 7, -5, 1, 0, -7,
					-- layer=2 filter=40 channel=21
					7, 10, 15, 2, -6, 5, 1, 10, 9,
					-- layer=2 filter=40 channel=22
					2, -8, 6, -1, -9, 1, 10, 5, 8,
					-- layer=2 filter=40 channel=23
					-8, 40, 15, -59, 9, -16, -45, -50, -26,
					-- layer=2 filter=40 channel=24
					0, 1, 22, 25, 30, 35, -3, 1, 0,
					-- layer=2 filter=40 channel=25
					-2, 17, 9, 16, 34, 19, -7, 20, 26,
					-- layer=2 filter=40 channel=26
					0, 1, -8, 7, -10, -7, -5, -1, -2,
					-- layer=2 filter=40 channel=27
					-35, -17, -42, -33, -37, -44, 1, -8, -21,
					-- layer=2 filter=40 channel=28
					4, 5, -1, 7, 25, 59, 63, -6, -5,
					-- layer=2 filter=40 channel=29
					-2, 3, -6, 0, -5, 4, -11, 8, 7,
					-- layer=2 filter=40 channel=30
					13, -6, -19, -81, -67, -47, -29, -42, -46,
					-- layer=2 filter=40 channel=31
					17, -6, 40, 16, 35, -7, 46, 66, 13,
					-- layer=2 filter=40 channel=32
					6, 4, 0, -1, 4, -9, -4, -6, -7,
					-- layer=2 filter=40 channel=33
					43, 5, 28, 29, -22, -37, -14, -31, 18,
					-- layer=2 filter=40 channel=34
					26, -35, 0, 10, 17, -37, -5, -63, 0,
					-- layer=2 filter=40 channel=35
					-11, -3, -6, 5, 9, -15, 20, -26, -17,
					-- layer=2 filter=40 channel=36
					16, 4, 11, 4, 9, 18, -6, 8, 19,
					-- layer=2 filter=40 channel=37
					9, 7, -9, 18, -4, -13, 14, 10, 4,
					-- layer=2 filter=40 channel=38
					-2, -17, -24, -47, -38, -72, 6, 8, -38,
					-- layer=2 filter=40 channel=39
					-16, 5, 17, -25, -28, -34, -69, -20, 0,
					-- layer=2 filter=40 channel=40
					-17, -20, -21, 7, 42, -26, 66, -24, -4,
					-- layer=2 filter=40 channel=41
					7, -2, 3, -1, 9, -1, 8, 0, -3,
					-- layer=2 filter=40 channel=42
					0, 39, 19, -59, 12, -2, -14, 14, -33,
					-- layer=2 filter=40 channel=43
					-8, -22, -15, 23, 7, -22, 24, -4, -30,
					-- layer=2 filter=40 channel=44
					-10, -7, -1, -7, 3, 9, -9, 8, -3,
					-- layer=2 filter=40 channel=45
					-21, -47, -15, 11, 16, -28, -86, -37, -61,
					-- layer=2 filter=40 channel=46
					-9, -17, -30, -18, -4, -34, -14, -10, -20,
					-- layer=2 filter=40 channel=47
					-30, 15, 28, 28, 22, 6, 24, 27, 5,
					-- layer=2 filter=40 channel=48
					7, 0, -6, -5, -7, 7, 0, -3, 6,
					-- layer=2 filter=40 channel=49
					-16, -18, -42, -26, -33, -45, -28, -18, -46,
					-- layer=2 filter=40 channel=50
					-16, -9, -6, 13, 6, -1, 18, 26, 11,
					-- layer=2 filter=40 channel=51
					-2, 8, -6, 8, 3, 11, 8, 22, -7,
					-- layer=2 filter=40 channel=52
					19, -2, 3, 33, 0, -27, 32, 15, 14,
					-- layer=2 filter=40 channel=53
					-29, -25, -12, -48, -27, -32, -16, -52, 10,
					-- layer=2 filter=40 channel=54
					-20, 11, 0, 20, -14, 9, 20, 22, 23,
					-- layer=2 filter=40 channel=55
					-3, -2, -5, 1, -4, -10, -3, -8, 7,
					-- layer=2 filter=40 channel=56
					0, -5, -6, -3, -7, 5, 7, 1, 4,
					-- layer=2 filter=40 channel=57
					-9, 6, -7, 4, -15, -6, -10, 8, 3,
					-- layer=2 filter=40 channel=58
					2, -2, 2, 25, 0, -6, 29, 30, 28,
					-- layer=2 filter=40 channel=59
					-3, -21, -49, -11, -16, -104, -25, 3, -19,
					-- layer=2 filter=40 channel=60
					-30, 0, -1, 5, -60, -29, 25, 39, 0,
					-- layer=2 filter=40 channel=61
					-47, 3, 26, -29, -71, 21, -6, 9, -20,
					-- layer=2 filter=40 channel=62
					18, 0, -43, -23, 6, -16, -11, -8, -16,
					-- layer=2 filter=40 channel=63
					-25, 20, 3, -36, -30, -30, -26, -9, -7,
					-- layer=2 filter=40 channel=64
					2, 22, 26, -44, -4, 0, -44, -2, 6,
					-- layer=2 filter=40 channel=65
					-20, 14, -18, -53, -22, 25, 25, 10, 7,
					-- layer=2 filter=40 channel=66
					-5, 7, 3, 9, -19, -32, -3, -10, -9,
					-- layer=2 filter=40 channel=67
					-39, -25, -14, -55, -6, -18, -59, -23, -24,
					-- layer=2 filter=40 channel=68
					-2, 1, -11, -6, -11, -9, -9, 2, -8,
					-- layer=2 filter=40 channel=69
					32, 57, 41, -63, -7, -15, -74, 22, -14,
					-- layer=2 filter=40 channel=70
					-11, -18, -2, 0, 17, 27, 62, 9, 18,
					-- layer=2 filter=40 channel=71
					-53, -9, -14, -28, -17, -16, -12, -13, -21,
					-- layer=2 filter=40 channel=72
					49, 21, 44, 3, -7, 26, 41, -13, 40,
					-- layer=2 filter=40 channel=73
					36, 19, 57, 39, 10, 35, -28, 25, -1,
					-- layer=2 filter=40 channel=74
					-32, -2, 28, -65, -56, -40, -44, -21, -35,
					-- layer=2 filter=40 channel=75
					-45, -28, -39, 49, -7, 32, -26, -39, -3,
					-- layer=2 filter=40 channel=76
					-15, 10, 18, 53, 22, -38, -28, 16, -33,
					-- layer=2 filter=40 channel=77
					7, 7, -3, 3, -2, -10, 3, -5, 1,
					-- layer=2 filter=40 channel=78
					-2, 0, -5, 39, 3, 10, 4, 21, 17,
					-- layer=2 filter=40 channel=79
					-3, 7, 3, -11, -8, 5, -1, -4, -1,
					-- layer=2 filter=40 channel=80
					-13, -11, 2, -15, 0, -33, -72, -37, -13,
					-- layer=2 filter=40 channel=81
					-3, -17, -4, -13, -15, -7, -7, -7, -5,
					-- layer=2 filter=40 channel=82
					-5, -7, -5, 4, 6, 7, -7, 9, 10,
					-- layer=2 filter=40 channel=83
					-42, 19, -23, -79, 10, -6, -23, -66, -11,
					-- layer=2 filter=40 channel=84
					1, -3, -5, 3, 3, 8, 7, -6, 8,
					-- layer=2 filter=40 channel=85
					0, 0, -9, -2, 0, -4, -11, -14, 0,
					-- layer=2 filter=40 channel=86
					3, 0, 2, 4, -11, -10, 1, 3, 9,
					-- layer=2 filter=40 channel=87
					-7, 21, -33, -21, -9, -48, 13, -38, -33,
					-- layer=2 filter=40 channel=88
					29, 26, 24, -74, -46, -24, -36, -55, -29,
					-- layer=2 filter=40 channel=89
					20, 20, 9, -14, -28, -24, -8, 11, -1,
					-- layer=2 filter=40 channel=90
					10, -5, -3, 1, -7, -6, 9, -10, 8,
					-- layer=2 filter=40 channel=91
					-8, -14, 5, 11, -14, 9, 3, -12, 24,
					-- layer=2 filter=40 channel=92
					7, 14, 17, -28, -24, -10, 4, -2, -4,
					-- layer=2 filter=40 channel=93
					31, 65, -21, -37, 20, -4, 7, 45, 26,
					-- layer=2 filter=40 channel=94
					3, -7, 16, -13, -58, 19, 54, 24, 0,
					-- layer=2 filter=40 channel=95
					-11, -19, -22, -18, 5, -12, 7, -12, -13,
					-- layer=2 filter=40 channel=96
					25, 18, 10, 14, -31, -25, 14, -31, -11,
					-- layer=2 filter=40 channel=97
					10, 2, -30, 22, -11, 6, 0, 14, -11,
					-- layer=2 filter=40 channel=98
					-28, 0, 21, 35, 14, 27, 48, 13, 11,
					-- layer=2 filter=40 channel=99
					-6, 10, -2, 51, -22, 23, 5, 24, 5,
					-- layer=2 filter=40 channel=100
					-14, 22, 20, 10, 9, 0, 19, 23, -22,
					-- layer=2 filter=40 channel=101
					-30, -18, 4, -4, 12, -2, -7, 7, 9,
					-- layer=2 filter=40 channel=102
					0, -2, -56, -33, -18, -80, -20, -8, -32,
					-- layer=2 filter=40 channel=103
					-54, -53, 7, -30, 36, 33, -2, 0, 23,
					-- layer=2 filter=40 channel=104
					-8, -57, -25, -28, -62, -48, -3, -61, -46,
					-- layer=2 filter=40 channel=105
					-31, -18, -39, 27, 2, -42, -40, 40, -31,
					-- layer=2 filter=40 channel=106
					-19, -19, -3, 3, 2, -1, -22, 18, 17,
					-- layer=2 filter=40 channel=107
					32, -4, 45, 8, 61, 13, -60, 14, -36,
					-- layer=2 filter=40 channel=108
					-25, -16, -31, -39, -51, -72, -13, 3, -23,
					-- layer=2 filter=40 channel=109
					10, 6, -4, 19, -1, -9, 20, 3, -1,
					-- layer=2 filter=40 channel=110
					-8, 23, 16, -56, 2, 13, -48, -33, 0,
					-- layer=2 filter=40 channel=111
					-14, 3, 0, 1, -5, 5, 10, -5, -5,
					-- layer=2 filter=40 channel=112
					-12, 19, 2, -7, 2, 21, 8, 26, 24,
					-- layer=2 filter=40 channel=113
					-19, -34, -3, -106, -42, -46, -14, -49, -16,
					-- layer=2 filter=40 channel=114
					-19, -16, 0, -8, 1, -12, -18, -5, -14,
					-- layer=2 filter=40 channel=115
					-5, 2, 7, -3, 2, -6, 9, 10, 5,
					-- layer=2 filter=40 channel=116
					2, 9, -29, -23, -31, -43, 29, -26, -14,
					-- layer=2 filter=40 channel=117
					9, 14, 40, 22, 4, 21, -27, -4, 27,
					-- layer=2 filter=40 channel=118
					-4, 0, 2, 35, 29, 28, -8, -5, -20,
					-- layer=2 filter=40 channel=119
					0, -30, -62, -45, 0, -29, -26, -49, -74,
					-- layer=2 filter=40 channel=120
					7, 4, -4, -7, -5, 1, -6, 0, 7,
					-- layer=2 filter=40 channel=121
					0, -5, -5, 9, 2, -7, -2, 11, 7,
					-- layer=2 filter=40 channel=122
					-15, 6, 5, -1, -4, -8, -14, 2, 2,
					-- layer=2 filter=40 channel=123
					31, 63, 56, 44, 11, 15, 17, 24, 25,
					-- layer=2 filter=40 channel=124
					34, 41, -5, 24, 7, -31, -9, 11, -22,
					-- layer=2 filter=40 channel=125
					0, 1, -2, -3, -2, 0, -5, 10, -4,
					-- layer=2 filter=40 channel=126
					15, -35, 22, -5, -38, -34, -39, -63, -39,
					-- layer=2 filter=40 channel=127
					35, 14, 19, -69, -39, -62, -15, -37, 8,
					-- layer=2 filter=41 channel=0
					-23, 0, -24, -7, 17, -24, 24, -1, -4,
					-- layer=2 filter=41 channel=1
					-10, 7, -16, -14, 6, -32, -2, -9, -4,
					-- layer=2 filter=41 channel=2
					1, 3, -1, 8, 4, 8, 7, -4, 6,
					-- layer=2 filter=41 channel=3
					12, 0, -13, -6, 20, -16, -8, 41, 41,
					-- layer=2 filter=41 channel=4
					23, 5, -8, -23, 7, -7, -16, -51, -34,
					-- layer=2 filter=41 channel=5
					-11, -30, -29, -12, -39, -24, 4, -63, -22,
					-- layer=2 filter=41 channel=6
					-66, 13, 5, -9, 48, 12, -4, 43, 47,
					-- layer=2 filter=41 channel=7
					32, 41, -6, 29, 15, -3, -14, -93, -32,
					-- layer=2 filter=41 channel=8
					-2, 5, 6, -4, 8, -9, 9, 1, -4,
					-- layer=2 filter=41 channel=9
					-36, -58, -20, 1, -16, -20, -7, 5, -8,
					-- layer=2 filter=41 channel=10
					0, -20, -24, 23, 4, -7, 2, -3, 6,
					-- layer=2 filter=41 channel=11
					3, -33, -18, -26, -54, -54, -4, -18, -18,
					-- layer=2 filter=41 channel=12
					15, 19, -27, 10, 35, -12, -42, -23, 9,
					-- layer=2 filter=41 channel=13
					9, -8, 0, 4, -5, 3, 0, 6, 3,
					-- layer=2 filter=41 channel=14
					7, 29, -3, -5, 3, -23, 10, -6, -1,
					-- layer=2 filter=41 channel=15
					12, -2, -34, 25, 25, -34, 45, -78, -47,
					-- layer=2 filter=41 channel=16
					-23, -38, 2, 12, 19, 38, -3, 0, 56,
					-- layer=2 filter=41 channel=17
					-3, -7, -8, 9, 3, 5, 1, -10, 0,
					-- layer=2 filter=41 channel=18
					4, 6, -36, -24, 6, -9, 12, 17, -27,
					-- layer=2 filter=41 channel=19
					-16, 21, -2, 0, 29, -7, 17, -9, -3,
					-- layer=2 filter=41 channel=20
					7, -7, 0, -10, 7, 2, 0, 0, 0,
					-- layer=2 filter=41 channel=21
					-2, -1, 10, -7, -13, 0, -14, -8, 9,
					-- layer=2 filter=41 channel=22
					10, -9, -2, -4, 1, -8, -3, -5, -1,
					-- layer=2 filter=41 channel=23
					-3, 5, 1, 31, 12, 40, 19, -11, 9,
					-- layer=2 filter=41 channel=24
					-18, -21, -5, -16, 24, 1, 0, 34, 40,
					-- layer=2 filter=41 channel=25
					-10, -9, 1, -31, 21, 2, -3, 46, 25,
					-- layer=2 filter=41 channel=26
					1, -5, -5, -4, 0, -1, 4, 9, 4,
					-- layer=2 filter=41 channel=27
					-14, -8, 51, -36, -68, 26, -52, -91, -32,
					-- layer=2 filter=41 channel=28
					-7, -13, 8, -3, 31, 2, -63, 13, -8,
					-- layer=2 filter=41 channel=29
					-5, 3, 8, 11, 9, 3, -3, 2, 7,
					-- layer=2 filter=41 channel=30
					-17, 0, -11, -7, 0, 17, 17, -34, 2,
					-- layer=2 filter=41 channel=31
					28, 51, -15, 56, -13, -47, 28, -71, 36,
					-- layer=2 filter=41 channel=32
					-5, -8, -7, 8, -7, 10, -3, -1, -3,
					-- layer=2 filter=41 channel=33
					-32, 19, -5, -57, -16, -22, -37, -15, -63,
					-- layer=2 filter=41 channel=34
					-35, -27, -40, -16, -28, -10, 11, 10, -50,
					-- layer=2 filter=41 channel=35
					-26, -5, 3, 32, 34, 26, -40, -29, -35,
					-- layer=2 filter=41 channel=36
					-7, 1, 9, -6, -6, 11, -14, -12, -5,
					-- layer=2 filter=41 channel=37
					0, -24, 0, -7, -47, -40, 8, -44, -26,
					-- layer=2 filter=41 channel=38
					-3, -7, 27, -1, -53, 2, 24, -6, -22,
					-- layer=2 filter=41 channel=39
					29, 1, -15, -19, -6, -31, 6, -26, 24,
					-- layer=2 filter=41 channel=40
					95, 0, -29, 34, 33, -22, 31, 50, 4,
					-- layer=2 filter=41 channel=41
					0, -2, -11, -6, 1, -3, 4, -2, -4,
					-- layer=2 filter=41 channel=42
					23, -8, 24, 26, 24, 26, 11, 30, 51,
					-- layer=2 filter=41 channel=43
					-43, -13, -29, 0, 3, 20, -28, 3, 11,
					-- layer=2 filter=41 channel=44
					-6, -8, 4, 0, -9, 2, 3, 10, -8,
					-- layer=2 filter=41 channel=45
					5, 23, 31, -12, -34, -6, -22, -37, 44,
					-- layer=2 filter=41 channel=46
					-5, -24, -25, -34, -59, 11, -1, -22, 2,
					-- layer=2 filter=41 channel=47
					8, 6, 27, 27, 9, 3, -61, -32, -23,
					-- layer=2 filter=41 channel=48
					-2, 2, 4, -9, -9, 8, 11, -2, 8,
					-- layer=2 filter=41 channel=49
					5, 28, 46, -13, 15, 12, 25, 49, 65,
					-- layer=2 filter=41 channel=50
					15, -2, 14, 11, 0, -2, 10, 18, 11,
					-- layer=2 filter=41 channel=51
					-13, -20, -3, 7, -34, -42, -3, -9, -34,
					-- layer=2 filter=41 channel=52
					-22, -12, -48, -30, -26, -26, 28, -3, -89,
					-- layer=2 filter=41 channel=53
					-7, 10, 12, -14, -1, 0, 29, -41, 44,
					-- layer=2 filter=41 channel=54
					16, 24, -15, -2, 15, -14, 0, -25, -11,
					-- layer=2 filter=41 channel=55
					1, 0, -3, 2, -7, 0, -5, -8, 12,
					-- layer=2 filter=41 channel=56
					14, -12, -11, -13, -46, -52, -1, -15, -26,
					-- layer=2 filter=41 channel=57
					-3, -12, -5, -12, 14, -2, 0, -4, 17,
					-- layer=2 filter=41 channel=58
					5, 12, -5, 3, 20, -1, -46, -27, -1,
					-- layer=2 filter=41 channel=59
					3, 4, 11, -35, -4, 35, -14, -16, -16,
					-- layer=2 filter=41 channel=60
					20, 11, 4, 4, 3, -26, 5, 1, 11,
					-- layer=2 filter=41 channel=61
					-10, 48, 44, 5, 38, 21, 24, 58, 21,
					-- layer=2 filter=41 channel=62
					-37, -27, -13, -16, 3, -5, 13, 10, 13,
					-- layer=2 filter=41 channel=63
					36, -1, 4, -2, 16, 0, 1, -2, -24,
					-- layer=2 filter=41 channel=64
					-13, 6, -10, -4, 6, 8, 8, 11, 24,
					-- layer=2 filter=41 channel=65
					-40, -13, 28, -16, 14, -4, -2, 45, 9,
					-- layer=2 filter=41 channel=66
					-10, 40, 0, -22, 46, 41, 21, 13, 50,
					-- layer=2 filter=41 channel=67
					-12, -44, -44, -48, -70, -19, 27, -16, -4,
					-- layer=2 filter=41 channel=68
					5, 4, -1, -5, -9, 10, 6, -3, -5,
					-- layer=2 filter=41 channel=69
					1, -15, 3, -5, 27, 20, 18, 9, 53,
					-- layer=2 filter=41 channel=70
					-43, 13, -22, 1, 20, -4, -35, -12, -52,
					-- layer=2 filter=41 channel=71
					6, 24, 88, -23, -30, 104, -57, -72, 36,
					-- layer=2 filter=41 channel=72
					9, 44, 16, 28, 12, -7, 0, -11, -36,
					-- layer=2 filter=41 channel=73
					33, 30, -15, 27, -3, 50, 28, 33, 67,
					-- layer=2 filter=41 channel=74
					27, 1, -50, -7, -10, -27, 12, -3, -15,
					-- layer=2 filter=41 channel=75
					8, 38, 4, -17, -11, -4, 30, 35, -10,
					-- layer=2 filter=41 channel=76
					-3, -12, -37, 11, -53, -56, 35, -23, 13,
					-- layer=2 filter=41 channel=77
					5, 1, -12, -3, 4, 5, -3, 0, -6,
					-- layer=2 filter=41 channel=78
					-12, -18, -62, -19, -7, -45, -2, 11, -1,
					-- layer=2 filter=41 channel=79
					-4, -7, 6, -6, 3, 2, 4, -7, -2,
					-- layer=2 filter=41 channel=80
					18, 0, 4, -3, -7, -12, -14, 0, 24,
					-- layer=2 filter=41 channel=81
					2, 1, 4, 23, 8, -3, 13, -2, 0,
					-- layer=2 filter=41 channel=82
					5, -6, 2, 13, 2, 9, -4, -1, 0,
					-- layer=2 filter=41 channel=83
					-9, 2, -10, -10, 26, 31, -5, -22, 5,
					-- layer=2 filter=41 channel=84
					-3, 8, -5, 5, 0, 5, 0, -8, 11,
					-- layer=2 filter=41 channel=85
					5, -9, 14, 7, 10, 0, 3, -16, 0,
					-- layer=2 filter=41 channel=86
					7, -1, -5, 0, 0, -3, 13, 2, 11,
					-- layer=2 filter=41 channel=87
					-25, -23, -23, -11, -36, 20, -8, -49, -61,
					-- layer=2 filter=41 channel=88
					1, -12, -7, -19, 7, -13, 2, -13, -5,
					-- layer=2 filter=41 channel=89
					8, 15, -6, -4, 14, 9, -5, -34, 24,
					-- layer=2 filter=41 channel=90
					-10, -6, 0, -3, -10, 0, 6, -2, -7,
					-- layer=2 filter=41 channel=91
					-14, 18, -36, 0, 14, -12, -16, -5, 6,
					-- layer=2 filter=41 channel=92
					-7, 11, -23, -20, 6, -27, -34, -7, -4,
					-- layer=2 filter=41 channel=93
					-23, -49, -15, 16, -23, 1, -19, -27, -6,
					-- layer=2 filter=41 channel=94
					-17, 43, 36, -2, 55, 19, 4, 12, 41,
					-- layer=2 filter=41 channel=95
					-16, -12, 6, 10, -10, -7, 2, -10, -4,
					-- layer=2 filter=41 channel=96
					21, 2, 4, -1, 17, -16, 29, -3, -5,
					-- layer=2 filter=41 channel=97
					-33, -13, -36, -35, -12, -24, -4, 29, 7,
					-- layer=2 filter=41 channel=98
					0, 5, 2, 28, 22, -1, -22, -1, -38,
					-- layer=2 filter=41 channel=99
					-3, 12, 13, -20, -1, -10, -18, 7, 5,
					-- layer=2 filter=41 channel=100
					11, 10, -26, 0, -19, -12, 8, -24, -12,
					-- layer=2 filter=41 channel=101
					62, 30, 50, -31, -22, 29, -18, -20, -2,
					-- layer=2 filter=41 channel=102
					2, 10, 29, -23, 9, 14, -13, 9, 27,
					-- layer=2 filter=41 channel=103
					-42, -24, -6, 18, -10, -74, -40, 4, 11,
					-- layer=2 filter=41 channel=104
					15, -10, 1, -16, 23, -5, 5, -18, 4,
					-- layer=2 filter=41 channel=105
					-8, 2, 50, 53, 75, 11, 8, 36, -36,
					-- layer=2 filter=41 channel=106
					-23, -6, -16, -20, -34, -49, -23, -4, 8,
					-- layer=2 filter=41 channel=107
					-3, 14, -34, 35, 11, -48, -20, 41, -5,
					-- layer=2 filter=41 channel=108
					18, 2, 44, -8, -27, -27, -22, -65, -8,
					-- layer=2 filter=41 channel=109
					9, -14, 7, 12, 4, 4, 7, 0, 9,
					-- layer=2 filter=41 channel=110
					-16, 32, 15, -12, 39, 33, -3, 28, 31,
					-- layer=2 filter=41 channel=111
					5, -8, 6, 7, 7, 7, 7, -7, 9,
					-- layer=2 filter=41 channel=112
					4, -28, 42, 14, -1, 10, 10, 17, 31,
					-- layer=2 filter=41 channel=113
					18, 14, -8, 24, 26, 15, 4, 5, 21,
					-- layer=2 filter=41 channel=114
					-5, -5, -9, -3, 12, 6, 4, -17, 1,
					-- layer=2 filter=41 channel=115
					-9, 0, -4, 4, -4, 6, -4, 0, 9,
					-- layer=2 filter=41 channel=116
					-35, -24, -37, -17, -38, 23, -7, 0, -62,
					-- layer=2 filter=41 channel=117
					15, 25, -12, 27, 36, -29, 3, -24, -30,
					-- layer=2 filter=41 channel=118
					0, -29, -44, -37, -22, -16, 4, 5, 39,
					-- layer=2 filter=41 channel=119
					-23, 1, -1, -30, -11, -12, -26, -13, -5,
					-- layer=2 filter=41 channel=120
					-1, -7, -9, 5, -10, -9, 0, 2, 9,
					-- layer=2 filter=41 channel=121
					3, -12, -6, 1, 1, -2, 3, 7, -10,
					-- layer=2 filter=41 channel=122
					0, -8, 4, 5, 0, -3, 5, 0, 10,
					-- layer=2 filter=41 channel=123
					20, 10, -2, 17, 34, -15, 16, -16, -32,
					-- layer=2 filter=41 channel=124
					-13, -4, -32, 0, -7, 16, 41, -26, 23,
					-- layer=2 filter=41 channel=125
					6, 0, -6, -9, 8, -7, 3, 3, 6,
					-- layer=2 filter=41 channel=126
					-9, 23, 40, -12, 19, 2, -24, 31, 49,
					-- layer=2 filter=41 channel=127
					-6, -2, -6, -18, 4, -22, -13, -9, -1,
					-- layer=2 filter=42 channel=0
					-4, 9, -14, 56, 26, -21, 29, 26, -24,
					-- layer=2 filter=42 channel=1
					7, -11, 3, -20, -10, 15, 13, -12, 27,
					-- layer=2 filter=42 channel=2
					1, 4, -5, -7, 5, 10, 0, 0, -7,
					-- layer=2 filter=42 channel=3
					4, 16, 10, 9, -22, -13, -21, -32, -56,
					-- layer=2 filter=42 channel=4
					-13, -15, -16, -4, -6, -5, -35, -10, -4,
					-- layer=2 filter=42 channel=5
					11, 10, -25, 31, 25, -6, 6, 3, -19,
					-- layer=2 filter=42 channel=6
					5, -7, -58, 12, 3, -21, 0, -16, 14,
					-- layer=2 filter=42 channel=7
					-2, -6, 21, -32, -37, -23, 13, 19, 8,
					-- layer=2 filter=42 channel=8
					4, -5, 6, 3, 9, 6, -5, -7, 7,
					-- layer=2 filter=42 channel=9
					-2, 4, 38, -10, 27, 3, -28, -23, 33,
					-- layer=2 filter=42 channel=10
					13, 20, -2, 44, 40, 14, 1, 17, -15,
					-- layer=2 filter=42 channel=11
					-8, 15, -42, 16, 11, -47, 14, 2, -46,
					-- layer=2 filter=42 channel=12
					31, -7, -1, -25, -19, 3, 23, 6, -23,
					-- layer=2 filter=42 channel=13
					-5, 11, 5, -4, -5, 11, -4, -8, 0,
					-- layer=2 filter=42 channel=14
					16, 7, -7, -28, -12, -19, 0, -20, -12,
					-- layer=2 filter=42 channel=15
					11, -20, -32, 35, 41, -8, 42, 39, 26,
					-- layer=2 filter=42 channel=16
					-28, -42, 23, -54, -53, 30, -72, -25, 72,
					-- layer=2 filter=42 channel=17
					-6, 12, 0, 5, 3, -7, -5, 10, 7,
					-- layer=2 filter=42 channel=18
					-21, -6, 9, 6, 18, 7, -15, 2, -2,
					-- layer=2 filter=42 channel=19
					0, 1, 6, 1, 1, 17, -9, 30, 48,
					-- layer=2 filter=42 channel=20
					9, 1, -8, 2, -4, 1, 7, 0, 9,
					-- layer=2 filter=42 channel=21
					7, 14, -9, -2, -2, 0, 3, -15, 1,
					-- layer=2 filter=42 channel=22
					-4, -2, 9, -3, -11, 3, 4, 1, 10,
					-- layer=2 filter=42 channel=23
					-13, -22, 2, -8, -56, -19, -24, 11, 22,
					-- layer=2 filter=42 channel=24
					19, 13, -21, -4, -13, -22, -22, -64, -28,
					-- layer=2 filter=42 channel=25
					-16, 6, -102, -8, -9, -98, -15, -55, -99,
					-- layer=2 filter=42 channel=26
					-7, 5, -8, -6, -8, -3, 6, 6, 6,
					-- layer=2 filter=42 channel=27
					-12, 16, 3, 13, 25, 13, 13, 16, -23,
					-- layer=2 filter=42 channel=28
					14, -9, -25, 12, 14, -15, 11, 5, -1,
					-- layer=2 filter=42 channel=29
					-4, -10, -3, 1, -2, 0, -2, -3, 9,
					-- layer=2 filter=42 channel=30
					11, -32, 7, -24, 0, -8, 23, -39, 17,
					-- layer=2 filter=42 channel=31
					60, 8, 16, 94, 56, -13, 36, 26, 2,
					-- layer=2 filter=42 channel=32
					1, 7, -1, 2, 1, 10, -3, 7, 8,
					-- layer=2 filter=42 channel=33
					13, -6, -35, 13, -3, -16, 28, 7, -17,
					-- layer=2 filter=42 channel=34
					-25, 1, 40, -25, 35, -20, -3, 30, 20,
					-- layer=2 filter=42 channel=35
					7, -5, 21, 8, 23, 42, 7, 4, 20,
					-- layer=2 filter=42 channel=36
					5, -10, -1, 0, -5, 6, 5, -3, -12,
					-- layer=2 filter=42 channel=37
					-4, 19, -33, 22, 1, -26, 6, 5, -40,
					-- layer=2 filter=42 channel=38
					-1, 0, 1, 7, 4, 23, 22, 6, 8,
					-- layer=2 filter=42 channel=39
					-12, 9, 39, 5, -39, 17, -6, -15, 104,
					-- layer=2 filter=42 channel=40
					0, -3, 28, -1, 21, -50, 12, 14, 58,
					-- layer=2 filter=42 channel=41
					10, 0, 8, -1, -7, -3, 9, -6, -7,
					-- layer=2 filter=42 channel=42
					0, -39, 25, -29, -87, 28, -11, 5, 67,
					-- layer=2 filter=42 channel=43
					-19, 31, -18, -2, 28, -5, -18, 9, -27,
					-- layer=2 filter=42 channel=44
					8, 10, 2, 8, -8, 5, -11, -5, -5,
					-- layer=2 filter=42 channel=45
					8, 18, 17, -1, -11, 16, -5, 3, -36,
					-- layer=2 filter=42 channel=46
					14, -12, 20, 21, 17, 28, -10, 18, 22,
					-- layer=2 filter=42 channel=47
					-5, -18, -27, 1, 13, -46, 44, 5, -9,
					-- layer=2 filter=42 channel=48
					9, -7, -8, 8, 9, 0, 3, 10, 2,
					-- layer=2 filter=42 channel=49
					-26, 9, 29, -12, 1, 3, -29, -40, 25,
					-- layer=2 filter=42 channel=50
					-9, 2, -6, 14, -14, -2, 10, 12, 3,
					-- layer=2 filter=42 channel=51
					8, 4, -56, 33, 7, -37, 25, -4, -37,
					-- layer=2 filter=42 channel=52
					36, 3, -13, -20, 4, -21, -10, -9, 13,
					-- layer=2 filter=42 channel=53
					34, -8, 10, -14, -8, -37, 8, 22, 22,
					-- layer=2 filter=42 channel=54
					19, -8, -25, 14, -27, -13, 27, 9, -29,
					-- layer=2 filter=42 channel=55
					14, 9, -1, -9, 4, 13, 6, -4, -8,
					-- layer=2 filter=42 channel=56
					-13, 5, -40, 27, 24, -50, 15, 9, -58,
					-- layer=2 filter=42 channel=57
					-11, 8, 10, 0, -2, 8, 3, -1, 10,
					-- layer=2 filter=42 channel=58
					59, -5, 0, -8, 16, -9, 45, -1, -18,
					-- layer=2 filter=42 channel=59
					-11, 17, -5, -5, 11, 33, 29, 17, 19,
					-- layer=2 filter=42 channel=60
					7, 15, 30, 18, -9, 42, 35, 50, 31,
					-- layer=2 filter=42 channel=61
					5, 31, 28, -2, 15, 40, -3, 5, 33,
					-- layer=2 filter=42 channel=62
					-31, 20, -15, 0, -18, -25, -17, -7, 19,
					-- layer=2 filter=42 channel=63
					18, 7, 8, 30, -31, -7, 39, 11, 18,
					-- layer=2 filter=42 channel=64
					2, -20, 21, -17, -53, -8, -25, -33, 42,
					-- layer=2 filter=42 channel=65
					-2, -4, -5, 32, -4, 1, 0, 19, 26,
					-- layer=2 filter=42 channel=66
					-8, -7, -55, 38, 17, 21, 50, 1, 16,
					-- layer=2 filter=42 channel=67
					8, -12, -19, 1, -13, 1, 0, -6, 3,
					-- layer=2 filter=42 channel=68
					-6, -7, -7, -8, 11, -7, 8, -6, 8,
					-- layer=2 filter=42 channel=69
					-25, -11, 21, -35, -45, 17, -8, -8, 51,
					-- layer=2 filter=42 channel=70
					40, -8, 9, 22, 33, 31, 5, 11, 0,
					-- layer=2 filter=42 channel=71
					-10, 11, -9, -21, -13, -19, 3, 1, -49,
					-- layer=2 filter=42 channel=72
					29, 16, -26, 5, -22, -5, -1, 12, -11,
					-- layer=2 filter=42 channel=73
					15, 14, 62, -3, -4, 5, 32, 15, 29,
					-- layer=2 filter=42 channel=74
					28, -4, 7, 36, -4, 17, 28, 4, 31,
					-- layer=2 filter=42 channel=75
					3, -4, 10, 42, 60, 20, -28, -40, -41,
					-- layer=2 filter=42 channel=76
					31, -15, 6, -31, 26, 7, 3, 40, 17,
					-- layer=2 filter=42 channel=77
					-3, 10, -4, 0, -2, 3, -3, -6, -7,
					-- layer=2 filter=42 channel=78
					-18, 9, -57, 10, 20, -61, -24, -20, -37,
					-- layer=2 filter=42 channel=79
					1, -1, 7, -6, 10, 3, -6, 0, 6,
					-- layer=2 filter=42 channel=80
					23, -17, 14, -13, -5, 18, -47, -36, 45,
					-- layer=2 filter=42 channel=81
					-4, -14, 2, 0, 2, 0, 1, -6, -2,
					-- layer=2 filter=42 channel=82
					5, 2, 6, 12, 0, -4, 0, 7, -7,
					-- layer=2 filter=42 channel=83
					29, -13, 23, -21, -22, 0, -31, -34, 11,
					-- layer=2 filter=42 channel=84
					8, 11, -4, -3, -5, 8, -5, 3, 4,
					-- layer=2 filter=42 channel=85
					12, -3, 0, 1, 13, 5, -4, 9, -1,
					-- layer=2 filter=42 channel=86
					-9, 15, 10, 7, 2, 24, 7, 8, 1,
					-- layer=2 filter=42 channel=87
					-26, -15, 10, -32, 11, -18, 21, 28, 55,
					-- layer=2 filter=42 channel=88
					-19, -16, 13, 23, -19, 2, 12, 4, 23,
					-- layer=2 filter=42 channel=89
					-12, 5, -24, -22, -11, -21, -19, -21, -1,
					-- layer=2 filter=42 channel=90
					6, 1, -7, -1, 1, 5, 4, 2, 5,
					-- layer=2 filter=42 channel=91
					44, -19, 18, -22, 10, 35, 26, 22, 16,
					-- layer=2 filter=42 channel=92
					-7, -6, -9, -25, -36, 7, -17, 2, 30,
					-- layer=2 filter=42 channel=93
					35, 8, -47, 57, -5, -31, -33, -16, -32,
					-- layer=2 filter=42 channel=94
					4, 0, -23, -43, -4, -28, -25, -23, 34,
					-- layer=2 filter=42 channel=95
					-11, 3, -9, 1, -2, 3, 0, -3, -7,
					-- layer=2 filter=42 channel=96
					-2, 21, -31, -21, 34, -21, -1, -13, 6,
					-- layer=2 filter=42 channel=97
					19, -10, 9, 22, -30, -13, -5, -24, -24,
					-- layer=2 filter=42 channel=98
					4, -15, 3, 17, 9, -42, -5, 12, -4,
					-- layer=2 filter=42 channel=99
					11, -6, -12, -16, -17, -16, 8, 17, 21,
					-- layer=2 filter=42 channel=100
					20, -1, -6, 14, -9, 47, 6, 10, 37,
					-- layer=2 filter=42 channel=101
					0, 9, -40, 2, -26, -37, 7, 8, -69,
					-- layer=2 filter=42 channel=102
					-2, -7, 5, -15, 0, 29, -10, -15, 5,
					-- layer=2 filter=42 channel=103
					-32, -40, -7, 1, -11, 8, -11, 21, 7,
					-- layer=2 filter=42 channel=104
					-13, 30, 3, 0, 8, 0, 23, 15, 14,
					-- layer=2 filter=42 channel=105
					-16, 3, 23, -23, -14, 37, -1, 61, 45,
					-- layer=2 filter=42 channel=106
					23, 14, -30, 43, -15, -46, 28, 11, -31,
					-- layer=2 filter=42 channel=107
					-41, -46, 26, -4, -17, 57, 27, -7, 37,
					-- layer=2 filter=42 channel=108
					-6, 7, -15, -1, 19, -4, -19, -14, -2,
					-- layer=2 filter=42 channel=109
					-2, -7, -10, 2, -8, -2, -10, 2, -10,
					-- layer=2 filter=42 channel=110
					8, -32, -5, -1, -50, -35, -37, -13, 37,
					-- layer=2 filter=42 channel=111
					12, 8, 8, -3, -6, -7, -1, -2, -2,
					-- layer=2 filter=42 channel=112
					49, -7, -40, 53, 20, -8, 29, 6, -8,
					-- layer=2 filter=42 channel=113
					26, -41, 19, 20, -52, -4, 11, -12, 20,
					-- layer=2 filter=42 channel=114
					-1, -5, -5, 19, 4, 3, 9, 5, -3,
					-- layer=2 filter=42 channel=115
					-8, 3, 0, 5, -9, -1, -2, -3, -1,
					-- layer=2 filter=42 channel=116
					-7, -5, 14, 1, 23, -15, 22, 12, 37,
					-- layer=2 filter=42 channel=117
					-17, 11, 11, -65, -13, -3, 16, 17, 15,
					-- layer=2 filter=42 channel=118
					-5, -2, -3, 22, 32, -7, -24, -6, -11,
					-- layer=2 filter=42 channel=119
					-31, -20, 28, -15, -10, 57, -29, -50, 10,
					-- layer=2 filter=42 channel=120
					-2, 6, 1, -4, 3, 5, -1, 6, 8,
					-- layer=2 filter=42 channel=121
					-5, -3, 1, 10, -8, 0, 12, -8, 6,
					-- layer=2 filter=42 channel=122
					-4, 4, -2, 6, -1, -7, 5, 2, 16,
					-- layer=2 filter=42 channel=123
					38, 2, -17, -2, -32, -26, 21, 20, -3,
					-- layer=2 filter=42 channel=124
					23, -42, 2, -23, -25, 4, 0, -5, 65,
					-- layer=2 filter=42 channel=125
					8, 2, -1, 1, 8, 0, -8, 10, 9,
					-- layer=2 filter=42 channel=126
					-28, 17, -28, -28, -38, -7, 17, -28, -35,
					-- layer=2 filter=42 channel=127
					-11, -10, 10, -27, 17, 1, 10, 8, 8,
					-- layer=2 filter=43 channel=0
					26, -16, -14, 3, 11, 18, -20, 24, 27,
					-- layer=2 filter=43 channel=1
					3, 6, 16, 0, -7, 11, 7, -21, 9,
					-- layer=2 filter=43 channel=2
					-7, 4, -7, -4, 1, 1, 8, 10, 4,
					-- layer=2 filter=43 channel=3
					-11, -9, -2, 25, 0, -3, 41, 20, 18,
					-- layer=2 filter=43 channel=4
					11, -15, -1, -12, -52, -11, -31, -9, -30,
					-- layer=2 filter=43 channel=5
					-10, 13, 17, 0, 13, 31, -14, -14, 15,
					-- layer=2 filter=43 channel=6
					24, 22, -13, -18, 0, -22, -38, -20, 14,
					-- layer=2 filter=43 channel=7
					-29, -80, 55, -34, -41, -17, 12, 20, -14,
					-- layer=2 filter=43 channel=8
					8, 9, -3, -4, 3, 4, 11, -6, 6,
					-- layer=2 filter=43 channel=9
					-6, 13, 41, 26, 10, 8, 24, 27, -8,
					-- layer=2 filter=43 channel=10
					18, 12, 0, 11, 10, 13, 0, -3, -10,
					-- layer=2 filter=43 channel=11
					-2, -3, 5, -19, 7, 5, -18, 1, 23,
					-- layer=2 filter=43 channel=12
					-23, 6, 48, 11, -17, 15, 2, -17, 6,
					-- layer=2 filter=43 channel=13
					-4, -5, 1, -7, 9, -2, -8, 5, 7,
					-- layer=2 filter=43 channel=14
					-19, -10, 29, -8, -34, -15, -2, -41, 29,
					-- layer=2 filter=43 channel=15
					18, -14, -36, -60, -15, 4, 17, 67, 0,
					-- layer=2 filter=43 channel=16
					-16, -24, -48, -32, -27, -30, 23, 0, -18,
					-- layer=2 filter=43 channel=17
					0, -5, -10, -7, 5, 10, -10, 7, 0,
					-- layer=2 filter=43 channel=18
					18, 7, -21, -35, -25, 0, 34, -44, -19,
					-- layer=2 filter=43 channel=19
					16, 22, 18, -34, -16, -6, 58, 39, 45,
					-- layer=2 filter=43 channel=20
					-8, 5, -10, -8, -4, -2, 2, 7, -7,
					-- layer=2 filter=43 channel=21
					7, 6, 5, -3, 4, 4, -6, 1, 11,
					-- layer=2 filter=43 channel=22
					10, -6, 9, -8, 11, -4, -8, -9, -1,
					-- layer=2 filter=43 channel=23
					16, 10, 8, -12, -12, -1, 0, 0, -7,
					-- layer=2 filter=43 channel=24
					-7, 4, -16, 20, 29, 11, 31, 52, 42,
					-- layer=2 filter=43 channel=25
					-47, -24, -18, -6, 21, 9, 8, 25, 45,
					-- layer=2 filter=43 channel=26
					4, -5, 6, 9, -1, -3, 0, -8, 0,
					-- layer=2 filter=43 channel=27
					-1, 13, 52, -15, -15, 20, -23, -40, -9,
					-- layer=2 filter=43 channel=28
					-31, -90, -89, -21, -39, 12, -15, -12, 11,
					-- layer=2 filter=43 channel=29
					-5, 1, 1, 0, 0, -1, 0, 2, -9,
					-- layer=2 filter=43 channel=30
					0, 8, 11, 3, 8, -21, -28, -6, -14,
					-- layer=2 filter=43 channel=31
					-44, -41, 27, -15, -22, -5, -16, 63, 18,
					-- layer=2 filter=43 channel=32
					-9, -11, 0, -8, 4, 8, -3, 2, -10,
					-- layer=2 filter=43 channel=33
					-71, -63, 5, -90, -83, -37, 12, 12, -17,
					-- layer=2 filter=43 channel=34
					-17, 4, -4, -32, -126, 0, -62, -37, 11,
					-- layer=2 filter=43 channel=35
					-25, -82, -77, -57, -60, -12, -15, -11, -43,
					-- layer=2 filter=43 channel=36
					9, 6, -4, -8, -9, 7, 0, -6, 4,
					-- layer=2 filter=43 channel=37
					5, 20, 8, -26, -14, -5, -14, 0, 10,
					-- layer=2 filter=43 channel=38
					-5, 12, 42, 3, -11, 17, -15, -41, -6,
					-- layer=2 filter=43 channel=39
					25, 10, 4, 27, 8, 11, -25, -18, -50,
					-- layer=2 filter=43 channel=40
					-10, -22, -36, -66, 21, 24, -10, 12, -2,
					-- layer=2 filter=43 channel=41
					3, 1, -9, -5, -4, 2, -6, 6, -6,
					-- layer=2 filter=43 channel=42
					28, 24, 42, 24, 1, 12, 20, 30, -8,
					-- layer=2 filter=43 channel=43
					10, 31, 17, 18, 36, 1, -12, -13, -41,
					-- layer=2 filter=43 channel=44
					10, -2, -3, 2, -7, 0, 2, -6, -9,
					-- layer=2 filter=43 channel=45
					-41, -15, 21, -20, -5, 35, 36, 26, 52,
					-- layer=2 filter=43 channel=46
					6, -4, 2, 9, 0, -10, -10, 13, -40,
					-- layer=2 filter=43 channel=47
					-32, -23, -37, 9, -14, 51, -13, 9, 32,
					-- layer=2 filter=43 channel=48
					-3, 6, 0, 8, -4, 4, -8, 4, 7,
					-- layer=2 filter=43 channel=49
					-17, 53, 20, -33, 30, 24, 14, -16, 26,
					-- layer=2 filter=43 channel=50
					-2, 7, -8, 9, -1, -2, -19, -22, 2,
					-- layer=2 filter=43 channel=51
					11, -9, 1, 0, 14, 19, 15, 16, 27,
					-- layer=2 filter=43 channel=52
					-1, 3, 11, -22, 12, 10, -16, -3, -17,
					-- layer=2 filter=43 channel=53
					44, -12, -20, 17, 16, -33, 13, 0, 15,
					-- layer=2 filter=43 channel=54
					-52, -62, -75, -62, -76, -13, -8, -10, 19,
					-- layer=2 filter=43 channel=55
					-13, -4, -8, 2, 0, 8, 0, -5, -12,
					-- layer=2 filter=43 channel=56
					10, 14, 11, 14, 39, 12, -1, 13, 8,
					-- layer=2 filter=43 channel=57
					-7, 9, -9, -6, 15, -4, -2, 3, 4,
					-- layer=2 filter=43 channel=58
					-7, -15, 19, 19, -38, 9, 0, -30, -21,
					-- layer=2 filter=43 channel=59
					-14, -1, 45, -4, 2, -6, 3, -15, -18,
					-- layer=2 filter=43 channel=60
					25, 9, -61, 22, 5, -3, 3, -45, 12,
					-- layer=2 filter=43 channel=61
					47, 28, -60, 35, 17, -7, 10, 32, 31,
					-- layer=2 filter=43 channel=62
					13, 27, -18, -48, -34, -36, -32, -24, 3,
					-- layer=2 filter=43 channel=63
					10, 4, -4, 22, 2, -23, -25, -21, -29,
					-- layer=2 filter=43 channel=64
					18, 7, 21, 12, 1, -11, -1, -7, -11,
					-- layer=2 filter=43 channel=65
					47, 25, -33, 38, 3, -27, 8, -19, -1,
					-- layer=2 filter=43 channel=66
					16, -18, -12, 35, -33, 1, 59, 28, 53,
					-- layer=2 filter=43 channel=67
					0, 13, 6, 5, 35, 4, 10, 17, -16,
					-- layer=2 filter=43 channel=68
					6, -8, 11, -3, 7, 8, 8, -7, 9,
					-- layer=2 filter=43 channel=69
					29, 13, 11, 26, 8, 16, 7, -13, 0,
					-- layer=2 filter=43 channel=70
					-33, -68, -85, -55, -87, -14, -29, -24, -38,
					-- layer=2 filter=43 channel=71
					25, 27, 53, -10, -14, -6, -6, -21, 24,
					-- layer=2 filter=43 channel=72
					-71, 13, 0, -58, -30, 4, 9, 11, -5,
					-- layer=2 filter=43 channel=73
					-5, -2, -1, 7, 23, 35, 52, 79, 60,
					-- layer=2 filter=43 channel=74
					1, -2, 1, 20, 15, -9, -21, 5, -32,
					-- layer=2 filter=43 channel=75
					-35, -31, 3, -11, 18, 35, 11, -1, 40,
					-- layer=2 filter=43 channel=76
					44, -39, -4, 0, 12, 64, 12, -20, 1,
					-- layer=2 filter=43 channel=77
					-5, -10, -7, 2, 1, -8, -4, -8, 6,
					-- layer=2 filter=43 channel=78
					-7, 15, 7, -4, -1, -14, 15, 9, -4,
					-- layer=2 filter=43 channel=79
					7, -1, 11, 9, 9, -6, 2, -5, 11,
					-- layer=2 filter=43 channel=80
					18, 6, -1, 13, -11, 17, 1, 0, -18,
					-- layer=2 filter=43 channel=81
					0, 3, 5, 3, 0, 19, 8, 3, 11,
					-- layer=2 filter=43 channel=82
					6, 4, -7, -2, 8, 1, -6, 1, 3,
					-- layer=2 filter=43 channel=83
					12, -2, 10, -5, -13, -6, -1, -7, 4,
					-- layer=2 filter=43 channel=84
					5, 7, -4, 3, -9, -6, 7, 3, 11,
					-- layer=2 filter=43 channel=85
					-2, 12, 5, 11, 8, 11, 3, 17, 10,
					-- layer=2 filter=43 channel=86
					-23, 6, -11, -18, -2, -4, 8, -8, -10,
					-- layer=2 filter=43 channel=87
					-8, -77, -10, -27, -82, -10, -28, -2, -18,
					-- layer=2 filter=43 channel=88
					3, 6, 23, 16, 7, -9, -37, -16, -1,
					-- layer=2 filter=43 channel=89
					-25, -9, 26, -3, -6, 9, 23, -2, 43,
					-- layer=2 filter=43 channel=90
					0, -7, 6, -3, -5, 6, 5, 1, 2,
					-- layer=2 filter=43 channel=91
					-8, 15, 39, 3, -9, 26, 34, 9, 35,
					-- layer=2 filter=43 channel=92
					2, 7, 30, -21, -17, 7, 5, -22, 5,
					-- layer=2 filter=43 channel=93
					53, -16, 4, 56, -4, -36, 38, -46, -19,
					-- layer=2 filter=43 channel=94
					40, 14, -23, 16, -10, -35, -4, 21, -8,
					-- layer=2 filter=43 channel=95
					-4, -15, 1, -16, -3, -5, -8, -6, -17,
					-- layer=2 filter=43 channel=96
					-2, -4, -40, 22, 7, -41, 26, -16, 6,
					-- layer=2 filter=43 channel=97
					-24, 5, 29, 19, 12, 28, 39, 9, -7,
					-- layer=2 filter=43 channel=98
					-30, -73, -78, -36, -38, 17, -30, 14, -9,
					-- layer=2 filter=43 channel=99
					29, 7, 29, 2, 15, 0, 3, 22, 32,
					-- layer=2 filter=43 channel=100
					6, 38, 30, 0, -12, -5, -9, -16, -87,
					-- layer=2 filter=43 channel=101
					-16, -18, 12, -35, -19, -15, -40, -12, 35,
					-- layer=2 filter=43 channel=102
					-28, 14, -67, -8, -29, -13, 41, -52, 19,
					-- layer=2 filter=43 channel=103
					6, -8, 19, -24, 4, 15, -9, -57, -19,
					-- layer=2 filter=43 channel=104
					13, 12, 14, -2, 18, -23, -32, -43, 15,
					-- layer=2 filter=43 channel=105
					37, -51, -46, -55, -12, 30, -36, 40, -7,
					-- layer=2 filter=43 channel=106
					-45, -42, -39, -4, -19, -5, 1, -3, 31,
					-- layer=2 filter=43 channel=107
					0, 36, 0, -6, 40, 2, -61, -18, 10,
					-- layer=2 filter=43 channel=108
					-20, 42, 46, -5, -3, 7, 20, -30, 19,
					-- layer=2 filter=43 channel=109
					17, -6, -9, 11, 7, 9, 23, -1, 14,
					-- layer=2 filter=43 channel=110
					-20, -19, -20, 10, 13, -7, 21, 47, 23,
					-- layer=2 filter=43 channel=111
					-11, -8, 5, -9, -6, -4, 1, 0, -1,
					-- layer=2 filter=43 channel=112
					43, 0, -23, 32, 4, 39, 6, 29, 50,
					-- layer=2 filter=43 channel=113
					23, -1, -9, 21, -11, 1, -4, -6, -1,
					-- layer=2 filter=43 channel=114
					-14, 0, -1, -18, -20, -2, -8, 0, 1,
					-- layer=2 filter=43 channel=115
					-2, 5, -5, 9, 2, 8, -6, -4, 4,
					-- layer=2 filter=43 channel=116
					-22, -82, -43, -51, -83, -27, 23, -27, -13,
					-- layer=2 filter=43 channel=117
					-33, -52, -21, -87, -59, -55, 2, -2, 16,
					-- layer=2 filter=43 channel=118
					15, 13, 15, 8, 1, -14, 33, 14, -25,
					-- layer=2 filter=43 channel=119
					12, -5, -23, -13, -24, -18, 47, -41, -25,
					-- layer=2 filter=43 channel=120
					0, 3, -10, -2, 6, 3, 0, -6, -9,
					-- layer=2 filter=43 channel=121
					5, 0, -11, 10, -7, -4, 6, 4, -4,
					-- layer=2 filter=43 channel=122
					0, 10, 6, 8, -10, 14, 8, 10, 4,
					-- layer=2 filter=43 channel=123
					-58, -52, 13, -75, -52, 5, 1, 5, -36,
					-- layer=2 filter=43 channel=124
					-17, -65, -19, -52, 12, 33, 38, 58, -1,
					-- layer=2 filter=43 channel=125
					-7, 6, 7, -10, 2, 0, 0, -7, 8,
					-- layer=2 filter=43 channel=126
					10, 0, 48, 5, 45, -24, 8, 47, 8,
					-- layer=2 filter=43 channel=127
					8, 10, -3, -13, -26, -13, -21, -22, -7,
					-- layer=2 filter=44 channel=0
					7, 6, 10, 29, 17, -7, -9, -9, -11,
					-- layer=2 filter=44 channel=1
					-25, -31, 3, 2, -3, -1, -36, 11, 21,
					-- layer=2 filter=44 channel=2
					-5, 5, 2, 5, -3, 3, 4, -5, -7,
					-- layer=2 filter=44 channel=3
					-8, -23, 19, 5, 6, 25, 4, 8, -27,
					-- layer=2 filter=44 channel=4
					-13, -21, -38, -22, 1, 13, -46, -37, -9,
					-- layer=2 filter=44 channel=5
					13, 26, -8, 6, 9, -9, -6, 6, -2,
					-- layer=2 filter=44 channel=6
					25, -26, -52, -16, -28, -20, -93, -56, -2,
					-- layer=2 filter=44 channel=7
					24, 22, 17, 43, 31, 40, -22, 7, 30,
					-- layer=2 filter=44 channel=8
					-11, 3, -8, 2, -3, -11, -5, 4, 7,
					-- layer=2 filter=44 channel=9
					40, 6, 66, -4, 27, -6, -8, -11, -23,
					-- layer=2 filter=44 channel=10
					6, -5, 40, 11, 0, 15, -4, -10, -19,
					-- layer=2 filter=44 channel=11
					21, 14, 4, 2, 4, -32, -2, -17, -32,
					-- layer=2 filter=44 channel=12
					13, 1, -2, 44, 36, 32, 35, 37, 41,
					-- layer=2 filter=44 channel=13
					0, -3, -6, 1, 8, 10, 0, -3, 1,
					-- layer=2 filter=44 channel=14
					19, 22, 30, 13, 12, 6, 4, 17, 18,
					-- layer=2 filter=44 channel=15
					3, -50, -72, -40, 22, 20, 1, -28, 0,
					-- layer=2 filter=44 channel=16
					-61, -59, -75, -49, -46, -18, -43, -38, -34,
					-- layer=2 filter=44 channel=17
					4, 0, -10, 9, -6, -6, -6, -2, -5,
					-- layer=2 filter=44 channel=18
					-20, 29, -12, -7, 20, 3, 8, 11, -9,
					-- layer=2 filter=44 channel=19
					-42, -33, -7, -39, -46, 18, -45, -30, 33,
					-- layer=2 filter=44 channel=20
					7, 10, -10, 5, 6, 3, 2, -1, 9,
					-- layer=2 filter=44 channel=21
					-6, -13, 2, -10, -9, -4, -4, -8, -7,
					-- layer=2 filter=44 channel=22
					-8, 0, 7, -1, 2, -7, 1, -4, 3,
					-- layer=2 filter=44 channel=23
					18, 12, -39, -14, 3, 23, -8, 24, 20,
					-- layer=2 filter=44 channel=24
					-25, -41, -10, -6, -12, -13, 27, 9, 3,
					-- layer=2 filter=44 channel=25
					-32, -21, -6, -8, -19, -28, 4, 2, -13,
					-- layer=2 filter=44 channel=26
					-12, 1, 4, -10, 5, 5, -1, 3, -3,
					-- layer=2 filter=44 channel=27
					15, -4, -4, 7, 10, -7, 0, 27, -7,
					-- layer=2 filter=44 channel=28
					2, 21, 0, 23, 15, 17, 7, 23, 36,
					-- layer=2 filter=44 channel=29
					-4, 11, 7, 1, 6, -4, -2, 1, -2,
					-- layer=2 filter=44 channel=30
					25, -31, -3, 10, -10, 7, 3, 25, 13,
					-- layer=2 filter=44 channel=31
					-17, -9, 16, -17, -9, 20, -34, -34, 6,
					-- layer=2 filter=44 channel=32
					6, 2, 7, 5, -1, -3, 8, -8, 10,
					-- layer=2 filter=44 channel=33
					12, 15, -2, 4, 28, 0, -21, 2, -30,
					-- layer=2 filter=44 channel=34
					16, 30, -18, -49, -25, 20, -62, -53, -9,
					-- layer=2 filter=44 channel=35
					-23, 13, -1, 5, 23, 27, -18, 18, 21,
					-- layer=2 filter=44 channel=36
					8, 6, 12, 8, 8, 11, 7, -1, 3,
					-- layer=2 filter=44 channel=37
					19, 19, -4, 1, -7, -15, -5, 6, -21,
					-- layer=2 filter=44 channel=38
					10, 6, -10, 12, 10, 13, 8, 4, -7,
					-- layer=2 filter=44 channel=39
					6, -6, -16, 51, 11, 26, 12, 11, 10,
					-- layer=2 filter=44 channel=40
					-22, -11, -37, -61, 14, -53, -44, -101, 24,
					-- layer=2 filter=44 channel=41
					-4, 7, -7, -4, -8, 0, -6, -1, -9,
					-- layer=2 filter=44 channel=42
					-22, -24, -15, 0, 27, 2, 21, 21, 30,
					-- layer=2 filter=44 channel=43
					-20, -9, 4, 2, -24, -41, -21, -31, -77,
					-- layer=2 filter=44 channel=44
					0, -6, -9, -8, 8, 0, 10, -2, -2,
					-- layer=2 filter=44 channel=45
					-71, -52, -44, -22, -23, -4, 0, 32, -20,
					-- layer=2 filter=44 channel=46
					5, 11, 34, 25, 31, -2, -13, -26, -28,
					-- layer=2 filter=44 channel=47
					-44, -24, -15, 15, 16, -16, 10, 10, 10,
					-- layer=2 filter=44 channel=48
					7, 0, 0, 7, -7, -3, -3, 1, -1,
					-- layer=2 filter=44 channel=49
					-39, 8, -32, 1, -23, 22, 34, 53, 34,
					-- layer=2 filter=44 channel=50
					10, 12, 30, 3, 7, 10, 7, -7, 6,
					-- layer=2 filter=44 channel=51
					29, 25, 16, 4, -11, -21, 3, -18, -37,
					-- layer=2 filter=44 channel=52
					16, 43, -5, -32, 4, -53, -14, -34, -6,
					-- layer=2 filter=44 channel=53
					76, 49, 0, -31, -51, -39, 29, -79, -20,
					-- layer=2 filter=44 channel=54
					33, 12, 10, 2, 4, -1, -22, 7, 8,
					-- layer=2 filter=44 channel=55
					8, 12, 10, -5, 3, -2, -4, -3, -3,
					-- layer=2 filter=44 channel=56
					34, 38, -5, 22, -1, -24, 11, -12, -29,
					-- layer=2 filter=44 channel=57
					-6, -2, 0, -11, -4, 2, 3, 2, -9,
					-- layer=2 filter=44 channel=58
					13, 20, 3, 41, 34, 44, 36, 40, 36,
					-- layer=2 filter=44 channel=59
					10, -8, -17, 22, -26, 4, 0, 2, 22,
					-- layer=2 filter=44 channel=60
					17, 8, 24, 0, -11, 47, -31, 1, 41,
					-- layer=2 filter=44 channel=61
					62, -9, -7, 3, -22, 13, -25, -13, -7,
					-- layer=2 filter=44 channel=62
					-20, -7, -16, -43, -38, 9, -60, -44, 2,
					-- layer=2 filter=44 channel=63
					15, 26, -35, 23, -17, 1, -11, 7, -6,
					-- layer=2 filter=44 channel=64
					-11, -33, -19, 18, 12, 18, 13, 40, 48,
					-- layer=2 filter=44 channel=65
					47, 0, -24, 3, -53, -3, -20, -45, -36,
					-- layer=2 filter=44 channel=66
					-30, -4, -33, -9, -11, -5, 29, -32, -27,
					-- layer=2 filter=44 channel=67
					20, -9, 19, -10, -25, -40, -31, -34, -40,
					-- layer=2 filter=44 channel=68
					7, -4, 0, -5, -9, -1, 7, 7, -8,
					-- layer=2 filter=44 channel=69
					-2, -32, -25, 29, 16, 19, -1, 16, 24,
					-- layer=2 filter=44 channel=70
					22, 15, -12, -2, 16, 32, 5, 7, 10,
					-- layer=2 filter=44 channel=71
					31, 17, -25, 9, 11, -3, 22, 29, -8,
					-- layer=2 filter=44 channel=72
					16, 52, 11, 20, 8, -1, -6, -14, 8,
					-- layer=2 filter=44 channel=73
					-6, 48, 82, -23, -93, -33, 43, 43, 13,
					-- layer=2 filter=44 channel=74
					4, -14, 4, 8, -3, -8, 0, -2, 10,
					-- layer=2 filter=44 channel=75
					8, -5, -33, 14, 6, 59, -33, -9, 14,
					-- layer=2 filter=44 channel=76
					51, 2, 32, -55, -40, 70, -16, -87, -28,
					-- layer=2 filter=44 channel=77
					-5, -4, 2, 3, 0, 2, 7, -9, 2,
					-- layer=2 filter=44 channel=78
					6, 17, -22, 4, -19, -32, 27, -18, -35,
					-- layer=2 filter=44 channel=79
					8, 10, -7, 2, -11, 1, 6, 9, 3,
					-- layer=2 filter=44 channel=80
					-3, -12, -3, -6, 9, -2, -48, -17, -39,
					-- layer=2 filter=44 channel=81
					-3, 8, -9, 10, 11, -5, 9, -1, -1,
					-- layer=2 filter=44 channel=82
					-5, 0, -3, -2, -3, -7, 9, -2, -6,
					-- layer=2 filter=44 channel=83
					-10, -13, -52, -30, -21, 15, -39, -8, -5,
					-- layer=2 filter=44 channel=84
					-5, -7, -5, -4, -4, -1, 0, -4, 0,
					-- layer=2 filter=44 channel=85
					8, 8, 10, 4, 13, -5, 10, 0, 0,
					-- layer=2 filter=44 channel=86
					-12, -14, -10, -15, -2, 2, -12, -12, -3,
					-- layer=2 filter=44 channel=87
					4, -6, -7, -34, -4, 38, -57, -39, 26,
					-- layer=2 filter=44 channel=88
					-1, -8, 14, 16, -6, 0, -24, -9, 27,
					-- layer=2 filter=44 channel=89
					-26, -19, -7, 20, -12, -8, -13, 0, 15,
					-- layer=2 filter=44 channel=90
					8, -2, 0, -1, 9, 7, -6, -9, -7,
					-- layer=2 filter=44 channel=91
					10, 16, 8, 25, 14, 19, 21, 10, 28,
					-- layer=2 filter=44 channel=92
					-2, -23, 6, 31, 8, -1, 18, 17, 33,
					-- layer=2 filter=44 channel=93
					-4, -40, -2, -9, -28, 9, -58, -35, -13,
					-- layer=2 filter=44 channel=94
					47, -4, 14, -21, -26, -79, -87, -59, -35,
					-- layer=2 filter=44 channel=95
					11, 4, -1, -1, 6, 7, 0, -4, 0,
					-- layer=2 filter=44 channel=96
					-18, 109, -4, -14, -21, -25, -59, -60, 0,
					-- layer=2 filter=44 channel=97
					0, -29, -19, 15, 22, 0, 48, 31, 7,
					-- layer=2 filter=44 channel=98
					1, 5, 3, -15, 12, 34, -12, 25, 9,
					-- layer=2 filter=44 channel=99
					71, 36, 4, -43, -46, 13, -10, -58, 7,
					-- layer=2 filter=44 channel=100
					-8, 2, -12, 15, 18, 1, -31, 5, -1,
					-- layer=2 filter=44 channel=101
					33, 19, -8, 6, -21, -9, -5, 8, -10,
					-- layer=2 filter=44 channel=102
					19, 29, -10, 4, -20, 0, -24, -2, 13,
					-- layer=2 filter=44 channel=103
					-11, 4, 7, -22, -34, -23, -34, -30, -35,
					-- layer=2 filter=44 channel=104
					32, 41, -47, 1, 0, -17, 66, -54, -17,
					-- layer=2 filter=44 channel=105
					-9, 20, 37, -41, -27, 82, -47, 8, 0,
					-- layer=2 filter=44 channel=106
					-11, 3, 22, 19, 2, -10, 6, -7, 9,
					-- layer=2 filter=44 channel=107
					-23, -50, 42, 21, 12, -34, 0, -19, 16,
					-- layer=2 filter=44 channel=108
					-11, 14, -33, -38, 7, -10, -25, 21, -34,
					-- layer=2 filter=44 channel=109
					3, 6, -10, -3, -4, -5, 6, 0, 4,
					-- layer=2 filter=44 channel=110
					4, 14, -20, 6, -10, 1, -21, -3, 14,
					-- layer=2 filter=44 channel=111
					-13, -8, -6, -3, 1, -8, -4, 1, -7,
					-- layer=2 filter=44 channel=112
					8, -11, 0, 1, 3, 32, -1, -13, -15,
					-- layer=2 filter=44 channel=113
					24, 9, -14, 0, -36, 14, 33, 10, 13,
					-- layer=2 filter=44 channel=114
					17, 11, 12, 3, 0, 0, -8, -13, 8,
					-- layer=2 filter=44 channel=115
					9, 1, 8, -5, 0, 8, -4, -4, 7,
					-- layer=2 filter=44 channel=116
					-14, 3, -40, -33, 11, 32, -46, -47, 38,
					-- layer=2 filter=44 channel=117
					-6, -14, 6, 24, -2, -8, -8, -25, 3,
					-- layer=2 filter=44 channel=118
					7, 28, -14, -10, -2, -3, -15, -9, -40,
					-- layer=2 filter=44 channel=119
					-25, 0, -24, -25, -20, 13, -43, -27, 8,
					-- layer=2 filter=44 channel=120
					-10, -7, -2, 6, 5, 3, 4, -8, 8,
					-- layer=2 filter=44 channel=121
					-3, 0, -7, 0, 0, -4, 0, 10, -1,
					-- layer=2 filter=44 channel=122
					-13, -4, 5, -4, -2, -8, 0, -2, -4,
					-- layer=2 filter=44 channel=123
					3, 26, -33, 6, 14, 6, -10, 12, -7,
					-- layer=2 filter=44 channel=124
					-3, -92, -115, -49, 0, 0, -8, -18, 51,
					-- layer=2 filter=44 channel=125
					6, 0, -4, 3, -7, 4, -6, 10, 7,
					-- layer=2 filter=44 channel=126
					1, 102, -13, 25, -30, -52, -69, -22, 82,
					-- layer=2 filter=44 channel=127
					-20, 22, -34, -10, -22, -2, -12, 1, -7,
					-- layer=2 filter=45 channel=0
					5, 3, 11, -8, -5, -10, 2, -12, -4,
					-- layer=2 filter=45 channel=1
					-29, 32, 41, 13, -6, -13, -14, -26, -14,
					-- layer=2 filter=45 channel=2
					5, -4, -1, 9, -3, 6, 11, -3, 8,
					-- layer=2 filter=45 channel=3
					37, 3, -43, 9, 30, -25, 31, 28, 23,
					-- layer=2 filter=45 channel=4
					48, 13, 12, -24, 10, -45, -14, -10, -23,
					-- layer=2 filter=45 channel=5
					-4, 3, -2, -31, -13, 9, -21, 19, 8,
					-- layer=2 filter=45 channel=6
					15, 15, 15, 12, 25, 5, -19, 21, 41,
					-- layer=2 filter=45 channel=7
					20, 1, -43, -42, -14, 19, -8, -44, -14,
					-- layer=2 filter=45 channel=8
					-10, 5, 6, -10, 6, 1, 4, 1, 4,
					-- layer=2 filter=45 channel=9
					27, 13, 28, -16, -35, -23, -25, -13, -25,
					-- layer=2 filter=45 channel=10
					7, -8, -24, -7, -1, -7, 17, 2, 5,
					-- layer=2 filter=45 channel=11
					-37, 4, -5, -37, 5, 16, -24, -44, -2,
					-- layer=2 filter=45 channel=12
					-7, 6, 43, 25, -11, -7, -2, 38, 18,
					-- layer=2 filter=45 channel=13
					-7, 1, 3, -8, 5, 0, 0, -6, -9,
					-- layer=2 filter=45 channel=14
					3, 51, 71, 0, -11, -2, -25, 5, -8,
					-- layer=2 filter=45 channel=15
					18, -26, -31, -30, 1, -37, -58, -12, -52,
					-- layer=2 filter=45 channel=16
					42, 18, -50, -23, -48, -49, 19, -13, -12,
					-- layer=2 filter=45 channel=17
					-5, 3, 5, -9, 4, 6, -3, 1, 3,
					-- layer=2 filter=45 channel=18
					-5, 12, 39, 4, 6, 2, 14, -13, 14,
					-- layer=2 filter=45 channel=19
					-45, -52, -11, 21, 5, -4, -79, -43, -42,
					-- layer=2 filter=45 channel=20
					-2, 7, 5, 4, 0, 0, 1, -9, -2,
					-- layer=2 filter=45 channel=21
					15, 0, 18, -3, 11, 13, 2, 15, 10,
					-- layer=2 filter=45 channel=22
					1, 5, 3, -5, 3, -6, 5, 2, -6,
					-- layer=2 filter=45 channel=23
					14, -1, -12, -20, -16, -28, 2, 15, 15,
					-- layer=2 filter=45 channel=24
					31, -24, -1, 19, 5, -30, 28, 31, -2,
					-- layer=2 filter=45 channel=25
					14, -40, -11, 18, 9, 2, 10, 26, -7,
					-- layer=2 filter=45 channel=26
					1, 9, 12, -9, -4, 6, -9, -2, -3,
					-- layer=2 filter=45 channel=27
					-15, -9, -9, -32, 18, 3, -28, -59, -22,
					-- layer=2 filter=45 channel=28
					2, 0, -47, 5, -18, -20, 41, -15, -37,
					-- layer=2 filter=45 channel=29
					2, 1, 10, 4, 2, 7, 9, -7, 2,
					-- layer=2 filter=45 channel=30
					6, 7, 19, -1, 13, 0, -20, 21, -25,
					-- layer=2 filter=45 channel=31
					10, -38, 23, 73, -18, -22, -58, 36, -19,
					-- layer=2 filter=45 channel=32
					2, -4, 11, -5, 1, 4, -3, 4, -5,
					-- layer=2 filter=45 channel=33
					52, 72, 59, -26, 35, 26, 20, -36, -17,
					-- layer=2 filter=45 channel=34
					-33, 34, 12, -1, 5, 19, 0, -63, 23,
					-- layer=2 filter=45 channel=35
					-38, -14, -68, 0, 26, -21, 6, -15, 15,
					-- layer=2 filter=45 channel=36
					-11, -8, 5, 2, 0, -3, -1, -1, -4,
					-- layer=2 filter=45 channel=37
					-45, -2, 4, -50, -17, -2, -18, -23, -2,
					-- layer=2 filter=45 channel=38
					-4, 36, 29, 5, 1, -26, -17, -18, -24,
					-- layer=2 filter=45 channel=39
					57, 16, -16, -5, -54, -2, 25, 7, 8,
					-- layer=2 filter=45 channel=40
					14, 11, 8, -7, -32, 27, 2, 49, 9,
					-- layer=2 filter=45 channel=41
					2, 1, 4, -1, -1, 1, -6, -8, -7,
					-- layer=2 filter=45 channel=42
					0, -39, 19, -6, -14, -44, 17, 22, 9,
					-- layer=2 filter=45 channel=43
					-29, 6, -29, -37, 13, -45, 21, -20, -13,
					-- layer=2 filter=45 channel=44
					0, 2, -1, 7, -2, -3, 8, -6, 1,
					-- layer=2 filter=45 channel=45
					39, 49, -36, 9, -14, -11, -7, -15, 5,
					-- layer=2 filter=45 channel=46
					10, 17, 5, -12, -28, -30, -6, -11, -29,
					-- layer=2 filter=45 channel=47
					19, -24, -4, -23, -22, 15, 4, -68, -25,
					-- layer=2 filter=45 channel=48
					-10, -5, 2, -8, -5, -10, 6, -3, -4,
					-- layer=2 filter=45 channel=49
					-2, 12, 36, 0, 9, -6, -12, 18, -20,
					-- layer=2 filter=45 channel=50
					25, 11, 13, 0, 4, -16, -11, 0, -12,
					-- layer=2 filter=45 channel=51
					-4, 14, 27, -22, 17, 8, -16, -19, -2,
					-- layer=2 filter=45 channel=52
					-6, 13, 26, -46, 51, -14, -32, -41, -1,
					-- layer=2 filter=45 channel=53
					12, -52, 29, 11, -37, -23, -44, 31, -12,
					-- layer=2 filter=45 channel=54
					-23, -30, -14, -38, 17, -35, -35, -7, -9,
					-- layer=2 filter=45 channel=55
					-6, -5, 10, -10, 6, 4, -5, 1, 0,
					-- layer=2 filter=45 channel=56
					-19, 19, 7, -35, -20, 14, -23, -36, 8,
					-- layer=2 filter=45 channel=57
					-1, -8, -12, -6, -5, 10, 6, 13, -8,
					-- layer=2 filter=45 channel=58
					-33, 0, 16, 22, 11, 6, -29, 11, 46,
					-- layer=2 filter=45 channel=59
					-38, 45, -8, 15, 16, 13, 0, -41, 44,
					-- layer=2 filter=45 channel=60
					-26, -9, 35, 37, 4, 48, -28, -7, 17,
					-- layer=2 filter=45 channel=61
					-60, -20, 1, -11, -32, 21, -41, -64, 0,
					-- layer=2 filter=45 channel=62
					-11, 2, 11, -7, -2, -6, -44, -27, 10,
					-- layer=2 filter=45 channel=63
					19, 11, -5, 7, -10, 17, -5, -14, -3,
					-- layer=2 filter=45 channel=64
					16, -3, 5, -22, -4, -13, -4, 29, 21,
					-- layer=2 filter=45 channel=65
					-30, 0, 18, -7, 16, 15, -56, -34, -12,
					-- layer=2 filter=45 channel=66
					37, 19, 38, 47, -9, 13, -20, -1, 10,
					-- layer=2 filter=45 channel=67
					22, 5, 3, -10, -18, -39, -2, -26, -42,
					-- layer=2 filter=45 channel=68
					-6, 0, -4, -4, -3, 10, -9, 7, 2,
					-- layer=2 filter=45 channel=69
					18, 6, 12, -30, 5, -18, 11, 34, 22,
					-- layer=2 filter=45 channel=70
					-15, -8, -17, 5, 3, 9, -4, -2, 5,
					-- layer=2 filter=45 channel=71
					-5, 10, 30, 5, 51, 32, -16, -17, -25,
					-- layer=2 filter=45 channel=72
					1, 51, 28, -26, 4, 37, 5, -17, 9,
					-- layer=2 filter=45 channel=73
					7, -5, -59, 10, -64, 0, -28, -40, -91,
					-- layer=2 filter=45 channel=74
					8, 6, -5, -14, 6, -34, 18, -9, -1,
					-- layer=2 filter=45 channel=75
					-24, -18, -10, -34, -41, 3, 4, 81, -15,
					-- layer=2 filter=45 channel=76
					-2, -21, 8, 9, -5, -18, -33, -32, -52,
					-- layer=2 filter=45 channel=77
					-10, -9, 4, 7, -9, -1, 0, 6, 1,
					-- layer=2 filter=45 channel=78
					-8, 23, -25, -15, 11, 17, -8, -26, 33,
					-- layer=2 filter=45 channel=79
					-8, 1, -9, 5, 5, -4, -6, 5, 8,
					-- layer=2 filter=45 channel=80
					43, -2, -2, 23, -22, -41, -11, 3, -1,
					-- layer=2 filter=45 channel=81
					4, -11, -9, 6, -5, -10, -3, -6, -1,
					-- layer=2 filter=45 channel=82
					-4, -9, -7, -3, -6, -9, -4, 1, -4,
					-- layer=2 filter=45 channel=83
					39, -16, -2, -7, -16, -25, -8, 26, -18,
					-- layer=2 filter=45 channel=84
					-2, -2, 2, -5, 6, -7, 0, 5, 0,
					-- layer=2 filter=45 channel=85
					-15, 10, -9, 2, -7, -6, 0, 12, -7,
					-- layer=2 filter=45 channel=86
					-3, -8, 5, -18, 5, 7, -1, -9, -5,
					-- layer=2 filter=45 channel=87
					44, 20, 13, 26, 33, 37, 19, 29, 29,
					-- layer=2 filter=45 channel=88
					35, 26, 22, 8, 23, -32, -14, 0, -20,
					-- layer=2 filter=45 channel=89
					-36, 35, 38, 31, 7, 13, -8, 6, 20,
					-- layer=2 filter=45 channel=90
					0, 6, -6, 8, 3, 0, 0, 5, 1,
					-- layer=2 filter=45 channel=91
					6, -9, 10, 26, -18, -18, 15, 34, 32,
					-- layer=2 filter=45 channel=92
					0, 24, 31, 12, -4, -23, 11, 0, 27,
					-- layer=2 filter=45 channel=93
					-4, -36, -1, 42, 42, 19, -53, 1, 5,
					-- layer=2 filter=45 channel=94
					-53, -54, 15, -30, 11, 16, -71, -25, -30,
					-- layer=2 filter=45 channel=95
					3, 3, 3, 14, 10, 13, 5, 13, 3,
					-- layer=2 filter=45 channel=96
					-42, 58, 34, 22, 64, 44, -8, 33, 26,
					-- layer=2 filter=45 channel=97
					17, 2, -10, -5, 8, -40, -3, 29, 6,
					-- layer=2 filter=45 channel=98
					-9, -22, -14, -2, -19, -3, -6, -71, -15,
					-- layer=2 filter=45 channel=99
					-61, -33, -17, -19, 23, -28, -87, -57, -41,
					-- layer=2 filter=45 channel=100
					15, 4, 4, -9, 1, 7, -36, 28, 14,
					-- layer=2 filter=45 channel=101
					-13, -25, -7, 8, 17, 37, -17, -15, -7,
					-- layer=2 filter=45 channel=102
					-47, 41, 47, -20, 68, 32, -20, -12, 17,
					-- layer=2 filter=45 channel=103
					27, -22, 43, 45, 12, 3, 43, -5, 5,
					-- layer=2 filter=45 channel=104
					3, 4, 11, 2, 8, -18, -50, -4, 4,
					-- layer=2 filter=45 channel=105
					-29, -17, -49, -25, -14, -3, 39, -38, 43,
					-- layer=2 filter=45 channel=106
					27, -4, 29, 20, -7, 12, -11, 2, -19,
					-- layer=2 filter=45 channel=107
					-30, 2, 32, 30, 38, -17, 16, -23, 25,
					-- layer=2 filter=45 channel=108
					-23, 24, 24, -7, 15, 5, -53, -59, -32,
					-- layer=2 filter=45 channel=109
					-1, 1, -6, 6, 1, -9, 14, 0, -4,
					-- layer=2 filter=45 channel=110
					-25, -32, -32, -44, -33, -13, 0, 39, 51,
					-- layer=2 filter=45 channel=111
					-11, 5, -12, -12, 3, 3, 8, 1, 5,
					-- layer=2 filter=45 channel=112
					-14, -14, 11, 11, -4, 12, -32, -19, -38,
					-- layer=2 filter=45 channel=113
					-2, -3, 4, -5, -10, 15, -20, -5, -17,
					-- layer=2 filter=45 channel=114
					4, -12, 6, 7, 2, 2, 6, 0, -1,
					-- layer=2 filter=45 channel=115
					7, -1, -1, -2, -5, 5, -5, 6, 8,
					-- layer=2 filter=45 channel=116
					31, 20, 11, 9, 51, 25, 13, 16, 15,
					-- layer=2 filter=45 channel=117
					-3, 42, 0, -16, 26, 41, -34, -39, -82,
					-- layer=2 filter=45 channel=118
					7, 11, -43, -12, -41, -56, 20, -16, 25,
					-- layer=2 filter=45 channel=119
					-10, 4, 2, -3, -34, -41, 73, -6, -25,
					-- layer=2 filter=45 channel=120
					5, 9, -4, -9, -6, -9, 5, 3, 2,
					-- layer=2 filter=45 channel=121
					2, -5, -1, -1, -11, -1, -3, -6, 0,
					-- layer=2 filter=45 channel=122
					5, 6, -8, 4, -5, -5, 1, -5, -14,
					-- layer=2 filter=45 channel=123
					41, 30, 5, -14, -36, 38, -24, -40, -8,
					-- layer=2 filter=45 channel=124
					45, 26, -6, 11, 4, -42, -12, 37, 6,
					-- layer=2 filter=45 channel=125
					-4, 5, -8, 0, -4, 9, -4, 10, 3,
					-- layer=2 filter=45 channel=126
					-52, 57, 18, -44, 35, 12, 31, -10, 14,
					-- layer=2 filter=45 channel=127
					31, 30, 36, 19, -3, -23, -6, 13, 18,
					-- layer=2 filter=46 channel=0
					-11, -11, -9, -2, -10, -2, 5, 8, -13,
					-- layer=2 filter=46 channel=1
					-4, -20, -5, -8, -5, -5, -16, -22, -15,
					-- layer=2 filter=46 channel=2
					-1, -5, 8, -8, 0, -1, 10, -4, -3,
					-- layer=2 filter=46 channel=3
					12, 4, -5, -11, 0, -1, -10, -9, -3,
					-- layer=2 filter=46 channel=4
					5, 8, 2, -11, -12, 2, -6, -9, -13,
					-- layer=2 filter=46 channel=5
					-6, -7, -4, -2, -10, -15, -8, -5, -9,
					-- layer=2 filter=46 channel=6
					-5, -1, -5, -3, 11, -9, -2, 2, 8,
					-- layer=2 filter=46 channel=7
					3, 2, -2, -10, 1, -15, -12, -26, 0,
					-- layer=2 filter=46 channel=8
					-1, 4, -9, 2, 7, 6, -7, 4, -5,
					-- layer=2 filter=46 channel=9
					3, -13, -14, 10, -7, 5, -4, -10, -13,
					-- layer=2 filter=46 channel=10
					-7, -13, -14, -10, 7, -10, -6, -2, -11,
					-- layer=2 filter=46 channel=11
					-11, -13, -1, -11, -15, -2, -3, -7, -13,
					-- layer=2 filter=46 channel=12
					-4, -21, -3, -18, -8, 5, -5, -17, -7,
					-- layer=2 filter=46 channel=13
					3, 6, 3, -1, 0, 10, -1, 2, -1,
					-- layer=2 filter=46 channel=14
					-11, -4, -16, -12, -18, 1, 0, -10, -6,
					-- layer=2 filter=46 channel=15
					-8, 0, 9, -10, -24, -9, 0, -2, -8,
					-- layer=2 filter=46 channel=16
					18, -5, -5, 5, -12, -9, 9, -11, 0,
					-- layer=2 filter=46 channel=17
					-3, 0, -6, 11, 9, 2, 9, -6, 0,
					-- layer=2 filter=46 channel=18
					-21, -1, 8, -1, -1, 6, -25, 1, 9,
					-- layer=2 filter=46 channel=19
					-3, 4, -10, -13, -14, -7, -6, -11, -14,
					-- layer=2 filter=46 channel=20
					3, -6, 0, -3, 8, -2, 7, 5, 5,
					-- layer=2 filter=46 channel=21
					-11, -8, -6, -2, 0, -7, -1, -8, 7,
					-- layer=2 filter=46 channel=22
					8, -5, 10, -5, 6, 5, -1, 3, -4,
					-- layer=2 filter=46 channel=23
					-10, 0, -11, -3, 0, -10, -6, -12, -18,
					-- layer=2 filter=46 channel=24
					0, 0, -10, 0, -17, -18, 0, -12, -5,
					-- layer=2 filter=46 channel=25
					5, 5, 7, -23, -15, -12, -6, -18, -5,
					-- layer=2 filter=46 channel=26
					-10, -9, -5, 5, 0, -3, 1, -3, 9,
					-- layer=2 filter=46 channel=27
					-15, -11, -9, 1, -5, 2, -4, -5, 1,
					-- layer=2 filter=46 channel=28
					-9, 2, 1, -3, -11, -8, -4, -15, -7,
					-- layer=2 filter=46 channel=29
					2, 9, -3, 4, -9, 2, -1, 0, 9,
					-- layer=2 filter=46 channel=30
					7, -2, -2, 0, -17, -5, 8, -14, -6,
					-- layer=2 filter=46 channel=31
					8, 8, 16, -1, 1, 6, 2, 8, -1,
					-- layer=2 filter=46 channel=32
					4, -2, 5, -3, -4, -5, -6, 8, -1,
					-- layer=2 filter=46 channel=33
					-6, -4, -2, 12, 6, 3, -2, 3, 0,
					-- layer=2 filter=46 channel=34
					-24, -13, 3, 11, -29, -5, -13, -6, -2,
					-- layer=2 filter=46 channel=35
					-26, -22, -2, 7, -11, 1, -23, 0, 2,
					-- layer=2 filter=46 channel=36
					7, 1, -9, 1, 6, 10, -3, 0, 5,
					-- layer=2 filter=46 channel=37
					-4, -2, -11, -10, -1, -3, -11, 0, -12,
					-- layer=2 filter=46 channel=38
					-22, -19, -19, -5, -3, -5, 6, -4, -4,
					-- layer=2 filter=46 channel=39
					13, -5, 3, -10, -9, -18, 3, 2, -7,
					-- layer=2 filter=46 channel=40
					-11, -9, -5, 4, -16, 17, -1, 13, -4,
					-- layer=2 filter=46 channel=41
					-9, 8, 1, -2, 5, -2, 4, -3, -3,
					-- layer=2 filter=46 channel=42
					-7, -7, -4, 2, 0, -8, -4, -9, -16,
					-- layer=2 filter=46 channel=43
					-10, 5, 8, -13, -3, 7, -3, 4, 10,
					-- layer=2 filter=46 channel=44
					-7, -9, -4, 2, -1, -4, -7, -8, -7,
					-- layer=2 filter=46 channel=45
					5, -9, 2, -1, 2, -10, 3, 4, 18,
					-- layer=2 filter=46 channel=46
					-3, 4, 4, -10, -16, 6, -17, -3, -7,
					-- layer=2 filter=46 channel=47
					16, 2, 14, -9, -11, -2, 0, 3, 11,
					-- layer=2 filter=46 channel=48
					-7, -1, 4, -6, -3, 10, 10, 5, -9,
					-- layer=2 filter=46 channel=49
					-15, -2, 2, -21, -6, -5, -15, -8, 3,
					-- layer=2 filter=46 channel=50
					-1, 2, 0, -8, -1, -8, 7, -5, -5,
					-- layer=2 filter=46 channel=51
					-15, -11, -4, 2, -1, -5, -10, 6, -8,
					-- layer=2 filter=46 channel=52
					-9, 1, -15, 8, 3, 3, -25, 4, -16,
					-- layer=2 filter=46 channel=53
					7, 4, 14, 0, 0, -19, 4, -9, -19,
					-- layer=2 filter=46 channel=54
					0, -2, -3, 5, -11, -7, -14, -16, -13,
					-- layer=2 filter=46 channel=55
					1, -5, 2, 0, 3, -1, -5, 8, -2,
					-- layer=2 filter=46 channel=56
					-11, -13, -15, -11, -12, -18, 1, -9, -5,
					-- layer=2 filter=46 channel=57
					-5, -5, 9, -2, 10, 7, 10, 5, -10,
					-- layer=2 filter=46 channel=58
					-9, -15, 0, 1, 7, 0, -3, 0, -5,
					-- layer=2 filter=46 channel=59
					0, 2, -8, -2, -7, -6, 0, 1, -2,
					-- layer=2 filter=46 channel=60
					0, 2, -2, 0, -13, -12, 9, -19, 1,
					-- layer=2 filter=46 channel=61
					-8, 0, -4, 3, -6, -4, 4, -4, -14,
					-- layer=2 filter=46 channel=62
					-18, 1, -16, -22, -10, 3, -23, 5, 0,
					-- layer=2 filter=46 channel=63
					7, -9, -8, -11, -13, -18, -5, -7, -8,
					-- layer=2 filter=46 channel=64
					5, -9, -8, -1, 3, -11, -4, -6, -2,
					-- layer=2 filter=46 channel=65
					-7, 4, -1, -13, 8, -12, 0, 1, -9,
					-- layer=2 filter=46 channel=66
					9, -7, 3, -3, -1, 7, 3, -5, 0,
					-- layer=2 filter=46 channel=67
					12, 0, 3, 9, 1, -6, -8, -2, -7,
					-- layer=2 filter=46 channel=68
					4, 10, 0, 4, 7, 2, 6, 3, -3,
					-- layer=2 filter=46 channel=69
					6, 4, -4, -10, -8, -10, -11, -4, 3,
					-- layer=2 filter=46 channel=70
					-19, -23, -15, 6, -14, -6, -15, -18, -5,
					-- layer=2 filter=46 channel=71
					-13, -15, -14, -4, -2, -4, 1, -5, -1,
					-- layer=2 filter=46 channel=72
					-7, 4, -15, -1, -11, -4, -15, -24, -15,
					-- layer=2 filter=46 channel=73
					2, 2, 8, 10, -3, 5, -17, 1, 3,
					-- layer=2 filter=46 channel=74
					3, 11, 6, 6, -8, -10, -10, -11, -10,
					-- layer=2 filter=46 channel=75
					-13, -1, -13, -31, -22, -14, 0, -5, 5,
					-- layer=2 filter=46 channel=76
					23, 0, 16, -10, -14, 0, -19, -9, 0,
					-- layer=2 filter=46 channel=77
					10, 10, 5, -4, -7, -11, -1, -1, -10,
					-- layer=2 filter=46 channel=78
					5, -1, -7, -1, -14, -15, -4, -9, -13,
					-- layer=2 filter=46 channel=79
					-1, 12, -6, 0, 9, -5, -7, -4, 5,
					-- layer=2 filter=46 channel=80
					5, -3, -6, -11, 3, -15, -4, 7, -14,
					-- layer=2 filter=46 channel=81
					3, 2, 5, -7, 1, -8, -2, -9, -5,
					-- layer=2 filter=46 channel=82
					4, 4, -5, 2, -1, -1, -8, -5, 8,
					-- layer=2 filter=46 channel=83
					-8, -8, -10, -8, -12, 7, 11, -9, -2,
					-- layer=2 filter=46 channel=84
					0, 3, 3, -6, 2, -7, -10, 6, 9,
					-- layer=2 filter=46 channel=85
					11, -9, 4, -3, -1, 1, -7, 1, 9,
					-- layer=2 filter=46 channel=86
					-1, 1, 1, -5, 6, 6, 6, -6, 7,
					-- layer=2 filter=46 channel=87
					0, 7, 9, -12, -7, 16, -16, 5, -21,
					-- layer=2 filter=46 channel=88
					-7, 7, -6, -1, 5, -13, 7, -7, -12,
					-- layer=2 filter=46 channel=89
					-8, -17, -5, -10, -24, -6, -4, -14, -6,
					-- layer=2 filter=46 channel=90
					3, 1, 6, -3, 0, -4, 5, -4, -9,
					-- layer=2 filter=46 channel=91
					-1, -17, -10, -4, -19, 4, 0, -18, -13,
					-- layer=2 filter=46 channel=92
					-16, -17, -8, -12, -16, -11, -11, -14, -3,
					-- layer=2 filter=46 channel=93
					-11, 3, 5, 3, 3, 1, -14, -5, 0,
					-- layer=2 filter=46 channel=94
					-5, -10, -13, -18, 7, -10, -18, -6, -17,
					-- layer=2 filter=46 channel=95
					8, 6, 6, -3, 4, 3, 11, -6, 1,
					-- layer=2 filter=46 channel=96
					-3, 4, 5, -2, 3, -11, -8, 6, -18,
					-- layer=2 filter=46 channel=97
					0, -10, 5, -11, -12, -16, 4, -2, -9,
					-- layer=2 filter=46 channel=98
					3, -13, 6, -4, -21, 8, -17, 4, -11,
					-- layer=2 filter=46 channel=99
					4, -7, 2, 0, 0, 4, -3, -15, -8,
					-- layer=2 filter=46 channel=100
					-11, -10, -10, -10, -16, -12, 4, 0, 2,
					-- layer=2 filter=46 channel=101
					4, 0, -8, -4, -11, -11, -11, -16, -24,
					-- layer=2 filter=46 channel=102
					7, 0, -12, -8, -9, 5, -12, 10, 5,
					-- layer=2 filter=46 channel=103
					-4, 9, 11, 1, -6, 2, -6, 8, 0,
					-- layer=2 filter=46 channel=104
					-5, -1, -12, -11, 7, -18, -24, 15, -10,
					-- layer=2 filter=46 channel=105
					7, 0, 0, -10, -31, 8, -15, -7, -18,
					-- layer=2 filter=46 channel=106
					-4, 0, -14, -4, -8, -20, -12, -2, -10,
					-- layer=2 filter=46 channel=107
					-1, 8, -10, 6, -9, -3, -6, 2, 0,
					-- layer=2 filter=46 channel=108
					-11, -7, -23, 0, -10, 10, 14, -1, -1,
					-- layer=2 filter=46 channel=109
					5, -9, -10, 9, 9, -2, 3, 1, -3,
					-- layer=2 filter=46 channel=110
					-9, 2, -3, -15, -9, -11, -9, -10, 0,
					-- layer=2 filter=46 channel=111
					5, 1, -6, -7, 6, 5, -10, 0, -5,
					-- layer=2 filter=46 channel=112
					3, 6, -9, -7, -2, -10, 7, -10, -1,
					-- layer=2 filter=46 channel=113
					-9, -11, -19, 5, -11, -15, -4, -23, -10,
					-- layer=2 filter=46 channel=114
					6, 3, -6, 8, 0, -7, 1, 9, 0,
					-- layer=2 filter=46 channel=115
					-6, 2, -5, 3, 1, -7, -5, 10, 6,
					-- layer=2 filter=46 channel=116
					-10, -3, 0, 9, 0, 14, -21, 6, -7,
					-- layer=2 filter=46 channel=117
					7, 12, 3, -14, 0, -16, -4, -23, 4,
					-- layer=2 filter=46 channel=118
					5, 6, 6, -1, -1, 8, -5, 5, 12,
					-- layer=2 filter=46 channel=119
					-5, 2, -6, 2, -19, -5, -3, -4, -1,
					-- layer=2 filter=46 channel=120
					-8, 10, 6, 2, 1, 3, 0, -5, 6,
					-- layer=2 filter=46 channel=121
					-6, 0, 6, -7, 6, -4, -1, 1, -3,
					-- layer=2 filter=46 channel=122
					8, 2, 1, -7, 9, 0, -9, 8, -8,
					-- layer=2 filter=46 channel=123
					-4, 6, -3, -17, -18, 7, -25, -2, -8,
					-- layer=2 filter=46 channel=124
					-1, 1, 9, -19, -17, -4, -10, -10, -21,
					-- layer=2 filter=46 channel=125
					8, 7, 0, 3, 6, 3, 2, 3, -3,
					-- layer=2 filter=46 channel=126
					-8, 0, 8, -14, 5, -13, -12, 6, -6,
					-- layer=2 filter=46 channel=127
					-17, -4, -19, 3, -8, -11, 4, -20, -18,
					-- layer=2 filter=47 channel=0
					3, -4, 6, -10, 0, -2, -7, 0, -4,
					-- layer=2 filter=47 channel=1
					-12, -9, -1, 0, -13, -15, -3, -9, -11,
					-- layer=2 filter=47 channel=2
					7, -8, -11, 3, -8, -10, 4, 2, 7,
					-- layer=2 filter=47 channel=3
					-2, 9, -11, -7, -6, -14, -11, -9, 5,
					-- layer=2 filter=47 channel=4
					3, 1, -10, -11, -1, -8, -4, -4, 1,
					-- layer=2 filter=47 channel=5
					-18, 1, -14, -6, -12, -7, 2, -4, 0,
					-- layer=2 filter=47 channel=6
					5, -11, -9, -9, 0, 0, -10, -6, 4,
					-- layer=2 filter=47 channel=7
					2, -16, -5, -8, -6, -1, -10, -1, 12,
					-- layer=2 filter=47 channel=8
					-9, 1, -2, -8, 1, 0, 9, 4, -7,
					-- layer=2 filter=47 channel=9
					-4, 2, -6, -1, -9, -4, -11, 3, -7,
					-- layer=2 filter=47 channel=10
					2, -1, -14, -5, 3, -7, -2, 2, -4,
					-- layer=2 filter=47 channel=11
					0, -4, 1, -15, -4, -2, 3, 0, -4,
					-- layer=2 filter=47 channel=12
					-23, -10, -7, -1, 0, 7, 3, -4, -12,
					-- layer=2 filter=47 channel=13
					8, -1, -3, 0, -5, 2, -4, 1, -7,
					-- layer=2 filter=47 channel=14
					6, 5, -2, -12, -5, -3, -2, 2, -3,
					-- layer=2 filter=47 channel=15
					-5, 7, -10, -1, -10, -8, 6, 0, 8,
					-- layer=2 filter=47 channel=16
					0, 4, -11, -2, -9, 4, 6, -11, 0,
					-- layer=2 filter=47 channel=17
					-11, 5, -9, -4, 5, 5, -9, -4, 4,
					-- layer=2 filter=47 channel=18
					1, -18, -8, -6, -7, 0, 10, -8, 4,
					-- layer=2 filter=47 channel=19
					-4, -3, -10, -8, -16, -3, 1, -11, -15,
					-- layer=2 filter=47 channel=20
					7, 10, 5, 6, 5, 0, -6, 8, 8,
					-- layer=2 filter=47 channel=21
					7, -5, 9, 7, 7, -5, 8, -8, -10,
					-- layer=2 filter=47 channel=22
					0, -9, 8, 0, 2, 7, -3, -1, 3,
					-- layer=2 filter=47 channel=23
					8, 0, -2, 1, 8, -3, 3, 0, 0,
					-- layer=2 filter=47 channel=24
					3, -2, -12, -4, 0, -7, -3, -1, -9,
					-- layer=2 filter=47 channel=25
					-18, -3, -14, 2, 5, 8, -13, -12, 3,
					-- layer=2 filter=47 channel=26
					-9, 3, -4, 0, 9, 1, -2, -1, 0,
					-- layer=2 filter=47 channel=27
					0, -11, 0, -11, -8, 4, 2, -16, -10,
					-- layer=2 filter=47 channel=28
					0, -9, 3, -10, -12, 0, 0, -5, -6,
					-- layer=2 filter=47 channel=29
					-8, -9, 3, 3, -6, -2, -7, 3, -2,
					-- layer=2 filter=47 channel=30
					-12, -1, -10, 1, -4, 3, -5, 0, -4,
					-- layer=2 filter=47 channel=31
					-4, 5, 4, 7, -3, 3, 1, -2, 5,
					-- layer=2 filter=47 channel=32
					-9, -8, -4, -6, 7, -8, -7, 6, -10,
					-- layer=2 filter=47 channel=33
					-14, 3, 0, 0, -10, -9, -17, 0, -2,
					-- layer=2 filter=47 channel=34
					-10, -12, 0, -4, 3, -8, -7, 4, -7,
					-- layer=2 filter=47 channel=35
					2, -11, -10, -9, -4, 3, -4, -5, 0,
					-- layer=2 filter=47 channel=36
					9, 2, -8, -3, 0, 5, -6, -4, -2,
					-- layer=2 filter=47 channel=37
					-6, -1, -13, -2, -6, -12, -4, 5, 0,
					-- layer=2 filter=47 channel=38
					-16, -10, 0, 2, -1, 1, 3, 7, -2,
					-- layer=2 filter=47 channel=39
					-4, -3, -11, 3, -8, -1, -10, -11, -2,
					-- layer=2 filter=47 channel=40
					-5, -2, -8, -15, -2, 0, -9, 8, 0,
					-- layer=2 filter=47 channel=41
					3, 0, 3, 3, -11, -1, 0, -6, -9,
					-- layer=2 filter=47 channel=42
					-8, 0, 8, -11, -9, 7, -8, 0, -3,
					-- layer=2 filter=47 channel=43
					3, -1, -1, -7, 6, 0, 0, 0, -7,
					-- layer=2 filter=47 channel=44
					2, -8, 0, -10, -6, 9, 7, -5, -8,
					-- layer=2 filter=47 channel=45
					-1, 9, 1, 3, -7, -8, 5, -3, -4,
					-- layer=2 filter=47 channel=46
					-9, 6, 4, -6, 0, 4, 2, 0, -8,
					-- layer=2 filter=47 channel=47
					-4, 4, -11, 0, 5, -6, -9, -10, 2,
					-- layer=2 filter=47 channel=48
					3, -7, 6, -2, -4, -6, 0, -6, 11,
					-- layer=2 filter=47 channel=49
					-2, -4, 2, -13, -21, 1, -3, -19, -6,
					-- layer=2 filter=47 channel=50
					-9, -8, 10, 0, 0, -5, 4, 8, -9,
					-- layer=2 filter=47 channel=51
					3, -3, -10, 0, -10, 4, -3, -3, -5,
					-- layer=2 filter=47 channel=52
					-9, -6, -14, 3, 0, -2, 3, -5, -11,
					-- layer=2 filter=47 channel=53
					-3, -9, -13, -14, 0, -16, 11, -1, 0,
					-- layer=2 filter=47 channel=54
					-3, -9, -10, -14, 1, -3, 0, 0, -5,
					-- layer=2 filter=47 channel=55
					-6, -3, 0, 0, -8, -7, 0, -10, 4,
					-- layer=2 filter=47 channel=56
					0, 4, -5, -1, -1, -9, -2, -3, -6,
					-- layer=2 filter=47 channel=57
					-6, -5, 6, -4, -4, 7, 5, -5, 0,
					-- layer=2 filter=47 channel=58
					-7, -2, -10, -7, 1, -6, -8, 9, 5,
					-- layer=2 filter=47 channel=59
					0, -18, -8, 2, -5, -14, 5, -8, -13,
					-- layer=2 filter=47 channel=60
					-7, 7, -6, -10, 0, 3, -1, -6, 6,
					-- layer=2 filter=47 channel=61
					4, -6, 2, 1, -11, 3, -8, -7, 3,
					-- layer=2 filter=47 channel=62
					5, 2, 8, -17, -4, -2, -9, -5, -3,
					-- layer=2 filter=47 channel=63
					-5, 10, 2, 2, -2, -3, -4, -7, -13,
					-- layer=2 filter=47 channel=64
					6, -12, 4, -8, 0, -6, 8, -6, 6,
					-- layer=2 filter=47 channel=65
					-3, -10, -1, -3, -7, -1, -11, 0, 2,
					-- layer=2 filter=47 channel=66
					-5, -10, -6, 8, 8, -6, 6, -3, -8,
					-- layer=2 filter=47 channel=67
					-6, -5, 1, -12, 0, -6, -6, -8, 0,
					-- layer=2 filter=47 channel=68
					-9, 7, -11, 0, -9, 6, 7, 4, -5,
					-- layer=2 filter=47 channel=69
					3, -5, 4, 6, -10, 0, 4, -5, 1,
					-- layer=2 filter=47 channel=70
					-1, 2, -9, -10, 4, 0, -6, -11, 12,
					-- layer=2 filter=47 channel=71
					-7, 3, 7, -8, -10, -2, 2, -4, -6,
					-- layer=2 filter=47 channel=72
					14, 1, -13, -9, -3, 7, -11, -13, 4,
					-- layer=2 filter=47 channel=73
					-15, 2, 8, -2, 6, -8, -5, -6, -7,
					-- layer=2 filter=47 channel=74
					0, 0, -5, 3, -10, -10, -1, 5, -13,
					-- layer=2 filter=47 channel=75
					5, -3, -8, -3, -9, 6, -2, -2, -1,
					-- layer=2 filter=47 channel=76
					-7, -9, -8, 0, 1, 7, 10, -3, -1,
					-- layer=2 filter=47 channel=77
					4, -10, 0, 4, 3, 1, -5, -5, -9,
					-- layer=2 filter=47 channel=78
					1, 7, -11, -11, 5, -5, 0, 2, 0,
					-- layer=2 filter=47 channel=79
					-8, 3, -4, 1, -2, -6, 6, 0, 1,
					-- layer=2 filter=47 channel=80
					0, 5, -8, -11, -5, 5, -1, -5, 1,
					-- layer=2 filter=47 channel=81
					6, 1, 8, 4, -1, -11, 3, -6, 5,
					-- layer=2 filter=47 channel=82
					-6, 5, 4, -7, -7, 0, 6, 1, -9,
					-- layer=2 filter=47 channel=83
					4, -4, -7, -8, -2, -7, 2, -9, 0,
					-- layer=2 filter=47 channel=84
					0, 0, 2, 6, 5, 2, -9, -7, -11,
					-- layer=2 filter=47 channel=85
					6, -6, 1, 10, 1, 1, 0, 7, -5,
					-- layer=2 filter=47 channel=86
					-1, -2, -7, -5, 11, 8, -3, -5, -5,
					-- layer=2 filter=47 channel=87
					-9, 0, 4, 6, 2, 5, -3, 5, 7,
					-- layer=2 filter=47 channel=88
					1, 5, 7, 0, -1, -2, -9, -3, -7,
					-- layer=2 filter=47 channel=89
					-8, -17, -12, -10, 7, -1, -6, -5, -6,
					-- layer=2 filter=47 channel=90
					6, -5, -9, -5, 6, -6, -3, 0, 0,
					-- layer=2 filter=47 channel=91
					3, 4, -1, -15, -4, 6, 0, 0, -2,
					-- layer=2 filter=47 channel=92
					0, -11, 0, -14, -9, -7, -4, -4, -4,
					-- layer=2 filter=47 channel=93
					-10, 0, 0, -7, 1, -5, -7, 7, 8,
					-- layer=2 filter=47 channel=94
					-6, -8, 2, 4, -7, -2, -12, -1, 0,
					-- layer=2 filter=47 channel=95
					0, 0, 3, -3, 4, -1, 6, 0, -1,
					-- layer=2 filter=47 channel=96
					-1, 0, -3, -4, -10, -6, 1, 2, 0,
					-- layer=2 filter=47 channel=97
					-10, -1, 0, -11, 0, -11, 6, -10, -3,
					-- layer=2 filter=47 channel=98
					9, 3, 0, -4, -11, 2, -11, 3, 4,
					-- layer=2 filter=47 channel=99
					-14, -1, 0, -5, 0, -11, 3, -13, -16,
					-- layer=2 filter=47 channel=100
					-6, -2, -1, 2, -4, 0, -12, -11, 4,
					-- layer=2 filter=47 channel=101
					-12, 0, 3, -11, 10, 11, -13, -9, 0,
					-- layer=2 filter=47 channel=102
					-10, -15, -4, -2, -15, -3, -6, 2, 2,
					-- layer=2 filter=47 channel=103
					-11, -10, -3, 9, -11, -6, 3, -10, 8,
					-- layer=2 filter=47 channel=104
					-5, 3, -5, 1, -13, -12, 10, -9, -10,
					-- layer=2 filter=47 channel=105
					6, 2, -6, -2, 0, 7, -10, -7, 0,
					-- layer=2 filter=47 channel=106
					0, -18, -9, -9, -8, -1, -15, -13, 6,
					-- layer=2 filter=47 channel=107
					0, 0, -4, 0, -1, 2, 6, 3, -8,
					-- layer=2 filter=47 channel=108
					-3, -1, -1, 2, 5, -13, 9, -2, 2,
					-- layer=2 filter=47 channel=109
					7, -5, 5, 4, -8, -4, -11, -6, -4,
					-- layer=2 filter=47 channel=110
					9, 0, -2, -4, -3, 0, 4, -4, 3,
					-- layer=2 filter=47 channel=111
					0, 2, -8, -3, -5, 6, -11, 2, 2,
					-- layer=2 filter=47 channel=112
					-2, 0, -1, -6, -2, -2, -8, 1, 0,
					-- layer=2 filter=47 channel=113
					-3, -8, -5, -3, -2, 3, 5, -9, -3,
					-- layer=2 filter=47 channel=114
					-8, -8, 5, 7, 2, 3, 6, 7, -10,
					-- layer=2 filter=47 channel=115
					9, -6, 6, -8, -2, -2, -3, 6, 2,
					-- layer=2 filter=47 channel=116
					0, -2, 0, -11, 0, 4, 3, -9, 4,
					-- layer=2 filter=47 channel=117
					-3, -5, -1, -15, 6, 10, -9, -8, -5,
					-- layer=2 filter=47 channel=118
					6, 7, -2, -11, -9, 0, -5, -8, 0,
					-- layer=2 filter=47 channel=119
					-6, 3, -3, -5, -8, -12, -11, -3, -3,
					-- layer=2 filter=47 channel=120
					9, 10, -9, 3, -3, 2, -9, -6, -8,
					-- layer=2 filter=47 channel=121
					-5, 0, 5, 0, -9, 5, -9, -3, 1,
					-- layer=2 filter=47 channel=122
					-9, -4, -9, -1, -7, -7, -5, 3, -3,
					-- layer=2 filter=47 channel=123
					9, 13, 2, 0, -2, 3, -14, 0, -15,
					-- layer=2 filter=47 channel=124
					-1, 4, -11, 0, -6, -3, 8, -10, 4,
					-- layer=2 filter=47 channel=125
					8, -1, 1, 7, -3, 5, 5, 5, -1,
					-- layer=2 filter=47 channel=126
					-10, 8, 4, 8, 2, 7, 2, -3, 6,
					-- layer=2 filter=47 channel=127
					-2, -7, 9, 5, 0, 6, 3, 0, 1,
					-- layer=2 filter=48 channel=0
					-20, -8, -12, -12, -7, -12, -24, -6, -14,
					-- layer=2 filter=48 channel=1
					3, -3, -11, -20, -2, -23, 9, -9, -19,
					-- layer=2 filter=48 channel=2
					4, 0, -6, -10, -3, -4, 11, -1, 4,
					-- layer=2 filter=48 channel=3
					0, -14, -4, 0, 0, -4, -24, -18, -22,
					-- layer=2 filter=48 channel=4
					-23, -6, -28, -12, 0, -6, -15, -13, -5,
					-- layer=2 filter=48 channel=5
					-10, -27, -24, -17, -7, -14, -4, -19, 0,
					-- layer=2 filter=48 channel=6
					-20, -22, 7, 13, 5, 11, 3, -15, -7,
					-- layer=2 filter=48 channel=7
					8, -4, 13, 5, -18, 6, -18, -12, 7,
					-- layer=2 filter=48 channel=8
					0, -6, -4, 9, -1, -1, 4, -10, 4,
					-- layer=2 filter=48 channel=9
					-24, -18, -13, -23, -5, -12, -16, -6, -11,
					-- layer=2 filter=48 channel=10
					-21, -12, -22, -15, -23, -12, -21, -20, -19,
					-- layer=2 filter=48 channel=11
					-10, 2, -13, -2, -11, 0, -10, -4, -5,
					-- layer=2 filter=48 channel=12
					-4, -1, 7, -5, -1, -5, 6, 0, 0,
					-- layer=2 filter=48 channel=13
					9, 10, 8, 3, 0, 4, -1, 8, 1,
					-- layer=2 filter=48 channel=14
					1, -17, -1, -6, -17, -23, 9, -8, -4,
					-- layer=2 filter=48 channel=15
					0, 7, -8, 2, -6, 18, -3, 16, -4,
					-- layer=2 filter=48 channel=16
					-3, -9, -18, -20, -13, -6, -13, -7, 15,
					-- layer=2 filter=48 channel=17
					0, 5, 8, 0, 2, 5, -9, 5, 7,
					-- layer=2 filter=48 channel=18
					-45, 5, -20, -23, 12, -14, -2, -20, 0,
					-- layer=2 filter=48 channel=19
					0, -1, 6, -6, -7, -19, 6, -3, -20,
					-- layer=2 filter=48 channel=20
					-7, 10, 7, 12, 6, 6, 1, 0, 6,
					-- layer=2 filter=48 channel=21
					-10, -10, -8, 7, 0, -6, -12, -10, 1,
					-- layer=2 filter=48 channel=22
					-2, 7, -4, 6, 0, -7, 0, -6, -5,
					-- layer=2 filter=48 channel=23
					-21, -3, -12, -7, -3, -15, -13, -5, -11,
					-- layer=2 filter=48 channel=24
					4, -7, -2, -9, 0, 0, -20, -14, -14,
					-- layer=2 filter=48 channel=25
					4, -5, -1, -1, -1, 10, -16, -6, -2,
					-- layer=2 filter=48 channel=26
					6, -5, 1, 7, 0, 2, -5, 4, 6,
					-- layer=2 filter=48 channel=27
					-10, -19, -16, -7, 2, -15, 4, 6, 12,
					-- layer=2 filter=48 channel=28
					-22, -2, 24, 1, -15, 13, -13, -26, -6,
					-- layer=2 filter=48 channel=29
					7, -3, -9, 6, -9, 4, -1, -3, -7,
					-- layer=2 filter=48 channel=30
					-8, -30, -17, -7, -5, -3, -2, -14, -10,
					-- layer=2 filter=48 channel=31
					5, 4, 7, -9, 0, 12, -1, -5, -3,
					-- layer=2 filter=48 channel=32
					10, -3, 3, -8, 0, -9, -1, -6, -2,
					-- layer=2 filter=48 channel=33
					-3, 5, -7, -12, -14, -6, -30, 2, -8,
					-- layer=2 filter=48 channel=34
					-15, 1, 2, 5, 0, -11, 18, -29, 0,
					-- layer=2 filter=48 channel=35
					-8, 6, 4, 11, -2, -5, -8, -27, -1,
					-- layer=2 filter=48 channel=36
					-3, -6, -2, 6, -8, 3, -5, 1, 8,
					-- layer=2 filter=48 channel=37
					-16, -10, -10, -17, -11, -24, -4, 7, 1,
					-- layer=2 filter=48 channel=38
					-3, -22, -21, -10, -14, -6, -16, -8, -7,
					-- layer=2 filter=48 channel=39
					8, -3, 12, 7, -5, -4, -16, 8, 3,
					-- layer=2 filter=48 channel=40
					-4, -3, 6, 2, -16, 23, 12, 13, 27,
					-- layer=2 filter=48 channel=41
					-3, -4, 6, -4, -1, -3, 4, -2, 7,
					-- layer=2 filter=48 channel=42
					-1, 5, -6, -1, 3, 9, -4, 2, -1,
					-- layer=2 filter=48 channel=43
					-17, -10, -7, 0, -4, -11, -15, -9, -2,
					-- layer=2 filter=48 channel=44
					-6, -1, 7, -2, -9, -3, -10, -7, -11,
					-- layer=2 filter=48 channel=45
					-1, 1, 0, -4, -11, 11, -13, 7, 6,
					-- layer=2 filter=48 channel=46
					-5, -30, -22, -14, -20, -6, -25, -1, -10,
					-- layer=2 filter=48 channel=47
					4, 1, 17, 18, 3, -1, -8, -26, 6,
					-- layer=2 filter=48 channel=48
					4, -6, 6, -9, 4, -4, 6, 8, 0,
					-- layer=2 filter=48 channel=49
					-31, -11, -27, -12, -1, -26, 2, -16, -9,
					-- layer=2 filter=48 channel=50
					-2, 3, 26, 11, 12, 3, 6, -8, 3,
					-- layer=2 filter=48 channel=51
					-8, -11, -4, 1, -26, -14, -14, -21, -13,
					-- layer=2 filter=48 channel=52
					-1, 3, -3, 0, -14, -11, -8, -10, -6,
					-- layer=2 filter=48 channel=53
					6, -31, -2, 1, -19, -3, -5, 5, 5,
					-- layer=2 filter=48 channel=54
					-4, 8, 5, 9, 9, 1, -13, -3, 1,
					-- layer=2 filter=48 channel=55
					-3, -2, 6, -5, 1, 2, -3, -5, -4,
					-- layer=2 filter=48 channel=56
					1, -3, -19, -10, -9, -21, -5, -14, 3,
					-- layer=2 filter=48 channel=57
					-2, 4, -1, 10, -6, 5, 6, 0, -4,
					-- layer=2 filter=48 channel=58
					9, -2, 5, -12, -14, -2, 19, 23, -15,
					-- layer=2 filter=48 channel=59
					6, -1, 4, -3, -19, 0, 12, 17, -8,
					-- layer=2 filter=48 channel=60
					6, 0, 8, 7, -14, -9, 6, 0, -6,
					-- layer=2 filter=48 channel=61
					-33, -29, -6, -2, 1, -3, -3, -15, -27,
					-- layer=2 filter=48 channel=62
					-12, -12, -18, -18, 4, -3, 7, -14, -1,
					-- layer=2 filter=48 channel=63
					-11, -18, -15, -7, 9, 0, -17, -15, -11,
					-- layer=2 filter=48 channel=64
					-2, 1, -7, -6, 6, 7, -3, -7, -12,
					-- layer=2 filter=48 channel=65
					-10, -23, 2, -7, -12, 4, -4, -18, -19,
					-- layer=2 filter=48 channel=66
					-1, -3, -1, -7, 2, 3, 3, -13, 0,
					-- layer=2 filter=48 channel=67
					-23, -29, -25, -22, -17, -21, -12, -4, -17,
					-- layer=2 filter=48 channel=68
					-4, -11, 5, 8, -8, -3, 6, -3, 9,
					-- layer=2 filter=48 channel=69
					3, -16, -5, -16, 0, 5, 6, 4, 8,
					-- layer=2 filter=48 channel=70
					-19, -6, 14, 3, 6, 0, -19, -18, 3,
					-- layer=2 filter=48 channel=71
					-1, -9, -7, -14, -12, -21, -2, 11, -7,
					-- layer=2 filter=48 channel=72
					4, 7, 4, -8, -7, -14, -21, -19, 0,
					-- layer=2 filter=48 channel=73
					15, -15, -7, -12, -10, -3, -8, 3, -20,
					-- layer=2 filter=48 channel=74
					1, -2, -10, -8, -16, -15, -7, -1, -17,
					-- layer=2 filter=48 channel=75
					-9, -5, 13, -31, -13, -5, 29, 16, 13,
					-- layer=2 filter=48 channel=76
					16, -5, 7, 17, -23, 7, -1, 8, 2,
					-- layer=2 filter=48 channel=77
					4, 9, 8, 7, -1, -1, -1, -12, 5,
					-- layer=2 filter=48 channel=78
					1, 7, -15, 0, -12, -12, -11, 4, 1,
					-- layer=2 filter=48 channel=79
					8, 5, 2, -1, -1, 3, 1, -4, -2,
					-- layer=2 filter=48 channel=80
					-7, -19, -23, -7, -9, -2, -18, -7, -6,
					-- layer=2 filter=48 channel=81
					7, 7, 5, 2, -11, 7, -11, -6, 0,
					-- layer=2 filter=48 channel=82
					1, -4, 10, 1, 0, 8, 6, 8, 8,
					-- layer=2 filter=48 channel=83
					-22, -30, -18, -17, -20, 0, 0, -3, -3,
					-- layer=2 filter=48 channel=84
					3, 3, -7, 5, -6, -3, 5, 1, 0,
					-- layer=2 filter=48 channel=85
					-1, 0, -4, 3, 11, 8, 4, -6, 7,
					-- layer=2 filter=48 channel=86
					1, -8, -5, 0, 6, 4, 9, 1, -4,
					-- layer=2 filter=48 channel=87
					-24, 6, -9, 10, -10, 10, 4, -3, -2,
					-- layer=2 filter=48 channel=88
					-14, 7, -1, -4, -12, -15, -5, -5, -12,
					-- layer=2 filter=48 channel=89
					4, -1, 9, -24, -8, -18, -5, -2, -4,
					-- layer=2 filter=48 channel=90
					1, -2, -4, 8, 4, -7, 3, -4, -5,
					-- layer=2 filter=48 channel=91
					24, 12, 1, -15, -8, -7, 19, -9, -7,
					-- layer=2 filter=48 channel=92
					-8, 0, 5, -4, -9, -14, 6, -5, -1,
					-- layer=2 filter=48 channel=93
					9, 8, 0, 4, 17, 10, 0, -5, -19,
					-- layer=2 filter=48 channel=94
					-25, -34, -3, 6, -18, -9, 7, 7, -10,
					-- layer=2 filter=48 channel=95
					4, -7, 6, 6, -4, 3, -11, -12, 6,
					-- layer=2 filter=48 channel=96
					-4, 10, -4, -12, -7, -14, -3, 7, -25,
					-- layer=2 filter=48 channel=97
					-8, -12, -16, -10, -2, -5, -16, -4, 0,
					-- layer=2 filter=48 channel=98
					-22, 6, 4, 0, -9, 2, -12, -23, -9,
					-- layer=2 filter=48 channel=99
					-6, 7, -4, -4, -20, -9, 7, -3, -6,
					-- layer=2 filter=48 channel=100
					-22, -12, -21, -9, -7, -18, -10, 11, -6,
					-- layer=2 filter=48 channel=101
					6, -10, -12, 1, -24, -17, -1, -20, -7,
					-- layer=2 filter=48 channel=102
					-16, 10, -13, -16, 9, -16, -7, -24, 7,
					-- layer=2 filter=48 channel=103
					-9, 6, -7, -4, -7, -11, -11, -21, -9,
					-- layer=2 filter=48 channel=104
					-22, -6, -20, 5, 0, -8, -1, -8, -4,
					-- layer=2 filter=48 channel=105
					5, 16, -6, -16, -9, 2, -18, 12, -15,
					-- layer=2 filter=48 channel=106
					17, 7, 11, 0, -9, -2, -7, -13, -9,
					-- layer=2 filter=48 channel=107
					-4, 12, -4, -1, -13, -7, 3, -4, 6,
					-- layer=2 filter=48 channel=108
					-12, -4, -11, -1, -8, -11, 3, -2, -9,
					-- layer=2 filter=48 channel=109
					-2, 8, -7, -4, 0, 0, 11, -4, 11,
					-- layer=2 filter=48 channel=110
					10, 11, 27, -1, 16, 16, -2, 5, 15,
					-- layer=2 filter=48 channel=111
					3, 2, 2, 4, -9, 11, -8, -6, -5,
					-- layer=2 filter=48 channel=112
					-11, -30, -27, -17, -15, -26, -20, -34, -8,
					-- layer=2 filter=48 channel=113
					-17, -24, -14, -8, -16, -3, -6, -11, -4,
					-- layer=2 filter=48 channel=114
					-7, 2, -5, -9, -8, -4, 8, -6, 7,
					-- layer=2 filter=48 channel=115
					2, 5, 6, 3, 8, 3, -11, -4, 3,
					-- layer=2 filter=48 channel=116
					-32, 4, -9, -2, -6, 2, 8, -11, -13,
					-- layer=2 filter=48 channel=117
					-3, -1, -4, 1, -6, 7, -3, -9, -16,
					-- layer=2 filter=48 channel=118
					-26, -16, -21, -17, -8, -6, -17, -17, -17,
					-- layer=2 filter=48 channel=119
					-26, -3, -21, 10, 13, -22, 5, -6, 11,
					-- layer=2 filter=48 channel=120
					-4, 2, 2, 0, -2, -4, 5, 9, -9,
					-- layer=2 filter=48 channel=121
					8, 10, 4, 9, 12, 1, 0, 3, 7,
					-- layer=2 filter=48 channel=122
					6, 3, -1, -2, 4, 0, 2, -7, 9,
					-- layer=2 filter=48 channel=123
					-1, 3, 16, 0, -13, 0, -4, 0, 12,
					-- layer=2 filter=48 channel=124
					-10, -5, 5, 0, -23, 12, -3, 6, -4,
					-- layer=2 filter=48 channel=125
					5, -7, 2, 8, -6, 1, 0, 0, -4,
					-- layer=2 filter=48 channel=126
					-4, -18, 10, 3, 9, -26, 15, 11, -4,
					-- layer=2 filter=48 channel=127
					-8, 0, -2, 0, -7, -6, -17, -2, -8,
					-- layer=2 filter=49 channel=0
					-5, -37, -11, -28, -29, -13, 0, 0, 21,
					-- layer=2 filter=49 channel=1
					-31, -53, -50, -18, -40, -6, 5, 8, -14,
					-- layer=2 filter=49 channel=2
					6, 3, -4, -3, 11, 3, 0, -2, 10,
					-- layer=2 filter=49 channel=3
					15, 11, -25, 1, -12, -7, 25, -9, 27,
					-- layer=2 filter=49 channel=4
					-2, -12, 0, -9, 10, 3, 14, 21, 0,
					-- layer=2 filter=49 channel=5
					-16, -28, -35, -7, -20, 8, -7, -15, 7,
					-- layer=2 filter=49 channel=6
					6, -10, -59, 0, 56, -32, 66, -90, 13,
					-- layer=2 filter=49 channel=7
					-4, -2, -29, -23, 1, 26, 16, 33, 22,
					-- layer=2 filter=49 channel=8
					6, 0, -1, 0, 7, 2, -2, -5, 3,
					-- layer=2 filter=49 channel=9
					4, -6, 18, -42, 5, 13, -22, -11, -22,
					-- layer=2 filter=49 channel=10
					14, -2, 13, 26, 4, 29, 10, 35, 26,
					-- layer=2 filter=49 channel=11
					-12, -42, -24, -43, -43, -34, 15, -23, 2,
					-- layer=2 filter=49 channel=12
					-29, -40, -59, 0, 0, 8, 0, 4, 16,
					-- layer=2 filter=49 channel=13
					8, -6, -6, -8, -6, 8, -11, -10, -3,
					-- layer=2 filter=49 channel=14
					-27, -81, -65, -24, -20, -11, -28, 2, 2,
					-- layer=2 filter=49 channel=15
					-49, -18, -35, -11, 62, -69, -57, -17, 28,
					-- layer=2 filter=49 channel=16
					2, -1, -9, 12, 38, 14, 38, 9, -13,
					-- layer=2 filter=49 channel=17
					7, -1, -4, -5, 7, 2, 8, 2, -8,
					-- layer=2 filter=49 channel=18
					-43, -23, -43, -40, -56, -16, -38, -16, -103,
					-- layer=2 filter=49 channel=19
					-10, -13, -26, 29, -18, -24, -18, -75, 2,
					-- layer=2 filter=49 channel=20
					-7, -8, 1, -3, -9, 0, 0, 5, -7,
					-- layer=2 filter=49 channel=21
					-6, 20, 14, -8, 13, 14, -21, 5, 14,
					-- layer=2 filter=49 channel=22
					-11, -1, -8, -10, 5, 0, 5, 4, 6,
					-- layer=2 filter=49 channel=23
					12, -7, 23, 24, 9, -3, 25, 24, 12,
					-- layer=2 filter=49 channel=24
					9, 1, -4, -14, 3, -20, 15, -30, -8,
					-- layer=2 filter=49 channel=25
					-26, -8, -5, -15, -15, -3, -7, -28, 4,
					-- layer=2 filter=49 channel=26
					7, -5, 9, 0, 4, -8, -5, -6, 10,
					-- layer=2 filter=49 channel=27
					-17, -35, -25, 6, -8, 24, -19, 2, -23,
					-- layer=2 filter=49 channel=28
					-32, -4, -21, 12, -43, -12, 18, 19, 20,
					-- layer=2 filter=49 channel=29
					9, 12, 2, 0, -5, 10, 0, 1, 0,
					-- layer=2 filter=49 channel=30
					9, 15, 15, 9, 6, 8, -12, 31, -1,
					-- layer=2 filter=49 channel=31
					-17, -13, -32, -29, 30, 2, -73, -29, 2,
					-- layer=2 filter=49 channel=32
					4, 0, -9, -10, 11, -2, 9, -7, 5,
					-- layer=2 filter=49 channel=33
					-24, 7, 5, -41, 29, -21, -7, -7, -29,
					-- layer=2 filter=49 channel=34
					15, 37, -13, 6, -15, 40, 50, 41, -35,
					-- layer=2 filter=49 channel=35
					-49, 0, -50, -13, -10, -3, 1, 26, 27,
					-- layer=2 filter=49 channel=36
					9, 1, 1, -7, 0, 0, -11, 4, 5,
					-- layer=2 filter=49 channel=37
					-31, -28, -37, -10, -61, -29, 17, -6, 2,
					-- layer=2 filter=49 channel=38
					-11, -49, -22, -19, 0, -2, 10, -6, -24,
					-- layer=2 filter=49 channel=39
					-15, 0, -3, -6, 12, 27, 8, 19, 4,
					-- layer=2 filter=49 channel=40
					-44, -43, -5, -18, 29, -52, 0, -35, -33,
					-- layer=2 filter=49 channel=41
					-1, 0, -9, 7, -8, 7, -1, -10, 1,
					-- layer=2 filter=49 channel=42
					7, 10, -2, 21, 20, -7, -2, 24, 20,
					-- layer=2 filter=49 channel=43
					-14, -13, -10, -6, -24, 18, 28, 1, 3,
					-- layer=2 filter=49 channel=44
					1, -2, 0, -3, 6, 4, 6, -8, 0,
					-- layer=2 filter=49 channel=45
					3, -48, -55, 5, -33, 22, -56, -16, 22,
					-- layer=2 filter=49 channel=46
					22, 5, -3, 17, -1, -13, 18, 29, -12,
					-- layer=2 filter=49 channel=47
					-21, -20, 6, -16, 3, 12, 26, 44, 12,
					-- layer=2 filter=49 channel=48
					5, 5, 7, -11, -4, 0, 0, -6, -2,
					-- layer=2 filter=49 channel=49
					19, -17, -28, 3, -32, 5, -21, -18, 11,
					-- layer=2 filter=49 channel=50
					14, -22, 17, 13, 8, 9, 9, 0, 13,
					-- layer=2 filter=49 channel=51
					-9, -43, -23, -34, -33, -1, 11, -4, 30,
					-- layer=2 filter=49 channel=52
					-18, -19, -55, -17, -23, -26, 58, 11, -5,
					-- layer=2 filter=49 channel=53
					21, -59, -114, 4, 4, -27, -13, -46, -29,
					-- layer=2 filter=49 channel=54
					-19, -2, -10, -31, -18, -5, 34, 21, 64,
					-- layer=2 filter=49 channel=55
					-2, -8, 0, 5, 0, -3, -10, 14, -5,
					-- layer=2 filter=49 channel=56
					-21, -28, -31, -7, -49, -17, -25, -22, -58,
					-- layer=2 filter=49 channel=57
					-2, -2, -8, 0, 6, -6, 1, 1, 3,
					-- layer=2 filter=49 channel=58
					-19, -18, -20, 2, 3, 20, 3, -30, 32,
					-- layer=2 filter=49 channel=59
					-19, -41, -26, 15, -6, -20, -26, -15, -49,
					-- layer=2 filter=49 channel=60
					-6, 3, 11, -3, -51, -27, 13, -21, 42,
					-- layer=2 filter=49 channel=61
					-10, -58, -15, -29, -15, -11, 17, 29, 7,
					-- layer=2 filter=49 channel=62
					14, -9, -44, 2, -2, -38, 31, -45, -55,
					-- layer=2 filter=49 channel=63
					-21, -17, -8, 5, -16, -7, 15, 20, 11,
					-- layer=2 filter=49 channel=64
					9, -4, 0, 6, 15, -15, 2, 16, 1,
					-- layer=2 filter=49 channel=65
					-6, -38, -28, 11, 36, -49, 32, 1, -15,
					-- layer=2 filter=49 channel=66
					14, 10, 6, 22, -29, 10, -18, 3, -9,
					-- layer=2 filter=49 channel=67
					24, 15, 19, -2, -17, -4, 4, -24, -36,
					-- layer=2 filter=49 channel=68
					-5, -2, 2, 8, 2, -7, 10, 5, -7,
					-- layer=2 filter=49 channel=69
					12, 11, 8, -1, 15, 0, 0, 24, 15,
					-- layer=2 filter=49 channel=70
					-19, 7, -34, -16, -31, -33, 21, 37, 49,
					-- layer=2 filter=49 channel=71
					-33, 2, 25, -59, -3, 20, -82, -22, -10,
					-- layer=2 filter=49 channel=72
					-70, 7, 0, -22, -16, -36, -27, -51, 0,
					-- layer=2 filter=49 channel=73
					9, -9, -6, 72, 14, 34, 62, 12, 33,
					-- layer=2 filter=49 channel=74
					14, -9, -16, 13, 0, -7, -12, 2, 1,
					-- layer=2 filter=49 channel=75
					2, -25, -78, -77, -78, 15, -46, 28, 16,
					-- layer=2 filter=49 channel=76
					25, -2, 9, -10, -44, -60, 17, -40, 3,
					-- layer=2 filter=49 channel=77
					-2, -6, -6, 10, -3, -2, 0, -7, 10,
					-- layer=2 filter=49 channel=78
					-26, -17, -20, -27, -18, -13, 2, 15, -27,
					-- layer=2 filter=49 channel=79
					-3, -8, 7, -6, -5, -2, 0, 0, 9,
					-- layer=2 filter=49 channel=80
					8, 14, -2, 25, 28, -5, 28, 6, -2,
					-- layer=2 filter=49 channel=81
					-3, -5, 0, -1, -1, 6, 11, 4, 0,
					-- layer=2 filter=49 channel=82
					0, 11, -5, 11, -6, -8, -6, -6, -2,
					-- layer=2 filter=49 channel=83
					-4, 0, 2, 28, 27, 13, 9, 33, 19,
					-- layer=2 filter=49 channel=84
					-8, 8, -7, -4, -8, 1, 0, -6, 7,
					-- layer=2 filter=49 channel=85
					11, 3, 12, -14, 1, 0, -18, 4, 0,
					-- layer=2 filter=49 channel=86
					16, -5, 4, 16, 2, -20, -13, 7, -6,
					-- layer=2 filter=49 channel=87
					48, 9, 14, -20, 19, -18, 11, 18, -45,
					-- layer=2 filter=49 channel=88
					0, -8, -12, -6, 4, 0, -3, 9, -6,
					-- layer=2 filter=49 channel=89
					1, -7, -30, -15, -14, -42, -8, -17, -4,
					-- layer=2 filter=49 channel=90
					3, -2, -8, 0, 8, -2, 5, 6, 1,
					-- layer=2 filter=49 channel=91
					-57, -31, -42, -22, -24, -24, 23, -23, 29,
					-- layer=2 filter=49 channel=92
					-46, -53, -31, -11, -11, -35, -16, -21, -2,
					-- layer=2 filter=49 channel=93
					68, 13, -38, 57, 26, -36, 18, -51, -45,
					-- layer=2 filter=49 channel=94
					-28, -14, 25, 0, 12, -1, 49, -30, 4,
					-- layer=2 filter=49 channel=95
					-15, -8, -9, -1, 3, -7, 2, 2, 5,
					-- layer=2 filter=49 channel=96
					31, -47, -14, 50, -64, 1, 66, -65, -15,
					-- layer=2 filter=49 channel=97
					10, -5, -12, -29, -25, -6, -34, -12, 16,
					-- layer=2 filter=49 channel=98
					-13, -6, 1, -41, -13, -5, 36, 53, 38,
					-- layer=2 filter=49 channel=99
					32, -31, 0, 9, -39, -8, 29, 15, 5,
					-- layer=2 filter=49 channel=100
					13, 13, 6, 3, 0, 22, 14, -15, 9,
					-- layer=2 filter=49 channel=101
					-32, -42, -23, -70, -56, -9, -52, -21, -7,
					-- layer=2 filter=49 channel=102
					-17, -21, 0, 8, -24, 16, 23, -28, -6,
					-- layer=2 filter=49 channel=103
					-29, 23, -42, -18, -39, -23, 59, -16, -11,
					-- layer=2 filter=49 channel=104
					14, 20, 26, 19, -20, -64, -8, -28, 0,
					-- layer=2 filter=49 channel=105
					81, -2, 24, -11, 43, -33, 42, -30, -31,
					-- layer=2 filter=49 channel=106
					-33, -51, -38, -21, -56, -9, -8, -48, -17,
					-- layer=2 filter=49 channel=107
					-30, 2, -34, 3, 14, -23, 2, -2, 18,
					-- layer=2 filter=49 channel=108
					-16, -77, -26, 4, -36, 37, 23, -31, 38,
					-- layer=2 filter=49 channel=109
					6, 0, 7, -1, -2, 8, 12, 0, 10,
					-- layer=2 filter=49 channel=110
					-17, 8, -19, -8, -8, -35, -37, 9, -16,
					-- layer=2 filter=49 channel=111
					-6, 3, 8, 2, 2, -7, -7, 0, 6,
					-- layer=2 filter=49 channel=112
					-9, -68, 17, 13, -23, 29, -6, 74, 37,
					-- layer=2 filter=49 channel=113
					-19, 3, 14, 24, 26, 3, 0, 26, 7,
					-- layer=2 filter=49 channel=114
					1, 8, 6, 14, 9, 10, -14, -5, 8,
					-- layer=2 filter=49 channel=115
					0, -2, -6, 8, 0, -4, -1, -5, 7,
					-- layer=2 filter=49 channel=116
					15, -7, -2, 17, -16, 2, 28, -7, -57,
					-- layer=2 filter=49 channel=117
					-10, -27, -5, -7, 6, 12, 1, -1, 10,
					-- layer=2 filter=49 channel=118
					11, 12, 5, 23, 4, 10, 67, 33, -2,
					-- layer=2 filter=49 channel=119
					-8, 15, -19, 0, 8, 6, 10, 15, 2,
					-- layer=2 filter=49 channel=120
					-8, -7, -3, 4, -5, 8, 5, -10, 10,
					-- layer=2 filter=49 channel=121
					-2, 11, 6, -8, 4, 0, -10, 4, -2,
					-- layer=2 filter=49 channel=122
					-10, -5, -10, -13, 2, 4, 4, -4, -4,
					-- layer=2 filter=49 channel=123
					-9, 7, 24, -24, 10, -11, 24, 4, 2,
					-- layer=2 filter=49 channel=124
					36, -15, -32, -25, 44, -65, -14, 0, -29,
					-- layer=2 filter=49 channel=125
					-7, -7, -4, 3, -2, 10, -6, -6, 4,
					-- layer=2 filter=49 channel=126
					8, 6, -45, -15, -26, -53, 13, -120, -16,
					-- layer=2 filter=49 channel=127
					7, -21, 10, -6, 3, -5, -27, 14, -9,
					-- layer=2 filter=50 channel=0
					-9, -18, 11, -14, -4, 10, 35, 13, 22,
					-- layer=2 filter=50 channel=1
					19, 29, 16, -12, 26, 27, -27, -62, -28,
					-- layer=2 filter=50 channel=2
					-8, 8, 9, 3, -4, -7, 0, -12, -2,
					-- layer=2 filter=50 channel=3
					-13, -32, -48, 22, -56, -34, 58, 55, 34,
					-- layer=2 filter=50 channel=4
					-27, 7, -14, 9, 5, -7, 47, 0, -10,
					-- layer=2 filter=50 channel=5
					-12, -5, 28, -24, -12, 15, 4, -4, -2,
					-- layer=2 filter=50 channel=6
					9, 19, 0, 34, 13, 58, -6, -11, 17,
					-- layer=2 filter=50 channel=7
					20, 27, 19, 50, 28, 18, -2, 21, 12,
					-- layer=2 filter=50 channel=8
					-3, 1, 9, 3, 0, 6, 9, 0, -2,
					-- layer=2 filter=50 channel=9
					-36, -10, 1, 28, 11, -30, 49, 70, 29,
					-- layer=2 filter=50 channel=10
					-24, -15, 0, 8, -12, -38, 54, 43, 14,
					-- layer=2 filter=50 channel=11
					-6, 15, 37, -14, -18, 12, 0, -6, 11,
					-- layer=2 filter=50 channel=12
					36, 14, 24, 22, 25, 47, -61, -83, -3,
					-- layer=2 filter=50 channel=13
					9, 11, 3, -7, 2, 4, -2, 5, -3,
					-- layer=2 filter=50 channel=14
					21, 32, 15, -32, -6, 7, -59, -84, -57,
					-- layer=2 filter=50 channel=15
					-56, 7, -15, -86, 11, 21, -60, 3, 19,
					-- layer=2 filter=50 channel=16
					-14, -5, 19, -25, -33, -16, -32, -39, -66,
					-- layer=2 filter=50 channel=17
					-10, -4, 10, 10, 8, 2, 10, 3, -5,
					-- layer=2 filter=50 channel=18
					-27, 2, -25, 10, -18, 1, 9, -28, 9,
					-- layer=2 filter=50 channel=19
					27, 31, 8, 6, 51, 20, -55, -18, 13,
					-- layer=2 filter=50 channel=20
					-5, 2, -5, -3, 0, -9, -7, 0, 5,
					-- layer=2 filter=50 channel=21
					-16, 4, -19, 1, 9, 9, -1, 5, 7,
					-- layer=2 filter=50 channel=22
					5, -3, 3, -6, -3, 7, 3, -8, -10,
					-- layer=2 filter=50 channel=23
					19, 15, -16, 29, 49, -3, 30, 5, -23,
					-- layer=2 filter=50 channel=24
					4, -8, 13, -25, -92, -78, 30, 10, 8,
					-- layer=2 filter=50 channel=25
					0, -8, 16, -26, -75, -23, 9, -19, 3,
					-- layer=2 filter=50 channel=26
					3, 5, 0, -4, -5, 2, 8, -9, 1,
					-- layer=2 filter=50 channel=27
					11, 32, 41, -45, -28, 13, -57, -56, -22,
					-- layer=2 filter=50 channel=28
					4, -18, -8, -11, 13, -13, 4, 22, 31,
					-- layer=2 filter=50 channel=29
					7, -1, -6, -3, 0, -9, 7, 1, -1,
					-- layer=2 filter=50 channel=30
					-50, -17, -7, -16, 3, 2, 1, 22, 4,
					-- layer=2 filter=50 channel=31
					-8, -19, -21, 1, -47, -4, -20, -7, 42,
					-- layer=2 filter=50 channel=32
					-8, -7, -2, 0, -6, 0, 8, -7, 6,
					-- layer=2 filter=50 channel=33
					-6, -18, -5, -29, -62, -24, -49, -37, 22,
					-- layer=2 filter=50 channel=34
					4, -9, -14, -12, 9, 26, 1, 17, 20,
					-- layer=2 filter=50 channel=35
					12, -22, -16, -34, -19, -29, -10, -2, -3,
					-- layer=2 filter=50 channel=36
					0, -8, -4, -1, 10, 3, -2, 3, 2,
					-- layer=2 filter=50 channel=37
					1, 5, 41, -13, -7, 16, -19, -12, 6,
					-- layer=2 filter=50 channel=38
					9, 27, 31, -20, -36, 0, -46, -30, -27,
					-- layer=2 filter=50 channel=39
					-66, -16, -11, 4, -35, -17, -3, 17, -69,
					-- layer=2 filter=50 channel=40
					17, 24, 52, 29, 8, 5, -21, -3, 30,
					-- layer=2 filter=50 channel=41
					-8, 0, 6, -5, -5, -8, -10, 2, 1,
					-- layer=2 filter=50 channel=42
					24, 36, 21, 34, 20, -12, -10, -4, -33,
					-- layer=2 filter=50 channel=43
					-17, 11, 25, -13, -40, -44, 59, 25, 10,
					-- layer=2 filter=50 channel=44
					8, 3, 5, 0, 1, 5, 12, 10, 6,
					-- layer=2 filter=50 channel=45
					2, -10, 30, -44, -69, -3, -41, -40, -51,
					-- layer=2 filter=50 channel=46
					-45, -4, -10, -2, 3, -48, 4, 15, -21,
					-- layer=2 filter=50 channel=47
					5, 19, 21, -15, -29, -9, 17, 5, 31,
					-- layer=2 filter=50 channel=48
					5, -5, -2, -7, 3, 2, 3, 10, -2,
					-- layer=2 filter=50 channel=49
					-34, -3, -32, -16, -33, -6, -17, 12, -33,
					-- layer=2 filter=50 channel=50
					5, 4, 24, 12, 10, -19, -10, 3, 5,
					-- layer=2 filter=50 channel=51
					3, 1, 21, -17, -9, 12, 17, 25, 11,
					-- layer=2 filter=50 channel=52
					-25, -9, 9, -43, 28, 8, 8, 3, 1,
					-- layer=2 filter=50 channel=53
					-25, 4, 21, 15, -9, 18, 19, -19, 26,
					-- layer=2 filter=50 channel=54
					-7, -19, -19, 6, 21, 9, -5, -1, 20,
					-- layer=2 filter=50 channel=55
					10, 6, 3, -2, 9, 0, 0, -10, -5,
					-- layer=2 filter=50 channel=56
					-14, 21, 22, -17, -25, 6, 6, -8, 8,
					-- layer=2 filter=50 channel=57
					-5, -11, 15, -10, 7, 13, -8, 5, 5,
					-- layer=2 filter=50 channel=58
					35, 42, 16, -1, 37, 65, -71, -98, -34,
					-- layer=2 filter=50 channel=59
					-4, 0, 21, -33, 3, 18, -32, -37, -2,
					-- layer=2 filter=50 channel=60
					22, 32, -19, -1, 19, 11, -38, -27, 6,
					-- layer=2 filter=50 channel=61
					-19, -21, -25, 1, 10, -6, 4, -15, 41,
					-- layer=2 filter=50 channel=62
					15, 21, -19, 29, 3, 32, -19, -34, 11,
					-- layer=2 filter=50 channel=63
					-42, -8, -15, -44, 0, -27, -4, 13, -5,
					-- layer=2 filter=50 channel=64
					-20, -1, -20, -8, -30, -34, -13, -34, -58,
					-- layer=2 filter=50 channel=65
					8, 13, 4, 14, 33, 16, 5, 8, 25,
					-- layer=2 filter=50 channel=66
					-10, -62, 9, -40, -16, -39, -20, 3, -34,
					-- layer=2 filter=50 channel=67
					-23, -27, 9, 51, 10, -2, 52, 43, 31,
					-- layer=2 filter=50 channel=68
					-7, 3, 2, 4, 0, -2, -6, 3, 7,
					-- layer=2 filter=50 channel=69
					-6, 40, -11, 2, 3, -18, 3, -3, -52,
					-- layer=2 filter=50 channel=70
					-7, -28, -13, -9, -13, -28, -9, 9, 2,
					-- layer=2 filter=50 channel=71
					-4, 14, 41, -26, -4, 14, -2, -25, 19,
					-- layer=2 filter=50 channel=72
					6, 36, 15, 10, 33, 1, -47, 1, 21,
					-- layer=2 filter=50 channel=73
					-38, 4, 1, 10, -3, -26, -21, -14, 0,
					-- layer=2 filter=50 channel=74
					-33, -17, 4, -15, -4, -17, 13, 9, -4,
					-- layer=2 filter=50 channel=75
					-13, 16, 25, -63, -4, -22, 2, -22, -6,
					-- layer=2 filter=50 channel=76
					-31, 20, -3, -20, -16, 31, -13, -6, 0,
					-- layer=2 filter=50 channel=77
					7, -11, -7, 0, -4, 0, -4, 1, -11,
					-- layer=2 filter=50 channel=78
					-6, 10, 1, -13, -16, -4, 25, -2, 16,
					-- layer=2 filter=50 channel=79
					0, -9, -8, -6, -2, 7, 0, -2, -11,
					-- layer=2 filter=50 channel=80
					-31, -15, 2, 0, -34, -25, 25, 15, -16,
					-- layer=2 filter=50 channel=81
					5, 9, 8, -1, 2, 6, -1, -5, -8,
					-- layer=2 filter=50 channel=82
					-3, 0, 1, 4, 7, -6, -11, 2, -8,
					-- layer=2 filter=50 channel=83
					-2, 2, 40, 7, 50, -3, -14, -13, -12,
					-- layer=2 filter=50 channel=84
					2, 2, -6, -6, -10, -2, 2, -4, -2,
					-- layer=2 filter=50 channel=85
					-9, -4, -16, -13, 7, -15, 2, 11, 1,
					-- layer=2 filter=50 channel=86
					-8, -10, -6, 0, 3, -8, -9, -1, -4,
					-- layer=2 filter=50 channel=87
					3, 22, -33, 5, 4, -27, 7, -7, -12,
					-- layer=2 filter=50 channel=88
					-2, -2, 24, -39, -6, 0, -23, 14, -42,
					-- layer=2 filter=50 channel=89
					37, 28, 16, -25, 18, 56, -69, -90, -8,
					-- layer=2 filter=50 channel=90
					4, 8, -3, 1, -5, 3, -2, 5, -7,
					-- layer=2 filter=50 channel=91
					27, 18, 8, 17, 31, 19, -43, -58, 22,
					-- layer=2 filter=50 channel=92
					22, 38, 10, 6, 34, 26, -52, -94, -35,
					-- layer=2 filter=50 channel=93
					4, 19, 13, 33, 16, -10, -11, 7, -14,
					-- layer=2 filter=50 channel=94
					-31, 0, -1, 30, 35, 20, 12, -39, 37,
					-- layer=2 filter=50 channel=95
					4, 14, 0, 0, 10, 15, 9, 14, 11,
					-- layer=2 filter=50 channel=96
					28, 25, 28, -5, 19, 34, -26, 1, -34,
					-- layer=2 filter=50 channel=97
					-15, 33, 18, 14, -54, -76, 52, 8, -12,
					-- layer=2 filter=50 channel=98
					37, -26, -32, -15, -4, -18, 0, 3, 18,
					-- layer=2 filter=50 channel=99
					-38, 24, 23, -25, 25, 39, 8, -24, 1,
					-- layer=2 filter=50 channel=100
					-26, -12, -2, -22, -9, 1, -3, -30, 4,
					-- layer=2 filter=50 channel=101
					19, 13, 38, -4, -57, -8, 16, -18, -10,
					-- layer=2 filter=50 channel=102
					0, -10, -3, -30, 4, -6, -1, -12, -25,
					-- layer=2 filter=50 channel=103
					21, 24, 15, 59, 45, -43, -49, 12, 86,
					-- layer=2 filter=50 channel=104
					18, 1, -28, -4, 0, -2, -51, -12, 16,
					-- layer=2 filter=50 channel=105
					20, -9, 0, 18, -15, 0, 10, -5, 17,
					-- layer=2 filter=50 channel=106
					27, 19, 14, -35, -77, -9, 14, -43, 3,
					-- layer=2 filter=50 channel=107
					-8, 15, 38, 3, -44, -12, 57, 92, 0,
					-- layer=2 filter=50 channel=108
					-14, 5, 35, -54, -6, 21, -22, -47, -35,
					-- layer=2 filter=50 channel=109
					-4, -7, 8, -3, 5, 2, -6, 4, 3,
					-- layer=2 filter=50 channel=110
					-8, 21, 43, 20, 14, 6, -50, -44, -35,
					-- layer=2 filter=50 channel=111
					-1, 3, 11, 5, -1, -4, 7, -7, 3,
					-- layer=2 filter=50 channel=112
					-4, 1, 13, -18, -23, -12, 25, 13, 29,
					-- layer=2 filter=50 channel=113
					-15, 12, -12, 4, 19, 0, -42, 23, -12,
					-- layer=2 filter=50 channel=114
					14, 0, 2, -5, -5, 7, -2, 3, -11,
					-- layer=2 filter=50 channel=115
					-4, 7, 4, 9, 0, -1, -6, 3, 6,
					-- layer=2 filter=50 channel=116
					-5, 24, -10, 7, 28, 6, -1, 4, 3,
					-- layer=2 filter=50 channel=117
					-6, -2, 16, 4, 44, 0, -5, 41, 46,
					-- layer=2 filter=50 channel=118
					7, -6, -8, 14, -12, 0, 56, 50, 18,
					-- layer=2 filter=50 channel=119
					-17, 2, 34, -13, -29, -22, 42, -27, 23,
					-- layer=2 filter=50 channel=120
					5, 7, 8, 0, 3, 5, -4, 0, 2,
					-- layer=2 filter=50 channel=121
					0, -2, -5, 9, -6, 5, -4, -6, 8,
					-- layer=2 filter=50 channel=122
					1, 3, 14, 3, -3, 10, -4, 10, 5,
					-- layer=2 filter=50 channel=123
					-9, -14, -7, 22, 26, 0, 0, 26, 9,
					-- layer=2 filter=50 channel=124
					9, 15, -20, 2, 58, 45, -22, 34, 20,
					-- layer=2 filter=50 channel=125
					2, 3, 0, 8, -7, -14, 1, 3, -12,
					-- layer=2 filter=50 channel=126
					-46, 3, 26, -36, -3, -4, 43, -11, -32,
					-- layer=2 filter=50 channel=127
					-1, 30, -23, -29, 2, -12, 13, 3, 3,
					-- layer=2 filter=51 channel=0
					1, 2, 14, -2, -3, -7, -24, 5, -21,
					-- layer=2 filter=51 channel=1
					17, 24, 14, 10, 3, 20, 18, 21, -24,
					-- layer=2 filter=51 channel=2
					-2, 9, 6, 0, -9, -6, -1, -9, 10,
					-- layer=2 filter=51 channel=3
					26, 6, -14, 4, 3, -10, 8, -18, -1,
					-- layer=2 filter=51 channel=4
					-33, 16, -23, -59, 1, -9, -19, -46, -24,
					-- layer=2 filter=51 channel=5
					12, 16, -9, 4, -7, 11, 14, 19, 19,
					-- layer=2 filter=51 channel=6
					-2, 0, 1, 9, 19, 2, -11, 3, 11,
					-- layer=2 filter=51 channel=7
					-19, 9, -36, 5, -20, -1, 25, 4, 24,
					-- layer=2 filter=51 channel=8
					-5, 1, -1, 10, -13, 8, 5, 4, -3,
					-- layer=2 filter=51 channel=9
					32, -5, 24, -4, 8, 44, -39, -39, 0,
					-- layer=2 filter=51 channel=10
					30, 3, 15, -3, 13, 23, -1, -12, -19,
					-- layer=2 filter=51 channel=11
					-2, 11, -5, 8, 1, 6, 9, 19, 22,
					-- layer=2 filter=51 channel=12
					6, 21, 9, 14, 11, 16, 31, 14, 34,
					-- layer=2 filter=51 channel=13
					-5, 5, 2, 2, 1, 1, -1, -8, -8,
					-- layer=2 filter=51 channel=14
					4, 15, 20, 24, 9, 38, 17, 27, 10,
					-- layer=2 filter=51 channel=15
					-4, -19, -2, -9, -5, 17, -12, 1, 2,
					-- layer=2 filter=51 channel=16
					16, 24, 96, 58, -85, -5, 9, -27, -29,
					-- layer=2 filter=51 channel=17
					-3, -8, -3, 6, -3, 2, 3, 7, 3,
					-- layer=2 filter=51 channel=18
					-21, 25, -28, -21, -19, -7, -37, 11, 28,
					-- layer=2 filter=51 channel=19
					30, -29, 19, 7, 21, 0, 16, -12, 1,
					-- layer=2 filter=51 channel=20
					1, -9, 3, 8, 7, 10, 0, 9, -6,
					-- layer=2 filter=51 channel=21
					17, 16, 17, 13, -4, 13, 14, -9, 5,
					-- layer=2 filter=51 channel=22
					0, -2, -4, 6, 8, 0, 4, 7, 0,
					-- layer=2 filter=51 channel=23
					-5, -7, 23, -43, -48, -9, -4, -59, -12,
					-- layer=2 filter=51 channel=24
					-7, 16, 24, -3, 0, 0, -18, -6, 10,
					-- layer=2 filter=51 channel=25
					27, 35, 20, -12, 2, 2, -5, 2, 17,
					-- layer=2 filter=51 channel=26
					2, 5, 13, -6, 0, -6, 6, -6, 7,
					-- layer=2 filter=51 channel=27
					0, 6, 15, 15, 9, 29, 34, -11, -3,
					-- layer=2 filter=51 channel=28
					-4, 0, 14, -19, -76, 1, 2, -15, 0,
					-- layer=2 filter=51 channel=29
					-2, -7, 0, -11, 0, -11, 1, 6, 1,
					-- layer=2 filter=51 channel=30
					-40, -16, 16, -16, -19, 15, -24, -51, -60,
					-- layer=2 filter=51 channel=31
					-38, -35, 34, -32, -24, -63, -41, -39, -49,
					-- layer=2 filter=51 channel=32
					0, 0, 2, -5, -1, -7, 7, 1, -4,
					-- layer=2 filter=51 channel=33
					-3, -30, -25, -14, -15, 33, 25, -38, -30,
					-- layer=2 filter=51 channel=34
					-12, -31, -14, -1, -45, -11, -30, -16, 0,
					-- layer=2 filter=51 channel=35
					10, 5, -1, 5, -67, -34, -45, -77, -21,
					-- layer=2 filter=51 channel=36
					-2, -4, 2, -5, 0, 5, 0, 0, 14,
					-- layer=2 filter=51 channel=37
					7, 6, 8, 0, 16, 10, 12, 27, 17,
					-- layer=2 filter=51 channel=38
					-10, -6, 0, -9, -21, -2, 11, -18, -6,
					-- layer=2 filter=51 channel=39
					-18, -66, 21, -68, -98, -83, 26, -30, -34,
					-- layer=2 filter=51 channel=40
					-7, -70, -40, -39, 0, 14, -68, 4, 30,
					-- layer=2 filter=51 channel=41
					3, -8, -1, 6, 8, 10, 1, -9, -2,
					-- layer=2 filter=51 channel=42
					22, 29, 33, 7, -24, -5, -12, -20, -62,
					-- layer=2 filter=51 channel=43
					-8, -12, -19, -40, 2, -26, -43, -28, 21,
					-- layer=2 filter=51 channel=44
					-9, 9, 2, 2, -9, 7, -7, 10, 6,
					-- layer=2 filter=51 channel=45
					26, 0, 33, -20, -2, -7, -42, -103, -74,
					-- layer=2 filter=51 channel=46
					-9, -59, 1, -36, -20, -6, -25, -47, -27,
					-- layer=2 filter=51 channel=47
					-28, -72, -2, -40, -48, -12, -13, -24, -10,
					-- layer=2 filter=51 channel=48
					0, 3, -5, -4, 0, -6, -8, -5, 0,
					-- layer=2 filter=51 channel=49
					58, 63, 20, 22, 13, 44, 6, 29, -2,
					-- layer=2 filter=51 channel=50
					-6, -10, -5, 4, -2, -13, -14, -17, -14,
					-- layer=2 filter=51 channel=51
					-6, 22, 5, -13, 17, 7, 3, 11, 12,
					-- layer=2 filter=51 channel=52
					-46, -9, 14, 17, 25, 17, 17, 10, 22,
					-- layer=2 filter=51 channel=53
					14, -24, 3, 31, -4, 20, 28, -30, -27,
					-- layer=2 filter=51 channel=54
					35, -6, -4, 24, -3, 10, 24, 13, 3,
					-- layer=2 filter=51 channel=55
					-1, 12, -8, 9, 12, -6, -4, -3, 5,
					-- layer=2 filter=51 channel=56
					-3, -10, 1, 6, 3, 10, 0, 21, 22,
					-- layer=2 filter=51 channel=57
					7, 0, 6, 8, 10, 15, 3, -9, -3,
					-- layer=2 filter=51 channel=58
					10, 20, -9, 31, 18, -4, 38, -5, 23,
					-- layer=2 filter=51 channel=59
					-26, -18, -17, -8, -2, 0, 0, 11, 19,
					-- layer=2 filter=51 channel=60
					11, 1, 22, 9, 3, 6, 7, 44, 24,
					-- layer=2 filter=51 channel=61
					11, 18, -22, 20, 2, -17, -33, -8, -16,
					-- layer=2 filter=51 channel=62
					-2, 3, -7, 21, 9, -3, -18, 1, 27,
					-- layer=2 filter=51 channel=63
					0, -7, -7, -9, -18, -28, -18, 6, -30,
					-- layer=2 filter=51 channel=64
					-1, 1, 51, -9, -32, -24, 14, -26, -13,
					-- layer=2 filter=51 channel=65
					-4, 10, 14, 7, 9, -33, 8, 10, -15,
					-- layer=2 filter=51 channel=66
					22, -40, 7, -36, -43, -31, 37, -3, -25,
					-- layer=2 filter=51 channel=67
					-25, -53, -9, -69, -32, -23, -38, -27, -11,
					-- layer=2 filter=51 channel=68
					5, -5, 12, -9, -1, 5, -1, 6, 0,
					-- layer=2 filter=51 channel=69
					14, 14, 35, -13, -20, -3, -6, -17, -22,
					-- layer=2 filter=51 channel=70
					26, 8, 27, 14, -34, 14, 24, 6, 0,
					-- layer=2 filter=51 channel=71
					-12, -8, -35, -8, -22, -3, -13, -32, -10,
					-- layer=2 filter=51 channel=72
					30, -13, 2, 25, 8, 39, 38, -16, 19,
					-- layer=2 filter=51 channel=73
					16, 0, 35, 25, -18, -16, 5, -50, -24,
					-- layer=2 filter=51 channel=74
					-6, -21, 11, -35, -17, -72, -38, -46, -35,
					-- layer=2 filter=51 channel=75
					-16, -4, -10, 13, -39, -27, -9, 12, 62,
					-- layer=2 filter=51 channel=76
					-29, -23, -2, -9, -41, 32, -9, -3, -36,
					-- layer=2 filter=51 channel=77
					5, -4, 9, -7, 5, 4, -2, -1, -3,
					-- layer=2 filter=51 channel=78
					20, 3, 0, 3, 2, -19, -25, 21, 31,
					-- layer=2 filter=51 channel=79
					5, 5, -10, 10, 2, -11, -4, 9, -2,
					-- layer=2 filter=51 channel=80
					-8, 22, 38, -31, 0, -56, -44, -26, -36,
					-- layer=2 filter=51 channel=81
					-6, 3, -5, 0, 2, -1, 8, -10, -5,
					-- layer=2 filter=51 channel=82
					-3, 2, -2, 1, -10, 4, 5, -1, 4,
					-- layer=2 filter=51 channel=83
					19, 40, 19, 18, -5, -3, -2, -14, -39,
					-- layer=2 filter=51 channel=84
					3, 1, -9, 8, 4, 1, -6, 3, 8,
					-- layer=2 filter=51 channel=85
					9, 12, 12, 17, 10, -4, -1, 25, 1,
					-- layer=2 filter=51 channel=86
					0, 0, 18, -12, -13, 0, -9, -9, 6,
					-- layer=2 filter=51 channel=87
					-33, -1, -2, -47, -29, -2, -33, -27, 46,
					-- layer=2 filter=51 channel=88
					-27, 1, 6, 0, 2, -7, -17, -99, -22,
					-- layer=2 filter=51 channel=89
					15, -6, -9, -11, 23, 17, 13, 21, 30,
					-- layer=2 filter=51 channel=90
					3, 0, 5, 9, 5, -3, -6, 0, -6,
					-- layer=2 filter=51 channel=91
					-32, -24, -7, 16, -9, -17, 9, -10, 16,
					-- layer=2 filter=51 channel=92
					29, 36, 3, 11, 22, 28, 33, 16, -6,
					-- layer=2 filter=51 channel=93
					-23, -22, 9, -22, 8, -47, -13, -32, 3,
					-- layer=2 filter=51 channel=94
					19, 8, -12, 31, 43, -7, -21, 32, -25,
					-- layer=2 filter=51 channel=95
					-6, -12, 0, -12, -9, 1, -5, -9, -7,
					-- layer=2 filter=51 channel=96
					44, 16, 28, 3, 29, 22, -46, 14, 14,
					-- layer=2 filter=51 channel=97
					13, 2, 42, -6, -10, -1, -17, 2, -3,
					-- layer=2 filter=51 channel=98
					20, -2, 37, 21, -18, 28, -1, -7, 34,
					-- layer=2 filter=51 channel=99
					-31, -13, -9, 6, 43, 3, 9, 14, 6,
					-- layer=2 filter=51 channel=100
					0, 5, 5, 11, -42, -3, -13, 10, -39,
					-- layer=2 filter=51 channel=101
					-24, 3, -13, -17, -44, -35, -16, -23, 9,
					-- layer=2 filter=51 channel=102
					-7, -3, 10, -43, -14, 4, -50, -16, -14,
					-- layer=2 filter=51 channel=103
					-69, -10, 1, -6, -2, -26, -41, 12, 2,
					-- layer=2 filter=51 channel=104
					17, 24, -7, 31, -3, 48, -5, 21, 0,
					-- layer=2 filter=51 channel=105
					17, -24, 4, -23, 37, 31, 2, -9, 10,
					-- layer=2 filter=51 channel=106
					18, 21, 14, -20, -15, -16, -20, -25, 7,
					-- layer=2 filter=51 channel=107
					-6, 24, 10, 21, 13, -16, 2, 7, -1,
					-- layer=2 filter=51 channel=108
					10, 1, 30, -16, -5, 20, 21, 0, -13,
					-- layer=2 filter=51 channel=109
					7, -5, -8, 3, 7, -8, 0, 4, 5,
					-- layer=2 filter=51 channel=110
					-5, -1, 38, 1, -9, 8, -18, -12, 9,
					-- layer=2 filter=51 channel=111
					-5, -8, 3, -8, 1, -2, -3, -11, -8,
					-- layer=2 filter=51 channel=112
					11, 1, -1, -6, -3, -17, -18, 11, 3,
					-- layer=2 filter=51 channel=113
					0, 14, 18, 0, -22, -8, 18, -30, -52,
					-- layer=2 filter=51 channel=114
					6, -4, -10, -7, -8, -13, 12, 5, -4,
					-- layer=2 filter=51 channel=115
					8, -12, 6, -9, 7, -8, 8, 4, 9,
					-- layer=2 filter=51 channel=116
					-4, 6, -17, -45, -42, -21, 3, -14, 15,
					-- layer=2 filter=51 channel=117
					26, 0, -12, -6, -26, 17, 13, -6, 1,
					-- layer=2 filter=51 channel=118
					12, 2, 6, 22, 18, 3, -9, -5, 29,
					-- layer=2 filter=51 channel=119
					-10, 9, 13, -14, -83, -11, -39, -48, -25,
					-- layer=2 filter=51 channel=120
					3, 6, -1, 8, 6, -9, -1, 7, -3,
					-- layer=2 filter=51 channel=121
					7, -1, -3, -1, 10, -4, -10, -4, 1,
					-- layer=2 filter=51 channel=122
					13, 15, -1, -7, -5, 4, 16, 4, 8,
					-- layer=2 filter=51 channel=123
					-23, -25, -12, -31, -35, 1, 44, -21, 16,
					-- layer=2 filter=51 channel=124
					-11, -27, -23, -17, -25, 0, 16, 15, -26,
					-- layer=2 filter=51 channel=125
					2, -6, 3, 6, -8, 4, 2, -5, -10,
					-- layer=2 filter=51 channel=126
					32, -31, -71, -46, -4, -130, -32, 0, -35,
					-- layer=2 filter=51 channel=127
					-4, -2, 18, 0, 27, -6, -18, 0, -39,
					-- layer=2 filter=52 channel=0
					1, -18, 16, -7, -6, -8, 11, 34, 39,
					-- layer=2 filter=52 channel=1
					16, 12, 8, 20, -9, 11, -1, -41, -12,
					-- layer=2 filter=52 channel=2
					-6, -5, 0, 9, 6, 3, 10, 9, 7,
					-- layer=2 filter=52 channel=3
					-30, -24, -28, 13, -20, -11, 29, 11, 30,
					-- layer=2 filter=52 channel=4
					-2, -17, 7, 1, -37, 16, -4, 12, -7,
					-- layer=2 filter=52 channel=5
					2, 14, -16, -26, 6, -7, -15, 30, 31,
					-- layer=2 filter=52 channel=6
					2, -19, 14, 14, 1, 25, -15, -4, 9,
					-- layer=2 filter=52 channel=7
					-7, -35, 18, 16, 3, 44, 20, 12, 21,
					-- layer=2 filter=52 channel=8
					6, -1, -10, 0, -4, 9, 3, 9, -2,
					-- layer=2 filter=52 channel=9
					-4, -30, -8, 22, -13, -4, -36, -7, 0,
					-- layer=2 filter=52 channel=10
					-20, -14, -3, 1, -12, -13, 21, 48, 38,
					-- layer=2 filter=52 channel=11
					6, -5, 3, 4, -2, 15, 6, 18, 21,
					-- layer=2 filter=52 channel=12
					-19, -20, 6, 32, 3, 29, 5, -4, 0,
					-- layer=2 filter=52 channel=13
					9, -1, -8, -6, -3, -10, -8, -7, -7,
					-- layer=2 filter=52 channel=14
					-5, -20, 5, 42, -4, 12, -20, -31, -2,
					-- layer=2 filter=52 channel=15
					10, -48, 36, -45, -29, -8, 6, -18, 7,
					-- layer=2 filter=52 channel=16
					37, 36, 44, -40, -13, 23, -54, -29, -36,
					-- layer=2 filter=52 channel=17
					0, -2, 5, -10, 0, -5, -5, 4, 10,
					-- layer=2 filter=52 channel=18
					3, -24, 20, -11, -24, 3, -22, -14, -27,
					-- layer=2 filter=52 channel=19
					24, 23, 24, 22, 16, 48, 3, -18, 22,
					-- layer=2 filter=52 channel=20
					-10, -8, 6, -1, -7, 0, 5, 0, 6,
					-- layer=2 filter=52 channel=21
					-6, -1, -4, -13, 9, 1, 9, -14, 6,
					-- layer=2 filter=52 channel=22
					-1, 8, 1, -6, -4, -8, -8, 0, 2,
					-- layer=2 filter=52 channel=23
					-2, 0, -1, -16, -6, -9, -5, -22, -5,
					-- layer=2 filter=52 channel=24
					-9, -25, -69, 15, -33, -53, 40, 15, -14,
					-- layer=2 filter=52 channel=25
					14, -5, -40, 31, -16, -45, 38, 25, -5,
					-- layer=2 filter=52 channel=26
					3, 6, -6, -10, -9, -8, 6, -1, 10,
					-- layer=2 filter=52 channel=27
					8, 0, 2, -31, -14, -15, -81, -31, -15,
					-- layer=2 filter=52 channel=28
					16, -53, -23, -30, -22, -22, 31, 19, 36,
					-- layer=2 filter=52 channel=29
					-2, 0, 10, -5, -5, -8, 9, 0, 5,
					-- layer=2 filter=52 channel=30
					-31, -14, -1, -22, -42, -33, -36, -32, -50,
					-- layer=2 filter=52 channel=31
					-20, -43, -15, -21, 16, 0, 47, 15, 37,
					-- layer=2 filter=52 channel=32
					-4, 0, 5, -1, -9, -8, -2, 5, 7,
					-- layer=2 filter=52 channel=33
					-6, -15, 0, 20, 0, 18, -14, -12, 24,
					-- layer=2 filter=52 channel=34
					56, 29, -5, 7, 10, 20, -50, -13, 0,
					-- layer=2 filter=52 channel=35
					35, -3, 0, -26, -3, -6, 11, 4, -3,
					-- layer=2 filter=52 channel=36
					-10, 13, 11, -13, 0, -10, 6, 19, 9,
					-- layer=2 filter=52 channel=37
					2, -1, -9, 3, 6, -9, -15, -8, 22,
					-- layer=2 filter=52 channel=38
					6, 13, -4, -29, -22, -20, -52, -45, -10,
					-- layer=2 filter=52 channel=39
					19, 19, -2, -45, -72, -7, -45, -15, -60,
					-- layer=2 filter=52 channel=40
					-18, -25, 42, -37, 21, -39, -16, -12, 0,
					-- layer=2 filter=52 channel=41
					-11, 3, -1, -3, -6, 4, -5, -9, 3,
					-- layer=2 filter=52 channel=42
					-5, 13, 5, -11, -15, -34, -34, -11, -46,
					-- layer=2 filter=52 channel=43
					15, -11, -41, -53, -28, -29, -8, 28, 10,
					-- layer=2 filter=52 channel=44
					-8, 5, -9, 6, -10, -10, -6, 7, 7,
					-- layer=2 filter=52 channel=45
					2, -58, -44, -40, -68, 10, -59, -53, -55,
					-- layer=2 filter=52 channel=46
					-40, -17, 18, -27, -40, -28, -20, -10, 0,
					-- layer=2 filter=52 channel=47
					-60, -41, -9, -34, -14, -13, 1, 11, 48,
					-- layer=2 filter=52 channel=48
					4, 6, -8, -1, 9, 8, -5, 1, -8,
					-- layer=2 filter=52 channel=49
					9, -18, 14, -5, -8, 8, -14, -24, -50,
					-- layer=2 filter=52 channel=50
					-25, 4, -2, -7, -9, 7, 0, 9, 1,
					-- layer=2 filter=52 channel=51
					7, -11, -5, 20, 0, 7, 21, 15, 15,
					-- layer=2 filter=52 channel=52
					-33, 5, 12, 12, -4, 11, 30, -17, -4,
					-- layer=2 filter=52 channel=53
					-43, 26, 22, 11, -45, 45, -9, 58, 21,
					-- layer=2 filter=52 channel=54
					-24, -13, -26, 10, 3, 25, 24, 26, 46,
					-- layer=2 filter=52 channel=55
					5, -2, -2, 13, -12, 3, 8, 7, 3,
					-- layer=2 filter=52 channel=56
					15, -22, 4, 5, 2, 13, 3, 5, 25,
					-- layer=2 filter=52 channel=57
					-6, -9, -1, 0, 11, 0, -3, 0, -9,
					-- layer=2 filter=52 channel=58
					-23, 0, -6, 9, -9, 8, -14, -14, -8,
					-- layer=2 filter=52 channel=59
					15, 39, -8, -8, 21, 22, -49, -7, -36,
					-- layer=2 filter=52 channel=60
					15, 45, 13, 0, 5, 30, 1, -29, -46,
					-- layer=2 filter=52 channel=61
					7, -25, 18, 6, -27, -38, 26, -32, -28,
					-- layer=2 filter=52 channel=62
					19, -20, -19, -2, 21, 0, -17, 16, -7,
					-- layer=2 filter=52 channel=63
					-30, 2, -4, -34, -43, 5, -34, 2, -7,
					-- layer=2 filter=52 channel=64
					1, 21, -1, -26, -31, -18, -12, -12, -23,
					-- layer=2 filter=52 channel=65
					-4, -27, -12, 1, -13, -23, 22, -21, -16,
					-- layer=2 filter=52 channel=66
					29, -38, -13, -52, -40, -31, -41, 50, -39,
					-- layer=2 filter=52 channel=67
					-10, 11, -3, -46, -21, -21, -36, -18, -3,
					-- layer=2 filter=52 channel=68
					-1, -9, 2, -5, -4, 3, 0, -4, -4,
					-- layer=2 filter=52 channel=69
					38, 50, 19, -12, -4, -10, -44, -14, -44,
					-- layer=2 filter=52 channel=70
					5, -25, 15, -23, -8, 7, -2, 19, 18,
					-- layer=2 filter=52 channel=71
					3, 6, -12, -23, 17, -32, -26, -14, -20,
					-- layer=2 filter=52 channel=72
					-24, -19, 39, 26, 3, 6, -30, 10, 2,
					-- layer=2 filter=52 channel=73
					-43, -22, -9, -20, 0, -1, -40, 6, -31,
					-- layer=2 filter=52 channel=74
					-26, -7, 0, -67, -26, -48, -34, -28, 1,
					-- layer=2 filter=52 channel=75
					18, -48, 12, -1, -10, -4, 49, 10, -16,
					-- layer=2 filter=52 channel=76
					23, 9, -2, 66, -18, 23, 10, 36, 1,
					-- layer=2 filter=52 channel=77
					-10, 1, 6, 7, -3, -5, 0, 7, 1,
					-- layer=2 filter=52 channel=78
					11, -11, -6, -3, 15, -6, 39, 31, 11,
					-- layer=2 filter=52 channel=79
					0, 0, 11, -5, 0, 0, -11, -10, -3,
					-- layer=2 filter=52 channel=80
					-18, 26, 28, -58, 5, -8, -4, 10, 7,
					-- layer=2 filter=52 channel=81
					-9, -2, -1, -12, 6, 3, 9, -9, 1,
					-- layer=2 filter=52 channel=82
					-7, 0, -6, -2, -2, -7, -2, -1, -4,
					-- layer=2 filter=52 channel=83
					45, 5, -9, -15, -64, -18, 5, -38, -7,
					-- layer=2 filter=52 channel=84
					5, -4, -8, 3, 5, 7, -7, -2, -7,
					-- layer=2 filter=52 channel=85
					-4, 14, 5, 6, -7, -2, -16, 9, 14,
					-- layer=2 filter=52 channel=86
					5, 3, -2, -15, 1, -11, 4, -6, -2,
					-- layer=2 filter=52 channel=87
					65, 4, 16, -1, 26, -13, -28, -48, -42,
					-- layer=2 filter=52 channel=88
					12, 0, -1, -23, -12, -6, -66, -54, -64,
					-- layer=2 filter=52 channel=89
					17, 4, 17, 31, 12, -3, -28, -12, -14,
					-- layer=2 filter=52 channel=90
					-5, 1, -9, -10, 7, -2, -3, 8, -7,
					-- layer=2 filter=52 channel=91
					-18, 13, -3, 29, 0, 10, 3, 30, -9,
					-- layer=2 filter=52 channel=92
					-11, 11, -4, 48, -7, 17, -25, 1, -23,
					-- layer=2 filter=52 channel=93
					-17, -16, -39, -31, 8, -11, -13, 20, 4,
					-- layer=2 filter=52 channel=94
					-15, -4, 20, 45, 18, 22, 3, -12, -5,
					-- layer=2 filter=52 channel=95
					-8, 8, -17, -1, 10, 14, -13, 0, -12,
					-- layer=2 filter=52 channel=96
					26, 34, 53, 27, 30, 7, 13, 7, 19,
					-- layer=2 filter=52 channel=97
					0, 12, 7, -37, -20, -40, 18, -13, 22,
					-- layer=2 filter=52 channel=98
					8, -43, 4, -17, 11, 8, 6, 6, 37,
					-- layer=2 filter=52 channel=99
					-17, 26, 17, 20, 28, 42, 26, -11, 13,
					-- layer=2 filter=52 channel=100
					-8, 23, -34, -50, -35, -47, -16, -15, -21,
					-- layer=2 filter=52 channel=101
					-25, -17, 4, 17, 14, -13, 42, 15, -20,
					-- layer=2 filter=52 channel=102
					-4, -21, 15, 6, -18, -37, 36, -23, -23,
					-- layer=2 filter=52 channel=103
					-15, 0, 20, 28, 27, -30, 37, 21, 21,
					-- layer=2 filter=52 channel=104
					10, -20, 19, -17, 12, 29, 6, -4, -12,
					-- layer=2 filter=52 channel=105
					53, 18, -21, -8, 7, 3, 12, -7, 0,
					-- layer=2 filter=52 channel=106
					10, -11, -38, 20, -28, -23, 32, 25, 7,
					-- layer=2 filter=52 channel=107
					9, 16, 15, 4, -6, -17, 29, 50, 2,
					-- layer=2 filter=52 channel=108
					5, -32, 14, 42, -48, 6, -9, -62, -10,
					-- layer=2 filter=52 channel=109
					-7, 18, 5, -1, 6, 12, 2, -1, 0,
					-- layer=2 filter=52 channel=110
					-1, -8, -9, 24, -28, -23, 2, -27, -63,
					-- layer=2 filter=52 channel=111
					6, 9, -7, 8, -8, 2, -3, 9, 9,
					-- layer=2 filter=52 channel=112
					5, 3, 15, 12, -16, -15, 13, 8, 14,
					-- layer=2 filter=52 channel=113
					-3, -18, -13, -29, -37, 30, -1, -1, -54,
					-- layer=2 filter=52 channel=114
					-3, -13, 8, -2, 9, 6, 8, -4, -4,
					-- layer=2 filter=52 channel=115
					10, 5, 0, 3, 4, 0, 3, 4, 7,
					-- layer=2 filter=52 channel=116
					46, 19, 11, -8, 0, 0, -18, -35, -14,
					-- layer=2 filter=52 channel=117
					-39, -35, 60, 36, 26, 24, -2, 12, 25,
					-- layer=2 filter=52 channel=118
					6, 4, 10, -13, 10, 19, 16, 23, 18,
					-- layer=2 filter=52 channel=119
					64, 9, -3, 16, -41, -22, -3, 11, -19,
					-- layer=2 filter=52 channel=120
					4, -3, 3, 10, 0, 0, -2, 9, 0,
					-- layer=2 filter=52 channel=121
					-2, 9, 2, 0, 7, -10, -1, 0, -3,
					-- layer=2 filter=52 channel=122
					2, 0, 6, -6, 11, 10, -5, 2, 3,
					-- layer=2 filter=52 channel=123
					-22, -5, 55, 20, 18, 32, -11, 1, 42,
					-- layer=2 filter=52 channel=124
					19, -6, 10, 16, 4, -10, 2, 24, -4,
					-- layer=2 filter=52 channel=125
					-5, 9, -6, 1, -6, 7, 0, -1, -5,
					-- layer=2 filter=52 channel=126
					20, 40, 25, 18, 29, -105, -3, 40, -42,
					-- layer=2 filter=52 channel=127
					24, 1, -4, -26, -8, -13, -41, -47, -3,
					-- layer=2 filter=53 channel=0
					6, 4, 23, 12, 12, -1, -4, -16, -19,
					-- layer=2 filter=53 channel=1
					-8, -25, 14, 9, 22, 20, 11, 4, -33,
					-- layer=2 filter=53 channel=2
					4, 2, -5, 4, -1, 5, 6, 3, -3,
					-- layer=2 filter=53 channel=3
					-21, 6, 14, -39, -10, -9, 6, 13, 9,
					-- layer=2 filter=53 channel=4
					8, 31, 23, 10, 10, 26, -11, -16, 15,
					-- layer=2 filter=53 channel=5
					29, 1, -3, 0, -16, -6, -1, -32, -42,
					-- layer=2 filter=53 channel=6
					-22, 14, 4, 16, -14, -13, 7, -4, -11,
					-- layer=2 filter=53 channel=7
					17, 19, 8, -3, 58, 52, 4, 56, 54,
					-- layer=2 filter=53 channel=8
					-7, 5, 1, 8, -7, -3, 5, 1, 11,
					-- layer=2 filter=53 channel=9
					-12, 30, 6, -39, -16, -23, -20, -12, -34,
					-- layer=2 filter=53 channel=10
					-6, 6, 10, -10, -4, -16, -12, -15, -2,
					-- layer=2 filter=53 channel=11
					7, 4, -1, -7, -11, -12, -19, -15, -22,
					-- layer=2 filter=53 channel=12
					31, 24, 21, -2, 38, 33, 23, 29, 12,
					-- layer=2 filter=53 channel=13
					-2, -4, 7, 6, -6, -2, 3, -6, 0,
					-- layer=2 filter=53 channel=14
					-8, 21, -1, -13, 1, 40, 2, 35, 0,
					-- layer=2 filter=53 channel=15
					8, -50, -38, -98, -40, 9, -121, -41, -1,
					-- layer=2 filter=53 channel=16
					-4, 23, 10, -23, 0, 16, -37, -27, -7,
					-- layer=2 filter=53 channel=17
					7, 10, 2, -7, -8, -4, -2, -7, 3,
					-- layer=2 filter=53 channel=18
					-16, -7, 16, -21, -64, -36, -11, -21, -6,
					-- layer=2 filter=53 channel=19
					-23, -22, -20, 15, 43, 9, 33, 5, 2,
					-- layer=2 filter=53 channel=20
					0, 2, 5, 8, -10, -7, 1, 0, -4,
					-- layer=2 filter=53 channel=21
					-14, -30, -17, -19, -9, 5, -9, 2, 4,
					-- layer=2 filter=53 channel=22
					6, 15, 0, 2, -8, 8, 11, 0, -8,
					-- layer=2 filter=53 channel=23
					-10, 26, 20, 1, 25, 34, 11, 10, 14,
					-- layer=2 filter=53 channel=24
					-11, -7, -3, -22, 27, -23, -5, 23, -4,
					-- layer=2 filter=53 channel=25
					-27, -11, -11, 0, 18, -1, -17, 16, 20,
					-- layer=2 filter=53 channel=26
					-8, -2, -3, -4, 5, -2, 7, 9, 0,
					-- layer=2 filter=53 channel=27
					-3, 13, -11, -11, 17, 23, -8, 8, -1,
					-- layer=2 filter=53 channel=28
					-44, 0, 7, 7, -22, 8, 0, 27, 23,
					-- layer=2 filter=53 channel=29
					-5, 6, 0, 0, 0, 2, 6, 6, -7,
					-- layer=2 filter=53 channel=30
					6, 31, 8, -12, 5, 7, 13, 29, 6,
					-- layer=2 filter=53 channel=31
					-52, -4, -38, -106, -18, -48, -67, -31, -76,
					-- layer=2 filter=53 channel=32
					4, 7, 6, -3, -3, -4, 0, -7, -5,
					-- layer=2 filter=53 channel=33
					-7, -5, 12, -57, -20, 24, -43, 4, 33,
					-- layer=2 filter=53 channel=34
					33, -18, 16, -36, -61, -74, -5, -16, -46,
					-- layer=2 filter=53 channel=35
					-21, -22, 8, -3, -17, -11, -47, 32, 27,
					-- layer=2 filter=53 channel=36
					1, 0, -6, 7, 3, 7, -2, 3, 5,
					-- layer=2 filter=53 channel=37
					9, -2, 0, -12, -12, -11, 3, -14, -18,
					-- layer=2 filter=53 channel=38
					0, -4, 4, 4, -5, 7, 4, -16, -10,
					-- layer=2 filter=53 channel=39
					-17, -24, 10, -62, 0, 9, -32, 17, -6,
					-- layer=2 filter=53 channel=40
					-13, -41, 10, -24, -35, -31, -62, -19, 35,
					-- layer=2 filter=53 channel=41
					0, -1, -1, -7, 1, -11, -6, 1, -3,
					-- layer=2 filter=53 channel=42
					-23, 23, 31, 2, 24, 16, -35, 8, 22,
					-- layer=2 filter=53 channel=43
					-7, -26, 2, -36, 9, -24, -5, 28, 17,
					-- layer=2 filter=53 channel=44
					11, -5, 4, -3, 6, 1, 3, -5, -6,
					-- layer=2 filter=53 channel=45
					-30, 3, -5, -38, 15, 29, -41, -2, 17,
					-- layer=2 filter=53 channel=46
					7, 0, 16, 22, 26, 0, -12, -6, -7,
					-- layer=2 filter=53 channel=47
					7, 41, 21, -12, 8, 23, -18, 0, 9,
					-- layer=2 filter=53 channel=48
					4, 2, -4, 7, 2, 7, 11, -9, -3,
					-- layer=2 filter=53 channel=49
					22, 13, -35, 3, -42, -7, 18, -21, -10,
					-- layer=2 filter=53 channel=50
					11, -3, 10, 7, 18, 15, -14, 14, 25,
					-- layer=2 filter=53 channel=51
					-1, 9, 7, -6, -3, -6, -5, -33, -19,
					-- layer=2 filter=53 channel=52
					3, 16, 32, 1, -19, -5, 31, 5, -14,
					-- layer=2 filter=53 channel=53
					-32, -46, -74, -24, -42, -75, 10, -40, -21,
					-- layer=2 filter=53 channel=54
					7, -14, 35, -13, 22, -14, -22, -11, -6,
					-- layer=2 filter=53 channel=55
					8, 6, -6, -2, 6, -1, -5, -10, -4,
					-- layer=2 filter=53 channel=56
					4, 15, 4, -16, 1, 0, -14, -25, -21,
					-- layer=2 filter=53 channel=57
					-2, -2, -1, 2, 0, -4, 1, 1, -6,
					-- layer=2 filter=53 channel=58
					5, 8, 1, -5, 17, 33, 0, 32, 21,
					-- layer=2 filter=53 channel=59
					0, -37, -14, 15, -7, -10, 34, -28, -31,
					-- layer=2 filter=53 channel=60
					-1, -28, 0, 26, -2, -40, 28, 0, -3,
					-- layer=2 filter=53 channel=61
					-24, -45, -6, 31, -20, -84, 21, 10, 25,
					-- layer=2 filter=53 channel=62
					26, 16, 27, 21, -3, -24, 28, -10, -16,
					-- layer=2 filter=53 channel=63
					12, -8, 12, 7, 20, 2, 1, 16, 15,
					-- layer=2 filter=53 channel=64
					-15, 10, 11, 5, 13, 13, 17, -12, 0,
					-- layer=2 filter=53 channel=65
					17, -12, -3, 33, -32, -67, 7, -9, 12,
					-- layer=2 filter=53 channel=66
					38, 94, 8, 3, 16, 57, 34, 10, 9,
					-- layer=2 filter=53 channel=67
					10, 7, -2, -19, -15, -33, 7, -17, -36,
					-- layer=2 filter=53 channel=68
					0, -4, -10, 0, -9, -11, 6, -9, 0,
					-- layer=2 filter=53 channel=69
					-3, 11, 9, -2, 1, 3, -8, -2, -12,
					-- layer=2 filter=53 channel=70
					-22, 7, 1, -2, -23, 16, -51, 6, 2,
					-- layer=2 filter=53 channel=71
					-20, 3, -20, 4, 29, 11, 1, 22, 19,
					-- layer=2 filter=53 channel=72
					4, -9, 5, -42, -15, 27, 9, 34, 30,
					-- layer=2 filter=53 channel=73
					4, -26, -54, 49, -13, -13, 9, 4, 5,
					-- layer=2 filter=53 channel=74
					3, -16, 3, -2, 10, 1, -5, 34, -6,
					-- layer=2 filter=53 channel=75
					-18, 22, 23, -28, 9, 9, 13, 59, 34,
					-- layer=2 filter=53 channel=76
					-54, 26, -63, -48, -68, -79, -36, -40, -24,
					-- layer=2 filter=53 channel=77
					2, 1, -3, 0, -10, 0, -6, -1, -6,
					-- layer=2 filter=53 channel=78
					-1, -37, -21, 2, -28, -42, -30, -14, -6,
					-- layer=2 filter=53 channel=79
					-7, -8, 2, -10, 4, -1, -1, 4, 0,
					-- layer=2 filter=53 channel=80
					-18, 5, 7, -15, 9, -11, 10, 3, 18,
					-- layer=2 filter=53 channel=81
					3, 2, 8, -3, -2, 7, 13, 3, -2,
					-- layer=2 filter=53 channel=82
					7, 7, 2, 2, -5, 4, 0, -2, 8,
					-- layer=2 filter=53 channel=83
					-31, -1, 8, 10, 15, 15, -8, 2, 0,
					-- layer=2 filter=53 channel=84
					6, -5, -10, 1, -10, -10, -10, 8, 0,
					-- layer=2 filter=53 channel=85
					3, 1, 18, 1, 11, 12, 12, -9, 12,
					-- layer=2 filter=53 channel=86
					-2, -5, 5, -21, -14, 9, -10, -3, 6,
					-- layer=2 filter=53 channel=87
					-20, -43, 18, -57, -75, -55, -71, -57, 0,
					-- layer=2 filter=53 channel=88
					13, -7, 14, 1, 0, 8, -4, 11, -25,
					-- layer=2 filter=53 channel=89
					1, -11, -11, -21, -8, 29, 10, 23, 29,
					-- layer=2 filter=53 channel=90
					0, 5, 7, 0, -5, 0, 3, -2, 5,
					-- layer=2 filter=53 channel=91
					-20, -19, 1, -37, -25, 16, -24, 23, 46,
					-- layer=2 filter=53 channel=92
					17, 8, 21, -9, 10, 28, -16, 27, 0,
					-- layer=2 filter=53 channel=93
					13, -9, -26, 57, -20, -34, 21, 22, -17,
					-- layer=2 filter=53 channel=94
					0, -31, -5, 8, 18, -75, 32, -1, -47,
					-- layer=2 filter=53 channel=95
					15, 12, 14, -8, 16, 0, 9, 11, -7,
					-- layer=2 filter=53 channel=96
					-3, 2, -8, 58, -6, -9, 61, 23, -53,
					-- layer=2 filter=53 channel=97
					-30, 7, 3, -38, 6, 11, -13, 5, 9,
					-- layer=2 filter=53 channel=98
					-1, 9, 10, -7, 5, -19, -14, 34, 30,
					-- layer=2 filter=53 channel=99
					-11, 21, -7, 6, 12, -61, 25, -2, 44,
					-- layer=2 filter=53 channel=100
					-17, -13, 8, -18, -15, -18, -25, -2, -19,
					-- layer=2 filter=53 channel=101
					16, 5, 6, 3, 16, 38, -4, 31, 61,
					-- layer=2 filter=53 channel=102
					10, 13, -6, 23, -9, 0, 23, -19, -9,
					-- layer=2 filter=53 channel=103
					-9, 3, -14, -50, -25, -10, -59, 3, -26,
					-- layer=2 filter=53 channel=104
					-4, -9, -44, -13, -35, -24, -22, -45, -32,
					-- layer=2 filter=53 channel=105
					23, 22, -32, -41, -15, 8, 3, 2, -3,
					-- layer=2 filter=53 channel=106
					-38, -26, -8, -38, 10, 28, -19, 37, 30,
					-- layer=2 filter=53 channel=107
					-51, 9, -13, -17, -4, -10, -32, -9, -31,
					-- layer=2 filter=53 channel=108
					-2, 4, -17, 4, 19, 6, 16, 7, -17,
					-- layer=2 filter=53 channel=109
					4, -8, -8, 8, 3, 1, 12, -9, -5,
					-- layer=2 filter=53 channel=110
					8, -2, 11, 5, 7, -13, 21, 18, -11,
					-- layer=2 filter=53 channel=111
					3, -5, 6, -4, 0, 2, -1, -8, -7,
					-- layer=2 filter=53 channel=112
					-21, 17, -13, 3, -21, -24, 4, -24, 30,
					-- layer=2 filter=53 channel=113
					-5, 24, 21, 14, 0, 0, -5, 20, 47,
					-- layer=2 filter=53 channel=114
					4, 5, 7, 0, -4, -1, 0, 10, 5,
					-- layer=2 filter=53 channel=115
					-3, 8, 0, 12, -3, -5, -4, 8, 4,
					-- layer=2 filter=53 channel=116
					-31, -20, 18, -44, -45, -18, -51, -43, -12,
					-- layer=2 filter=53 channel=117
					-4, -11, -26, -24, 9, 14, 15, 30, 30,
					-- layer=2 filter=53 channel=118
					15, 2, 12, -19, -20, -22, 13, -35, 17,
					-- layer=2 filter=53 channel=119
					-6, 3, 20, -3, 29, 0, 29, 13, 28,
					-- layer=2 filter=53 channel=120
					-3, -5, 7, -9, -5, -1, 0, 4, -6,
					-- layer=2 filter=53 channel=121
					-1, 10, -1, -10, 11, 11, 4, -6, 9,
					-- layer=2 filter=53 channel=122
					-19, -1, 5, 0, 8, -12, 2, -9, -9,
					-- layer=2 filter=53 channel=123
					-3, 18, 6, -19, 12, 5, 15, 1, 16,
					-- layer=2 filter=53 channel=124
					-3, -50, -31, -64, -47, 4, -59, -29, -14,
					-- layer=2 filter=53 channel=125
					9, 11, -4, 9, 2, 8, 1, 6, -11,
					-- layer=2 filter=53 channel=126
					-36, -26, 9, -16, 31, -14, -4, 56, -37,
					-- layer=2 filter=53 channel=127
					4, 13, 24, 22, 6, 11, 4, 2, -44,
					-- layer=2 filter=54 channel=0
					-2, -13, -6, -8, 4, -3, 1, -7, 1,
					-- layer=2 filter=54 channel=1
					-13, -6, -8, -3, -3, 0, 2, -2, -7,
					-- layer=2 filter=54 channel=2
					-1, 2, 5, -6, 4, -1, 0, -7, 6,
					-- layer=2 filter=54 channel=3
					4, -8, 6, -11, 6, -9, -7, 7, 1,
					-- layer=2 filter=54 channel=4
					3, -10, -9, -8, -4, -15, -3, -17, 3,
					-- layer=2 filter=54 channel=5
					0, -7, -10, -3, 0, -7, -2, -13, -1,
					-- layer=2 filter=54 channel=6
					5, -2, -2, -1, -4, -7, -2, -19, -1,
					-- layer=2 filter=54 channel=7
					-16, 2, 2, -10, 1, -8, 5, -5, -1,
					-- layer=2 filter=54 channel=8
					-2, 8, 8, -4, -9, -9, -7, 3, 10,
					-- layer=2 filter=54 channel=9
					2, -2, 4, -2, -9, 1, -8, -1, -1,
					-- layer=2 filter=54 channel=10
					-7, -13, -12, -5, 1, -10, 1, 4, -1,
					-- layer=2 filter=54 channel=11
					2, -5, -17, -4, -3, 3, -10, -6, 1,
					-- layer=2 filter=54 channel=12
					-14, -12, -2, -4, 8, 0, -12, -8, -13,
					-- layer=2 filter=54 channel=13
					4, 0, 0, -8, 3, -5, -7, 1, 9,
					-- layer=2 filter=54 channel=14
					-8, -10, 2, -5, -16, 0, -12, -10, -10,
					-- layer=2 filter=54 channel=15
					-8, -8, 6, -11, -10, -6, -12, 1, 8,
					-- layer=2 filter=54 channel=16
					8, 2, -6, 4, -14, -7, 7, -6, -14,
					-- layer=2 filter=54 channel=17
					10, 10, 6, -2, -2, 0, -1, -3, 2,
					-- layer=2 filter=54 channel=18
					4, -1, 9, 1, -11, -10, 1, 5, -12,
					-- layer=2 filter=54 channel=19
					-8, -1, -9, -4, -3, -9, -9, -9, -15,
					-- layer=2 filter=54 channel=20
					-5, 0, 9, 7, -7, -7, 5, -5, 1,
					-- layer=2 filter=54 channel=21
					7, 8, 5, 6, 6, -2, 2, -2, 7,
					-- layer=2 filter=54 channel=22
					-9, 0, -5, 2, -5, 8, 9, -3, 2,
					-- layer=2 filter=54 channel=23
					5, -15, -7, -9, 2, 2, 4, -5, -5,
					-- layer=2 filter=54 channel=24
					-12, -9, -8, -9, 1, -9, -10, -13, 4,
					-- layer=2 filter=54 channel=25
					0, 2, -13, -10, -1, -6, 1, 3, 10,
					-- layer=2 filter=54 channel=26
					3, -3, -8, -6, -6, 4, -10, -2, 2,
					-- layer=2 filter=54 channel=27
					-2, -1, -15, -11, 7, 6, 0, 0, -11,
					-- layer=2 filter=54 channel=28
					-13, -9, 1, -17, 9, 1, 1, -2, 4,
					-- layer=2 filter=54 channel=29
					0, 6, -10, 3, -9, 10, -3, -1, 4,
					-- layer=2 filter=54 channel=30
					2, 6, 1, 0, 9, -6, -10, -1, -7,
					-- layer=2 filter=54 channel=31
					7, -10, 1, -10, -5, 0, -10, -10, -8,
					-- layer=2 filter=54 channel=32
					-1, 2, -9, -2, 0, -4, -9, -3, 0,
					-- layer=2 filter=54 channel=33
					-15, -4, -4, -5, 4, -8, 0, 3, -1,
					-- layer=2 filter=54 channel=34
					-5, 5, -9, -6, 3, -17, 0, -7, -13,
					-- layer=2 filter=54 channel=35
					-8, -1, -5, 4, -1, 0, -12, 0, -14,
					-- layer=2 filter=54 channel=36
					8, -7, 0, -4, 1, 5, -9, -3, 4,
					-- layer=2 filter=54 channel=37
					9, -8, -9, -17, -11, 0, 2, 2, 3,
					-- layer=2 filter=54 channel=38
					2, 0, -13, -1, -12, -7, 2, 0, -6,
					-- layer=2 filter=54 channel=39
					-7, -10, -8, -2, -7, -3, 2, 1, -6,
					-- layer=2 filter=54 channel=40
					6, -5, 0, 6, -15, -5, -4, -3, 3,
					-- layer=2 filter=54 channel=41
					7, 6, 0, -7, 8, 1, -3, 0, -7,
					-- layer=2 filter=54 channel=42
					-13, -2, 1, -7, 0, 3, 5, -3, -7,
					-- layer=2 filter=54 channel=43
					7, 2, 1, -7, -9, -4, 1, 3, -12,
					-- layer=2 filter=54 channel=44
					0, 9, -10, 9, 0, -5, 3, -10, 7,
					-- layer=2 filter=54 channel=45
					0, -4, -12, -8, -10, -2, 0, 3, 1,
					-- layer=2 filter=54 channel=46
					-4, 5, -10, -16, 9, -2, -2, 7, -16,
					-- layer=2 filter=54 channel=47
					-6, -11, -5, -1, -10, -4, -14, 4, 5,
					-- layer=2 filter=54 channel=48
					9, 0, 4, 7, 8, -9, -6, 0, -8,
					-- layer=2 filter=54 channel=49
					3, -9, 12, 13, -6, -8, -10, -1, 5,
					-- layer=2 filter=54 channel=50
					7, 8, 1, 1, -9, 3, -10, -9, -1,
					-- layer=2 filter=54 channel=51
					0, 0, -2, -13, -7, -3, -3, -4, -10,
					-- layer=2 filter=54 channel=52
					2, -8, 2, -10, -3, 2, -9, -8, -12,
					-- layer=2 filter=54 channel=53
					2, -11, 7, 7, -6, 1, -2, -2, -3,
					-- layer=2 filter=54 channel=54
					-13, -2, -14, -5, -4, 2, -3, -8, 4,
					-- layer=2 filter=54 channel=55
					-9, 10, -2, -2, 7, 0, 2, -1, 1,
					-- layer=2 filter=54 channel=56
					4, -4, -11, -2, -10, -4, -4, -10, -13,
					-- layer=2 filter=54 channel=57
					-1, -5, -3, -2, 0, 8, -6, 1, -4,
					-- layer=2 filter=54 channel=58
					-10, -8, 5, -10, -5, -3, 1, -9, -4,
					-- layer=2 filter=54 channel=59
					-3, 2, -2, 4, 2, -1, -1, 3, -10,
					-- layer=2 filter=54 channel=60
					3, 0, -2, -4, 4, -7, -2, -2, -1,
					-- layer=2 filter=54 channel=61
					-1, -3, -9, 5, 6, -15, 1, -8, 4,
					-- layer=2 filter=54 channel=62
					0, -4, -5, 0, 3, -9, -7, -13, -14,
					-- layer=2 filter=54 channel=63
					-18, -10, 0, -15, -4, -4, -3, 9, -17,
					-- layer=2 filter=54 channel=64
					3, 2, 0, -8, -2, 7, -9, -10, -9,
					-- layer=2 filter=54 channel=65
					-3, -4, -1, -12, -11, -12, 7, -8, -1,
					-- layer=2 filter=54 channel=66
					9, -6, -2, -5, 7, 2, -11, 7, 1,
					-- layer=2 filter=54 channel=67
					-1, -3, 8, -2, -2, -13, -2, -6, -11,
					-- layer=2 filter=54 channel=68
					-9, 2, 8, -12, 2, 0, 8, 7, -3,
					-- layer=2 filter=54 channel=69
					-1, -13, 6, 0, -3, -12, -3, -2, -6,
					-- layer=2 filter=54 channel=70
					-11, -4, -9, -11, -5, 2, -13, -5, -12,
					-- layer=2 filter=54 channel=71
					-3, -12, -14, -11, 5, -11, 2, 9, -6,
					-- layer=2 filter=54 channel=72
					0, -4, -11, 3, -13, 4, 5, -12, -8,
					-- layer=2 filter=54 channel=73
					-12, 2, -11, 6, 2, 7, 7, -11, 9,
					-- layer=2 filter=54 channel=74
					-10, -3, -12, -1, -8, -7, 7, 0, -10,
					-- layer=2 filter=54 channel=75
					-7, -9, 0, -10, -5, -9, 3, -8, -3,
					-- layer=2 filter=54 channel=76
					4, -4, 1, 0, 0, -12, 9, 4, -4,
					-- layer=2 filter=54 channel=77
					1, -9, -1, 6, -2, 8, -11, -7, 8,
					-- layer=2 filter=54 channel=78
					-4, -14, 0, 1, -4, -14, 0, -1, 0,
					-- layer=2 filter=54 channel=79
					-11, 9, -8, 7, 8, 4, -4, -7, -4,
					-- layer=2 filter=54 channel=80
					-2, 6, -4, 0, -7, 7, -9, 2, -9,
					-- layer=2 filter=54 channel=81
					0, -4, -2, 8, 2, -11, -11, -1, 7,
					-- layer=2 filter=54 channel=82
					5, -3, 4, 1, 9, 2, 2, 5, -3,
					-- layer=2 filter=54 channel=83
					-3, -7, -8, -4, -1, -8, -9, 2, -11,
					-- layer=2 filter=54 channel=84
					-3, -7, -3, 1, 6, -4, 2, 5, -10,
					-- layer=2 filter=54 channel=85
					-5, -1, 9, 2, 0, -8, 4, 8, -8,
					-- layer=2 filter=54 channel=86
					1, 7, 7, -1, -4, -9, 5, 5, -10,
					-- layer=2 filter=54 channel=87
					1, -9, -3, -13, -13, 4, 3, -5, 7,
					-- layer=2 filter=54 channel=88
					-13, -3, -1, -3, -1, 0, -8, -9, 3,
					-- layer=2 filter=54 channel=89
					-10, -16, -8, 9, 0, 0, -16, -1, -5,
					-- layer=2 filter=54 channel=90
					2, -6, -8, 5, 3, 5, 10, 0, 0,
					-- layer=2 filter=54 channel=91
					-15, 0, -11, 0, -10, 5, -6, -7, 2,
					-- layer=2 filter=54 channel=92
					0, 3, -5, -1, -8, 8, -12, -4, -9,
					-- layer=2 filter=54 channel=93
					6, 1, -4, -9, 0, -6, 7, -10, -6,
					-- layer=2 filter=54 channel=94
					-16, 1, 4, 2, -1, -10, -4, -5, 0,
					-- layer=2 filter=54 channel=95
					3, -11, 0, -7, 7, -8, -11, 7, -9,
					-- layer=2 filter=54 channel=96
					0, -4, 7, -10, 3, 3, -9, -10, 10,
					-- layer=2 filter=54 channel=97
					-5, 1, -3, -2, -16, -4, -5, 3, -3,
					-- layer=2 filter=54 channel=98
					-8, -5, -15, -14, 5, 6, -8, -3, -9,
					-- layer=2 filter=54 channel=99
					-6, -4, -2, -14, 2, 9, 12, -8, -11,
					-- layer=2 filter=54 channel=100
					-11, -7, 8, -10, -5, -6, -10, -14, 0,
					-- layer=2 filter=54 channel=101
					-1, -7, -10, 0, -4, 5, -12, -2, -2,
					-- layer=2 filter=54 channel=102
					3, 3, -5, -3, 2, -1, -6, -5, 3,
					-- layer=2 filter=54 channel=103
					6, 9, 4, 0, -10, 3, 0, -5, 3,
					-- layer=2 filter=54 channel=104
					-6, 0, 5, -6, -9, -5, -10, -1, -1,
					-- layer=2 filter=54 channel=105
					-4, 9, 4, 1, -5, 5, -2, 5, 2,
					-- layer=2 filter=54 channel=106
					-5, -6, -1, -12, -2, 0, -9, -11, 0,
					-- layer=2 filter=54 channel=107
					-10, 8, 9, -2, -2, -2, 10, -1, 6,
					-- layer=2 filter=54 channel=108
					-7, 0, -8, -1, -9, -2, -22, 1, -10,
					-- layer=2 filter=54 channel=109
					-8, -10, -10, -5, -7, -9, -5, -10, 1,
					-- layer=2 filter=54 channel=110
					-13, -9, -16, 4, 3, 2, 1, 2, -9,
					-- layer=2 filter=54 channel=111
					-2, -1, 3, 5, -5, -8, 2, -8, 8,
					-- layer=2 filter=54 channel=112
					-6, 0, 0, -13, -3, -4, 0, -11, -2,
					-- layer=2 filter=54 channel=113
					1, -4, 0, 8, -3, 4, -9, -3, -8,
					-- layer=2 filter=54 channel=114
					8, 1, 8, -3, -3, -7, -8, 8, 8,
					-- layer=2 filter=54 channel=115
					0, -10, 9, -5, 2, 0, -9, 9, -1,
					-- layer=2 filter=54 channel=116
					4, -11, -4, -2, 0, 5, 7, 0, 1,
					-- layer=2 filter=54 channel=117
					-12, -13, -7, -6, 3, 1, 1, 2, -5,
					-- layer=2 filter=54 channel=118
					0, -3, -9, 0, -6, -10, -13, -4, -14,
					-- layer=2 filter=54 channel=119
					3, -12, 2, -18, -1, -16, -7, -13, -10,
					-- layer=2 filter=54 channel=120
					-1, -9, -5, 0, -7, 0, -6, 8, 3,
					-- layer=2 filter=54 channel=121
					-4, 1, 6, 10, 1, -4, -8, 4, -10,
					-- layer=2 filter=54 channel=122
					7, 1, 7, 5, 3, 0, 9, 7, -1,
					-- layer=2 filter=54 channel=123
					-1, 1, -2, 2, 7, -3, 2, -12, -8,
					-- layer=2 filter=54 channel=124
					-12, -16, 8, -10, -2, 4, 12, -13, 8,
					-- layer=2 filter=54 channel=125
					-10, 4, 10, 2, -8, -4, 6, 9, -2,
					-- layer=2 filter=54 channel=126
					1, -2, 2, 5, -1, -5, 0, -4, -5,
					-- layer=2 filter=54 channel=127
					0, -7, 6, -8, -5, 2, -2, 2, -12,
					-- layer=2 filter=55 channel=0
					-22, -4, -25, 7, -15, -10, -5, 36, 46,
					-- layer=2 filter=55 channel=1
					-19, -20, -1, -19, -12, -7, -14, -30, -26,
					-- layer=2 filter=55 channel=2
					2, -8, -7, -5, -6, 7, 4, -6, 4,
					-- layer=2 filter=55 channel=3
					-30, 7, -23, 3, 19, -9, 19, 38, 9,
					-- layer=2 filter=55 channel=4
					-19, 14, 11, -19, -23, 1, -22, -14, -15,
					-- layer=2 filter=55 channel=5
					-25, -9, -31, -6, 5, 23, 0, 0, 72,
					-- layer=2 filter=55 channel=6
					19, 12, -37, 5, 17, -20, 6, -52, -6,
					-- layer=2 filter=55 channel=7
					-19, -1, -10, -17, 6, -24, 13, 19, -13,
					-- layer=2 filter=55 channel=8
					4, -4, 2, 6, -3, -2, -9, -9, 4,
					-- layer=2 filter=55 channel=9
					-26, -17, -29, 12, 29, 25, -30, -7, -19,
					-- layer=2 filter=55 channel=10
					-17, 7, 0, -7, -15, 6, 1, -3, 25,
					-- layer=2 filter=55 channel=11
					-6, -11, -3, 2, 1, 1, 10, 6, 4,
					-- layer=2 filter=55 channel=12
					-27, -22, 7, 0, 16, 23, -11, -51, -29,
					-- layer=2 filter=55 channel=13
					-3, 5, 5, -7, -10, 9, -2, 3, 2,
					-- layer=2 filter=55 channel=14
					-38, -20, -14, 1, 17, 11, 10, -19, -14,
					-- layer=2 filter=55 channel=15
					-13, -5, 15, -27, 5, -25, -29, -17, -10,
					-- layer=2 filter=55 channel=16
					-27, -10, 9, -16, -24, -9, -7, -14, -24,
					-- layer=2 filter=55 channel=17
					1, -5, 4, 1, -2, -4, -2, -9, 2,
					-- layer=2 filter=55 channel=18
					-22, 2, 17, 1, -28, -11, 0, -22, -11,
					-- layer=2 filter=55 channel=19
					-2, -32, -53, -35, -22, -28, -24, -34, -18,
					-- layer=2 filter=55 channel=20
					-6, 6, -7, -6, 4, 0, -3, -10, -3,
					-- layer=2 filter=55 channel=21
					-5, -1, -3, -4, -10, -11, -4, -10, 0,
					-- layer=2 filter=55 channel=22
					2, 3, -6, -1, 5, 0, 10, -1, 2,
					-- layer=2 filter=55 channel=23
					-18, -25, -2, -22, -64, -57, -63, -45, -19,
					-- layer=2 filter=55 channel=24
					-22, 9, -6, -17, -6, -47, -19, -31, -30,
					-- layer=2 filter=55 channel=25
					8, 5, -7, -20, -19, -35, -11, -37, -34,
					-- layer=2 filter=55 channel=26
					-5, 4, -7, 0, -5, 10, 3, -6, 3,
					-- layer=2 filter=55 channel=27
					-21, -18, -10, 7, 4, 3, 6, 19, 18,
					-- layer=2 filter=55 channel=28
					40, 51, 26, -37, -35, -23, 18, 21, 12,
					-- layer=2 filter=55 channel=29
					4, -1, 0, -6, -11, -2, 4, 6, 8,
					-- layer=2 filter=55 channel=30
					-25, -32, -8, -11, -5, 23, -41, -11, 0,
					-- layer=2 filter=55 channel=31
					-7, -23, -11, 18, 2, -8, -8, -19, -6,
					-- layer=2 filter=55 channel=32
					-10, 7, -8, -8, 7, -7, 4, -1, -3,
					-- layer=2 filter=55 channel=33
					-16, -7, 24, -4, 11, -7, 27, 55, -27,
					-- layer=2 filter=55 channel=34
					19, 8, -7, 11, 7, 6, 4, 5, 5,
					-- layer=2 filter=55 channel=35
					-19, 32, 13, -64, -57, -20, 43, 40, -22,
					-- layer=2 filter=55 channel=36
					0, 0, 4, -5, -8, -4, -10, -7, -1,
					-- layer=2 filter=55 channel=37
					22, 6, 1, -1, 7, 13, 26, 14, 13,
					-- layer=2 filter=55 channel=38
					-31, -24, -11, 0, 2, 27, -10, -26, 21,
					-- layer=2 filter=55 channel=39
					-13, -34, -17, -39, -11, -2, -42, 2, -57,
					-- layer=2 filter=55 channel=40
					5, 28, 1, -20, -5, 5, 10, -24, -2,
					-- layer=2 filter=55 channel=41
					4, -5, 2, 2, 7, -2, 10, -9, 2,
					-- layer=2 filter=55 channel=42
					-5, -4, -6, -11, -8, -18, -44, -31, -29,
					-- layer=2 filter=55 channel=43
					-11, -9, 8, -28, -19, -8, 10, 18, 5,
					-- layer=2 filter=55 channel=44
					7, 4, 9, -5, 4, -3, -2, 5, -4,
					-- layer=2 filter=55 channel=45
					-50, -21, -8, -11, -25, 13, 7, -19, -28,
					-- layer=2 filter=55 channel=46
					-9, -28, -35, -16, -26, -2, -14, -35, -8,
					-- layer=2 filter=55 channel=47
					37, 41, 32, -11, -27, 10, 11, 40, 8,
					-- layer=2 filter=55 channel=48
					3, 6, -9, 9, -1, -5, -3, 8, -1,
					-- layer=2 filter=55 channel=49
					-28, -7, 0, 12, -24, -29, -3, -47, -11,
					-- layer=2 filter=55 channel=50
					-6, 7, 4, 0, 1, -2, -5, 8, 5,
					-- layer=2 filter=55 channel=51
					22, -23, 1, -16, 0, 0, -1, 14, 41,
					-- layer=2 filter=55 channel=52
					-21, 2, 42, 22, 10, -11, 0, 35, 12,
					-- layer=2 filter=55 channel=53
					-5, -29, -17, -18, -27, -45, -16, -64, -10,
					-- layer=2 filter=55 channel=54
					-14, -2, -6, -14, -14, -22, 1, -18, 14,
					-- layer=2 filter=55 channel=55
					6, -5, -9, 6, 2, 3, 1, 8, -5,
					-- layer=2 filter=55 channel=56
					-1, 5, -27, -5, 15, 2, 0, 11, 14,
					-- layer=2 filter=55 channel=57
					-2, 6, -5, -6, 2, 1, -10, 9, -6,
					-- layer=2 filter=55 channel=58
					-44, -46, -42, -10, 11, 10, 0, -35, -42,
					-- layer=2 filter=55 channel=59
					-19, -41, 19, -15, -20, 4, -2, -20, -43,
					-- layer=2 filter=55 channel=60
					-21, -28, -42, -37, -10, 7, -28, -25, -7,
					-- layer=2 filter=55 channel=61
					-16, -30, -20, -12, -45, -42, -17, 2, -42,
					-- layer=2 filter=55 channel=62
					26, -34, -45, 9, -15, -12, 14, -44, 3,
					-- layer=2 filter=55 channel=63
					-10, 11, 4, -27, -31, -7, -40, -7, -26,
					-- layer=2 filter=55 channel=64
					-19, 12, -8, 12, -10, 2, -16, -13, -21,
					-- layer=2 filter=55 channel=65
					13, -19, 3, -12, -3, -59, -17, -24, -23,
					-- layer=2 filter=55 channel=66
					8, 5, 2, -21, -26, -17, -19, -9, -29,
					-- layer=2 filter=55 channel=67
					-31, 4, -37, -9, 7, 0, -43, -64, -25,
					-- layer=2 filter=55 channel=68
					-9, -11, -1, -6, 5, -4, -9, 0, -5,
					-- layer=2 filter=55 channel=69
					-4, -25, 12, 11, 12, 17, 0, -24, -25,
					-- layer=2 filter=55 channel=70
					4, 18, 4, -48, -26, -23, 36, 21, -16,
					-- layer=2 filter=55 channel=71
					7, -5, -17, -5, -14, -1, 17, -10, 1,
					-- layer=2 filter=55 channel=72
					18, 19, 32, 12, -2, -11, 11, 33, 5,
					-- layer=2 filter=55 channel=73
					-20, -5, -31, -35, -27, -23, -6, -24, -39,
					-- layer=2 filter=55 channel=74
					-66, -14, -35, -16, 9, 18, -33, -40, -7,
					-- layer=2 filter=55 channel=75
					17, 35, 23, -6, 25, -7, 33, -25, -5,
					-- layer=2 filter=55 channel=76
					-32, 0, 20, -33, -3, -45, -17, -10, 0,
					-- layer=2 filter=55 channel=77
					-4, 0, -1, -1, 5, -8, -11, 1, -10,
					-- layer=2 filter=55 channel=78
					5, -6, 7, -30, -18, -20, 0, -3, -8,
					-- layer=2 filter=55 channel=79
					-1, 5, -5, 7, -6, -1, 3, -5, -8,
					-- layer=2 filter=55 channel=80
					7, 11, -18, -34, -18, -20, -52, -52, -39,
					-- layer=2 filter=55 channel=81
					-4, 5, 1, -9, 8, 0, 2, 1, -4,
					-- layer=2 filter=55 channel=82
					3, -8, -3, 1, 6, -8, -10, 0, 5,
					-- layer=2 filter=55 channel=83
					-18, -12, -15, -50, -30, -26, -3, -45, -45,
					-- layer=2 filter=55 channel=84
					-6, -10, 8, -2, -7, 7, -3, -7, 7,
					-- layer=2 filter=55 channel=85
					-2, 2, 10, -5, 0, 2, 0, 3, -4,
					-- layer=2 filter=55 channel=86
					-10, 5, 7, -3, -6, -1, -7, -9, -2,
					-- layer=2 filter=55 channel=87
					-32, 24, 17, -24, -26, -55, -41, 25, -16,
					-- layer=2 filter=55 channel=88
					-24, -34, -8, -2, 47, 52, -31, 1, -31,
					-- layer=2 filter=55 channel=89
					-15, -12, 9, -2, -9, 7, -22, -33, -19,
					-- layer=2 filter=55 channel=90
					-4, -4, 6, 2, 0, -5, -7, 10, -8,
					-- layer=2 filter=55 channel=91
					35, 14, 22, -13, -5, 16, -35, -8, -56,
					-- layer=2 filter=55 channel=92
					-20, -36, 2, 4, 0, 2, -31, -35, -24,
					-- layer=2 filter=55 channel=93
					50, 0, -10, 22, 4, -10, 18, -26, -4,
					-- layer=2 filter=55 channel=94
					18, -11, -54, -1, -24, -51, -17, -4, -5,
					-- layer=2 filter=55 channel=95
					-10, 0, -9, -4, 6, -8, 8, -6, 6,
					-- layer=2 filter=55 channel=96
					-34, -15, 0, -4, -22, 49, -36, 13, 22,
					-- layer=2 filter=55 channel=97
					-12, 28, 11, 32, 41, 13, -27, -28, -35,
					-- layer=2 filter=55 channel=98
					28, 34, 26, -33, -44, -20, 27, 34, -32,
					-- layer=2 filter=55 channel=99
					-16, -31, -36, -11, -17, -18, -22, -48, -33,
					-- layer=2 filter=55 channel=100
					-26, -11, -23, -56, -8, 17, 5, -3, 15,
					-- layer=2 filter=55 channel=101
					-18, -13, -12, -27, -6, -14, 9, -2, -32,
					-- layer=2 filter=55 channel=102
					-42, -18, -5, 3, -4, 28, -36, -27, 31,
					-- layer=2 filter=55 channel=103
					15, -10, 0, -16, -22, -3, 0, 12, 12,
					-- layer=2 filter=55 channel=104
					-35, -16, -4, -9, -39, -32, -16, -17, -13,
					-- layer=2 filter=55 channel=105
					2, 12, 22, -71, -28, -19, -40, -7, -15,
					-- layer=2 filter=55 channel=106
					18, 8, -12, -22, 0, 11, -22, -24, -29,
					-- layer=2 filter=55 channel=107
					-19, -25, -19, -17, -10, 5, 13, -13, 16,
					-- layer=2 filter=55 channel=108
					-20, -2, -25, 10, -23, 24, 11, -24, -4,
					-- layer=2 filter=55 channel=109
					5, 0, 1, 0, -2, 5, -4, 0, -6,
					-- layer=2 filter=55 channel=110
					-16, -25, -37, -7, -24, -25, -13, -23, -18,
					-- layer=2 filter=55 channel=111
					-5, 6, -6, 4, -4, 10, 4, 8, 2,
					-- layer=2 filter=55 channel=112
					-31, -29, -22, -24, -37, -12, 17, -16, -15,
					-- layer=2 filter=55 channel=113
					10, -25, 3, -34, -16, 7, 0, -22, -51,
					-- layer=2 filter=55 channel=114
					-4, 5, 0, -1, -9, 3, 7, -6, 6,
					-- layer=2 filter=55 channel=115
					-9, 9, 0, -4, 0, 3, 0, -3, 1,
					-- layer=2 filter=55 channel=116
					-41, 16, 18, -33, -35, -12, -53, 9, -10,
					-- layer=2 filter=55 channel=117
					-63, -22, -11, -13, -13, 19, -17, 10, 9,
					-- layer=2 filter=55 channel=118
					17, 3, 17, -12, -5, -29, 2, 13, -2,
					-- layer=2 filter=55 channel=119
					-7, 27, 15, 14, -41, -16, -5, -31, -27,
					-- layer=2 filter=55 channel=120
					1, 0, 6, 7, 2, -5, -1, 10, 0,
					-- layer=2 filter=55 channel=121
					-7, -4, -6, -6, -2, -7, -8, 0, -8,
					-- layer=2 filter=55 channel=122
					1, 4, -5, -9, -8, 6, -8, 0, 1,
					-- layer=2 filter=55 channel=123
					22, 16, 22, 15, -8, -32, 4, 10, -30,
					-- layer=2 filter=55 channel=124
					-43, -26, 4, -6, 4, -9, 4, 0, 23,
					-- layer=2 filter=55 channel=125
					-10, -2, 0, -9, 1, 3, -5, -1, -3,
					-- layer=2 filter=55 channel=126
					-39, -27, -8, 0, -20, -10, -43, -8, -11,
					-- layer=2 filter=55 channel=127
					-13, -24, 1, -44, 1, -4, -14, -29, -16,
					-- layer=2 filter=56 channel=0
					-2, -6, 19, 26, 4, 11, 15, 34, 4,
					-- layer=2 filter=56 channel=1
					-2, 13, -7, 2, -5, -15, -28, -19, 16,
					-- layer=2 filter=56 channel=2
					8, 10, 11, -3, -6, 6, 7, -1, 8,
					-- layer=2 filter=56 channel=3
					-31, -15, 41, 13, -7, 31, -7, 36, 63,
					-- layer=2 filter=56 channel=4
					-5, -25, -27, -9, 3, -31, 0, -25, -15,
					-- layer=2 filter=56 channel=5
					5, 0, 16, 15, 28, -2, 5, 5, -18,
					-- layer=2 filter=56 channel=6
					20, 27, -31, 32, 35, 12, 15, -2, 34,
					-- layer=2 filter=56 channel=7
					7, -27, 8, -20, -60, 70, -67, -3, 36,
					-- layer=2 filter=56 channel=8
					1, 0, -3, -3, 1, -1, 5, 3, -4,
					-- layer=2 filter=56 channel=9
					27, 31, 0, 24, 0, 3, 27, 0, -11,
					-- layer=2 filter=56 channel=10
					2, -2, 22, 15, 18, 0, 10, 8, 22,
					-- layer=2 filter=56 channel=11
					30, 26, -7, 6, 13, -26, 12, -19, -39,
					-- layer=2 filter=56 channel=12
					25, 8, 13, -39, -13, 23, -17, -13, 37,
					-- layer=2 filter=56 channel=13
					-3, -8, 2, -1, 3, -8, -1, 3, 2,
					-- layer=2 filter=56 channel=14
					27, 24, 2, -35, -29, -15, -15, -24, 2,
					-- layer=2 filter=56 channel=15
					22, -52, -82, -49, -53, -27, -39, -4, 5,
					-- layer=2 filter=56 channel=16
					0, -19, 11, -55, -12, -8, -15, -8, 8,
					-- layer=2 filter=56 channel=17
					-9, -3, 7, 4, -1, 11, 8, 9, 5,
					-- layer=2 filter=56 channel=18
					12, 5, -44, -35, -1, -59, 10, -22, -85,
					-- layer=2 filter=56 channel=19
					10, -50, -43, 8, -29, -12, -11, -37, 14,
					-- layer=2 filter=56 channel=20
					-5, -7, -4, 8, -8, 2, 5, -2, -1,
					-- layer=2 filter=56 channel=21
					-7, -13, -5, -9, -13, -19, 0, -8, -14,
					-- layer=2 filter=56 channel=22
					-5, -8, -3, -11, -10, -1, 6, -7, -2,
					-- layer=2 filter=56 channel=23
					15, -11, 6, 0, -8, -14, -12, 9, 6,
					-- layer=2 filter=56 channel=24
					9, -4, 21, -27, -27, -7, 1, 14, 18,
					-- layer=2 filter=56 channel=25
					-41, -11, 38, -48, -37, 4, 0, -6, 17,
					-- layer=2 filter=56 channel=26
					-3, -3, 8, -6, 1, -8, -10, 0, -3,
					-- layer=2 filter=56 channel=27
					13, -6, -36, 45, 19, -26, 37, -5, -32,
					-- layer=2 filter=56 channel=28
					-13, -6, 50, 11, -1, -23, -3, -4, 1,
					-- layer=2 filter=56 channel=29
					-7, 1, 5, 8, 3, 2, 10, -3, 1,
					-- layer=2 filter=56 channel=30
					0, 7, -25, -11, -12, -56, 38, -28, 8,
					-- layer=2 filter=56 channel=31
					-2, -20, -2, 14, -72, -22, 39, 1, -13,
					-- layer=2 filter=56 channel=32
					6, 6, -3, 0, -4, 0, -4, -5, 1,
					-- layer=2 filter=56 channel=33
					18, 13, 35, -14, -21, 47, -23, -19, 61,
					-- layer=2 filter=56 channel=34
					-15, -3, -7, -39, -21, -20, 18, -48, -50,
					-- layer=2 filter=56 channel=35
					-51, -41, -16, 9, 13, -5, -5, -15, 1,
					-- layer=2 filter=56 channel=36
					-9, -2, -3, 5, -8, 5, 1, 0, -6,
					-- layer=2 filter=56 channel=37
					15, 24, 2, 10, 30, -27, -5, -8, -41,
					-- layer=2 filter=56 channel=38
					13, 16, -21, 1, 21, -33, 10, 15, -14,
					-- layer=2 filter=56 channel=39
					-9, 2, 20, 12, -22, 9, -46, -1, 9,
					-- layer=2 filter=56 channel=40
					20, -10, -49, -19, 15, -11, -40, -10, -12,
					-- layer=2 filter=56 channel=41
					-11, -7, -3, 0, -1, -10, 0, -1, -9,
					-- layer=2 filter=56 channel=42
					12, -12, 21, -3, -6, 63, -43, 22, 44,
					-- layer=2 filter=56 channel=43
					-10, -40, -27, 17, 0, -16, 32, -6, 42,
					-- layer=2 filter=56 channel=44
					-4, -6, 8, 6, -1, 4, 2, 6, -4,
					-- layer=2 filter=56 channel=45
					-48, -28, 22, -23, -44, -11, -2, -28, -1,
					-- layer=2 filter=56 channel=46
					-8, -7, -15, -8, -6, -29, 26, -3, 4,
					-- layer=2 filter=56 channel=47
					-7, 0, 26, 8, -25, -5, 52, -43, -10,
					-- layer=2 filter=56 channel=48
					-12, 3, -10, -3, 6, 5, -4, -4, -10,
					-- layer=2 filter=56 channel=49
					8, 42, -24, -26, 2, -35, -15, -36, -26,
					-- layer=2 filter=56 channel=50
					-3, -17, 8, -6, 14, 7, -17, -24, 0,
					-- layer=2 filter=56 channel=51
					13, 28, 5, 5, 33, -18, 12, -2, -4,
					-- layer=2 filter=56 channel=52
					38, 59, 15, 16, 19, -25, 3, -46, -2,
					-- layer=2 filter=56 channel=53
					23, 8, 2, -9, -51, 34, -6, -21, 52,
					-- layer=2 filter=56 channel=54
					23, 0, 0, -12, -21, 1, -52, -21, -13,
					-- layer=2 filter=56 channel=55
					0, 4, -2, 4, 3, -11, -2, -1, -7,
					-- layer=2 filter=56 channel=56
					13, 22, 0, 31, 19, -25, 6, -7, -24,
					-- layer=2 filter=56 channel=57
					11, -4, -7, -16, -9, -16, 5, 14, 9,
					-- layer=2 filter=56 channel=58
					23, 0, 30, -10, 5, 1, 5, -15, 23,
					-- layer=2 filter=56 channel=59
					1, -9, 5, -9, -31, -6, -9, -7, -3,
					-- layer=2 filter=56 channel=60
					-22, 4, -2, -44, -5, 8, -35, -3, -15,
					-- layer=2 filter=56 channel=61
					11, 34, -4, 11, -5, 17, -14, -40, 3,
					-- layer=2 filter=56 channel=62
					12, 10, -49, 2, 0, -15, -1, -39, -24,
					-- layer=2 filter=56 channel=63
					25, -10, 37, 18, -34, 2, 28, 25, 23,
					-- layer=2 filter=56 channel=64
					-7, -11, -12, 13, 1, -15, 9, -3, 11,
					-- layer=2 filter=56 channel=65
					24, 37, -3, 35, 50, -6, 0, -30, 16,
					-- layer=2 filter=56 channel=66
					4, 29, 33, 22, -29, -19, 64, 22, 21,
					-- layer=2 filter=56 channel=67
					27, -10, -20, 28, -13, -30, 50, 14, -33,
					-- layer=2 filter=56 channel=68
					-6, 5, 0, -8, -10, 8, 9, 11, 0,
					-- layer=2 filter=56 channel=69
					-8, 0, 5, 11, -15, 5, 14, 8, 18,
					-- layer=2 filter=56 channel=70
					-29, -39, 13, 6, 15, -3, -16, 4, -10,
					-- layer=2 filter=56 channel=71
					7, -9, -7, 19, -2, -37, 45, 16, -27,
					-- layer=2 filter=56 channel=72
					2, 7, 15, -49, 19, 31, -60, -52, 28,
					-- layer=2 filter=56 channel=73
					1, -2, -5, 20, -68, 41, 3, -6, -20,
					-- layer=2 filter=56 channel=74
					16, 14, -13, 12, 15, 12, 34, 34, -3,
					-- layer=2 filter=56 channel=75
					37, 21, 54, -18, -10, 3, 41, 2, -6,
					-- layer=2 filter=56 channel=76
					71, 36, 30, -5, -27, -9, 30, -30, -60,
					-- layer=2 filter=56 channel=77
					5, 7, 8, -8, -2, -11, 6, 5, -6,
					-- layer=2 filter=56 channel=78
					-27, -3, -29, -4, 15, -33, 12, 1, -24,
					-- layer=2 filter=56 channel=79
					-1, -1, 9, 10, 0, 8, 12, 8, 3,
					-- layer=2 filter=56 channel=80
					-13, -27, 8, 3, -3, 0, -13, 3, 9,
					-- layer=2 filter=56 channel=81
					-5, 1, -18, 2, -7, 4, 2, 10, 11,
					-- layer=2 filter=56 channel=82
					12, -12, -8, 7, -2, -8, -4, -4, -3,
					-- layer=2 filter=56 channel=83
					-18, -27, -17, -19, -38, -45, -2, -25, 1,
					-- layer=2 filter=56 channel=84
					-4, -8, 11, 2, 1, 2, -4, -8, 8,
					-- layer=2 filter=56 channel=85
					1, -6, 3, 2, -17, -3, 2, -5, 8,
					-- layer=2 filter=56 channel=86
					-8, 4, -7, -14, 17, -8, -2, 8, 1,
					-- layer=2 filter=56 channel=87
					18, 0, -81, -24, -19, -47, -34, 19, -68,
					-- layer=2 filter=56 channel=88
					4, -4, -31, -10, -21, -13, 3, 11, 14,
					-- layer=2 filter=56 channel=89
					-4, -26, 12, -19, -19, -24, -17, -20, 7,
					-- layer=2 filter=56 channel=90
					-1, -6, -10, -4, -4, -6, -3, 4, -3,
					-- layer=2 filter=56 channel=91
					-3, -3, 55, -28, -14, 24, 13, 10, 40,
					-- layer=2 filter=56 channel=92
					-1, -20, 2, -24, -23, -1, -33, -7, 22,
					-- layer=2 filter=56 channel=93
					12, -1, -45, 30, 16, -5, 19, 4, 64,
					-- layer=2 filter=56 channel=94
					10, 0, 35, 1, -31, 28, 2, -36, 13,
					-- layer=2 filter=56 channel=95
					-10, -5, 0, 3, 0, 7, 2, -11, -7,
					-- layer=2 filter=56 channel=96
					33, 41, 38, 90, 44, 43, 40, 47, -18,
					-- layer=2 filter=56 channel=97
					-2, 26, 28, -18, -26, 21, 12, 10, 27,
					-- layer=2 filter=56 channel=98
					-25, -11, 26, -2, 9, 0, -31, -41, -32,
					-- layer=2 filter=56 channel=99
					31, 32, -8, 70, -6, -4, 25, -12, -25,
					-- layer=2 filter=56 channel=100
					10, -35, 9, -4, -2, -5, -13, 2, -30,
					-- layer=2 filter=56 channel=101
					0, -23, 43, 0, 7, 15, 15, 19, 9,
					-- layer=2 filter=56 channel=102
					7, 25, -4, 52, 51, -3, 44, -21, -47,
					-- layer=2 filter=56 channel=103
					-7, -4, 23, 5, 42, 55, -33, -3, -51,
					-- layer=2 filter=56 channel=104
					25, 27, -11, 0, 0, 2, -13, -10, -10,
					-- layer=2 filter=56 channel=105
					-1, 23, 21, -22, -45, 29, -15, -22, -49,
					-- layer=2 filter=56 channel=106
					1, 0, 62, -23, -12, 34, 2, 23, 23,
					-- layer=2 filter=56 channel=107
					8, 48, 1, 3, 14, 38, -47, -4, 11,
					-- layer=2 filter=56 channel=108
					-4, -8, -22, 36, 8, -17, 26, -18, -49,
					-- layer=2 filter=56 channel=109
					-6, 4, -9, 3, 0, 4, -3, 8, 8,
					-- layer=2 filter=56 channel=110
					8, -38, -7, -10, -15, -16, -2, -1, 42,
					-- layer=2 filter=56 channel=111
					-3, 4, -10, -6, 6, -3, 5, -1, -6,
					-- layer=2 filter=56 channel=112
					13, 2, -27, 25, 3, 0, -5, 1, 5,
					-- layer=2 filter=56 channel=113
					-24, -1, 18, -9, -22, -59, 18, -16, 13,
					-- layer=2 filter=56 channel=114
					7, 17, 7, 3, 11, 12, 0, 9, -9,
					-- layer=2 filter=56 channel=115
					2, 8, 4, 10, 3, -7, 7, 0, -9,
					-- layer=2 filter=56 channel=116
					40, 30, -39, -14, 19, -30, -3, -1, -41,
					-- layer=2 filter=56 channel=117
					23, -11, -2, 18, -3, 16, 0, -43, 12,
					-- layer=2 filter=56 channel=118
					-29, -17, -2, -3, -6, -7, 8, 21, 23,
					-- layer=2 filter=56 channel=119
					21, -5, 18, -12, -1, -12, 6, -3, 1,
					-- layer=2 filter=56 channel=120
					-6, 7, 10, -5, 9, -5, -3, -3, 5,
					-- layer=2 filter=56 channel=121
					-9, 0, -2, 6, 0, -1, 3, 0, -5,
					-- layer=2 filter=56 channel=122
					7, -2, 0, 0, -10, -5, 0, -1, 3,
					-- layer=2 filter=56 channel=123
					-14, -5, 26, -33, -27, 8, -46, -42, 14,
					-- layer=2 filter=56 channel=124
					-35, -76, -76, -30, -54, -7, -35, -12, -19,
					-- layer=2 filter=56 channel=125
					9, 2, -8, -11, 0, 10, 6, 9, 0,
					-- layer=2 filter=56 channel=126
					-4, -64, 0, -21, 0, 0, -3, 13, 40,
					-- layer=2 filter=56 channel=127
					1, 7, 20, -6, -44, -58, -20, -8, -1,
					-- layer=2 filter=57 channel=0
					3, 0, -10, -8, 1, -10, -10, -11, -1,
					-- layer=2 filter=57 channel=1
					7, -4, -8, -12, 1, -4, -3, 5, -3,
					-- layer=2 filter=57 channel=2
					0, -9, 8, -4, -2, -11, 4, 7, -3,
					-- layer=2 filter=57 channel=3
					-5, -4, 7, -8, 9, -11, 7, 4, -10,
					-- layer=2 filter=57 channel=4
					-11, -10, 5, -5, 3, 0, 9, 2, -2,
					-- layer=2 filter=57 channel=5
					-3, -5, -3, 4, -8, 5, 1, -1, 5,
					-- layer=2 filter=57 channel=6
					-11, 1, 0, -10, 0, -7, 7, 5, -7,
					-- layer=2 filter=57 channel=7
					0, 0, 1, 2, -4, -9, 3, -2, -2,
					-- layer=2 filter=57 channel=8
					1, 9, -6, 2, -1, 0, 2, -6, -8,
					-- layer=2 filter=57 channel=9
					-2, -8, -5, -2, 6, -5, -5, -7, -11,
					-- layer=2 filter=57 channel=10
					2, -9, 4, 5, 2, -1, -6, -1, -7,
					-- layer=2 filter=57 channel=11
					-8, 6, -7, -2, -2, -1, -1, -2, -5,
					-- layer=2 filter=57 channel=12
					6, -2, -3, -6, 2, -4, -4, 0, 2,
					-- layer=2 filter=57 channel=13
					-6, 9, 11, 4, -2, 5, 3, 0, 2,
					-- layer=2 filter=57 channel=14
					0, -11, -11, -8, 1, 8, 6, 6, -4,
					-- layer=2 filter=57 channel=15
					-6, 2, 5, 2, 3, 1, -8, 8, -7,
					-- layer=2 filter=57 channel=16
					0, -8, 7, -3, 1, -4, -6, -7, -2,
					-- layer=2 filter=57 channel=17
					-8, 0, -2, -11, 0, -8, -4, 10, -7,
					-- layer=2 filter=57 channel=18
					-1, 7, 3, 6, -14, 6, 5, -12, 8,
					-- layer=2 filter=57 channel=19
					-2, -13, -3, 0, -6, -1, -6, -3, -8,
					-- layer=2 filter=57 channel=20
					-6, 5, 3, 8, -7, 3, -2, 11, -3,
					-- layer=2 filter=57 channel=21
					6, -5, 4, -3, 10, 2, 8, 3, 6,
					-- layer=2 filter=57 channel=22
					-6, 0, 2, -6, 4, -7, -10, 10, 9,
					-- layer=2 filter=57 channel=23
					-5, 4, -13, 2, -1, 5, 2, -3, 0,
					-- layer=2 filter=57 channel=24
					4, -8, -1, 3, -5, -2, 0, -11, -10,
					-- layer=2 filter=57 channel=25
					6, -4, 3, -10, -1, 0, 5, 5, -2,
					-- layer=2 filter=57 channel=26
					-5, 2, -5, 5, 0, 8, 2, -7, -5,
					-- layer=2 filter=57 channel=27
					-4, -3, -2, -10, 5, -4, 3, 2, -14,
					-- layer=2 filter=57 channel=28
					3, -12, -5, -10, 2, 6, -12, -4, -8,
					-- layer=2 filter=57 channel=29
					-10, -4, -10, 1, -6, -6, 5, -7, 0,
					-- layer=2 filter=57 channel=30
					0, 1, -7, 0, 0, 5, -7, 0, -4,
					-- layer=2 filter=57 channel=31
					-4, -4, 5, -9, 7, 0, -5, 7, -7,
					-- layer=2 filter=57 channel=32
					-2, -3, 2, -11, -4, 6, 11, 3, -1,
					-- layer=2 filter=57 channel=33
					-6, -7, -2, 6, -1, -6, -12, 3, -2,
					-- layer=2 filter=57 channel=34
					0, 4, -4, -5, 5, 7, -11, 4, -1,
					-- layer=2 filter=57 channel=35
					-4, -2, 4, -2, 0, 1, -8, -8, -4,
					-- layer=2 filter=57 channel=36
					2, -7, -12, -6, -11, 3, 1, -3, 0,
					-- layer=2 filter=57 channel=37
					5, 6, -5, 3, -4, -13, -6, -5, -3,
					-- layer=2 filter=57 channel=38
					-6, -2, 5, -3, -1, 3, -8, 2, 0,
					-- layer=2 filter=57 channel=39
					-8, -5, -6, -6, -11, 0, 6, -1, 2,
					-- layer=2 filter=57 channel=40
					-10, -10, 4, -5, 3, 6, 5, 7, -3,
					-- layer=2 filter=57 channel=41
					5, -5, -11, -11, -12, 10, -3, -2, -6,
					-- layer=2 filter=57 channel=42
					-11, -6, -5, 4, -3, -7, -8, 8, -5,
					-- layer=2 filter=57 channel=43
					3, 6, -6, 0, -8, -8, -5, -9, -10,
					-- layer=2 filter=57 channel=44
					-5, -3, 7, 6, -3, -10, -2, -7, 10,
					-- layer=2 filter=57 channel=45
					-4, 5, 0, 1, 0, 8, -8, -9, 1,
					-- layer=2 filter=57 channel=46
					0, -9, 8, 7, -5, -9, 2, -1, -6,
					-- layer=2 filter=57 channel=47
					0, -3, 5, 7, 2, -4, 4, 3, 0,
					-- layer=2 filter=57 channel=48
					3, 10, -8, 4, -7, 10, 0, 10, 10,
					-- layer=2 filter=57 channel=49
					-8, -9, 4, -11, 5, 2, 2, -3, 6,
					-- layer=2 filter=57 channel=50
					-1, 10, 5, -2, 1, 9, 2, 2, 7,
					-- layer=2 filter=57 channel=51
					-5, 2, 0, -7, -4, 0, 5, -2, -12,
					-- layer=2 filter=57 channel=52
					-12, 2, -7, 0, -10, 6, -6, 7, -7,
					-- layer=2 filter=57 channel=53
					-3, 10, 3, -7, 3, -2, 10, 2, 5,
					-- layer=2 filter=57 channel=54
					-12, -12, -14, 2, -14, 1, -1, -7, -2,
					-- layer=2 filter=57 channel=55
					-6, 4, 3, 5, -2, 0, -11, 1, 9,
					-- layer=2 filter=57 channel=56
					0, -7, -5, 5, 3, 6, -4, 4, -7,
					-- layer=2 filter=57 channel=57
					-1, 4, 6, -5, -3, -2, 4, -3, -10,
					-- layer=2 filter=57 channel=58
					6, -6, 7, 4, -7, 3, -10, -4, 6,
					-- layer=2 filter=57 channel=59
					7, 3, -11, 3, -7, 5, -3, -9, 0,
					-- layer=2 filter=57 channel=60
					3, 0, -3, -1, -6, -1, -3, -3, 0,
					-- layer=2 filter=57 channel=61
					-5, 0, -7, -8, 7, -4, -8, -8, -8,
					-- layer=2 filter=57 channel=62
					0, -3, 0, -7, -9, 2, 0, 5, 4,
					-- layer=2 filter=57 channel=63
					6, -7, -5, -4, 5, -8, -1, -10, -9,
					-- layer=2 filter=57 channel=64
					7, -11, -3, -10, -3, 4, -4, 2, -9,
					-- layer=2 filter=57 channel=65
					0, -11, 3, 4, -12, 6, -5, -11, 2,
					-- layer=2 filter=57 channel=66
					-8, 6, -6, 4, -2, 8, -2, 6, 2,
					-- layer=2 filter=57 channel=67
					5, -2, -6, -8, -5, -10, -3, -8, 6,
					-- layer=2 filter=57 channel=68
					3, 4, 8, 0, 0, -10, 4, 1, 3,
					-- layer=2 filter=57 channel=69
					-13, 8, -4, 0, -6, 3, -12, -12, 11,
					-- layer=2 filter=57 channel=70
					-2, -11, 1, 3, -15, -10, 2, 5, 1,
					-- layer=2 filter=57 channel=71
					-4, -2, 9, -7, 6, -7, 3, 10, 5,
					-- layer=2 filter=57 channel=72
					7, 0, 1, 5, -9, 10, 2, -13, -9,
					-- layer=2 filter=57 channel=73
					-9, -6, 5, -6, -5, 1, -2, 4, 0,
					-- layer=2 filter=57 channel=74
					2, -3, -4, 6, 3, 0, -8, 2, 1,
					-- layer=2 filter=57 channel=75
					-6, 0, 1, -5, -3, 0, 8, -2, 5,
					-- layer=2 filter=57 channel=76
					-4, -10, -9, 4, 5, 4, 1, -5, -6,
					-- layer=2 filter=57 channel=77
					-2, 8, -6, 4, 8, -2, -5, -2, 7,
					-- layer=2 filter=57 channel=78
					8, -2, -10, -3, 2, 7, 1, -2, 3,
					-- layer=2 filter=57 channel=79
					-9, -5, -3, -4, -1, 0, 8, 5, 5,
					-- layer=2 filter=57 channel=80
					7, 3, 0, -3, -3, 1, -11, -11, 3,
					-- layer=2 filter=57 channel=81
					2, 5, -3, 8, 1, 8, 4, -7, -6,
					-- layer=2 filter=57 channel=82
					0, -4, 3, -5, -4, 10, 5, 2, -7,
					-- layer=2 filter=57 channel=83
					-11, 4, 6, -2, 2, -6, 7, 6, -1,
					-- layer=2 filter=57 channel=84
					-2, 5, 5, -9, 4, 6, -7, 4, -3,
					-- layer=2 filter=57 channel=85
					3, 8, -9, -5, 8, 0, -8, 5, -2,
					-- layer=2 filter=57 channel=86
					-3, -6, 0, -3, 7, 11, -9, 10, -6,
					-- layer=2 filter=57 channel=87
					2, 0, 0, 6, 7, -6, -2, -5, 5,
					-- layer=2 filter=57 channel=88
					-7, 0, 0, -7, 0, 3, -12, -6, 5,
					-- layer=2 filter=57 channel=89
					-4, -7, 0, -3, 1, 1, -5, 3, -8,
					-- layer=2 filter=57 channel=90
					-1, -3, 3, 7, -7, 0, 7, 0, -3,
					-- layer=2 filter=57 channel=91
					-6, -8, -8, 0, -5, -8, -8, -14, -6,
					-- layer=2 filter=57 channel=92
					1, -10, 2, 6, 0, 6, -9, -2, 5,
					-- layer=2 filter=57 channel=93
					3, -7, 0, -7, 8, -3, 6, 2, -8,
					-- layer=2 filter=57 channel=94
					2, -4, -1, -2, 7, -2, -8, -8, -1,
					-- layer=2 filter=57 channel=95
					-4, 4, -1, 3, 4, 3, -1, -8, 0,
					-- layer=2 filter=57 channel=96
					1, -2, 1, -7, -1, -2, -6, 7, 1,
					-- layer=2 filter=57 channel=97
					2, -11, -11, -3, 7, -1, 7, -3, 0,
					-- layer=2 filter=57 channel=98
					-10, -5, 5, -3, -12, -11, -3, 1, -7,
					-- layer=2 filter=57 channel=99
					-10, -8, 8, -12, -4, -3, -1, 2, 5,
					-- layer=2 filter=57 channel=100
					-9, -10, 6, 2, 0, -8, 8, 3, 2,
					-- layer=2 filter=57 channel=101
					-7, 0, 0, -6, 0, 0, 6, -12, -4,
					-- layer=2 filter=57 channel=102
					-2, -6, -9, 2, -11, 4, -1, -6, -10,
					-- layer=2 filter=57 channel=103
					-7, -5, 1, 0, 7, -6, -10, 1, 3,
					-- layer=2 filter=57 channel=104
					-6, 7, 2, -2, -10, -4, -3, -1, 5,
					-- layer=2 filter=57 channel=105
					6, 8, -6, -1, -3, -7, -1, -8, 9,
					-- layer=2 filter=57 channel=106
					3, -11, 7, -8, 0, -8, 6, -4, 8,
					-- layer=2 filter=57 channel=107
					0, 10, -5, 0, 1, 1, -11, 1, 5,
					-- layer=2 filter=57 channel=108
					3, 3, -10, -3, -3, -7, -2, 6, 6,
					-- layer=2 filter=57 channel=109
					-3, -4, 0, 2, -3, 0, -9, -11, -2,
					-- layer=2 filter=57 channel=110
					-10, 0, -5, -9, -5, 3, -2, -3, -8,
					-- layer=2 filter=57 channel=111
					-3, -2, 8, -3, -8, -4, -6, -3, -9,
					-- layer=2 filter=57 channel=112
					1, -8, 0, -6, -8, 2, -10, -11, 5,
					-- layer=2 filter=57 channel=113
					-7, 6, 1, -9, -12, -5, -4, 5, 6,
					-- layer=2 filter=57 channel=114
					-11, 0, -3, 1, -11, -2, -4, -3, 6,
					-- layer=2 filter=57 channel=115
					9, -4, 5, 3, 2, -2, 6, -9, -4,
					-- layer=2 filter=57 channel=116
					-6, -11, -6, -5, -2, 5, -7, 0, -5,
					-- layer=2 filter=57 channel=117
					-8, 6, 0, 4, 0, 2, 0, -3, -3,
					-- layer=2 filter=57 channel=118
					6, -10, -1, -5, 6, 4, -8, -9, -3,
					-- layer=2 filter=57 channel=119
					2, -10, -5, -10, -11, 4, -3, -9, 8,
					-- layer=2 filter=57 channel=120
					2, -3, 0, -8, -3, 0, 6, -1, -4,
					-- layer=2 filter=57 channel=121
					-1, -2, 0, -4, 5, 6, 7, -5, 8,
					-- layer=2 filter=57 channel=122
					6, -8, -9, -1, -1, -6, -7, -3, -3,
					-- layer=2 filter=57 channel=123
					-1, -8, 2, -10, 3, -7, 5, 6, -11,
					-- layer=2 filter=57 channel=124
					8, -6, -10, 4, -4, -5, -10, 7, 0,
					-- layer=2 filter=57 channel=125
					-10, 4, 0, -7, -8, 10, 3, 7, 1,
					-- layer=2 filter=57 channel=126
					0, -12, -6, 1, 7, 7, -8, -7, -2,
					-- layer=2 filter=57 channel=127
					-3, 6, -2, 2, -9, 1, -2, 3, -6,
					-- layer=2 filter=58 channel=0
					2, 0, -8, 1, -2, -11, 0, -3, -10,
					-- layer=2 filter=58 channel=1
					3, 7, 3, -12, 0, 0, -8, -11, 4,
					-- layer=2 filter=58 channel=2
					2, 2, -3, 4, -7, 5, -4, 6, 0,
					-- layer=2 filter=58 channel=3
					-4, -2, 0, 0, -7, -9, 5, 0, 2,
					-- layer=2 filter=58 channel=4
					0, 2, 2, 5, -7, -10, 0, 2, -9,
					-- layer=2 filter=58 channel=5
					3, -9, -8, 7, 4, -9, 2, 2, 0,
					-- layer=2 filter=58 channel=6
					-7, -6, -2, -9, 0, 4, -11, -3, 7,
					-- layer=2 filter=58 channel=7
					-7, 6, 0, 1, 4, 7, -6, -5, -5,
					-- layer=2 filter=58 channel=8
					1, 1, 8, -1, 2, 6, -11, -9, -2,
					-- layer=2 filter=58 channel=9
					-9, 6, -3, -7, -1, -5, -1, -5, 6,
					-- layer=2 filter=58 channel=10
					-11, 2, 7, 2, -8, 1, -6, -7, 0,
					-- layer=2 filter=58 channel=11
					-4, -2, 4, 2, 1, -10, -11, 0, -14,
					-- layer=2 filter=58 channel=12
					-7, -3, 0, -1, 6, -2, -7, -1, -11,
					-- layer=2 filter=58 channel=13
					-7, 4, 0, 0, -8, -6, -4, 6, 8,
					-- layer=2 filter=58 channel=14
					-9, -3, 2, 1, -6, -4, -12, 4, -14,
					-- layer=2 filter=58 channel=15
					-4, -8, 7, 6, 2, 4, -7, -6, 4,
					-- layer=2 filter=58 channel=16
					-2, 6, 0, -11, 4, 7, -7, -4, 2,
					-- layer=2 filter=58 channel=17
					7, -3, -7, 9, -6, -6, 9, 8, 2,
					-- layer=2 filter=58 channel=18
					3, 3, 3, -7, -10, 7, 0, 7, 0,
					-- layer=2 filter=58 channel=19
					-14, -9, -10, 0, 0, -5, -12, 1, -13,
					-- layer=2 filter=58 channel=20
					-2, -10, 8, 0, 7, -2, 8, 4, 2,
					-- layer=2 filter=58 channel=21
					-1, -10, -5, 4, 5, -2, -3, 3, 9,
					-- layer=2 filter=58 channel=22
					3, 1, -10, 1, -3, 4, 0, 4, -3,
					-- layer=2 filter=58 channel=23
					-12, 1, -5, 7, -3, -7, -7, 8, -3,
					-- layer=2 filter=58 channel=24
					-4, -5, -8, -10, -12, -9, 7, 3, 5,
					-- layer=2 filter=58 channel=25
					-9, -2, -5, 0, -10, 0, -10, -12, 6,
					-- layer=2 filter=58 channel=26
					2, -6, 5, 3, -3, 1, 9, -5, -10,
					-- layer=2 filter=58 channel=27
					8, -8, 0, -3, -8, 0, -5, -8, 6,
					-- layer=2 filter=58 channel=28
					-1, -11, 5, 3, -3, 4, 5, -13, 4,
					-- layer=2 filter=58 channel=29
					0, -9, -3, -1, -5, 0, 1, 0, -9,
					-- layer=2 filter=58 channel=30
					-1, -10, -8, -3, -1, 4, -10, 1, -6,
					-- layer=2 filter=58 channel=31
					2, -6, 2, 0, 2, -4, -5, -9, -5,
					-- layer=2 filter=58 channel=32
					4, -4, -5, -3, -3, 5, -5, -5, -2,
					-- layer=2 filter=58 channel=33
					-2, 1, -5, -2, -8, -6, 5, 8, -3,
					-- layer=2 filter=58 channel=34
					1, 7, -2, -9, -5, 0, 7, -1, -2,
					-- layer=2 filter=58 channel=35
					-9, -8, 3, -5, 5, -2, 1, 7, -7,
					-- layer=2 filter=58 channel=36
					8, 0, -3, 3, 4, 7, -4, 3, -3,
					-- layer=2 filter=58 channel=37
					-10, -5, -5, -5, -1, -13, -4, 3, -7,
					-- layer=2 filter=58 channel=38
					4, -9, 0, -7, -1, -3, -6, -1, -9,
					-- layer=2 filter=58 channel=39
					-8, 0, 0, 7, 0, -5, 3, -8, -6,
					-- layer=2 filter=58 channel=40
					4, 8, -6, -15, -3, -5, -4, 7, -12,
					-- layer=2 filter=58 channel=41
					4, -1, 4, -8, -2, 5, -2, -3, 10,
					-- layer=2 filter=58 channel=42
					-4, -12, -6, -9, 0, -7, -6, 1, 4,
					-- layer=2 filter=58 channel=43
					3, -6, -7, -4, -8, -1, -10, -10, 4,
					-- layer=2 filter=58 channel=44
					8, 9, 10, 3, 2, 0, -5, 4, -3,
					-- layer=2 filter=58 channel=45
					-8, 0, 4, -7, -7, 1, -10, -2, 3,
					-- layer=2 filter=58 channel=46
					-5, 0, -8, -9, 1, -10, -2, 7, 5,
					-- layer=2 filter=58 channel=47
					-6, 0, -9, -8, 7, -1, -2, -1, -7,
					-- layer=2 filter=58 channel=48
					10, 4, -11, 2, 4, 2, -1, 0, -10,
					-- layer=2 filter=58 channel=49
					6, 1, -3, -13, -9, -4, -3, -14, 1,
					-- layer=2 filter=58 channel=50
					-4, -6, 6, 8, 9, 3, -8, 6, -9,
					-- layer=2 filter=58 channel=51
					-6, -8, 4, 8, -3, -10, -9, -6, -1,
					-- layer=2 filter=58 channel=52
					7, 6, -14, -9, 5, -13, -8, 7, 0,
					-- layer=2 filter=58 channel=53
					2, 0, -8, -9, 5, -1, 0, -7, 8,
					-- layer=2 filter=58 channel=54
					-3, 3, -11, -5, 2, -12, -11, 1, 6,
					-- layer=2 filter=58 channel=55
					-2, 2, 9, 10, -2, -6, 9, -5, 5,
					-- layer=2 filter=58 channel=56
					0, 2, -5, 1, 4, -9, 7, -10, -8,
					-- layer=2 filter=58 channel=57
					0, 5, -10, -3, 0, -8, 0, 6, -7,
					-- layer=2 filter=58 channel=58
					1, 4, -6, 9, -1, 1, 0, -5, -12,
					-- layer=2 filter=58 channel=59
					-2, -5, 0, -4, -9, -2, 4, 4, -2,
					-- layer=2 filter=58 channel=60
					7, 10, 6, -6, 4, -7, -7, -13, 0,
					-- layer=2 filter=58 channel=61
					-3, -5, 3, -2, -1, -4, 0, 6, -6,
					-- layer=2 filter=58 channel=62
					-5, -4, -6, -13, 4, -2, 0, -6, 0,
					-- layer=2 filter=58 channel=63
					9, -1, -12, 4, -11, -2, -3, -10, 0,
					-- layer=2 filter=58 channel=64
					2, -6, -7, -8, -10, -3, -11, -8, 4,
					-- layer=2 filter=58 channel=65
					3, -5, 5, 5, -7, 6, -9, 4, -9,
					-- layer=2 filter=58 channel=66
					-7, -7, 6, -5, 2, 2, -4, 7, 2,
					-- layer=2 filter=58 channel=67
					-3, -6, 4, -9, 2, -11, -4, -1, 0,
					-- layer=2 filter=58 channel=68
					1, -8, 0, 0, 1, 0, 5, -9, 3,
					-- layer=2 filter=58 channel=69
					0, 3, 2, -6, -5, -3, -8, 2, -12,
					-- layer=2 filter=58 channel=70
					9, 2, -3, 2, 6, 3, -12, 2, -13,
					-- layer=2 filter=58 channel=71
					3, -10, -10, -7, -6, -4, 1, -3, 5,
					-- layer=2 filter=58 channel=72
					-1, 8, -5, -7, -8, -9, 4, -1, -3,
					-- layer=2 filter=58 channel=73
					-10, -2, 7, 5, 1, -3, -11, 3, -9,
					-- layer=2 filter=58 channel=74
					-3, -4, 1, 1, 5, -1, -3, -10, -4,
					-- layer=2 filter=58 channel=75
					-1, -3, -1, 1, -11, -4, 8, -11, -7,
					-- layer=2 filter=58 channel=76
					0, -9, 5, 9, 1, -14, -9, -11, 2,
					-- layer=2 filter=58 channel=77
					-3, 3, -5, 4, 6, 7, 6, 6, 0,
					-- layer=2 filter=58 channel=78
					3, 6, 0, -12, -7, -9, -8, -9, -1,
					-- layer=2 filter=58 channel=79
					8, 10, 2, 3, -8, 1, -6, 4, -7,
					-- layer=2 filter=58 channel=80
					4, -3, -3, 6, 4, 5, -7, -1, -8,
					-- layer=2 filter=58 channel=81
					-8, -5, 4, -2, 3, -5, 2, -9, 7,
					-- layer=2 filter=58 channel=82
					0, -1, -9, 5, -10, 7, 8, 7, 5,
					-- layer=2 filter=58 channel=83
					-8, 2, 4, -7, -2, 5, -8, 5, 0,
					-- layer=2 filter=58 channel=84
					3, 4, 6, -2, 1, 5, 5, -4, 8,
					-- layer=2 filter=58 channel=85
					-6, 7, 6, 9, -8, 8, 7, -7, -1,
					-- layer=2 filter=58 channel=86
					4, -7, -11, 3, 7, -7, -9, -5, -5,
					-- layer=2 filter=58 channel=87
					-3, -6, -3, 8, 0, -12, -4, -11, 1,
					-- layer=2 filter=58 channel=88
					-9, 8, 4, -8, 0, -7, 8, 3, -4,
					-- layer=2 filter=58 channel=89
					4, -8, 6, 0, -6, -9, -1, 3, 2,
					-- layer=2 filter=58 channel=90
					-5, 1, -2, -4, 0, 9, -5, 0, -4,
					-- layer=2 filter=58 channel=91
					-9, 3, 1, -4, -13, -1, 2, -4, -7,
					-- layer=2 filter=58 channel=92
					-14, -4, 2, -1, -9, 5, -1, 3, -12,
					-- layer=2 filter=58 channel=93
					-2, -3, 1, -4, 0, -6, -7, 3, -4,
					-- layer=2 filter=58 channel=94
					-14, 0, -2, -3, -9, 5, 3, -8, -1,
					-- layer=2 filter=58 channel=95
					6, -2, -1, 1, 5, -5, 0, -5, 3,
					-- layer=2 filter=58 channel=96
					0, 0, -15, -3, 4, -5, 6, 6, 0,
					-- layer=2 filter=58 channel=97
					2, 6, 5, 1, -2, -4, 5, -10, 0,
					-- layer=2 filter=58 channel=98
					-10, 1, -11, -4, -6, -8, -7, 0, 0,
					-- layer=2 filter=58 channel=99
					-7, -11, -7, 9, -1, 0, -5, 0, 4,
					-- layer=2 filter=58 channel=100
					6, 1, -7, -12, -4, 0, -8, 3, -11,
					-- layer=2 filter=58 channel=101
					4, -1, -6, -10, 10, 9, -4, -10, -2,
					-- layer=2 filter=58 channel=102
					0, 6, -10, -5, 3, -1, -8, 4, 0,
					-- layer=2 filter=58 channel=103
					5, -5, 3, -10, 7, -11, -11, -9, 6,
					-- layer=2 filter=58 channel=104
					8, -8, -8, -4, -4, 2, 7, -8, -5,
					-- layer=2 filter=58 channel=105
					0, 0, 7, -1, -11, -2, -3, 8, -7,
					-- layer=2 filter=58 channel=106
					4, -2, 4, 1, -7, -1, 0, -3, 2,
					-- layer=2 filter=58 channel=107
					6, -9, -1, -1, -9, -8, -5, 4, -10,
					-- layer=2 filter=58 channel=108
					-9, 6, -4, 6, 1, 0, -4, -9, -4,
					-- layer=2 filter=58 channel=109
					4, -12, -2, 0, -2, 7, 4, -1, -3,
					-- layer=2 filter=58 channel=110
					4, 1, -9, 2, -1, -3, -6, -5, -1,
					-- layer=2 filter=58 channel=111
					1, 1, -8, 10, -10, 9, 6, -4, 11,
					-- layer=2 filter=58 channel=112
					2, 2, 0, 7, -12, 4, -4, 0, -5,
					-- layer=2 filter=58 channel=113
					-1, 4, -2, -10, -10, -4, 4, 5, 0,
					-- layer=2 filter=58 channel=114
					2, 0, 8, 2, -2, -3, -3, 0, -6,
					-- layer=2 filter=58 channel=115
					-10, -3, 9, 4, -7, -6, 9, 9, 9,
					-- layer=2 filter=58 channel=116
					-4, 11, 5, 4, -8, 1, -8, -5, 2,
					-- layer=2 filter=58 channel=117
					1, 4, -4, -6, 9, 2, 8, 0, -8,
					-- layer=2 filter=58 channel=118
					-8, 3, -8, 3, 3, 5, -8, -7, 3,
					-- layer=2 filter=58 channel=119
					-2, -7, -13, -3, 1, 5, -9, -11, -15,
					-- layer=2 filter=58 channel=120
					8, -3, 5, -1, 3, 0, -8, 3, -8,
					-- layer=2 filter=58 channel=121
					-3, 4, -4, 6, -10, 6, 7, 7, 0,
					-- layer=2 filter=58 channel=122
					8, 7, -2, 5, 9, 8, -9, 0, 7,
					-- layer=2 filter=58 channel=123
					-3, -1, -12, 0, 0, 4, -5, -4, 2,
					-- layer=2 filter=58 channel=124
					7, -6, -4, -3, -9, -6, -1, -8, -11,
					-- layer=2 filter=58 channel=125
					-10, -2, 9, 6, 2, 2, 7, -8, -7,
					-- layer=2 filter=58 channel=126
					3, -7, 4, -9, 6, 7, 4, 3, 7,
					-- layer=2 filter=58 channel=127
					-10, 0, 2, -6, -4, 2, 0, 4, 5,
					-- layer=2 filter=59 channel=0
					-21, -14, 11, 0, -32, 31, -2, -24, 8,
					-- layer=2 filter=59 channel=1
					-23, -14, 9, -9, 25, 24, 28, 32, 25,
					-- layer=2 filter=59 channel=2
					-8, 5, -8, -8, -11, 5, -8, -2, -6,
					-- layer=2 filter=59 channel=3
					-18, 5, -4, -42, -66, -57, 21, 5, 13,
					-- layer=2 filter=59 channel=4
					-9, 9, -38, -4, -21, -29, -29, -21, 14,
					-- layer=2 filter=59 channel=5
					-7, -10, 33, -17, -2, 38, -15, -46, -2,
					-- layer=2 filter=59 channel=6
					5, -4, 28, 24, 26, 26, -20, 8, 31,
					-- layer=2 filter=59 channel=7
					17, -11, -5, -2, -45, -26, 32, 28, 11,
					-- layer=2 filter=59 channel=8
					-9, 9, 1, 8, 4, 8, -6, 4, 4,
					-- layer=2 filter=59 channel=9
					-53, -19, -60, -18, 2, -64, -38, -32, -54,
					-- layer=2 filter=59 channel=10
					-35, -13, -9, -23, -12, -25, 9, -12, 14,
					-- layer=2 filter=59 channel=11
					-47, -9, 3, -19, -26, 6, 0, -27, -6,
					-- layer=2 filter=59 channel=12
					-41, -25, 18, 15, 31, 37, 21, 32, 22,
					-- layer=2 filter=59 channel=13
					9, 3, 5, -2, -5, 5, -3, -10, 0,
					-- layer=2 filter=59 channel=14
					-19, -29, -15, 4, 4, -2, 34, 15, 14,
					-- layer=2 filter=59 channel=15
					41, -20, -54, 18, 20, -25, -9, 5, 45,
					-- layer=2 filter=59 channel=16
					61, 45, 17, 11, 16, 1, -20, -17, -8,
					-- layer=2 filter=59 channel=17
					2, 5, 9, 1, 10, 7, 8, -5, 1,
					-- layer=2 filter=59 channel=18
					-30, 4, -47, -11, -26, -10, 21, 25, 23,
					-- layer=2 filter=59 channel=19
					-8, 33, 15, -16, 14, 6, 22, 27, 39,
					-- layer=2 filter=59 channel=20
					-1, -7, 11, -6, 0, 0, 9, -2, 2,
					-- layer=2 filter=59 channel=21
					-12, 5, -12, -12, -2, -4, -6, -10, -18,
					-- layer=2 filter=59 channel=22
					4, -3, -7, 10, 2, 1, -1, 1, 6,
					-- layer=2 filter=59 channel=23
					2, 31, 8, -16, -2, -3, -18, -22, 10,
					-- layer=2 filter=59 channel=24
					5, 34, 22, -2, -20, -69, -19, -35, -85,
					-- layer=2 filter=59 channel=25
					44, 35, 39, -12, -12, -15, -26, -32, -49,
					-- layer=2 filter=59 channel=26
					-11, 10, -8, 4, 9, -8, -12, 2, -2,
					-- layer=2 filter=59 channel=27
					-6, 10, 26, -11, 9, 10, -27, -23, -10,
					-- layer=2 filter=59 channel=28
					-6, -7, -61, -55, -28, -29, -7, 28, 26,
					-- layer=2 filter=59 channel=29
					-6, 7, 8, 7, 1, 4, -5, 10, 1,
					-- layer=2 filter=59 channel=30
					30, -5, -11, 10, 25, -24, 2, -12, -25,
					-- layer=2 filter=59 channel=31
					17, 24, -23, 2, 39, -23, -29, -23, -39,
					-- layer=2 filter=59 channel=32
					9, -1, 0, -8, 4, 13, -7, -4, 1,
					-- layer=2 filter=59 channel=33
					13, -16, -38, -1, -23, 30, -33, -6, 56,
					-- layer=2 filter=59 channel=34
					6, 2, -22, -22, -33, -9, -28, -19, 16,
					-- layer=2 filter=59 channel=35
					5, -22, 14, -7, -35, -20, -32, 19, 18,
					-- layer=2 filter=59 channel=36
					-1, 4, 11, 5, -6, 13, -2, 3, 9,
					-- layer=2 filter=59 channel=37
					-19, 9, 24, -13, 0, 21, -26, -8, 17,
					-- layer=2 filter=59 channel=38
					-25, -4, 9, 12, 11, 30, -17, -32, -22,
					-- layer=2 filter=59 channel=39
					-4, 17, 21, -35, -16, 2, -17, -28, -57,
					-- layer=2 filter=59 channel=40
					58, 14, -19, -5, -25, -17, -41, -20, -17,
					-- layer=2 filter=59 channel=41
					-4, 9, -6, 3, -10, 6, 2, 9, 5,
					-- layer=2 filter=59 channel=42
					7, -11, 1, 2, -1, -11, -25, -7, -21,
					-- layer=2 filter=59 channel=43
					-13, 5, -20, -49, -32, -54, -47, -15, 61,
					-- layer=2 filter=59 channel=44
					8, 9, 9, 5, 10, 1, -7, -5, 0,
					-- layer=2 filter=59 channel=45
					40, 11, -16, 13, 1, 11, -16, -13, 13,
					-- layer=2 filter=59 channel=46
					-17, -15, -25, -6, 0, 12, 56, -2, -28,
					-- layer=2 filter=59 channel=47
					7, 1, -36, -27, -35, -43, -10, 6, 19,
					-- layer=2 filter=59 channel=48
					-4, 1, -4, 7, 10, -3, -7, 9, 3,
					-- layer=2 filter=59 channel=49
					32, 21, -31, 37, 20, -8, 41, 16, 2,
					-- layer=2 filter=59 channel=50
					36, 3, -11, 17, 24, 22, 21, 2, 6,
					-- layer=2 filter=59 channel=51
					-26, -16, 25, -27, -27, 20, -22, -26, -10,
					-- layer=2 filter=59 channel=52
					-14, 16, 29, 17, 6, 1, -31, 0, -6,
					-- layer=2 filter=59 channel=53
					38, -31, 9, 21, 51, -28, -3, 14, 5,
					-- layer=2 filter=59 channel=54
					4, -9, -5, -5, -42, 7, 22, 18, 32,
					-- layer=2 filter=59 channel=55
					9, 2, 2, 0, 3, 2, 4, -9, 14,
					-- layer=2 filter=59 channel=56
					-39, 9, 21, -53, -35, 13, -7, -62, -18,
					-- layer=2 filter=59 channel=57
					4, 0, -2, -12, -7, 2, 8, -6, -4,
					-- layer=2 filter=59 channel=58
					-12, -31, 2, 13, 29, 30, 18, 31, 44,
					-- layer=2 filter=59 channel=59
					-41, -12, 8, 0, 3, 16, -20, -12, 27,
					-- layer=2 filter=59 channel=60
					-29, -17, -3, -7, 4, 35, 42, 30, 1,
					-- layer=2 filter=59 channel=61
					-37, -9, 6, 31, -24, -7, 57, 3, -10,
					-- layer=2 filter=59 channel=62
					5, 22, -31, 11, 22, 14, 24, 18, 47,
					-- layer=2 filter=59 channel=63
					-4, 37, -13, -4, 2, -23, -3, -25, -44,
					-- layer=2 filter=59 channel=64
					45, 35, 14, 0, 15, -45, -19, -9, -30,
					-- layer=2 filter=59 channel=65
					-66, 9, 1, 32, -10, 30, 22, 12, -9,
					-- layer=2 filter=59 channel=66
					35, -62, 23, -18, -30, 37, 51, 9, -41,
					-- layer=2 filter=59 channel=67
					-82, -57, -56, -64, -37, -44, -28, -30, -21,
					-- layer=2 filter=59 channel=68
					10, 10, 9, 0, -7, -8, -3, 3, 0,
					-- layer=2 filter=59 channel=69
					19, 27, -12, 19, 0, -23, 16, -6, -12,
					-- layer=2 filter=59 channel=70
					12, -7, 22, -25, -25, 5, -8, 25, 28,
					-- layer=2 filter=59 channel=71
					-18, -4, 15, -15, -1, -18, -27, -38, -5,
					-- layer=2 filter=59 channel=72
					8, 12, -24, 19, -42, -50, 12, 8, 0,
					-- layer=2 filter=59 channel=73
					39, -65, -34, 12, -8, -5, 0, 16, -42,
					-- layer=2 filter=59 channel=74
					-21, -34, -37, -31, -9, -16, -3, -23, 0,
					-- layer=2 filter=59 channel=75
					21, -15, -27, 25, 13, -8, 74, 29, 24,
					-- layer=2 filter=59 channel=76
					5, -12, -21, -20, 6, 30, -41, 6, 3,
					-- layer=2 filter=59 channel=77
					7, 4, 2, 4, 2, -4, -2, 9, -11,
					-- layer=2 filter=59 channel=78
					0, 3, 5, 25, -11, 0, -2, -28, 5,
					-- layer=2 filter=59 channel=79
					-5, -7, 6, -5, 1, 10, -8, 1, -6,
					-- layer=2 filter=59 channel=80
					11, 28, 0, -32, 19, -3, -22, 16, -3,
					-- layer=2 filter=59 channel=81
					1, -3, -3, 3, -5, -12, -12, 1, -12,
					-- layer=2 filter=59 channel=82
					-4, 5, 4, 13, -8, 8, 6, 6, 0,
					-- layer=2 filter=59 channel=83
					15, 15, 24, 7, 30, -1, -18, 16, -3,
					-- layer=2 filter=59 channel=84
					-2, -5, -12, -1, 7, -1, -4, 2, -11,
					-- layer=2 filter=59 channel=85
					-12, 9, 16, -5, 8, 2, -10, 2, -6,
					-- layer=2 filter=59 channel=86
					-12, 18, 13, 4, 2, -1, 0, 13, 0,
					-- layer=2 filter=59 channel=87
					-24, 13, -54, 18, -3, 3, -3, 20, 50,
					-- layer=2 filter=59 channel=88
					-8, 35, -14, -5, 43, -9, -35, -12, -33,
					-- layer=2 filter=59 channel=89
					-8, -33, 12, 1, 19, -11, 3, 16, 29,
					-- layer=2 filter=59 channel=90
					5, -10, -7, -3, -2, -5, -4, 0, 6,
					-- layer=2 filter=59 channel=91
					-31, 1, 6, 14, 15, 11, 14, 41, -8,
					-- layer=2 filter=59 channel=92
					-11, 14, -1, -1, 26, 40, 3, 11, 0,
					-- layer=2 filter=59 channel=93
					-34, 44, 47, -17, 35, -2, 0, -10, 34,
					-- layer=2 filter=59 channel=94
					0, -9, 1, 48, 30, -30, 53, 19, 60,
					-- layer=2 filter=59 channel=95
					-16, -6, 0, -11, -15, 3, 0, -9, -9,
					-- layer=2 filter=59 channel=96
					-7, 57, 61, 6, 31, 4, 37, 48, 15,
					-- layer=2 filter=59 channel=97
					1, -16, -29, -58, -40, -65, -9, 0, -27,
					-- layer=2 filter=59 channel=98
					7, -9, -27, 7, -36, -23, 18, 12, 16,
					-- layer=2 filter=59 channel=99
					-27, -4, 29, 5, 2, 3, 36, 70, 7,
					-- layer=2 filter=59 channel=100
					-40, -5, 1, -6, 13, 0, -6, -11, -6,
					-- layer=2 filter=59 channel=101
					-20, -19, 14, -54, -36, 1, -42, -27, -12,
					-- layer=2 filter=59 channel=102
					1, 44, -3, 23, 16, -4, 24, 43, -3,
					-- layer=2 filter=59 channel=103
					-16, 43, -16, -23, 54, 49, 7, 0, 8,
					-- layer=2 filter=59 channel=104
					11, 21, -4, 20, 33, 4, 36, 13, 3,
					-- layer=2 filter=59 channel=105
					-8, 8, -34, 18, -20, -8, 41, -20, 29,
					-- layer=2 filter=59 channel=106
					-9, -9, -20, -14, -8, 23, -40, 3, -37,
					-- layer=2 filter=59 channel=107
					1, 45, -34, 11, 12, -32, 19, 30, -36,
					-- layer=2 filter=59 channel=108
					1, 8, 4, 9, 27, 3, -6, -19, 0,
					-- layer=2 filter=59 channel=109
					-3, 12, -15, 5, 0, 6, -11, 19, 7,
					-- layer=2 filter=59 channel=110
					13, 56, 30, -12, 14, -8, -25, -39, -70,
					-- layer=2 filter=59 channel=111
					2, -11, 3, 4, -8, 8, 6, 5, -10,
					-- layer=2 filter=59 channel=112
					-23, -46, 34, 8, -84, -4, 48, -4, -39,
					-- layer=2 filter=59 channel=113
					6, 29, -1, 16, 6, 10, 4, -19, -92,
					-- layer=2 filter=59 channel=114
					-8, 5, -1, -4, 7, 0, -7, -11, -5,
					-- layer=2 filter=59 channel=115
					8, -1, -1, -6, -3, -6, -11, 10, 3,
					-- layer=2 filter=59 channel=116
					-24, 32, -9, 16, 14, 6, 3, 46, 12,
					-- layer=2 filter=59 channel=117
					-36, -73, -11, 16, -36, -73, 22, 21, -9,
					-- layer=2 filter=59 channel=118
					18, 17, -22, -25, 2, -28, -20, 9, 23,
					-- layer=2 filter=59 channel=119
					11, 23, -26, -8, 1, -28, 1, 7, 37,
					-- layer=2 filter=59 channel=120
					-2, 7, -1, -4, 8, 4, 10, -8, 8,
					-- layer=2 filter=59 channel=121
					2, 4, -1, 3, 0, -4, -7, 0, 9,
					-- layer=2 filter=59 channel=122
					5, 3, 6, 20, -14, -11, -12, -10, -5,
					-- layer=2 filter=59 channel=123
					-6, -25, -24, -21, -38, -14, 20, 10, 10,
					-- layer=2 filter=59 channel=124
					35, -9, -54, 22, -13, 3, -6, 41, 61,
					-- layer=2 filter=59 channel=125
					8, -6, 5, 6, 5, 4, -4, -3, 0,
					-- layer=2 filter=59 channel=126
					32, 123, 2, -50, 34, -16, 35, -7, 33,
					-- layer=2 filter=59 channel=127
					0, 3, 8, 7, -4, -3, 1, 4, -21,
					-- layer=2 filter=60 channel=0
					-20, -27, -8, -5, 2, -8, -31, -14, 34,
					-- layer=2 filter=60 channel=1
					-20, 3, 3, 17, 8, 7, -39, 36, 16,
					-- layer=2 filter=60 channel=2
					11, 9, -4, -5, 6, 4, 4, 8, -4,
					-- layer=2 filter=60 channel=3
					-36, 1, 24, -45, -38, -23, -25, -25, -33,
					-- layer=2 filter=60 channel=4
					-5, 9, -12, -6, 5, -8, 24, 2, 6,
					-- layer=2 filter=60 channel=5
					-12, 0, -27, -11, -18, -22, -53, -7, 24,
					-- layer=2 filter=60 channel=6
					43, -27, -24, -27, -54, 31, -39, -105, 22,
					-- layer=2 filter=60 channel=7
					-21, 7, 44, -25, -21, -38, -3, 16, 11,
					-- layer=2 filter=60 channel=8
					10, 5, -5, -7, 6, 8, 9, 8, 7,
					-- layer=2 filter=60 channel=9
					-8, -43, 21, 12, -3, 6, 7, 24, -13,
					-- layer=2 filter=60 channel=10
					-27, -12, -11, -26, -12, 5, -14, -16, 21,
					-- layer=2 filter=60 channel=11
					12, -34, -8, -39, 1, 3, -23, 1, -12,
					-- layer=2 filter=60 channel=12
					10, -24, -32, 29, -26, -6, -64, 11, -8,
					-- layer=2 filter=60 channel=13
					-6, -3, 9, 9, -3, 1, 7, 4, 5,
					-- layer=2 filter=60 channel=14
					12, -7, -2, 3, -4, -6, -56, 9, -21,
					-- layer=2 filter=60 channel=15
					39, 16, -28, 20, -2, -14, 6, 32, 9,
					-- layer=2 filter=60 channel=16
					-43, -16, 10, 5, -23, -4, 23, 22, 1,
					-- layer=2 filter=60 channel=17
					0, -6, -5, -3, -1, -6, -3, 6, -5,
					-- layer=2 filter=60 channel=18
					0, -17, -55, 10, -55, -39, -30, -1, -17,
					-- layer=2 filter=60 channel=19
					-65, 16, -3, 12, 30, 16, 0, 38, 9,
					-- layer=2 filter=60 channel=20
					-7, -6, 2, 8, -4, 9, -7, 12, 7,
					-- layer=2 filter=60 channel=21
					-8, -15, -18, -2, -5, -4, -14, -16, -4,
					-- layer=2 filter=60 channel=22
					3, 4, 3, 2, 4, 3, 6, -9, 4,
					-- layer=2 filter=60 channel=23
					39, 28, 21, 26, 31, 3, 3, 16, 11,
					-- layer=2 filter=60 channel=24
					-26, -24, 0, -30, -51, -7, -14, -13, 2,
					-- layer=2 filter=60 channel=25
					45, 26, -4, -47, -50, -27, 1, -31, 33,
					-- layer=2 filter=60 channel=26
					10, -7, -8, 4, 5, -3, -8, 1, -10,
					-- layer=2 filter=60 channel=27
					-111, -62, -19, -20, 27, 34, -18, 2, 10,
					-- layer=2 filter=60 channel=28
					4, -18, -1, -4, -21, -29, -79, -35, -4,
					-- layer=2 filter=60 channel=29
					-8, 2, 7, -2, 0, 8, 5, -2, -10,
					-- layer=2 filter=60 channel=30
					1, 10, -15, 0, 25, -24, -9, 5, 3,
					-- layer=2 filter=60 channel=31
					-15, 4, 28, 35, 24, 1, 27, 37, -2,
					-- layer=2 filter=60 channel=32
					-2, -2, -5, 2, -1, -8, -10, -9, 2,
					-- layer=2 filter=60 channel=33
					8, 4, 74, -52, -12, -44, -16, -12, 32,
					-- layer=2 filter=60 channel=34
					28, 35, -2, 67, -20, -11, 36, 7, 45,
					-- layer=2 filter=60 channel=35
					11, 13, 11, 24, -10, -2, -51, -22, -3,
					-- layer=2 filter=60 channel=36
					0, 0, 11, -7, -4, 0, -1, 0, -2,
					-- layer=2 filter=60 channel=37
					-25, -13, -35, -23, 0, -4, -24, 18, -4,
					-- layer=2 filter=60 channel=38
					-45, 11, -24, 0, -4, 39, -18, -26, 0,
					-- layer=2 filter=60 channel=39
					-26, 18, 34, -7, 18, 0, 9, 25, 2,
					-- layer=2 filter=60 channel=40
					-36, 14, 23, 32, 53, 24, 15, -5, 17,
					-- layer=2 filter=60 channel=41
					2, -6, -1, -6, -1, -9, 7, -1, -7,
					-- layer=2 filter=60 channel=42
					-3, 3, 25, 20, 16, 9, 16, 2, -5,
					-- layer=2 filter=60 channel=43
					-13, -6, -39, -41, -23, 5, -23, -22, -33,
					-- layer=2 filter=60 channel=44
					3, 0, 0, -1, -7, 8, -4, 1, 3,
					-- layer=2 filter=60 channel=45
					-92, -82, -60, -21, -21, 0, 19, 0, 1,
					-- layer=2 filter=60 channel=46
					-12, 11, -17, 2, -6, -3, 46, 14, 17,
					-- layer=2 filter=60 channel=47
					-41, -50, -17, -43, -6, -19, 8, -9, 17,
					-- layer=2 filter=60 channel=48
					-8, 8, 2, 0, -7, 7, -11, 1, -9,
					-- layer=2 filter=60 channel=49
					14, -7, -36, 49, -54, 18, 1, 26, 0,
					-- layer=2 filter=60 channel=50
					-10, 1, 11, -13, -6, -3, -23, 1, -15,
					-- layer=2 filter=60 channel=51
					-16, -30, -23, -18, -39, -4, -54, -2, -7,
					-- layer=2 filter=60 channel=52
					13, -52, -51, 0, 5, -11, 13, 3, -20,
					-- layer=2 filter=60 channel=53
					3, -62, -6, -4, 20, 6, 55, -26, 42,
					-- layer=2 filter=60 channel=54
					28, -7, -23, -9, -50, -18, -8, 6, 28,
					-- layer=2 filter=60 channel=55
					12, 0, 11, -1, 16, -2, 7, 4, 1,
					-- layer=2 filter=60 channel=56
					-10, -16, 0, -18, 7, -13, -30, -17, -12,
					-- layer=2 filter=60 channel=57
					1, -4, -1, 2, -6, -1, -7, -7, 0,
					-- layer=2 filter=60 channel=58
					27, 5, -4, -10, -22, -4, -50, -27, 21,
					-- layer=2 filter=60 channel=59
					-10, -23, 0, -21, 55, -17, -30, 12, 17,
					-- layer=2 filter=60 channel=60
					0, 50, -58, -22, -20, 7, -39, -20, -8,
					-- layer=2 filter=60 channel=61
					-4, -44, -35, -33, -35, -6, -52, -43, 15,
					-- layer=2 filter=60 channel=62
					45, -18, 10, 7, -37, 4, -1, -17, 10,
					-- layer=2 filter=60 channel=63
					1, 14, 14, 11, 40, 21, -11, 18, 13,
					-- layer=2 filter=60 channel=64
					2, 6, 19, 19, 29, 5, 36, 25, -4,
					-- layer=2 filter=60 channel=65
					30, 0, -48, -44, -52, 6, -23, -68, 20,
					-- layer=2 filter=60 channel=66
					5, -12, 24, -1, 8, -2, -14, -17, -67,
					-- layer=2 filter=60 channel=67
					-19, 3, 0, 2, 16, -10, 33, 20, -25,
					-- layer=2 filter=60 channel=68
					1, 1, -6, 5, -7, 8, -3, -1, 1,
					-- layer=2 filter=60 channel=69
					11, 12, 19, 11, 12, 17, 12, 35, -10,
					-- layer=2 filter=60 channel=70
					13, -3, 6, -3, -20, -39, -23, -20, 10,
					-- layer=2 filter=60 channel=71
					-32, -2, 0, -9, 0, 0, 7, 12, 27,
					-- layer=2 filter=60 channel=72
					-54, -29, 28, -18, -24, -22, -22, -16, -22,
					-- layer=2 filter=60 channel=73
					8, -28, -24, 71, 30, -7, 96, 28, 35,
					-- layer=2 filter=60 channel=74
					-3, 7, -1, 24, 34, -10, 10, 29, -9,
					-- layer=2 filter=60 channel=75
					6, -6, 3, -8, -42, 19, -52, -18, 24,
					-- layer=2 filter=60 channel=76
					49, -16, -8, -1, -33, 5, 37, 8, 39,
					-- layer=2 filter=60 channel=77
					-2, -8, 3, 3, 5, 0, -9, 10, -2,
					-- layer=2 filter=60 channel=78
					18, -27, -50, -14, -23, -30, -7, 7, -24,
					-- layer=2 filter=60 channel=79
					4, -2, 0, -2, 0, 4, 6, -5, 2,
					-- layer=2 filter=60 channel=80
					-9, 1, 11, 0, 17, 1, 18, 15, -1,
					-- layer=2 filter=60 channel=81
					10, 10, 7, 9, 9, -2, 0, -7, 0,
					-- layer=2 filter=60 channel=82
					0, -8, 1, -10, 9, 6, -1, 0, -4,
					-- layer=2 filter=60 channel=83
					-17, -2, -17, 4, 9, -21, -1, 18, 0,
					-- layer=2 filter=60 channel=84
					-2, 9, 6, -1, -2, -5, 2, 2, -5,
					-- layer=2 filter=60 channel=85
					-2, 0, 1, 9, -4, -2, -3, 5, 10,
					-- layer=2 filter=60 channel=86
					15, 0, 2, 5, 1, -1, 9, 15, -15,
					-- layer=2 filter=60 channel=87
					56, 15, -33, 35, -13, 7, -11, 2, 42,
					-- layer=2 filter=60 channel=88
					-18, 2, 0, 9, 24, 17, -9, 11, -2,
					-- layer=2 filter=60 channel=89
					28, 2, 25, 35, 22, 7, -32, 21, -3,
					-- layer=2 filter=60 channel=90
					6, 7, -3, -6, 7, 0, 4, 8, 8,
					-- layer=2 filter=60 channel=91
					-34, -29, -6, 22, -12, -5, -46, -2, -43,
					-- layer=2 filter=60 channel=92
					-1, -14, -7, 15, 0, 15, -40, 22, -10,
					-- layer=2 filter=60 channel=93
					38, 30, 22, -14, -34, 12, 10, -35, 23,
					-- layer=2 filter=60 channel=94
					29, -71, -24, 0, -4, 18, -8, -54, 41,
					-- layer=2 filter=60 channel=95
					2, -16, -4, 0, 0, -7, 1, 2, -6,
					-- layer=2 filter=60 channel=96
					15, -51, 1, 30, -21, 36, -32, -24, 35,
					-- layer=2 filter=60 channel=97
					-19, -16, 20, -23, -29, -3, -5, 7, -2,
					-- layer=2 filter=60 channel=98
					-34, -56, -24, -29, -40, -41, -14, -14, 6,
					-- layer=2 filter=60 channel=99
					-38, -31, -32, 20, 38, -57, 0, 9, 22,
					-- layer=2 filter=60 channel=100
					-17, -10, -1, -2, 25, 6, 28, -23, -18,
					-- layer=2 filter=60 channel=101
					29, -4, -18, 30, -33, -36, 0, -32, -6,
					-- layer=2 filter=60 channel=102
					11, -26, -39, 42, -33, 2, -15, -8, -19,
					-- layer=2 filter=60 channel=103
					-4, -21, -2, 26, 13, 29, -15, -18, 6,
					-- layer=2 filter=60 channel=104
					24, -62, -34, 7, -45, 27, -17, 35, 24,
					-- layer=2 filter=60 channel=105
					60, -26, -5, -5, 22, 12, 39, 26, 19,
					-- layer=2 filter=60 channel=106
					45, 12, 14, -22, -41, 7, -53, -35, 12,
					-- layer=2 filter=60 channel=107
					50, 53, -3, 0, -21, -19, -6, 5, -33,
					-- layer=2 filter=60 channel=108
					-15, -34, -31, 23, 34, 20, -29, 68, 11,
					-- layer=2 filter=60 channel=109
					1, -1, 16, -5, 11, 3, 3, -4, 3,
					-- layer=2 filter=60 channel=110
					-21, 2, -11, 16, 14, -21, 4, 18, 3,
					-- layer=2 filter=60 channel=111
					8, -2, 9, -8, -6, -5, 5, 0, -8,
					-- layer=2 filter=60 channel=112
					-43, -36, -33, -44, -77, -25, -40, -48, 28,
					-- layer=2 filter=60 channel=113
					15, 23, -18, 15, 39, 0, 8, -2, 12,
					-- layer=2 filter=60 channel=114
					-9, 6, 5, 3, -6, 2, 0, 11, 7,
					-- layer=2 filter=60 channel=115
					7, 2, 0, -9, -1, 4, 0, -9, 3,
					-- layer=2 filter=60 channel=116
					26, 0, -83, 47, -18, -1, 9, -40, 20,
					-- layer=2 filter=60 channel=117
					-3, -32, -23, 15, 54, 9, -10, 1, 1,
					-- layer=2 filter=60 channel=118
					-3, -14, 0, -33, -25, 0, -20, -17, -1,
					-- layer=2 filter=60 channel=119
					29, -14, 7, -1, -6, -9, 13, -12, -25,
					-- layer=2 filter=60 channel=120
					2, 9, 0, 5, 8, 0, 7, 3, -6,
					-- layer=2 filter=60 channel=121
					-2, 3, -3, 6, 11, -4, -4, 0, 0,
					-- layer=2 filter=60 channel=122
					8, -1, 6, 7, 6, 7, -7, 4, 2,
					-- layer=2 filter=60 channel=123
					-23, -4, 23, -47, -30, -21, -4, 6, 16,
					-- layer=2 filter=60 channel=124
					67, 44, 26, -1, -31, -2, 32, 75, 28,
					-- layer=2 filter=60 channel=125
					-5, -8, 4, -5, -8, 4, 8, 9, 7,
					-- layer=2 filter=60 channel=126
					51, 11, 51, 27, 69, 24, -16, -30, 27,
					-- layer=2 filter=60 channel=127
					14, -1, 18, 33, 18, 17, 7, 17, -7,
					-- layer=2 filter=61 channel=0
					17, 9, -6, 3, 11, 7, 0, 9, 7,
					-- layer=2 filter=61 channel=1
					-33, -25, 6, 19, -40, -11, -16, -23, -24,
					-- layer=2 filter=61 channel=2
					-5, -5, -8, 4, -1, -5, -3, -2, 2,
					-- layer=2 filter=61 channel=3
					9, 29, -8, 32, 8, 0, -9, -4, -4,
					-- layer=2 filter=61 channel=4
					-19, 4, -5, -7, -29, 40, 31, -19, -19,
					-- layer=2 filter=61 channel=5
					9, 22, -4, -17, 12, 7, 12, 4, -1,
					-- layer=2 filter=61 channel=6
					-19, -10, 11, -34, 9, -64, 35, 5, -22,
					-- layer=2 filter=61 channel=7
					-32, -49, -57, -13, -15, 10, -4, -4, -32,
					-- layer=2 filter=61 channel=8
					-1, -10, -4, -4, 8, 3, 8, -4, 3,
					-- layer=2 filter=61 channel=9
					-19, 0, -7, -23, -11, 6, -36, -23, 2,
					-- layer=2 filter=61 channel=10
					24, 16, 9, 21, 20, 19, 3, -3, 31,
					-- layer=2 filter=61 channel=11
					11, 2, -34, 29, 13, -19, 16, 19, 0,
					-- layer=2 filter=61 channel=12
					-7, 1, -4, 31, -21, -25, 1, -28, -64,
					-- layer=2 filter=61 channel=13
					-1, 2, 1, -8, 3, 1, 7, -1, -3,
					-- layer=2 filter=61 channel=14
					-9, -11, -37, 41, -2, -22, 12, 0, -28,
					-- layer=2 filter=61 channel=15
					38, 0, 12, 18, 10, -28, 4, -12, -26,
					-- layer=2 filter=61 channel=16
					-13, -28, 3, 5, -5, 31, 23, -3, 18,
					-- layer=2 filter=61 channel=17
					6, -10, 8, -8, 0, -8, 7, 8, 9,
					-- layer=2 filter=61 channel=18
					9, 26, 1, 3, -42, 33, 30, 11, -35,
					-- layer=2 filter=61 channel=19
					-24, -48, 13, -36, -26, -14, -25, -40, -29,
					-- layer=2 filter=61 channel=20
					-3, -1, 5, -7, -9, 1, 5, 8, -9,
					-- layer=2 filter=61 channel=21
					-10, 5, -9, -8, -3, -3, 5, -7, 1,
					-- layer=2 filter=61 channel=22
					8, -10, -1, -4, -6, -8, -4, -11, -11,
					-- layer=2 filter=61 channel=23
					6, -5, -14, 18, 16, 3, -10, 7, 1,
					-- layer=2 filter=61 channel=24
					-7, 24, -1, 7, 30, 4, 10, 2, 18,
					-- layer=2 filter=61 channel=25
					0, -13, -23, -4, 14, 1, 16, 23, 10,
					-- layer=2 filter=61 channel=26
					5, 0, 1, 2, 10, 3, -3, -3, -5,
					-- layer=2 filter=61 channel=27
					-9, 31, 42, 2, 18, 27, 5, -12, 9,
					-- layer=2 filter=61 channel=28
					-16, -18, -63, 5, -33, -3, -6, -14, -12,
					-- layer=2 filter=61 channel=29
					-9, -11, 2, -7, -1, 4, 0, -7, -6,
					-- layer=2 filter=61 channel=30
					-7, -44, 19, 0, -9, 0, -6, 8, 17,
					-- layer=2 filter=61 channel=31
					-2, -27, -80, -21, -19, 96, -7, 45, 41,
					-- layer=2 filter=61 channel=32
					-3, -2, 7, -7, -5, 2, 4, -11, 3,
					-- layer=2 filter=61 channel=33
					-28, 36, -27, 13, 22, 22, -17, -1, -23,
					-- layer=2 filter=61 channel=34
					48, 31, 74, 36, 0, 29, 28, 37, 55,
					-- layer=2 filter=61 channel=35
					-10, 7, 2, 8, 1, 19, 45, 38, 10,
					-- layer=2 filter=61 channel=36
					-2, 10, 0, -10, -2, -9, 1, -4, 3,
					-- layer=2 filter=61 channel=37
					-1, -8, -17, 13, 7, 8, 17, 15, 10,
					-- layer=2 filter=61 channel=38
					-6, 4, 23, -1, 48, 1, 20, 1, -2,
					-- layer=2 filter=61 channel=39
					-47, -24, -11, 3, 16, 63, -1, 6, -9,
					-- layer=2 filter=61 channel=40
					5, -21, 4, -23, 0, -34, -12, -28, -38,
					-- layer=2 filter=61 channel=41
					-1, 5, -5, 1, 8, 10, 4, -2, 4,
					-- layer=2 filter=61 channel=42
					6, -1, 29, 10, 1, -1, 50, -12, 5,
					-- layer=2 filter=61 channel=43
					-30, -31, 16, -21, -11, 18, -6, 20, -18,
					-- layer=2 filter=61 channel=44
					-4, -7, 3, -8, -5, 6, -2, -8, 0,
					-- layer=2 filter=61 channel=45
					4, 23, -30, -43, -32, 15, 8, -64, -16,
					-- layer=2 filter=61 channel=46
					6, -2, -5, -14, -16, -12, 0, -13, -6,
					-- layer=2 filter=61 channel=47
					-31, -11, -40, -30, 0, -19, -41, -50, -7,
					-- layer=2 filter=61 channel=48
					-2, -7, -1, 7, 8, 0, -3, 2, 2,
					-- layer=2 filter=61 channel=49
					-3, -4, -22, 12, -38, 0, -7, -14, -29,
					-- layer=2 filter=61 channel=50
					15, 14, 8, 24, 25, 23, 21, 3, -2,
					-- layer=2 filter=61 channel=51
					10, -11, -14, 21, 16, -1, 22, 30, 4,
					-- layer=2 filter=61 channel=52
					11, -16, -2, 10, -34, -5, -2, 16, 0,
					-- layer=2 filter=61 channel=53
					-11, -34, -24, -15, -74, -52, -48, -8, -38,
					-- layer=2 filter=61 channel=54
					27, 8, -20, 15, 4, -2, 8, 5, 0,
					-- layer=2 filter=61 channel=55
					1, 10, 11, -2, -8, -7, 9, -9, -9,
					-- layer=2 filter=61 channel=56
					-1, 3, -27, 29, 12, -1, 20, 17, -1,
					-- layer=2 filter=61 channel=57
					11, -2, -16, 5, 10, -5, -8, 3, -4,
					-- layer=2 filter=61 channel=58
					-17, 14, 22, -1, -3, -2, -6, -25, -22,
					-- layer=2 filter=61 channel=59
					19, 42, 22, 5, -12, 38, 11, 35, 23,
					-- layer=2 filter=61 channel=60
					-4, 27, 58, 4, 36, 36, -5, -10, 56,
					-- layer=2 filter=61 channel=61
					0, 13, 24, -27, -1, 5, -33, 3, 19,
					-- layer=2 filter=61 channel=62
					0, -15, 1, 11, -24, -49, 17, 21, -12,
					-- layer=2 filter=61 channel=63
					-2, -21, 0, -8, 2, 18, 3, -8, 22,
					-- layer=2 filter=61 channel=64
					-1, 4, 13, 4, 7, -2, 23, 14, 5,
					-- layer=2 filter=61 channel=65
					-37, 0, 20, -1, -2, -29, 15, 17, 6,
					-- layer=2 filter=61 channel=66
					-7, -61, -25, -44, -14, 5, -20, 22, 3,
					-- layer=2 filter=61 channel=67
					-13, -20, -32, -36, -36, -22, -23, -56, -23,
					-- layer=2 filter=61 channel=68
					-8, -1, -6, 6, 8, 0, 1, 10, 5,
					-- layer=2 filter=61 channel=69
					-25, -18, 7, 16, 3, 18, 30, 15, 13,
					-- layer=2 filter=61 channel=70
					5, 21, 18, 10, 11, 17, 20, 2, 5,
					-- layer=2 filter=61 channel=71
					-49, -20, 0, 8, -28, -11, -47, -13, -13,
					-- layer=2 filter=61 channel=72
					2, 51, 2, 27, 6, 12, 9, 8, -24,
					-- layer=2 filter=61 channel=73
					-26, -46, -29, -69, -24, 22, -54, -24, 12,
					-- layer=2 filter=61 channel=74
					5, -4, -12, -30, -2, -31, 6, -20, -2,
					-- layer=2 filter=61 channel=75
					0, -4, -59, 38, -60, -129, -82, -52, -42,
					-- layer=2 filter=61 channel=76
					18, -21, 5, 2, 23, -16, -67, -58, -55,
					-- layer=2 filter=61 channel=77
					-10, 6, 0, 4, 5, 3, 0, 3, -7,
					-- layer=2 filter=61 channel=78
					3, -10, -32, 12, -22, -21, 14, 34, -12,
					-- layer=2 filter=61 channel=79
					-6, -1, 2, -2, -1, -8, 10, 1, 0,
					-- layer=2 filter=61 channel=80
					-28, -1, 7, -5, -7, 1, -3, -24, 8,
					-- layer=2 filter=61 channel=81
					-3, -12, 0, 8, 10, -3, -2, 8, -4,
					-- layer=2 filter=61 channel=82
					-7, 0, 4, -7, -4, -6, 2, -1, 9,
					-- layer=2 filter=61 channel=83
					-6, -12, 19, -25, -21, 6, 6, 4, -5,
					-- layer=2 filter=61 channel=84
					8, -5, 5, 6, 5, -1, -5, 6, -10,
					-- layer=2 filter=61 channel=85
					7, -2, -5, -7, -7, -11, -16, -3, 11,
					-- layer=2 filter=61 channel=86
					-11, -7, -22, -1, -9, 7, 3, 2, -20,
					-- layer=2 filter=61 channel=87
					11, 49, 64, 30, 24, -2, 14, 64, 20,
					-- layer=2 filter=61 channel=88
					-29, -14, -10, -34, -12, -6, 3, -3, -13,
					-- layer=2 filter=61 channel=89
					-7, -10, -6, 15, -23, -26, 0, 12, -43,
					-- layer=2 filter=61 channel=90
					-3, -5, 10, -7, 4, -8, 6, -3, -10,
					-- layer=2 filter=61 channel=91
					-6, 37, 30, 15, 6, 4, -22, -25, -19,
					-- layer=2 filter=61 channel=92
					-40, 7, 28, 16, -13, -3, 14, -21, -54,
					-- layer=2 filter=61 channel=93
					-37, -78, 75, -4, -43, -20, -4, -37, -39,
					-- layer=2 filter=61 channel=94
					-60, -41, -17, -18, -48, -54, -55, -3, -36,
					-- layer=2 filter=61 channel=95
					-13, -2, -2, 3, 8, -1, 9, -2, -3,
					-- layer=2 filter=61 channel=96
					22, -10, 7, 15, -23, -4, -14, 34, 0,
					-- layer=2 filter=61 channel=97
					-1, 35, -19, 16, 18, 23, -6, -4, 16,
					-- layer=2 filter=61 channel=98
					-9, 7, -1, 26, 14, 2, 1, 9, -8,
					-- layer=2 filter=61 channel=99
					-19, -43, -1, -37, -37, -33, -33, -15, 1,
					-- layer=2 filter=61 channel=100
					-9, 16, 24, -14, 33, 11, 7, -12, 16,
					-- layer=2 filter=61 channel=101
					-35, -54, -30, -3, -21, -30, -26, -2, -55,
					-- layer=2 filter=61 channel=102
					9, -19, -5, 3, -65, 14, 6, -12, -10,
					-- layer=2 filter=61 channel=103
					-74, -36, -18, -49, -62, -55, 67, 71, -15,
					-- layer=2 filter=61 channel=104
					-24, 33, -22, 24, -55, -34, -13, -1, -42,
					-- layer=2 filter=61 channel=105
					-18, -26, -66, -26, -23, -26, -33, -28, -57,
					-- layer=2 filter=61 channel=106
					-12, -5, -12, 22, 19, 7, 8, -18, 5,
					-- layer=2 filter=61 channel=107
					-41, -62, 56, -13, -6, -65, 38, 3, 27,
					-- layer=2 filter=61 channel=108
					-4, -19, -1, 21, -25, -15, -16, -20, -13,
					-- layer=2 filter=61 channel=109
					-5, 10, -4, -4, 10, -19, 5, -6, 2,
					-- layer=2 filter=61 channel=110
					-19, -7, 27, -5, 3, 32, 13, 29, 5,
					-- layer=2 filter=61 channel=111
					6, 2, 9, -1, 3, 7, 3, -4, 9,
					-- layer=2 filter=61 channel=112
					6, 10, -5, -28, -1, -5, -9, -17, 7,
					-- layer=2 filter=61 channel=113
					1, -25, 28, 8, 0, 17, -17, 27, 23,
					-- layer=2 filter=61 channel=114
					-10, -25, 0, 4, -3, -13, -5, -14, -5,
					-- layer=2 filter=61 channel=115
					-4, 9, 5, -2, -7, -5, -10, 6, -5,
					-- layer=2 filter=61 channel=116
					-7, 43, 31, 4, 5, -13, 14, 26, 1,
					-- layer=2 filter=61 channel=117
					-20, -40, -36, -32, -74, -42, -10, -30, -38,
					-- layer=2 filter=61 channel=118
					-36, 14, 3, -5, -6, -12, 2, -4, 8,
					-- layer=2 filter=61 channel=119
					-15, -23, -11, -8, -26, 19, 31, -2, -13,
					-- layer=2 filter=61 channel=120
					-1, 0, 2, 6, 8, 0, -5, 0, 9,
					-- layer=2 filter=61 channel=121
					-6, -5, -5, -4, -6, -3, -10, -10, 0,
					-- layer=2 filter=61 channel=122
					14, 15, 5, 0, -1, 2, -5, 10, -6,
					-- layer=2 filter=61 channel=123
					-16, 13, -22, 20, 0, 6, -4, 0, -6,
					-- layer=2 filter=61 channel=124
					35, -3, -25, 7, 8, -25, 0, 8, -19,
					-- layer=2 filter=61 channel=125
					-2, -8, 0, -2, -1, -10, 4, 3, 6,
					-- layer=2 filter=61 channel=126
					-3, -5, 37, -33, -25, 64, 5, 0, 7,
					-- layer=2 filter=61 channel=127
					0, -27, -3, 25, -18, 15, -1, -9, 16,
					-- layer=2 filter=62 channel=0
					-3, 8, -9, 3, 1, -5, 0, -1, -11,
					-- layer=2 filter=62 channel=1
					1, 5, 0, -13, -9, -1, -7, -2, 4,
					-- layer=2 filter=62 channel=2
					-6, 0, 5, 0, 8, -4, 0, 2, 8,
					-- layer=2 filter=62 channel=3
					-3, -7, 7, -9, 2, 5, 3, 0, 1,
					-- layer=2 filter=62 channel=4
					6, 5, 0, 4, 6, -5, 0, -2, 4,
					-- layer=2 filter=62 channel=5
					0, 7, -5, -3, 6, -12, -6, -7, 4,
					-- layer=2 filter=62 channel=6
					1, -8, 5, 0, 3, 0, -11, 7, 4,
					-- layer=2 filter=62 channel=7
					-7, 1, -2, -16, -3, -3, -15, -4, -14,
					-- layer=2 filter=62 channel=8
					-5, 4, 6, -3, 4, -9, -3, 2, 6,
					-- layer=2 filter=62 channel=9
					-10, 0, 1, -8, -10, -11, 8, -11, 6,
					-- layer=2 filter=62 channel=10
					-10, -6, 6, 1, -2, 6, -5, 7, 6,
					-- layer=2 filter=62 channel=11
					7, 9, 7, -8, -2, 0, 3, 3, 8,
					-- layer=2 filter=62 channel=12
					2, -15, -16, -4, -7, -2, -10, -13, 0,
					-- layer=2 filter=62 channel=13
					7, -6, -3, 7, -11, 5, -9, -1, -5,
					-- layer=2 filter=62 channel=14
					0, -7, 5, 0, -1, -2, -7, -2, 0,
					-- layer=2 filter=62 channel=15
					-11, -8, 4, 3, -12, 5, 4, 2, 2,
					-- layer=2 filter=62 channel=16
					9, 0, -6, 6, 3, -10, 2, 3, -12,
					-- layer=2 filter=62 channel=17
					-5, 8, -8, -9, -3, 8, 4, 11, -4,
					-- layer=2 filter=62 channel=18
					-9, 0, -4, -4, -7, -6, 1, 5, -5,
					-- layer=2 filter=62 channel=19
					2, 9, 7, -11, -3, 1, -8, -7, -6,
					-- layer=2 filter=62 channel=20
					-2, -4, 0, -11, -3, 6, 3, 5, -1,
					-- layer=2 filter=62 channel=21
					0, 6, -10, -2, -2, 3, -4, 3, -7,
					-- layer=2 filter=62 channel=22
					6, -9, -6, -9, -2, 2, -10, 9, -4,
					-- layer=2 filter=62 channel=23
					3, -8, -5, -6, 6, -15, 3, -13, -7,
					-- layer=2 filter=62 channel=24
					3, -8, -3, -8, 5, 5, -3, -2, -10,
					-- layer=2 filter=62 channel=25
					7, -9, 0, -5, -3, 2, -14, -1, 0,
					-- layer=2 filter=62 channel=26
					0, 5, 3, 2, -10, 1, -6, 2, 7,
					-- layer=2 filter=62 channel=27
					-9, 0, -2, 4, 5, 7, 4, 6, 1,
					-- layer=2 filter=62 channel=28
					6, -12, -9, 0, -10, -3, -5, 0, 4,
					-- layer=2 filter=62 channel=29
					-9, 0, -4, -12, -10, -9, -2, -8, -4,
					-- layer=2 filter=62 channel=30
					-4, -7, 0, -1, -9, 3, -5, 5, 6,
					-- layer=2 filter=62 channel=31
					-11, 4, 6, 8, -2, -3, -10, 6, -2,
					-- layer=2 filter=62 channel=32
					-10, 5, -10, -8, -4, 6, 9, 6, 3,
					-- layer=2 filter=62 channel=33
					5, 8, 0, 4, 7, -6, -5, -10, 2,
					-- layer=2 filter=62 channel=34
					5, -7, -11, -11, 4, 0, -5, -8, 3,
					-- layer=2 filter=62 channel=35
					0, -7, 5, 1, -5, 0, -5, -12, -14,
					-- layer=2 filter=62 channel=36
					-7, -7, 3, 0, 0, -11, -11, -11, -10,
					-- layer=2 filter=62 channel=37
					-10, -1, -1, -1, 10, -9, -10, 2, 0,
					-- layer=2 filter=62 channel=38
					2, -5, -9, -11, -10, -8, 0, -4, 4,
					-- layer=2 filter=62 channel=39
					-1, -11, 7, 0, -10, -6, -5, 1, -4,
					-- layer=2 filter=62 channel=40
					-3, -3, 1, 5, -1, -9, 8, 8, 8,
					-- layer=2 filter=62 channel=41
					-8, 3, 0, 3, -3, 3, -1, 0, 1,
					-- layer=2 filter=62 channel=42
					-9, 6, -4, 5, -2, -4, 4, -6, 0,
					-- layer=2 filter=62 channel=43
					0, 4, -4, -10, -2, -4, -8, -7, -11,
					-- layer=2 filter=62 channel=44
					6, -9, 7, 0, -5, -10, -8, 0, -4,
					-- layer=2 filter=62 channel=45
					4, 7, -5, 3, -1, 1, 4, -2, 8,
					-- layer=2 filter=62 channel=46
					-5, -4, -1, -1, -8, -2, -12, 7, -10,
					-- layer=2 filter=62 channel=47
					0, 5, -1, 1, -6, -12, 5, -11, -1,
					-- layer=2 filter=62 channel=48
					-6, -2, -3, -4, -10, -3, -4, 8, -7,
					-- layer=2 filter=62 channel=49
					7, -9, -15, 0, 3, -13, -4, -6, 3,
					-- layer=2 filter=62 channel=50
					5, 0, -5, 0, 0, -2, -6, -1, 0,
					-- layer=2 filter=62 channel=51
					-3, -6, -1, -7, 7, 0, -6, -9, -2,
					-- layer=2 filter=62 channel=52
					1, 0, -6, 0, 3, 3, 8, 1, -2,
					-- layer=2 filter=62 channel=53
					-5, -12, -3, 1, -5, 6, -9, -12, -11,
					-- layer=2 filter=62 channel=54
					-10, 4, -3, 5, -6, -9, 5, -8, -7,
					-- layer=2 filter=62 channel=55
					-11, -6, 5, 8, -4, 2, -10, 7, -8,
					-- layer=2 filter=62 channel=56
					2, -6, 9, -6, -6, 3, -3, -6, -2,
					-- layer=2 filter=62 channel=57
					0, 0, -9, -1, 4, 3, 5, -3, -8,
					-- layer=2 filter=62 channel=58
					-3, -8, -8, -8, 7, 3, 5, 6, -10,
					-- layer=2 filter=62 channel=59
					3, -9, -11, -10, -15, -1, 4, -6, -5,
					-- layer=2 filter=62 channel=60
					-2, -10, -13, -2, -7, -7, 4, 6, -5,
					-- layer=2 filter=62 channel=61
					-14, -6, -11, 4, -2, -9, 4, -5, 2,
					-- layer=2 filter=62 channel=62
					-9, 6, -7, -9, -5, -5, -8, -12, -7,
					-- layer=2 filter=62 channel=63
					0, 0, 8, -3, -9, 6, -5, -4, 0,
					-- layer=2 filter=62 channel=64
					0, 5, -5, -1, 1, 6, -12, 1, -4,
					-- layer=2 filter=62 channel=65
					-6, -9, 0, -9, 8, 6, -3, -8, 4,
					-- layer=2 filter=62 channel=66
					-2, 8, -2, 4, -9, -10, -3, -1, -7,
					-- layer=2 filter=62 channel=67
					-6, 0, -3, 1, -3, 1, 0, -7, -10,
					-- layer=2 filter=62 channel=68
					4, 5, -2, -8, -10, 5, -12, 6, 2,
					-- layer=2 filter=62 channel=69
					-2, 2, -8, 2, 5, 7, -13, 5, 1,
					-- layer=2 filter=62 channel=70
					9, 3, 5, 3, -4, 2, -1, 0, -11,
					-- layer=2 filter=62 channel=71
					0, -9, -1, 0, -8, -3, 1, -9, 5,
					-- layer=2 filter=62 channel=72
					-13, -7, -2, -3, -1, -1, -10, -9, -7,
					-- layer=2 filter=62 channel=73
					-11, -7, 0, -1, -5, 2, -11, -3, -8,
					-- layer=2 filter=62 channel=74
					7, -9, 6, -1, -4, -3, 0, -1, 1,
					-- layer=2 filter=62 channel=75
					5, 0, 8, -12, -6, 1, -11, -3, -7,
					-- layer=2 filter=62 channel=76
					-6, -9, -11, 4, 4, -11, 7, 5, -5,
					-- layer=2 filter=62 channel=77
					-8, -10, 6, 8, -3, 4, -5, -7, -3,
					-- layer=2 filter=62 channel=78
					-2, 4, -12, -5, -2, 4, -1, -8, -1,
					-- layer=2 filter=62 channel=79
					-5, -6, 0, 8, -11, 0, 2, -12, -10,
					-- layer=2 filter=62 channel=80
					-8, -1, 7, 8, 2, -3, -11, 3, -3,
					-- layer=2 filter=62 channel=81
					-3, -11, -3, 8, -6, -7, 4, 7, -6,
					-- layer=2 filter=62 channel=82
					-4, 5, 1, -6, 7, 4, 1, -6, -5,
					-- layer=2 filter=62 channel=83
					-6, -10, -2, -3, -7, -10, 0, -6, -9,
					-- layer=2 filter=62 channel=84
					-8, -9, 5, 5, -9, -9, -1, -7, -9,
					-- layer=2 filter=62 channel=85
					-2, -2, 8, -7, -3, -10, 2, -9, -5,
					-- layer=2 filter=62 channel=86
					-7, 5, 12, -5, -1, -1, -2, -3, -7,
					-- layer=2 filter=62 channel=87
					3, 1, -1, 0, 0, 6, -6, -5, -5,
					-- layer=2 filter=62 channel=88
					-2, -8, -1, 4, -11, 3, -2, -5, 7,
					-- layer=2 filter=62 channel=89
					-6, -2, 0, -6, -8, -9, 0, -6, -14,
					-- layer=2 filter=62 channel=90
					-1, 2, -3, -2, 1, 4, 10, 11, -2,
					-- layer=2 filter=62 channel=91
					-14, 1, -4, -12, -4, -13, 0, -16, 4,
					-- layer=2 filter=62 channel=92
					0, -9, -5, -15, -1, 3, 9, 1, -15,
					-- layer=2 filter=62 channel=93
					8, 0, -3, -3, 1, 3, -9, 0, -1,
					-- layer=2 filter=62 channel=94
					-8, -3, 0, 2, -9, -5, -4, -14, -13,
					-- layer=2 filter=62 channel=95
					1, 0, 3, -7, -6, 6, -6, -9, 0,
					-- layer=2 filter=62 channel=96
					-2, 4, 2, -5, -1, 3, 9, 4, -12,
					-- layer=2 filter=62 channel=97
					0, -5, 4, 7, 6, 3, 0, -5, -9,
					-- layer=2 filter=62 channel=98
					-9, 1, 4, -12, -3, 11, -14, 2, -13,
					-- layer=2 filter=62 channel=99
					1, 2, 7, 3, 10, -2, -13, -14, -1,
					-- layer=2 filter=62 channel=100
					-4, -8, 4, -9, -4, -7, -1, 7, -10,
					-- layer=2 filter=62 channel=101
					-5, 6, -9, -7, 4, -4, -3, -7, -11,
					-- layer=2 filter=62 channel=102
					9, -12, 4, -12, -6, -5, 5, -3, -13,
					-- layer=2 filter=62 channel=103
					8, 1, 1, 6, 1, 3, -3, -6, -1,
					-- layer=2 filter=62 channel=104
					-3, -5, 0, 6, -1, 0, -12, -10, -15,
					-- layer=2 filter=62 channel=105
					3, -1, -3, 3, 4, 0, 7, 5, -3,
					-- layer=2 filter=62 channel=106
					0, -6, -4, 7, 3, 7, 11, -10, -5,
					-- layer=2 filter=62 channel=107
					-10, -6, -5, 1, -5, 1, 3, -12, -4,
					-- layer=2 filter=62 channel=108
					0, 4, -10, 3, 7, 0, 6, 1, -11,
					-- layer=2 filter=62 channel=109
					3, -2, 2, 5, -10, -2, 0, 0, -1,
					-- layer=2 filter=62 channel=110
					-1, 6, -12, -12, 2, -2, -5, -2, -11,
					-- layer=2 filter=62 channel=111
					-3, 2, -5, 2, -10, -8, 6, -8, 8,
					-- layer=2 filter=62 channel=112
					5, 0, -5, -11, -1, -7, -3, 0, -12,
					-- layer=2 filter=62 channel=113
					-8, 3, 5, 8, -3, 3, -8, -8, 2,
					-- layer=2 filter=62 channel=114
					-9, 3, -4, 4, 10, 8, -8, -3, 9,
					-- layer=2 filter=62 channel=115
					9, 7, -4, -7, -4, 8, 0, 4, 4,
					-- layer=2 filter=62 channel=116
					-6, -7, 0, -1, -5, -1, 3, -3, -7,
					-- layer=2 filter=62 channel=117
					6, 1, 0, -3, 0, -11, -1, -1, 4,
					-- layer=2 filter=62 channel=118
					1, -1, 9, 2, 7, 4, -1, 5, 5,
					-- layer=2 filter=62 channel=119
					7, -6, -3, 1, -1, -12, 5, -8, -13,
					-- layer=2 filter=62 channel=120
					-4, 3, -3, 4, 0, 8, -6, 1, 0,
					-- layer=2 filter=62 channel=121
					-7, -10, -3, -5, 4, 1, -11, 10, -5,
					-- layer=2 filter=62 channel=122
					0, 0, -2, -10, 0, 8, -7, 4, -10,
					-- layer=2 filter=62 channel=123
					5, -4, -5, 1, -5, 2, -16, 0, -14,
					-- layer=2 filter=62 channel=124
					-4, 5, 9, 6, -1, 0, -3, 2, -12,
					-- layer=2 filter=62 channel=125
					-10, 7, -3, 6, -7, 4, 6, 9, 7,
					-- layer=2 filter=62 channel=126
					-5, -1, -6, -2, 3, -3, -3, 5, -1,
					-- layer=2 filter=62 channel=127
					0, -9, -5, 8, 7, -2, 3, -11, 7,
					-- layer=2 filter=63 channel=0
					-17, 6, 9, -17, -4, 14, -6, 26, -14,
					-- layer=2 filter=63 channel=1
					-18, 15, -12, -8, -13, 4, 1, -15, 15,
					-- layer=2 filter=63 channel=2
					0, -3, -1, 4, 6, -4, 9, -6, -1,
					-- layer=2 filter=63 channel=3
					10, 26, 19, 44, 49, 18, -1, -7, -8,
					-- layer=2 filter=63 channel=4
					-10, -13, -29, -43, -12, -4, -8, 39, -1,
					-- layer=2 filter=63 channel=5
					12, 12, 4, -13, 11, 2, 1, 5, -1,
					-- layer=2 filter=63 channel=6
					12, 10, -20, 40, 11, 9, 10, 16, -34,
					-- layer=2 filter=63 channel=7
					-6, 38, 36, 30, 16, 2, 62, 39, 32,
					-- layer=2 filter=63 channel=8
					-4, 4, 5, -11, -3, -3, -1, -6, -4,
					-- layer=2 filter=63 channel=9
					-2, 10, -12, 6, 29, 43, -2, -6, 3,
					-- layer=2 filter=63 channel=10
					-2, 36, 28, -12, 13, 30, 21, 12, -4,
					-- layer=2 filter=63 channel=11
					3, -5, 12, 19, -2, 9, 5, 11, -1,
					-- layer=2 filter=63 channel=12
					-5, 35, -17, 17, 30, 20, -5, -10, 32,
					-- layer=2 filter=63 channel=13
					-5, 7, 0, -1, -2, -11, -11, 9, -3,
					-- layer=2 filter=63 channel=14
					8, 13, -18, 8, 18, 29, 5, -7, 28,
					-- layer=2 filter=63 channel=15
					-10, -25, -23, -10, -27, -27, 28, -21, 1,
					-- layer=2 filter=63 channel=16
					8, 7, 18, 24, 23, 11, 12, -2, 9,
					-- layer=2 filter=63 channel=17
					8, 8, -6, 0, -7, -6, 6, -9, -2,
					-- layer=2 filter=63 channel=18
					5, -31, -49, -55, -41, -39, -48, -49, -50,
					-- layer=2 filter=63 channel=19
					-13, 6, 34, -4, -20, -14, 31, 14, -9,
					-- layer=2 filter=63 channel=20
					-8, 9, -7, -6, 0, 9, 9, 1, -8,
					-- layer=2 filter=63 channel=21
					5, -5, 2, 9, 18, 15, -13, -2, -1,
					-- layer=2 filter=63 channel=22
					-11, -9, 0, -4, -10, 8, 0, 6, 1,
					-- layer=2 filter=63 channel=23
					-4, -7, 20, 28, -1, 6, -6, -25, -43,
					-- layer=2 filter=63 channel=24
					-19, 2, -9, 20, 34, 25, -26, 3, -4,
					-- layer=2 filter=63 channel=25
					9, 5, 12, 15, 13, 18, -21, 15, 21,
					-- layer=2 filter=63 channel=26
					-5, -3, 8, 1, -10, 10, 6, -5, -8,
					-- layer=2 filter=63 channel=27
					-3, -9, 0, -13, 3, 19, 13, 20, 41,
					-- layer=2 filter=63 channel=28
					-7, 12, 33, 7, -18, -14, -5, -23, 23,
					-- layer=2 filter=63 channel=29
					2, 3, 4, 1, 2, -3, -3, 2, 7,
					-- layer=2 filter=63 channel=30
					-34, -11, -5, -73, 11, 38, -59, -72, -71,
					-- layer=2 filter=63 channel=31
					-32, 11, 31, -3, 30, -16, -17, 18, -22,
					-- layer=2 filter=63 channel=32
					7, 4, 6, 4, -2, 8, 5, 2, 8,
					-- layer=2 filter=63 channel=33
					-7, 5, 0, 16, -13, -6, 31, 1, 54,
					-- layer=2 filter=63 channel=34
					-1, 28, 37, 16, 17, 0, -53, 2, -7,
					-- layer=2 filter=63 channel=35
					-9, 5, 36, -2, -28, -27, 7, -45, -24,
					-- layer=2 filter=63 channel=36
					4, -1, -5, -8, 1, -2, -13, -12, -9,
					-- layer=2 filter=63 channel=37
					20, -3, 12, 12, -3, 8, -3, -5, 5,
					-- layer=2 filter=63 channel=38
					0, -10, 20, 0, -24, -2, 4, 10, 26,
					-- layer=2 filter=63 channel=39
					-24, 17, 15, -44, -1, -28, -8, -25, -62,
					-- layer=2 filter=63 channel=40
					25, -32, -13, -40, 11, 4, 2, -34, -12,
					-- layer=2 filter=63 channel=41
					-7, 0, 7, 0, 7, 4, 11, -5, -5,
					-- layer=2 filter=63 channel=42
					7, 31, 11, -2, 19, 6, 3, -17, -36,
					-- layer=2 filter=63 channel=43
					9, 3, 13, -14, -2, 5, 15, -26, -31,
					-- layer=2 filter=63 channel=44
					7, -8, 10, -4, -6, 8, 3, 10, -3,
					-- layer=2 filter=63 channel=45
					-28, 13, -11, -45, -45, 16, -34, -18, 24,
					-- layer=2 filter=63 channel=46
					-28, 6, 1, -40, 20, 5, 6, 27, 2,
					-- layer=2 filter=63 channel=47
					-15, 54, 27, -3, 4, 0, -11, -20, 3,
					-- layer=2 filter=63 channel=48
					8, 0, -6, 7, 8, -8, -3, 6, -4,
					-- layer=2 filter=63 channel=49
					17, -43, -28, -31, -13, 21, -19, -41, -40,
					-- layer=2 filter=63 channel=50
					-8, 4, 10, 24, 1, 7, -3, -2, 7,
					-- layer=2 filter=63 channel=51
					14, 6, 5, 20, 23, 2, 13, 1, 3,
					-- layer=2 filter=63 channel=52
					-6, -19, 32, 22, 1, 17, 0, -3, 16,
					-- layer=2 filter=63 channel=53
					-74, 19, 14, 15, 35, -6, -4, 6, 28,
					-- layer=2 filter=63 channel=54
					11, 15, 1, 8, 6, 8, 19, 20, 11,
					-- layer=2 filter=63 channel=55
					4, 7, 0, -8, -10, -8, 0, -5, 0,
					-- layer=2 filter=63 channel=56
					12, -3, 10, 7, -9, -1, -10, -5, 1,
					-- layer=2 filter=63 channel=57
					13, 1, 8, 5, 0, -6, 2, 2, -2,
					-- layer=2 filter=63 channel=58
					0, 25, -2, 17, 8, 31, -11, 3, 13,
					-- layer=2 filter=63 channel=59
					-1, 14, 14, -34, -27, -30, -14, 30, 14,
					-- layer=2 filter=63 channel=60
					20, -20, -9, 0, -26, -46, -5, -14, -20,
					-- layer=2 filter=63 channel=61
					-30, -21, -27, -42, -26, -48, -28, -7, -66,
					-- layer=2 filter=63 channel=62
					28, -4, -22, 38, 0, -18, -22, 1, -46,
					-- layer=2 filter=63 channel=63
					-34, -12, -44, -18, -45, -61, -36, -1, -51,
					-- layer=2 filter=63 channel=64
					-14, 4, 14, 10, 13, 29, -29, -17, -27,
					-- layer=2 filter=63 channel=65
					-11, -33, -8, 4, -14, -38, 9, 11, -20,
					-- layer=2 filter=63 channel=66
					0, -17, -23, -27, -32, -22, -32, 20, -4,
					-- layer=2 filter=63 channel=67
					-33, 2, 5, -37, 9, 15, -60, -25, -11,
					-- layer=2 filter=63 channel=68
					-11, -10, -4, -5, -5, 5, 7, 5, 0,
					-- layer=2 filter=63 channel=69
					17, 20, -6, 0, -1, 24, -4, 15, -11,
					-- layer=2 filter=63 channel=70
					-37, -29, 49, -39, -31, 11, 30, -2, 16,
					-- layer=2 filter=63 channel=71
					2, 0, -12, 22, -3, 34, 10, 13, 37,
					-- layer=2 filter=63 channel=72
					-2, 28, 21, 19, -11, -11, 41, 12, 35,
					-- layer=2 filter=63 channel=73
					2, -12, 32, 16, -13, 7, -27, 17, 2,
					-- layer=2 filter=63 channel=74
					-19, 22, 48, -60, 7, 8, -41, -31, -14,
					-- layer=2 filter=63 channel=75
					-11, 1, -43, 24, 18, 15, -28, -16, 12,
					-- layer=2 filter=63 channel=76
					30, 27, -4, 10, -20, -28, -54, 26, -53,
					-- layer=2 filter=63 channel=77
					5, -8, 3, 6, -5, -7, -3, 5, -6,
					-- layer=2 filter=63 channel=78
					22, -6, -5, 30, -4, -5, 1, 10, -4,
					-- layer=2 filter=63 channel=79
					7, -3, -8, 0, 0, 3, -6, 4, 3,
					-- layer=2 filter=63 channel=80
					9, 26, 6, -16, 49, 3, 0, -7, -42,
					-- layer=2 filter=63 channel=81
					0, 0, -5, 5, 11, 9, 11, -4, -8,
					-- layer=2 filter=63 channel=82
					3, -3, 3, -4, 0, 7, 9, -6, -9,
					-- layer=2 filter=63 channel=83
					-12, -10, -13, -17, -8, -3, 17, -4, -7,
					-- layer=2 filter=63 channel=84
					11, 10, -7, -8, 6, -1, 5, -5, 7,
					-- layer=2 filter=63 channel=85
					1, -3, 15, 14, -11, -6, 10, -7, 4,
					-- layer=2 filter=63 channel=86
					9, -9, 21, 10, -12, 0, 2, -10, 15,
					-- layer=2 filter=63 channel=87
					-9, -7, -6, 21, -3, 1, -42, -34, -20,
					-- layer=2 filter=63 channel=88
					-23, 17, -7, -39, -5, -2, -53, -37, 4,
					-- layer=2 filter=63 channel=89
					9, 22, 3, -16, 0, -4, -12, -13, 25,
					-- layer=2 filter=63 channel=90
					-9, -4, -1, -9, 1, 0, 0, 5, -3,
					-- layer=2 filter=63 channel=91
					-16, 18, 17, 21, 4, -3, -18, -48, 23,
					-- layer=2 filter=63 channel=92
					-12, 26, 3, -7, -1, 10, 6, -5, 8,
					-- layer=2 filter=63 channel=93
					-37, -8, -24, 0, 21, -6, 7, 31, -15,
					-- layer=2 filter=63 channel=94
					19, -5, 3, 0, 25, -23, -9, 44, -75,
					-- layer=2 filter=63 channel=95
					-6, -5, -12, -16, -20, -11, -4, 1, -5,
					-- layer=2 filter=63 channel=96
					34, 3, 3, 7, 54, 27, -29, 22, 32,
					-- layer=2 filter=63 channel=97
					-7, 11, -17, -18, 15, 26, -27, 6, 10,
					-- layer=2 filter=63 channel=98
					-9, 46, 35, 32, -18, 0, -1, -11, 20,
					-- layer=2 filter=63 channel=99
					-11, -21, 44, -4, 9, 23, -12, 28, -4,
					-- layer=2 filter=63 channel=100
					-26, -11, -2, -37, 6, -12, 24, -42, -2,
					-- layer=2 filter=63 channel=101
					0, 6, 4, 19, 0, 17, 16, 10, 42,
					-- layer=2 filter=63 channel=102
					51, -8, -7, -8, 5, 1, -26, -48, -28,
					-- layer=2 filter=63 channel=103
					-21, -2, -10, 7, 1, 29, 18, 12, 37,
					-- layer=2 filter=63 channel=104
					-6, -50, -52, -33, 7, 6, -43, -27, -61,
					-- layer=2 filter=63 channel=105
					-9, 23, 12, -4, -25, -42, -50, -2, -24,
					-- layer=2 filter=63 channel=106
					6, 16, 4, 29, 3, 10, -14, 1, 13,
					-- layer=2 filter=63 channel=107
					28, 35, -15, -19, 9, 9, 23, -16, 3,
					-- layer=2 filter=63 channel=108
					24, -33, -7, 7, 0, 20, 2, -6, 30,
					-- layer=2 filter=63 channel=109
					7, 0, -6, 5, 8, 0, 6, -3, -4,
					-- layer=2 filter=63 channel=110
					-29, 29, -19, -9, 5, -14, -55, -23, 5,
					-- layer=2 filter=63 channel=111
					-6, 7, 0, 0, 6, 3, -7, 1, 5,
					-- layer=2 filter=63 channel=112
					6, -8, -8, 6, 18, 0, 26, 16, 3,
					-- layer=2 filter=63 channel=113
					-55, -73, -20, -29, -53, -7, -61, -20, -34,
					-- layer=2 filter=63 channel=114
					-1, -19, 0, 7, -18, 1, 13, -11, 21,
					-- layer=2 filter=63 channel=115
					9, -4, -3, 9, -6, -11, 6, 5, 0,
					-- layer=2 filter=63 channel=116
					4, -22, 0, 4, 7, -1, -43, 1, -6,
					-- layer=2 filter=63 channel=117
					-2, 29, -2, 5, -4, 27, 25, 18, 14,
					-- layer=2 filter=63 channel=118
					26, 26, 16, 45, 27, 32, 15, -17, -20,
					-- layer=2 filter=63 channel=119
					3, -26, -32, -65, -55, -75, -51, -78, -60,
					-- layer=2 filter=63 channel=120
					4, 9, 9, -8, -1, -1, -5, 2, -9,
					-- layer=2 filter=63 channel=121
					8, 0, -4, 1, 7, 0, -4, 0, -6,
					-- layer=2 filter=63 channel=122
					6, 9, -5, 8, 3, -10, 8, 3, 14,
					-- layer=2 filter=63 channel=123
					5, 30, 19, 22, -34, -5, 17, -2, -5,
					-- layer=2 filter=63 channel=124
					23, 13, -11, -15, -28, -23, -10, -4, -22,
					-- layer=2 filter=63 channel=125
					-8, -5, -1, -4, -4, 3, -2, 6, -2,
					-- layer=2 filter=63 channel=126
					2, 9, -22, -81, 22, -24, -61, 0, -13,
					-- layer=2 filter=63 channel=127
					12, -15, 12, -16, -2, -24, -10, -12, 13,
					-- layer=2 filter=64 channel=0
					-14, -30, -16, -25, -14, -56, -34, -57, -36,
					-- layer=2 filter=64 channel=1
					-43, -30, 28, -10, 3, -25, 17, -6, 37,
					-- layer=2 filter=64 channel=2
					-7, -4, 1, -1, -11, 1, 5, 1, 1,
					-- layer=2 filter=64 channel=3
					-31, -35, -52, -31, -44, -1, -15, -27, -22,
					-- layer=2 filter=64 channel=4
					-3, -34, -40, -9, -43, -13, -28, -18, -16,
					-- layer=2 filter=64 channel=5
					-1, -30, -18, -19, -14, -36, -2, -11, -15,
					-- layer=2 filter=64 channel=6
					-44, -63, 4, -8, 8, -19, -12, -6, 13,
					-- layer=2 filter=64 channel=7
					-45, 2, -57, -65, -14, -36, -14, 2, 46,
					-- layer=2 filter=64 channel=8
					3, 4, -2, 4, -9, -4, -1, 1, -5,
					-- layer=2 filter=64 channel=9
					-9, -46, -28, -1, -15, -27, 5, -19, -24,
					-- layer=2 filter=64 channel=10
					-20, -50, -17, -37, -14, -28, -20, -36, -21,
					-- layer=2 filter=64 channel=11
					-8, -17, -25, 2, 2, -4, -7, -5, -26,
					-- layer=2 filter=64 channel=12
					-66, -34, -9, -27, -3, -67, 19, -2, 78,
					-- layer=2 filter=64 channel=13
					3, -11, 0, -6, 0, -8, -5, 0, -1,
					-- layer=2 filter=64 channel=14
					-36, -4, 3, -8, 3, -28, -1, 5, 27,
					-- layer=2 filter=64 channel=15
					-16, -34, 2, 35, -41, 45, 16, 15, -28,
					-- layer=2 filter=64 channel=16
					26, 23, 38, -81, -36, 52, -40, -69, 7,
					-- layer=2 filter=64 channel=17
					-9, 5, 1, 2, -3, 10, -5, 0, -6,
					-- layer=2 filter=64 channel=18
					-13, -43, -53, -6, -76, 8, 3, -11, -17,
					-- layer=2 filter=64 channel=19
					-11, 4, 35, 8, 10, -1, 25, -4, 39,
					-- layer=2 filter=64 channel=20
					9, -7, 6, 8, 1, -5, -3, -3, 4,
					-- layer=2 filter=64 channel=21
					-7, -2, -13, -26, -21, -4, -16, -28, -3,
					-- layer=2 filter=64 channel=22
					5, 7, -5, 1, 2, -8, -3, 5, -4,
					-- layer=2 filter=64 channel=23
					-16, -16, -41, -21, 15, 1, -24, 16, 43,
					-- layer=2 filter=64 channel=24
					-27, -23, -31, -40, -32, -58, -15, -37, -55,
					-- layer=2 filter=64 channel=25
					-43, -26, -28, -36, -40, -23, -46, -12, -44,
					-- layer=2 filter=64 channel=26
					-1, 0, 1, 6, -3, -3, 3, -6, 10,
					-- layer=2 filter=64 channel=27
					19, 20, 17, 29, 10, -6, 3, 12, -18,
					-- layer=2 filter=64 channel=28
					25, 10, -1, -2, -21, 2, -42, 17, -19,
					-- layer=2 filter=64 channel=29
					-11, 3, -11, -6, 8, -7, 2, 4, -6,
					-- layer=2 filter=64 channel=30
					-27, -31, -15, 31, 29, -3, 4, -16, -5,
					-- layer=2 filter=64 channel=31
					44, -23, 42, -63, -49, -39, -73, 3, -7,
					-- layer=2 filter=64 channel=32
					-2, -4, 8, -11, -5, 1, 6, -4, 7,
					-- layer=2 filter=64 channel=33
					-21, -33, -30, -28, -17, -19, -11, -52, -22,
					-- layer=2 filter=64 channel=34
					-26, 0, -33, 70, -8, 14, 42, -23, 5,
					-- layer=2 filter=64 channel=35
					-11, -5, -16, 11, 2, 46, -61, -9, 15,
					-- layer=2 filter=64 channel=36
					2, 3, -9, 4, 9, 0, 6, -5, -3,
					-- layer=2 filter=64 channel=37
					-5, -11, 7, 10, 2, -19, -5, -13, -33,
					-- layer=2 filter=64 channel=38
					4, -13, 17, 20, 11, -2, 9, -18, -32,
					-- layer=2 filter=64 channel=39
					-27, 19, -51, -45, 25, 0, -3, 4, 49,
					-- layer=2 filter=64 channel=40
					-3, 20, -45, 9, -47, 52, 46, 21, -23,
					-- layer=2 filter=64 channel=41
					-7, -7, 3, -3, -11, -3, -7, -9, -8,
					-- layer=2 filter=64 channel=42
					-17, -13, -80, -41, -45, -17, -4, 5, 52,
					-- layer=2 filter=64 channel=43
					7, 0, -24, -15, -18, 16, 3, -39, -46,
					-- layer=2 filter=64 channel=44
					3, 3, -6, 8, -4, 0, 11, -6, -2,
					-- layer=2 filter=64 channel=45
					14, 11, 12, 20, 2, -21, 4, -35, -43,
					-- layer=2 filter=64 channel=46
					-8, -21, -6, -7, -15, -8, -23, -10, -36,
					-- layer=2 filter=64 channel=47
					-3, -21, -29, -44, -31, -20, -78, -30, -73,
					-- layer=2 filter=64 channel=48
					-6, 0, -4, -2, -7, -9, -11, 8, 3,
					-- layer=2 filter=64 channel=49
					-40, -34, -32, 7, -99, 21, 0, -20, -16,
					-- layer=2 filter=64 channel=50
					-1, -9, 1, -2, -17, -2, -1, -17, -3,
					-- layer=2 filter=64 channel=51
					12, -17, -25, -2, 2, -14, -32, -13, -27,
					-- layer=2 filter=64 channel=52
					-10, -20, -42, 36, -8, 14, 0, -25, -21,
					-- layer=2 filter=64 channel=53
					-10, -16, 30, -19, 13, -18, -55, 7, -2,
					-- layer=2 filter=64 channel=54
					-19, -32, -2, -20, -34, -37, -38, -31, 16,
					-- layer=2 filter=64 channel=55
					8, -7, -6, -7, -3, -1, -9, 0, -6,
					-- layer=2 filter=64 channel=56
					-5, -4, -18, -20, 9, -19, -26, -8, -18,
					-- layer=2 filter=64 channel=57
					-9, 3, 6, 1, -10, -4, 1, -5, -7,
					-- layer=2 filter=64 channel=58
					-29, -18, 2, -20, 23, -61, 13, 10, 69,
					-- layer=2 filter=64 channel=59
					-30, 12, 19, -2, 21, -8, 11, -4, 39,
					-- layer=2 filter=64 channel=60
					25, 10, 59, 21, 23, -8, 6, 9, 96,
					-- layer=2 filter=64 channel=61
					28, 21, -9, 9, 14, 23, -5, -26, 5,
					-- layer=2 filter=64 channel=62
					-57, -47, -24, 13, 0, -17, -11, -4, 11,
					-- layer=2 filter=64 channel=63
					-63, 4, -51, -1, -11, 0, -25, -34, 4,
					-- layer=2 filter=64 channel=64
					-33, -28, -52, -20, -7, -17, 21, 20, 65,
					-- layer=2 filter=64 channel=65
					-35, -24, -6, -4, -7, -42, -25, -36, 4,
					-- layer=2 filter=64 channel=66
					-6, 51, 7, 25, -12, -8, 23, -31, 3,
					-- layer=2 filter=64 channel=67
					-1, 7, -12, 4, -16, 20, 6, 12, 7,
					-- layer=2 filter=64 channel=68
					-11, -2, -5, -5, 0, 4, 6, -9, -4,
					-- layer=2 filter=64 channel=69
					-85, -47, -55, -50, -52, -17, -18, -15, 58,
					-- layer=2 filter=64 channel=70
					0, -4, -7, 6, -10, -12, -8, -2, 5,
					-- layer=2 filter=64 channel=71
					21, 33, 18, 31, 14, 13, 20, 11, 5,
					-- layer=2 filter=64 channel=72
					-53, 5, -12, -34, -33, -11, -3, 3, -18,
					-- layer=2 filter=64 channel=73
					64, 53, 37, -35, 24, -2, -70, -33, -11,
					-- layer=2 filter=64 channel=74
					-18, -14, -58, -2, -17, 0, -15, -31, 28,
					-- layer=2 filter=64 channel=75
					-49, -33, 18, -20, -29, -47, 18, 65, 66,
					-- layer=2 filter=64 channel=76
					1, -28, -16, -18, 20, 28, -54, 48, 25,
					-- layer=2 filter=64 channel=77
					-9, -9, 6, -5, -4, 6, 5, 2, -7,
					-- layer=2 filter=64 channel=78
					-48, -47, -51, -7, -14, -19, -25, 0, 2,
					-- layer=2 filter=64 channel=79
					-6, 0, 0, 10, 6, 6, 7, 3, 2,
					-- layer=2 filter=64 channel=80
					-10, -14, -31, -9, -32, 14, 13, 16, 23,
					-- layer=2 filter=64 channel=81
					7, -3, -7, -14, -13, -4, -11, 0, 4,
					-- layer=2 filter=64 channel=82
					-10, 5, -3, -5, -4, -6, 6, 0, 10,
					-- layer=2 filter=64 channel=83
					-21, -15, 20, 39, -25, -9, 38, -2, 11,
					-- layer=2 filter=64 channel=84
					3, 4, -9, -6, -6, -7, 7, -8, 0,
					-- layer=2 filter=64 channel=85
					-7, 1, 4, 6, -10, 6, 1, -4, -3,
					-- layer=2 filter=64 channel=86
					5, 6, -5, 0, -1, 8, -7, -1, -2,
					-- layer=2 filter=64 channel=87
					-35, -19, -65, 24, -43, 42, -4, 31, -28,
					-- layer=2 filter=64 channel=88
					-60, -38, -79, 14, 4, -11, 25, -45, -32,
					-- layer=2 filter=64 channel=89
					-51, -31, 9, -27, -1, -35, 21, 49, 82,
					-- layer=2 filter=64 channel=90
					-1, 11, -11, -6, -6, -6, -10, 0, 3,
					-- layer=2 filter=64 channel=91
					-38, -24, 28, -46, -1, -35, -5, 27, 101,
					-- layer=2 filter=64 channel=92
					-22, -25, 0, -42, -6, -19, 10, 6, 44,
					-- layer=2 filter=64 channel=93
					-88, -51, 50, 70, -28, -9, 2, 19, 53,
					-- layer=2 filter=64 channel=94
					-36, -10, 0, -13, 32, -17, -24, -35, 31,
					-- layer=2 filter=64 channel=95
					-19, -5, -10, 4, 9, -5, -4, -6, -17,
					-- layer=2 filter=64 channel=96
					19, 3, 23, 6, -2, 26, -56, 15, 36,
					-- layer=2 filter=64 channel=97
					-15, -35, -28, -53, -43, -23, -18, -7, 0,
					-- layer=2 filter=64 channel=98
					18, 15, -30, -15, 2, 17, -8, 8, -25,
					-- layer=2 filter=64 channel=99
					35, 22, 40, 19, 40, 44, 24, 11, 61,
					-- layer=2 filter=64 channel=100
					-10, -4, -3, 17, -5, -35, 19, -8, 48,
					-- layer=2 filter=64 channel=101
					19, 50, 7, 14, 9, -20, -2, 24, 20,
					-- layer=2 filter=64 channel=102
					14, -19, 47, -6, -32, 17, -16, -32, 33,
					-- layer=2 filter=64 channel=103
					15, -3, 4, -29, -9, -5, 45, 36, 70,
					-- layer=2 filter=64 channel=104
					-10, -31, 0, 28, -47, -6, -11, -22, -22,
					-- layer=2 filter=64 channel=105
					38, 14, -4, -44, 50, 42, 50, -10, 70,
					-- layer=2 filter=64 channel=106
					17, -2, -10, -51, -16, -69, -50, 7, 14,
					-- layer=2 filter=64 channel=107
					58, 2, 14, -14, -35, -10, -37, -32, 11,
					-- layer=2 filter=64 channel=108
					3, 4, 15, 39, 0, -1, 38, 10, 4,
					-- layer=2 filter=64 channel=109
					0, 6, -5, -8, 4, -14, -2, -9, -10,
					-- layer=2 filter=64 channel=110
					3, 18, -5, 22, -17, 46, 14, 21, 54,
					-- layer=2 filter=64 channel=111
					6, 7, 7, -7, -6, -6, 0, -7, 8,
					-- layer=2 filter=64 channel=112
					34, 8, 9, -11, 5, -13, -18, -23, 4,
					-- layer=2 filter=64 channel=113
					-8, 35, -38, 24, -22, 0, 0, -27, 4,
					-- layer=2 filter=64 channel=114
					9, 12, -3, 13, 0, 2, 2, 2, 1,
					-- layer=2 filter=64 channel=115
					-8, -9, -5, 9, -4, -6, 5, -9, -1,
					-- layer=2 filter=64 channel=116
					-44, -34, -21, 33, -90, 35, 1, 12, -37,
					-- layer=2 filter=64 channel=117
					0, 31, 15, -47, -8, 34, -36, -53, 35,
					-- layer=2 filter=64 channel=118
					0, -13, -63, -4, -7, 10, -19, -47, -31,
					-- layer=2 filter=64 channel=119
					28, -34, -25, -15, -21, -19, -43, -57, -38,
					-- layer=2 filter=64 channel=120
					-8, -3, -8, -2, -6, -4, 0, 0, 5,
					-- layer=2 filter=64 channel=121
					7, -3, 1, -7, 0, -2, 6, 0, -2,
					-- layer=2 filter=64 channel=122
					0, 2, 7, -11, 0, 2, -6, -2, -8,
					-- layer=2 filter=64 channel=123
					-40, 7, -9, 2, -2, -21, -17, -21, 1,
					-- layer=2 filter=64 channel=124
					-4, 0, -7, -88, -29, 18, -41, -25, 32,
					-- layer=2 filter=64 channel=125
					5, -7, 4, 3, -7, -4, -3, 8, 1,
					-- layer=2 filter=64 channel=126
					-7, 27, -20, 12, 6, -9, 13, 0, -26,
					-- layer=2 filter=64 channel=127
					-39, -34, 0, 21, 5, -15, -3, -38, -34,
					-- layer=2 filter=65 channel=0
					-6, -6, -7, -5, -8, 8, -8, 3, 2,
					-- layer=2 filter=65 channel=1
					4, -3, 0, 2, -8, -2, 0, -12, 3,
					-- layer=2 filter=65 channel=2
					0, 6, -12, 8, -11, -6, -1, -8, 0,
					-- layer=2 filter=65 channel=3
					5, -8, 0, 3, -9, -9, 0, -13, 8,
					-- layer=2 filter=65 channel=4
					7, -3, -2, 0, -6, 3, -2, -4, -6,
					-- layer=2 filter=65 channel=5
					-9, 8, 8, -10, 3, 3, -7, 7, -6,
					-- layer=2 filter=65 channel=6
					4, 4, 0, -3, 7, -3, 0, 5, 3,
					-- layer=2 filter=65 channel=7
					3, -10, -11, 0, -11, 7, -12, -5, 0,
					-- layer=2 filter=65 channel=8
					7, 3, 3, -5, -1, 0, 4, -3, -7,
					-- layer=2 filter=65 channel=9
					2, -6, -9, 4, -5, -2, 8, 1, -3,
					-- layer=2 filter=65 channel=10
					-9, -1, 4, 8, 0, 3, 0, 0, -5,
					-- layer=2 filter=65 channel=11
					-8, -4, -10, 5, 0, -5, 9, -10, -10,
					-- layer=2 filter=65 channel=12
					7, -9, -13, 1, 7, -11, -4, 0, -7,
					-- layer=2 filter=65 channel=13
					-10, -8, -7, 1, 0, -10, -3, -3, -9,
					-- layer=2 filter=65 channel=14
					-4, 7, 3, -11, -8, 0, -7, -6, 0,
					-- layer=2 filter=65 channel=15
					7, -5, 0, 2, -8, -7, 1, -7, -7,
					-- layer=2 filter=65 channel=16
					-6, -5, 7, -2, 0, 8, 3, 2, 6,
					-- layer=2 filter=65 channel=17
					-11, 0, 0, -6, 1, 9, 9, -2, 0,
					-- layer=2 filter=65 channel=18
					8, 3, -2, -2, 0, -11, -6, -7, 0,
					-- layer=2 filter=65 channel=19
					1, -14, 1, 1, -3, 0, -6, -2, -1,
					-- layer=2 filter=65 channel=20
					-6, 2, 5, 5, 4, -3, -6, 1, 3,
					-- layer=2 filter=65 channel=21
					-6, 1, 7, 0, 6, 0, 1, -8, -9,
					-- layer=2 filter=65 channel=22
					-4, 3, -3, 2, -2, 10, 6, -2, -4,
					-- layer=2 filter=65 channel=23
					-4, -3, -10, -7, -15, -8, 6, -4, 0,
					-- layer=2 filter=65 channel=24
					-7, -8, -1, 6, 4, -11, -5, 7, -4,
					-- layer=2 filter=65 channel=25
					-5, 10, 0, 3, 4, -10, -9, 4, 5,
					-- layer=2 filter=65 channel=26
					9, 1, 9, 9, 3, 3, -3, 5, -7,
					-- layer=2 filter=65 channel=27
					6, 3, -3, -6, -11, -7, 5, -11, 1,
					-- layer=2 filter=65 channel=28
					7, -3, -5, 2, 1, -13, -9, -8, -11,
					-- layer=2 filter=65 channel=29
					3, 0, -9, 6, -4, 1, 7, -12, 3,
					-- layer=2 filter=65 channel=30
					-9, -4, -8, 7, 1, -10, 0, -9, 2,
					-- layer=2 filter=65 channel=31
					-10, -2, 0, -8, 0, -11, -8, -3, -8,
					-- layer=2 filter=65 channel=32
					-1, -11, -7, 5, 2, -1, -5, -2, 2,
					-- layer=2 filter=65 channel=33
					0, -10, 6, -6, 5, 5, 2, -2, -4,
					-- layer=2 filter=65 channel=34
					-10, 7, 3, 1, -7, 3, -11, -6, 0,
					-- layer=2 filter=65 channel=35
					4, -8, 4, -13, -7, 1, 2, 4, -10,
					-- layer=2 filter=65 channel=36
					-3, -12, -8, -4, 5, -8, -10, -4, -12,
					-- layer=2 filter=65 channel=37
					-14, -12, -3, 9, 7, 2, -5, -4, -8,
					-- layer=2 filter=65 channel=38
					-8, -1, -11, -6, -1, 8, -1, 0, 0,
					-- layer=2 filter=65 channel=39
					-11, -3, 4, 0, 3, -4, 5, 1, 3,
					-- layer=2 filter=65 channel=40
					-1, -13, 5, -11, 0, 3, -8, 1, -6,
					-- layer=2 filter=65 channel=41
					-3, -11, -6, -7, -9, -7, 11, 6, 0,
					-- layer=2 filter=65 channel=42
					-10, 4, 6, 5, -3, 3, -11, 0, -11,
					-- layer=2 filter=65 channel=43
					-6, -1, -4, -11, -12, -2, 8, -7, -3,
					-- layer=2 filter=65 channel=44
					7, -6, -9, -9, 4, -4, -11, -7, 6,
					-- layer=2 filter=65 channel=45
					3, -3, 7, 8, 1, 3, -5, 4, 1,
					-- layer=2 filter=65 channel=46
					-4, 7, 3, -12, 1, -2, 7, -13, -12,
					-- layer=2 filter=65 channel=47
					-1, 8, -7, -3, 1, 3, 7, 0, -3,
					-- layer=2 filter=65 channel=48
					7, 8, 3, -1, -1, 7, -7, 5, 6,
					-- layer=2 filter=65 channel=49
					2, 2, -5, 0, -10, -3, 1, 7, -5,
					-- layer=2 filter=65 channel=50
					-10, 5, 9, 7, 9, -1, -2, 3, 0,
					-- layer=2 filter=65 channel=51
					-10, 4, 2, 4, -12, -10, -1, 6, -7,
					-- layer=2 filter=65 channel=52
					-3, 5, -1, -11, -6, -1, 5, -6, -1,
					-- layer=2 filter=65 channel=53
					-3, -4, -3, 6, -10, -7, -3, -6, 5,
					-- layer=2 filter=65 channel=54
					1, -5, -8, -8, -12, -6, -2, -11, -8,
					-- layer=2 filter=65 channel=55
					-9, 5, -2, 0, 7, 5, 0, -4, -11,
					-- layer=2 filter=65 channel=56
					-4, -6, -12, -5, -3, -3, 7, -6, -4,
					-- layer=2 filter=65 channel=57
					-8, 0, 9, 4, 0, 0, 3, 5, 2,
					-- layer=2 filter=65 channel=58
					4, 7, -7, 0, 6, -8, -3, -16, 6,
					-- layer=2 filter=65 channel=59
					-9, -11, -1, 1, -6, -1, -9, 3, 0,
					-- layer=2 filter=65 channel=60
					-9, -9, -3, -4, -12, 3, -7, -10, 4,
					-- layer=2 filter=65 channel=61
					4, 1, -8, -8, 6, -9, 0, 9, -16,
					-- layer=2 filter=65 channel=62
					-1, -7, -14, 4, -10, 1, -13, 1, 4,
					-- layer=2 filter=65 channel=63
					0, 7, -10, -5, -10, -6, 0, -2, 5,
					-- layer=2 filter=65 channel=64
					5, -9, -2, -12, -2, 3, -8, 0, -10,
					-- layer=2 filter=65 channel=65
					-2, 3, -1, -2, -6, -7, 4, 6, -8,
					-- layer=2 filter=65 channel=66
					2, -2, 2, 7, -11, 4, -12, 1, 3,
					-- layer=2 filter=65 channel=67
					-4, -11, -3, -1, 6, -8, -10, 1, -8,
					-- layer=2 filter=65 channel=68
					6, -6, 8, -12, 6, -7, -3, 2, 2,
					-- layer=2 filter=65 channel=69
					3, 0, -2, -14, -13, -7, -13, -12, 4,
					-- layer=2 filter=65 channel=70
					1, 2, -7, -4, 3, -14, 2, 9, 1,
					-- layer=2 filter=65 channel=71
					-6, 0, -11, -10, -1, -1, 4, -6, -10,
					-- layer=2 filter=65 channel=72
					-5, -4, -5, -10, -11, -7, 0, -14, -4,
					-- layer=2 filter=65 channel=73
					3, -16, 3, 3, -9, 7, 6, -1, 6,
					-- layer=2 filter=65 channel=74
					-1, -10, -1, -3, -2, 4, 0, -6, -1,
					-- layer=2 filter=65 channel=75
					-9, 2, -11, -8, -11, 7, -12, -6, 2,
					-- layer=2 filter=65 channel=76
					1, -5, 0, -10, -10, 3, -5, -3, -2,
					-- layer=2 filter=65 channel=77
					8, -4, -5, 0, -10, 1, 1, 0, 7,
					-- layer=2 filter=65 channel=78
					-8, 7, 0, -8, 0, -11, 1, -12, -4,
					-- layer=2 filter=65 channel=79
					1, 8, -9, 3, -5, -6, 3, 4, -2,
					-- layer=2 filter=65 channel=80
					-7, 5, 0, 2, 0, -9, -7, -1, 7,
					-- layer=2 filter=65 channel=81
					-9, -8, 6, -2, -2, -7, -6, -5, 0,
					-- layer=2 filter=65 channel=82
					-3, 1, 4, -2, -8, -1, -2, -6, -5,
					-- layer=2 filter=65 channel=83
					5, -1, -5, 0, -2, -5, 1, -2, -6,
					-- layer=2 filter=65 channel=84
					7, -7, -2, -8, 7, -10, 7, -1, 5,
					-- layer=2 filter=65 channel=85
					-8, 2, 8, 3, 5, -6, 7, 2, -11,
					-- layer=2 filter=65 channel=86
					-6, 0, 4, -6, 9, 6, 9, 8, 7,
					-- layer=2 filter=65 channel=87
					-5, 0, 3, 0, 4, -3, -6, -4, -10,
					-- layer=2 filter=65 channel=88
					7, 6, -8, 0, -1, -1, -1, 1, -5,
					-- layer=2 filter=65 channel=89
					-10, -12, -1, 4, 4, -10, -4, 2, 0,
					-- layer=2 filter=65 channel=90
					7, 7, 4, 0, -10, -8, 4, 7, -5,
					-- layer=2 filter=65 channel=91
					-12, -2, -5, 0, -12, -14, -7, -16, -5,
					-- layer=2 filter=65 channel=92
					-6, -1, -13, -6, -2, 1, -7, -15, -6,
					-- layer=2 filter=65 channel=93
					5, 0, -2, -10, 2, -6, 8, 5, 5,
					-- layer=2 filter=65 channel=94
					-12, -4, 3, 7, 1, -2, -5, 3, -8,
					-- layer=2 filter=65 channel=95
					-1, 0, 0, -12, 3, -10, -10, -8, 3,
					-- layer=2 filter=65 channel=96
					-2, 0, -3, -10, -9, -3, -1, -1, -3,
					-- layer=2 filter=65 channel=97
					2, -12, 0, -8, 0, 6, -1, -10, 5,
					-- layer=2 filter=65 channel=98
					-11, -4, -10, 0, 4, -12, 0, -8, 7,
					-- layer=2 filter=65 channel=99
					4, -4, -1, -9, 7, -4, -7, -4, 0,
					-- layer=2 filter=65 channel=100
					5, -2, -10, 1, -6, -4, -7, -13, 0,
					-- layer=2 filter=65 channel=101
					-3, 3, 9, -9, -4, 2, -6, 7, 0,
					-- layer=2 filter=65 channel=102
					0, 3, -10, -11, -6, 5, -12, 0, 4,
					-- layer=2 filter=65 channel=103
					-11, 3, 4, -5, -1, 6, 7, 1, 5,
					-- layer=2 filter=65 channel=104
					-7, -3, 7, -5, 4, -10, 2, -6, -10,
					-- layer=2 filter=65 channel=105
					2, -12, -9, 0, 7, -8, -4, -4, 0,
					-- layer=2 filter=65 channel=106
					-5, 8, 9, 2, -2, -5, -9, 3, -1,
					-- layer=2 filter=65 channel=107
					2, -2, -8, 0, 0, 0, -4, -3, 2,
					-- layer=2 filter=65 channel=108
					8, 0, -4, 8, -2, 1, -10, 0, 1,
					-- layer=2 filter=65 channel=109
					3, 7, -6, -5, -10, 1, 5, -3, -10,
					-- layer=2 filter=65 channel=110
					-13, 2, 5, -4, -11, 0, -12, 6, -5,
					-- layer=2 filter=65 channel=111
					7, -5, -4, 8, -9, 6, 1, 11, 1,
					-- layer=2 filter=65 channel=112
					-2, 5, -6, 3, 0, -12, -6, 5, -9,
					-- layer=2 filter=65 channel=113
					-1, 1, 1, 6, 7, 0, 6, 5, -9,
					-- layer=2 filter=65 channel=114
					-2, -2, -9, -9, -1, -7, -2, 8, -4,
					-- layer=2 filter=65 channel=115
					2, 5, 5, 10, 3, 9, 5, 0, 8,
					-- layer=2 filter=65 channel=116
					-2, -11, 7, 0, -10, 0, 3, -1, 2,
					-- layer=2 filter=65 channel=117
					-11, -14, -15, -4, 4, 6, -5, 6, -14,
					-- layer=2 filter=65 channel=118
					4, -8, -3, 2, 6, -8, -10, 1, 6,
					-- layer=2 filter=65 channel=119
					-6, -5, -10, -9, 2, -1, 3, -9, -3,
					-- layer=2 filter=65 channel=120
					-6, 4, 9, -7, -9, -4, 9, 1, 2,
					-- layer=2 filter=65 channel=121
					0, 11, -7, -1, 7, -1, 0, -3, 0,
					-- layer=2 filter=65 channel=122
					-6, 8, 2, 6, 5, -2, 3, 7, 8,
					-- layer=2 filter=65 channel=123
					-10, -11, -16, -1, -9, -13, -12, 4, 2,
					-- layer=2 filter=65 channel=124
					-6, -6, -5, 3, 1, 0, -3, -5, 6,
					-- layer=2 filter=65 channel=125
					4, 9, -4, 6, 8, -5, -6, 7, 0,
					-- layer=2 filter=65 channel=126
					0, -9, 0, 0, 6, -9, -7, -12, 3,
					-- layer=2 filter=65 channel=127
					-1, 0, -5, -6, -7, -10, -8, -4, -14,
					-- layer=2 filter=66 channel=0
					-9, -9, -14, -20, -26, -37, -2, 4, 0,
					-- layer=2 filter=66 channel=1
					-1, 2, -2, 6, -1, 21, -6, 31, -7,
					-- layer=2 filter=66 channel=2
					2, 7, -9, -3, 0, -7, -9, 9, 2,
					-- layer=2 filter=66 channel=3
					2, -10, -7, -39, -10, -8, -20, 31, 54,
					-- layer=2 filter=66 channel=4
					-15, 2, 59, -13, 12, 7, -2, 3, 0,
					-- layer=2 filter=66 channel=5
					-28, -46, -35, -18, -50, 3, -12, -24, -6,
					-- layer=2 filter=66 channel=6
					22, -39, -23, -14, -103, -52, 0, -69, -47,
					-- layer=2 filter=66 channel=7
					45, -7, 42, 40, 48, 41, 28, 39, 17,
					-- layer=2 filter=66 channel=8
					10, 7, 5, 10, 8, 2, -1, 7, 2,
					-- layer=2 filter=66 channel=9
					-8, -8, 6, -20, -27, -42, -8, -36, -8,
					-- layer=2 filter=66 channel=10
					9, 30, -15, -13, -6, -8, 19, 4, 3,
					-- layer=2 filter=66 channel=11
					-32, -69, -45, -17, -50, -17, -19, -31, -4,
					-- layer=2 filter=66 channel=12
					12, 8, 21, 24, -7, 22, -44, -13, -1,
					-- layer=2 filter=66 channel=13
					8, 0, -8, -7, 3, -1, -4, -11, 10,
					-- layer=2 filter=66 channel=14
					12, -19, 1, 27, -9, 39, -17, 19, 14,
					-- layer=2 filter=66 channel=15
					7, 7, -29, 19, -7, -36, 7, 33, 35,
					-- layer=2 filter=66 channel=16
					-24, -19, -47, 7, 0, -17, 18, 15, 3,
					-- layer=2 filter=66 channel=17
					5, 4, 9, 7, 2, 0, -8, -4, -10,
					-- layer=2 filter=66 channel=18
					-64, 19, 5, 22, 27, -6, -13, 4, 9,
					-- layer=2 filter=66 channel=19
					7, -19, -30, -2, 7, -5, -15, -14, -50,
					-- layer=2 filter=66 channel=20
					8, -1, 0, 0, 1, 12, 2, -6, -6,
					-- layer=2 filter=66 channel=21
					0, 12, 11, 14, 8, 15, -8, 8, 20,
					-- layer=2 filter=66 channel=22
					-4, 2, 2, 7, 3, 3, 0, 4, -7,
					-- layer=2 filter=66 channel=23
					-24, -27, 2, -17, 40, 7, 22, -6, -2,
					-- layer=2 filter=66 channel=24
					-18, -24, -16, -1, 15, 14, 6, 56, 77,
					-- layer=2 filter=66 channel=25
					-8, -26, -11, -14, 0, 41, 17, 24, 57,
					-- layer=2 filter=66 channel=26
					9, -5, 7, -5, -4, 0, -4, -3, -3,
					-- layer=2 filter=66 channel=27
					8, -55, -18, 6, -8, -2, -19, -24, -25,
					-- layer=2 filter=66 channel=28
					-41, -4, -9, -19, 0, 20, 41, 16, 19,
					-- layer=2 filter=66 channel=29
					-2, 1, -8, -1, 2, 5, -7, -2, -3,
					-- layer=2 filter=66 channel=30
					-1, -22, -13, -23, 15, -27, -18, 5, -20,
					-- layer=2 filter=66 channel=31
					-39, 14, 1, -52, 21, -21, 46, -24, -59,
					-- layer=2 filter=66 channel=32
					-4, 3, 0, 0, 9, -11, 3, 4, 7,
					-- layer=2 filter=66 channel=33
					22, 4, 53, 5, -2, 47, -28, 12, 0,
					-- layer=2 filter=66 channel=34
					-32, -38, -23, -31, 7, 17, -10, -13, -7,
					-- layer=2 filter=66 channel=35
					-22, -15, -43, -1, 17, 40, 44, 18, 13,
					-- layer=2 filter=66 channel=36
					-10, -7, 8, -2, 0, -6, -10, 1, -4,
					-- layer=2 filter=66 channel=37
					-43, -72, -64, -43, -49, -42, -18, -33, -20,
					-- layer=2 filter=66 channel=38
					4, -37, -63, -5, -5, 14, -45, -4, 6,
					-- layer=2 filter=66 channel=39
					20, 6, -9, -21, 6, -19, 1, 3, 8,
					-- layer=2 filter=66 channel=40
					-5, 32, -31, -21, 30, 8, -10, 29, 38,
					-- layer=2 filter=66 channel=41
					4, -6, 10, 7, -4, -3, -11, 7, -4,
					-- layer=2 filter=66 channel=42
					-8, 10, 15, 13, 20, -2, 17, 12, 19,
					-- layer=2 filter=66 channel=43
					1, -35, -31, -17, -3, 23, -49, -23, 31,
					-- layer=2 filter=66 channel=44
					10, -3, -2, 8, 3, -4, 10, -6, -8,
					-- layer=2 filter=66 channel=45
					1, -25, -71, 30, 4, 13, -3, -20, 9,
					-- layer=2 filter=66 channel=46
					12, 19, -16, -29, -32, -35, 0, -17, -47,
					-- layer=2 filter=66 channel=47
					-40, 6, 11, 23, 7, 13, 23, 34, 25,
					-- layer=2 filter=66 channel=48
					-8, 10, -6, 6, -10, -4, 2, 0, 5,
					-- layer=2 filter=66 channel=49
					-43, 21, 29, 48, 19, -24, -16, 19, -18,
					-- layer=2 filter=66 channel=50
					10, -5, 16, 8, 7, 8, -7, 11, 0,
					-- layer=2 filter=66 channel=51
					-49, -81, -53, -26, -51, -12, -8, -12, 0,
					-- layer=2 filter=66 channel=52
					-37, -29, -20, -16, -25, -7, -24, -38, -29,
					-- layer=2 filter=66 channel=53
					40, -46, -26, -13, 12, -40, -18, -33, -27,
					-- layer=2 filter=66 channel=54
					-41, -9, -1, 0, 17, 33, 1, 21, 22,
					-- layer=2 filter=66 channel=55
					8, 2, 1, 10, 7, 4, -1, 3, -8,
					-- layer=2 filter=66 channel=56
					-20, -53, -12, -12, -35, -57, -8, -29, 5,
					-- layer=2 filter=66 channel=57
					6, -5, 2, 4, 0, -2, 6, -3, -7,
					-- layer=2 filter=66 channel=58
					39, -4, 4, 25, -26, 16, -51, -14, 10,
					-- layer=2 filter=66 channel=59
					33, -28, 38, -19, -12, 1, -41, -23, -62,
					-- layer=2 filter=66 channel=60
					9, -13, -26, -9, -6, -20, 5, 12, -46,
					-- layer=2 filter=66 channel=61
					12, -56, -40, 14, 22, -47, 9, 25, -37,
					-- layer=2 filter=66 channel=62
					16, -7, 3, -15, -1, -3, -36, -26, -18,
					-- layer=2 filter=66 channel=63
					10, -7, -9, -7, 1, -24, -10, -13, -8,
					-- layer=2 filter=66 channel=64
					-13, 14, 5, -17, 29, -4, 8, 26, 17,
					-- layer=2 filter=66 channel=65
					-6, -59, -23, 10, -53, -57, -20, -27, -89,
					-- layer=2 filter=66 channel=66
					-16, -6, -33, -7, 0, 13, 6, 15, 32,
					-- layer=2 filter=66 channel=67
					21, 41, -22, -37, -50, -6, -7, 4, -19,
					-- layer=2 filter=66 channel=68
					1, 0, 6, 7, 0, 1, -2, 7, -11,
					-- layer=2 filter=66 channel=69
					16, 4, 17, -10, 11, -6, 7, 5, 21,
					-- layer=2 filter=66 channel=70
					-48, -68, -68, -5, 6, 20, 22, 4, 2,
					-- layer=2 filter=66 channel=71
					27, -27, 1, 7, -8, 17, -36, -3, -24,
					-- layer=2 filter=66 channel=72
					-43, -26, 19, -5, -16, 3, 29, -11, 29,
					-- layer=2 filter=66 channel=73
					48, 0, -9, 35, 57, 3, 17, 28, -20,
					-- layer=2 filter=66 channel=74
					41, 19, -7, -23, -22, -20, 4, -6, 0,
					-- layer=2 filter=66 channel=75
					17, -14, 21, 13, -35, 23, -13, 22, 38,
					-- layer=2 filter=66 channel=76
					52, -18, -22, -53, 40, -53, 14, -7, -18,
					-- layer=2 filter=66 channel=77
					2, -2, 2, -1, 10, -9, 2, -8, 2,
					-- layer=2 filter=66 channel=78
					-76, -56, 0, -44, -8, 6, -4, 3, 37,
					-- layer=2 filter=66 channel=79
					1, -7, -7, 9, 11, 6, 5, -6, 0,
					-- layer=2 filter=66 channel=80
					4, 16, 20, -14, 1, -16, -3, 3, -13,
					-- layer=2 filter=66 channel=81
					5, 1, -8, -6, 2, 5, -10, -11, -10,
					-- layer=2 filter=66 channel=82
					0, 7, -7, -6, -5, 3, -3, 0, 8,
					-- layer=2 filter=66 channel=83
					-18, 0, -6, -4, 9, -12, 12, -4, -6,
					-- layer=2 filter=66 channel=84
					5, 2, 10, -7, 0, -12, -9, -3, 0,
					-- layer=2 filter=66 channel=85
					-10, 8, -8, -5, -9, -19, 0, 3, 4,
					-- layer=2 filter=66 channel=86
					-1, 8, 3, 0, -18, -1, 18, 7, 10,
					-- layer=2 filter=66 channel=87
					-16, 15, 24, -4, 38, -2, 38, 0, 53,
					-- layer=2 filter=66 channel=88
					21, -1, -8, -4, 8, -26, -8, 1, 10,
					-- layer=2 filter=66 channel=89
					32, 0, 15, -11, -10, 27, -9, -12, -16,
					-- layer=2 filter=66 channel=90
					-4, 4, 7, 5, -9, -6, -1, 1, 2,
					-- layer=2 filter=66 channel=91
					30, -8, 13, 5, -14, 6, -14, 6, -11,
					-- layer=2 filter=66 channel=92
					10, 0, 11, 7, -14, 28, -39, 0, -7,
					-- layer=2 filter=66 channel=93
					69, 13, 16, -13, -57, -41, -26, -36, -44,
					-- layer=2 filter=66 channel=94
					13, -84, 2, 16, 7, -47, 20, -18, -36,
					-- layer=2 filter=66 channel=95
					-8, 9, -7, -6, 7, -3, -2, 0, -4,
					-- layer=2 filter=66 channel=96
					8, -22, 32, -31, -58, -8, -1, -18, -36,
					-- layer=2 filter=66 channel=97
					-6, 15, 25, -40, -20, 20, -6, 21, 58,
					-- layer=2 filter=66 channel=98
					-33, 24, -15, 14, 12, 9, 44, -1, 19,
					-- layer=2 filter=66 channel=99
					44, -56, 1, -25, -40, -27, 20, -34, -52,
					-- layer=2 filter=66 channel=100
					-23, -16, -26, -1, -14, 12, -1, 21, 10,
					-- layer=2 filter=66 channel=101
					27, -20, -20, 8, -63, -22, -31, -17, -31,
					-- layer=2 filter=66 channel=102
					-12, -14, 6, 0, -47, -33, -32, 0, -37,
					-- layer=2 filter=66 channel=103
					-48, 23, 18, 32, 12, 19, 8, 15, 4,
					-- layer=2 filter=66 channel=104
					-55, -18, 1, 41, -26, -52, -17, -12, -12,
					-- layer=2 filter=66 channel=105
					20, -83, 15, -8, 68, -24, 15, -47, 25,
					-- layer=2 filter=66 channel=106
					45, -18, -11, -3, -25, -1, -6, 26, -1,
					-- layer=2 filter=66 channel=107
					-32, 24, -37, 64, 8, -29, -35, -8, -38,
					-- layer=2 filter=66 channel=108
					-2, 0, -18, 3, -26, -48, -35, 13, -29,
					-- layer=2 filter=66 channel=109
					23, 1, -7, 15, 6, 4, 0, 7, -6,
					-- layer=2 filter=66 channel=110
					-16, -27, -2, -43, 20, 17, 27, 2, 22,
					-- layer=2 filter=66 channel=111
					-5, -4, 5, -3, 1, 8, -6, 5, -6,
					-- layer=2 filter=66 channel=112
					-38, -59, -86, -1, -10, -26, -14, 31, -18,
					-- layer=2 filter=66 channel=113
					-5, -31, -46, 3, 0, -3, 1, -32, -18,
					-- layer=2 filter=66 channel=114
					-5, 3, 4, 3, -5, 11, 5, 2, 11,
					-- layer=2 filter=66 channel=115
					0, -4, 7, 8, -5, 7, -9, 4, -1,
					-- layer=2 filter=66 channel=116
					-22, 24, 6, -15, 0, -2, -11, 8, 40,
					-- layer=2 filter=66 channel=117
					1, -23, -9, 36, -8, 11, 20, 2, 0,
					-- layer=2 filter=66 channel=118
					-2, 3, 6, -41, 0, -9, -24, -9, 23,
					-- layer=2 filter=66 channel=119
					-23, -3, 14, 2, 12, -7, -4, 21, 7,
					-- layer=2 filter=66 channel=120
					3, 7, 5, 0, 0, -3, -5, -10, -2,
					-- layer=2 filter=66 channel=121
					-8, 3, 0, -7, 6, -12, 5, 7, -6,
					-- layer=2 filter=66 channel=122
					8, -3, -8, -5, 7, 6, 12, 15, 3,
					-- layer=2 filter=66 channel=123
					-10, -22, 38, 12, 26, 32, 3, -1, 17,
					-- layer=2 filter=66 channel=124
					12, 37, 58, 0, 41, 30, 34, 3, -7,
					-- layer=2 filter=66 channel=125
					5, 3, -6, 1, -3, 10, 6, 1, 2,
					-- layer=2 filter=66 channel=126
					58, 4, 67, 5, 27, 35, -16, -35, 12,
					-- layer=2 filter=66 channel=127
					-9, -54, 16, -13, -3, 51, -11, -13, 19,
					-- layer=2 filter=67 channel=0
					25, -17, -10, 1, -5, -7, -21, -1, -24,
					-- layer=2 filter=67 channel=1
					-2, -62, -11, 19, -32, -26, -34, 10, 0,
					-- layer=2 filter=67 channel=2
					-7, 4, -8, -2, 2, 4, -2, -5, 3,
					-- layer=2 filter=67 channel=3
					-2, 10, 11, 12, -4, 9, -24, -27, -21,
					-- layer=2 filter=67 channel=4
					9, -2, -11, -95, -33, -17, -33, -29, -63,
					-- layer=2 filter=67 channel=5
					-5, -8, -9, -15, 18, 23, -8, -11, -16,
					-- layer=2 filter=67 channel=6
					45, -14, -12, 27, -24, 17, -7, 1, -6,
					-- layer=2 filter=67 channel=7
					-25, 42, 19, -48, -14, -37, 64, 13, -5,
					-- layer=2 filter=67 channel=8
					3, -3, -3, -6, -5, 0, 9, -6, -8,
					-- layer=2 filter=67 channel=9
					-60, -35, -27, 26, 47, 18, -10, 19, -31,
					-- layer=2 filter=67 channel=10
					3, -16, 1, -14, -39, -6, -43, -26, -28,
					-- layer=2 filter=67 channel=11
					-7, 10, -5, 15, 14, -4, 4, 5, -4,
					-- layer=2 filter=67 channel=12
					-28, -63, -74, 4, -13, -4, -32, -15, -38,
					-- layer=2 filter=67 channel=13
					-9, 6, 7, -5, -11, 7, 3, 6, 4,
					-- layer=2 filter=67 channel=14
					-46, -34, -35, 19, 23, 0, -16, 10, 15,
					-- layer=2 filter=67 channel=15
					25, 14, 32, -11, -22, -7, 54, -20, 69,
					-- layer=2 filter=67 channel=16
					52, 32, 27, 13, 60, -2, 7, -50, -23,
					-- layer=2 filter=67 channel=17
					-6, 10, 0, -7, 5, 6, 4, 5, 9,
					-- layer=2 filter=67 channel=18
					-38, 9, 32, -41, 17, 11, -21, -5, -8,
					-- layer=2 filter=67 channel=19
					10, 8, 28, -5, -24, -11, -13, 50, 31,
					-- layer=2 filter=67 channel=20
					-3, -5, 9, 10, 2, -8, -6, 11, -3,
					-- layer=2 filter=67 channel=21
					-5, 8, -14, 5, -4, -3, -10, 1, 2,
					-- layer=2 filter=67 channel=22
					11, 4, 11, -9, 8, -2, -4, -5, -8,
					-- layer=2 filter=67 channel=23
					14, 8, -33, -47, -42, -47, -2, -27, -26,
					-- layer=2 filter=67 channel=24
					0, -14, -6, 22, 10, 12, -5, -15, 0,
					-- layer=2 filter=67 channel=25
					-24, -6, 3, 22, 7, 1, 22, 8, 7,
					-- layer=2 filter=67 channel=26
					-8, 7, 0, 10, -5, 4, 5, -4, -6,
					-- layer=2 filter=67 channel=27
					6, 13, 12, 3, 29, 11, -19, 17, 25,
					-- layer=2 filter=67 channel=28
					-11, 38, 32, -52, -35, -1, -42, -5, -22,
					-- layer=2 filter=67 channel=29
					-9, 7, -8, 4, 7, -7, 6, 8, 1,
					-- layer=2 filter=67 channel=30
					14, -4, -6, -4, 29, -17, -75, -39, -12,
					-- layer=2 filter=67 channel=31
					21, 54, 0, -28, -32, -40, -24, -8, -27,
					-- layer=2 filter=67 channel=32
					0, -1, -8, 5, 3, 8, -12, -10, 10,
					-- layer=2 filter=67 channel=33
					-2, 60, 18, -31, -42, -66, 20, -2, 5,
					-- layer=2 filter=67 channel=34
					-22, 56, 27, 7, -39, -13, -32, -2, 59,
					-- layer=2 filter=67 channel=35
					-14, 22, 13, -47, -58, -71, -10, -30, -66,
					-- layer=2 filter=67 channel=36
					-1, 7, 4, 0, 4, -1, -2, 3, 7,
					-- layer=2 filter=67 channel=37
					-5, -6, 0, -14, 14, 11, -1, 9, 17,
					-- layer=2 filter=67 channel=38
					4, -15, -28, 21, 30, 35, -21, -3, 11,
					-- layer=2 filter=67 channel=39
					49, 2, 14, -13, 30, 11, -1, -30, -19,
					-- layer=2 filter=67 channel=40
					31, 60, 46, -15, 8, 17, -10, -44, 30,
					-- layer=2 filter=67 channel=41
					-5, 11, 8, 6, -6, -8, -7, 9, -8,
					-- layer=2 filter=67 channel=42
					20, 35, -28, -35, -58, -69, 8, -48, -50,
					-- layer=2 filter=67 channel=43
					-43, 16, 54, -1, 60, 8, -25, -2, -34,
					-- layer=2 filter=67 channel=44
					4, -9, 10, 2, 8, -1, -1, -5, 6,
					-- layer=2 filter=67 channel=45
					23, 33, 3, -5, -31, -5, -5, -14, 14,
					-- layer=2 filter=67 channel=46
					32, -47, -29, -25, -4, 12, -4, -40, -14,
					-- layer=2 filter=67 channel=47
					27, 58, 39, -51, -54, -38, 11, -2, -16,
					-- layer=2 filter=67 channel=48
					-4, 0, -2, -5, 0, 1, -1, 1, 7,
					-- layer=2 filter=67 channel=49
					-23, 7, 11, 2, 12, -7, 16, 31, -22,
					-- layer=2 filter=67 channel=50
					0, 12, 1, -5, 11, 10, -5, -13, -11,
					-- layer=2 filter=67 channel=51
					-5, 0, -11, 13, 10, 9, -2, 7, -10,
					-- layer=2 filter=67 channel=52
					13, 17, 4, 5, 60, -5, 18, -1, 10,
					-- layer=2 filter=67 channel=53
					-12, 26, 5, 39, -25, -56, -19, 27, -7,
					-- layer=2 filter=67 channel=54
					34, 15, 6, -20, -14, -6, 5, -7, -9,
					-- layer=2 filter=67 channel=55
					-13, 10, 5, -6, -2, -5, -9, 8, -9,
					-- layer=2 filter=67 channel=56
					-24, 8, 17, 1, 26, 17, -8, 14, -4,
					-- layer=2 filter=67 channel=57
					0, 3, 3, -6, 3, 5, -3, 4, 2,
					-- layer=2 filter=67 channel=58
					-11, -41, -50, -16, 3, 14, -43, -17, -41,
					-- layer=2 filter=67 channel=59
					31, 19, -38, -1, -5, -16, -40, 9, 20,
					-- layer=2 filter=67 channel=60
					12, -12, 12, -86, -29, 45, -47, 7, 30,
					-- layer=2 filter=67 channel=61
					36, -1, 9, 7, -41, -1, -29, -11, 3,
					-- layer=2 filter=67 channel=62
					1, 19, 14, 0, -33, -1, 0, 34, 8,
					-- layer=2 filter=67 channel=63
					46, 47, 6, -50, -57, -35, -55, -39, -22,
					-- layer=2 filter=67 channel=64
					30, 14, -34, -14, 4, -31, -17, -40, -26,
					-- layer=2 filter=67 channel=65
					32, -25, -20, 25, -26, 50, 13, -36, 5,
					-- layer=2 filter=67 channel=66
					11, 7, -19, 34, -19, -13, -6, 4, -38,
					-- layer=2 filter=67 channel=67
					-1, -15, -20, 18, 27, 37, -12, -13, 24,
					-- layer=2 filter=67 channel=68
					-3, -10, -5, 3, 0, -10, 1, -9, 8,
					-- layer=2 filter=67 channel=69
					60, 19, 5, 23, -4, -29, -13, -12, -67,
					-- layer=2 filter=67 channel=70
					-15, 2, -2, -38, -14, -6, -16, -17, -35,
					-- layer=2 filter=67 channel=71
					-7, 18, -6, 3, 44, 10, 23, 31, 24,
					-- layer=2 filter=67 channel=72
					-44, 0, 17, -66, -39, -32, 5, 6, 40,
					-- layer=2 filter=67 channel=73
					42, 31, 20, 35, -10, -62, 26, 5, -20,
					-- layer=2 filter=67 channel=74
					30, 1, -30, -19, -23, -9, -89, -76, -66,
					-- layer=2 filter=67 channel=75
					5, 5, -42, 18, -6, 30, -29, 0, 6,
					-- layer=2 filter=67 channel=76
					33, 24, 12, 1, -34, -62, -56, 43, -34,
					-- layer=2 filter=67 channel=77
					-5, 0, -8, 2, 3, 2, -6, -5, 2,
					-- layer=2 filter=67 channel=78
					-16, -12, 3, -1, 4, -12, 7, 13, 6,
					-- layer=2 filter=67 channel=79
					-7, -6, 10, 2, 1, -10, 3, 0, 11,
					-- layer=2 filter=67 channel=80
					27, 63, 11, -40, 0, 13, -17, -53, -44,
					-- layer=2 filter=67 channel=81
					-2, -1, 8, 0, 1, 3, 3, -10, -1,
					-- layer=2 filter=67 channel=82
					0, 11, 10, -3, -7, -7, -12, 0, 9,
					-- layer=2 filter=67 channel=83
					-14, 19, -26, -22, 13, 9, -7, 20, -5,
					-- layer=2 filter=67 channel=84
					9, -4, -7, -8, 6, 1, 10, -7, 0,
					-- layer=2 filter=67 channel=85
					-1, 1, -12, -1, 4, -1, 0, -11, 4,
					-- layer=2 filter=67 channel=86
					3, 8, -9, -8, 3, 3, 2, -6, 3,
					-- layer=2 filter=67 channel=87
					-6, -30, 23, -2, -36, 13, -8, -21, 9,
					-- layer=2 filter=67 channel=88
					-8, -14, -51, -35, 6, -49, -107, -88, -65,
					-- layer=2 filter=67 channel=89
					-10, -32, -28, -9, 12, -13, -3, 23, -1,
					-- layer=2 filter=67 channel=90
					-7, 4, -11, 2, 0, 5, 10, 0, 3,
					-- layer=2 filter=67 channel=91
					7, -30, 20, -27, -23, 3, -47, 22, -8,
					-- layer=2 filter=67 channel=92
					-8, -50, -55, -7, -19, -11, -20, -5, -25,
					-- layer=2 filter=67 channel=93
					10, 54, 40, -12, -16, 36, -1, -28, 36,
					-- layer=2 filter=67 channel=94
					42, -11, 0, 33, 0, 5, -4, -9, -31,
					-- layer=2 filter=67 channel=95
					-7, 0, 4, 4, 0, 1, 10, 6, 11,
					-- layer=2 filter=67 channel=96
					3, 6, -6, 29, -12, -5, -18, 1, 0,
					-- layer=2 filter=67 channel=97
					-3, 3, -12, -6, 4, -3, -40, -19, -26,
					-- layer=2 filter=67 channel=98
					24, 45, 35, -56, -59, -38, 16, 29, 7,
					-- layer=2 filter=67 channel=99
					26, 26, -16, -18, -18, 4, 0, 22, 16,
					-- layer=2 filter=67 channel=100
					-38, -15, -16, -35, -9, 38, -52, -57, -37,
					-- layer=2 filter=67 channel=101
					-5, 11, 25, 34, 19, 19, 30, 11, 11,
					-- layer=2 filter=67 channel=102
					-7, -20, 11, 1, 9, -6, -1, -15, 4,
					-- layer=2 filter=67 channel=103
					-38, 3, -57, 1, -32, 8, 6, 30, -29,
					-- layer=2 filter=67 channel=104
					-14, -2, 10, 16, 15, -5, 4, 17, -21,
					-- layer=2 filter=67 channel=105
					-23, 39, 31, -76, 0, -35, 42, 30, -14,
					-- layer=2 filter=67 channel=106
					0, -25, 21, 18, 11, 28, 1, 9, 16,
					-- layer=2 filter=67 channel=107
					3, -3, -36, 16, -41, -4, 87, 1, -3,
					-- layer=2 filter=67 channel=108
					-17, 0, -7, 1, 32, -4, -7, 26, 46,
					-- layer=2 filter=67 channel=109
					-4, -3, -6, 1, -6, 0, 10, 0, -5,
					-- layer=2 filter=67 channel=110
					-33, 42, -12, -35, -29, -49, -34, -22, -17,
					-- layer=2 filter=67 channel=111
					-3, -4, -9, 3, 6, -11, -2, 1, 3,
					-- layer=2 filter=67 channel=112
					22, 2, 1, 4, -27, -8, 32, 14, 37,
					-- layer=2 filter=67 channel=113
					6, 12, -90, -77, -31, -44, -87, -91, -62,
					-- layer=2 filter=67 channel=114
					8, -1, 22, 8, 8, 25, 7, 6, 20,
					-- layer=2 filter=67 channel=115
					0, -4, -7, 1, -3, 0, 9, -6, 1,
					-- layer=2 filter=67 channel=116
					26, 6, 41, 7, 12, 14, 34, -29, 29,
					-- layer=2 filter=67 channel=117
					-2, 9, 10, -56, -71, -14, 38, 28, -28,
					-- layer=2 filter=67 channel=118
					1, 13, 27, -12, 36, 16, -14, 0, -30,
					-- layer=2 filter=67 channel=119
					0, -3, -9, -49, -56, -51, -91, -58, -63,
					-- layer=2 filter=67 channel=120
					-1, 6, 5, -3, -1, -7, 4, -4, -10,
					-- layer=2 filter=67 channel=121
					11, -5, -9, 2, 5, 0, 1, 1, -2,
					-- layer=2 filter=67 channel=122
					-4, 10, 4, 7, -2, -9, 0, 4, 0,
					-- layer=2 filter=67 channel=123
					13, 47, 18, -71, -15, -39, 31, -8, -13,
					-- layer=2 filter=67 channel=124
					39, 25, 3, -25, -40, -14, -26, -16, 1,
					-- layer=2 filter=67 channel=125
					-4, 8, -1, 0, -12, -5, 10, -8, 2,
					-- layer=2 filter=67 channel=126
					34, -14, 27, 23, 28, 13, -30, 46, -11,
					-- layer=2 filter=67 channel=127
					23, -33, -27, -30, 15, -44, -68, -14, -6,
					-- layer=2 filter=68 channel=0
					-22, -7, -5, -11, -18, -13, -23, -9, -12,
					-- layer=2 filter=68 channel=1
					5, 4, -17, 0, -10, -10, 4, -12, -17,
					-- layer=2 filter=68 channel=2
					-5, -4, -11, -11, 0, -3, -1, -5, -9,
					-- layer=2 filter=68 channel=3
					-17, -5, -24, -10, -6, -9, -7, -11, -3,
					-- layer=2 filter=68 channel=4
					-12, -8, -6, -2, 3, 0, -9, 0, -5,
					-- layer=2 filter=68 channel=5
					-10, -12, -18, -14, -2, -9, -15, -20, -2,
					-- layer=2 filter=68 channel=6
					1, -19, 13, -10, -16, 3, -10, 1, -8,
					-- layer=2 filter=68 channel=7
					1, -9, -14, -7, -17, -10, -5, 0, -13,
					-- layer=2 filter=68 channel=8
					3, -6, -2, -1, -7, 10, 0, 0, 8,
					-- layer=2 filter=68 channel=9
					-11, -2, -3, 0, -15, -11, -20, 1, -1,
					-- layer=2 filter=68 channel=10
					-21, -9, 0, -21, -18, -18, -23, -9, 2,
					-- layer=2 filter=68 channel=11
					-15, -10, -4, -9, -3, -14, -3, -8, -8,
					-- layer=2 filter=68 channel=12
					-1, -11, -5, 4, 4, -15, -10, -3, -9,
					-- layer=2 filter=68 channel=13
					-10, 7, 4, -7, 10, 6, -9, -4, -9,
					-- layer=2 filter=68 channel=14
					-6, -1, -18, -10, -11, -12, 7, -1, -18,
					-- layer=2 filter=68 channel=15
					-9, -10, 5, -14, -18, -5, -3, -10, 3,
					-- layer=2 filter=68 channel=16
					-2, 5, 12, 4, 0, 11, 8, -7, -11,
					-- layer=2 filter=68 channel=17
					4, -11, 8, 2, -7, 1, 8, 1, -1,
					-- layer=2 filter=68 channel=18
					-15, 2, -21, 2, -13, -6, -22, -6, 4,
					-- layer=2 filter=68 channel=19
					-7, -9, 2, -1, -20, -17, -2, -8, -7,
					-- layer=2 filter=68 channel=20
					3, 6, -5, -9, -11, -9, 0, 6, 3,
					-- layer=2 filter=68 channel=21
					3, 2, 2, 10, 9, 6, 5, -4, -3,
					-- layer=2 filter=68 channel=22
					2, -3, 3, -7, 11, 7, -3, 10, 9,
					-- layer=2 filter=68 channel=23
					6, 7, 15, -11, -6, 6, -15, -5, -12,
					-- layer=2 filter=68 channel=24
					-1, -8, -4, -14, -10, 5, -12, 3, -14,
					-- layer=2 filter=68 channel=25
					-8, -11, -24, -15, -15, -8, -3, 1, -4,
					-- layer=2 filter=68 channel=26
					-5, 6, -1, -3, 3, 6, 8, -2, 0,
					-- layer=2 filter=68 channel=27
					-8, -20, -11, -10, -6, -20, -4, -13, -17,
					-- layer=2 filter=68 channel=28
					-23, -18, -10, -10, -11, -15, 2, 7, -4,
					-- layer=2 filter=68 channel=29
					-10, -8, -6, -9, -9, -6, -5, -3, -2,
					-- layer=2 filter=68 channel=30
					-16, 0, 1, -16, -5, -7, -4, -18, -14,
					-- layer=2 filter=68 channel=31
					-10, -14, 5, -12, -8, -2, 5, -8, -5,
					-- layer=2 filter=68 channel=32
					0, -5, 0, 3, 5, 8, 0, 0, 5,
					-- layer=2 filter=68 channel=33
					-5, -11, -8, 1, -8, 1, 4, 8, -9,
					-- layer=2 filter=68 channel=34
					-11, -5, -6, -5, -2, -16, -16, -3, -9,
					-- layer=2 filter=68 channel=35
					-14, -10, -5, -15, -16, -6, -10, 1, -6,
					-- layer=2 filter=68 channel=36
					-3, 2, -8, -2, -11, -10, -8, -6, 7,
					-- layer=2 filter=68 channel=37
					-14, -14, -11, -14, -4, -20, 0, -18, 0,
					-- layer=2 filter=68 channel=38
					-2, -16, -14, -8, -4, -20, 1, -20, -9,
					-- layer=2 filter=68 channel=39
					-3, -5, -8, -3, -9, 4, -7, -14, -5,
					-- layer=2 filter=68 channel=40
					-9, -19, -4, 7, -13, 17, -15, -12, 0,
					-- layer=2 filter=68 channel=41
					0, 2, 0, 1, 0, -9, 7, -7, -5,
					-- layer=2 filter=68 channel=42
					0, 16, 3, 10, 2, -6, -5, -2, 5,
					-- layer=2 filter=68 channel=43
					0, -11, -15, -13, 1, 3, 7, -6, -6,
					-- layer=2 filter=68 channel=44
					9, 11, 10, 6, 6, 5, 7, -10, -5,
					-- layer=2 filter=68 channel=45
					-3, -17, -15, 4, 9, -3, -5, -11, 4,
					-- layer=2 filter=68 channel=46
					-15, -1, -13, -22, -8, -14, -14, -22, -14,
					-- layer=2 filter=68 channel=47
					-12, -11, -10, 8, 4, -3, -10, -1, 1,
					-- layer=2 filter=68 channel=48
					-7, -1, 5, 7, 7, 0, 0, 6, -7,
					-- layer=2 filter=68 channel=49
					0, -7, -1, -4, -8, -16, -15, -11, -8,
					-- layer=2 filter=68 channel=50
					-8, 0, 3, 10, -6, -2, 5, 3, 8,
					-- layer=2 filter=68 channel=51
					-3, -2, -9, -4, -13, -12, -4, -1, -1,
					-- layer=2 filter=68 channel=52
					-15, -4, -9, -1, -5, -6, 2, -11, 8,
					-- layer=2 filter=68 channel=53
					11, 3, 1, 1, 8, -11, -18, -3, -2,
					-- layer=2 filter=68 channel=54
					-14, -7, -16, -6, 0, -16, -20, -4, -5,
					-- layer=2 filter=68 channel=55
					-2, 2, -5, -6, 5, 7, 8, 0, 7,
					-- layer=2 filter=68 channel=56
					-4, -13, -15, -2, -21, -12, -7, -11, -8,
					-- layer=2 filter=68 channel=57
					-8, -3, -10, -2, 10, -2, -8, 4, -8,
					-- layer=2 filter=68 channel=58
					-5, 1, -10, 4, -2, -9, 5, -1, -14,
					-- layer=2 filter=68 channel=59
					-3, -6, 0, -7, 2, -10, -10, 0, -3,
					-- layer=2 filter=68 channel=60
					-24, -4, -3, -13, -14, -6, -5, -10, -3,
					-- layer=2 filter=68 channel=61
					-5, -5, -1, -2, -8, -14, -16, -10, -8,
					-- layer=2 filter=68 channel=62
					-5, -16, 0, -4, -7, -13, -9, -5, 5,
					-- layer=2 filter=68 channel=63
					0, 2, -5, 0, -14, 2, -3, -7, 4,
					-- layer=2 filter=68 channel=64
					-4, 4, 11, 4, 0, 4, -2, -16, 0,
					-- layer=2 filter=68 channel=65
					-16, -10, 16, -13, -9, 0, -14, -4, -20,
					-- layer=2 filter=68 channel=66
					7, 4, -3, -7, 0, -2, -7, 0, -6,
					-- layer=2 filter=68 channel=67
					-4, 0, -8, -14, -17, -3, -12, -22, -11,
					-- layer=2 filter=68 channel=68
					0, 4, 0, 3, 0, 0, 8, 7, 8,
					-- layer=2 filter=68 channel=69
					2, 0, 13, -9, -7, -1, 3, 0, 8,
					-- layer=2 filter=68 channel=70
					-3, 1, 3, -18, -23, -24, -8, -6, -13,
					-- layer=2 filter=68 channel=71
					3, -1, 8, -5, -13, -6, -10, -17, -8,
					-- layer=2 filter=68 channel=72
					-9, -7, -19, -17, -5, 0, -12, -15, -24,
					-- layer=2 filter=68 channel=73
					7, -15, 7, -4, -4, 6, -13, 16, -5,
					-- layer=2 filter=68 channel=74
					-9, 1, -1, -6, -4, -8, -17, -13, -1,
					-- layer=2 filter=68 channel=75
					-13, -14, 2, -17, -17, -3, 4, 0, -3,
					-- layer=2 filter=68 channel=76
					6, -10, -12, 2, 4, 10, 2, 8, 6,
					-- layer=2 filter=68 channel=77
					-1, -5, -6, -8, 7, -6, -4, 7, -5,
					-- layer=2 filter=68 channel=78
					-6, -9, -6, -10, -3, -9, -18, -9, 2,
					-- layer=2 filter=68 channel=79
					-2, 6, -3, 2, 6, 5, 2, 5, 4,
					-- layer=2 filter=68 channel=80
					-5, -2, 9, 2, -11, -5, -14, -2, -3,
					-- layer=2 filter=68 channel=81
					7, 1, 4, 7, 7, -4, 2, -4, -2,
					-- layer=2 filter=68 channel=82
					-1, 9, -11, -5, 7, 4, 1, 6, 1,
					-- layer=2 filter=68 channel=83
					3, 2, -1, -2, -4, -10, -5, 1, -7,
					-- layer=2 filter=68 channel=84
					4, 3, 6, -2, 0, 6, 7, -4, 5,
					-- layer=2 filter=68 channel=85
					0, -9, 5, -5, 9, -2, -2, 4, 5,
					-- layer=2 filter=68 channel=86
					1, -3, 4, 0, -7, -4, -7, -9, 8,
					-- layer=2 filter=68 channel=87
					-23, -12, -3, -6, -19, 12, -13, -3, -12,
					-- layer=2 filter=68 channel=88
					-5, 7, 1, -14, -5, -11, -17, -6, 2,
					-- layer=2 filter=68 channel=89
					-2, -13, -16, 3, -11, -9, -3, -3, -6,
					-- layer=2 filter=68 channel=90
					0, -4, 1, 2, -4, 0, -5, -10, -3,
					-- layer=2 filter=68 channel=91
					-15, 6, -6, 1, -10, -9, 0, -9, -14,
					-- layer=2 filter=68 channel=92
					-8, 8, 0, -1, -7, -14, 8, -7, -24,
					-- layer=2 filter=68 channel=93
					-6, 8, 0, 0, 7, 3, -2, -10, -16,
					-- layer=2 filter=68 channel=94
					-3, -8, 12, -1, 3, 5, -12, 0, -10,
					-- layer=2 filter=68 channel=95
					-12, 1, 4, 3, -7, 0, -1, -4, 8,
					-- layer=2 filter=68 channel=96
					1, -5, 7, 4, 3, 5, 1, 3, 0,
					-- layer=2 filter=68 channel=97
					5, -14, -3, -5, 2, -8, -18, -12, -1,
					-- layer=2 filter=68 channel=98
					-14, -15, -3, 1, -9, -21, -8, 4, -9,
					-- layer=2 filter=68 channel=99
					-7, 0, -12, -6, -4, -9, 5, -14, 3,
					-- layer=2 filter=68 channel=100
					-1, -13, -4, -18, -18, -12, 0, -23, 0,
					-- layer=2 filter=68 channel=101
					-10, 7, -2, -3, -19, 1, -4, -5, -26,
					-- layer=2 filter=68 channel=102
					11, 7, -17, -5, 2, 2, -8, 8, 4,
					-- layer=2 filter=68 channel=103
					-2, -7, -10, -5, -4, -11, 7, -8, 4,
					-- layer=2 filter=68 channel=104
					-14, -1, 10, -6, 5, -8, -22, 13, -15,
					-- layer=2 filter=68 channel=105
					4, -1, -9, -2, -1, 0, 3, 6, 0,
					-- layer=2 filter=68 channel=106
					-19, -6, -9, -5, -11, -11, -17, 7, -19,
					-- layer=2 filter=68 channel=107
					-4, 7, 6, 6, -6, 8, -3, -9, -3,
					-- layer=2 filter=68 channel=108
					4, 0, -18, 0, -2, -8, 12, -3, -10,
					-- layer=2 filter=68 channel=109
					-7, 0, 4, -1, 8, 8, 3, 4, 4,
					-- layer=2 filter=68 channel=110
					1, 0, 12, -9, -7, 3, -3, -12, -1,
					-- layer=2 filter=68 channel=111
					3, 4, 8, -6, 0, -11, 6, 0, 0,
					-- layer=2 filter=68 channel=112
					-22, -15, -13, -18, -15, -6, -6, -12, -17,
					-- layer=2 filter=68 channel=113
					0, 6, -4, -18, -5, -24, -9, -11, -4,
					-- layer=2 filter=68 channel=114
					11, -1, 6, -5, -4, -10, -9, -6, -5,
					-- layer=2 filter=68 channel=115
					8, 10, -6, 6, 3, 2, 4, -4, -4,
					-- layer=2 filter=68 channel=116
					-7, -15, 0, -11, -15, 0, -23, 0, -13,
					-- layer=2 filter=68 channel=117
					0, -15, -7, 10, -18, 4, -20, -3, -20,
					-- layer=2 filter=68 channel=118
					-22, -16, -19, -25, -5, -5, -26, -17, -9,
					-- layer=2 filter=68 channel=119
					-2, 6, -22, -3, -17, -19, -4, -19, -9,
					-- layer=2 filter=68 channel=120
					7, 1, 2, -8, -6, -9, 9, 4, 1,
					-- layer=2 filter=68 channel=121
					1, 8, -5, 4, 2, -5, -5, -10, 6,
					-- layer=2 filter=68 channel=122
					0, 9, -9, 9, 6, 7, 9, 6, -3,
					-- layer=2 filter=68 channel=123
					-15, -13, -21, 1, -15, -10, -6, -10, -11,
					-- layer=2 filter=68 channel=124
					-16, -2, 1, -5, -11, -6, -7, -6, -15,
					-- layer=2 filter=68 channel=125
					10, -7, 0, 5, -7, 3, 8, 7, 0,
					-- layer=2 filter=68 channel=126
					6, -12, 2, 3, -8, 3, -1, 0, 11,
					-- layer=2 filter=68 channel=127
					-15, -2, -4, -1, 3, 8, -15, -9, -6,
					-- layer=2 filter=69 channel=0
					-6, -7, -13, -15, 4, -1, -3, -21, -20,
					-- layer=2 filter=69 channel=1
					-7, -8, -12, 0, -22, -2, -4, -1, 7,
					-- layer=2 filter=69 channel=2
					-6, 6, -5, -11, 9, -2, 0, -10, 0,
					-- layer=2 filter=69 channel=3
					-7, -12, 0, 3, 2, -7, -17, -5, -4,
					-- layer=2 filter=69 channel=4
					0, 5, -8, -7, -17, -5, 2, -2, -7,
					-- layer=2 filter=69 channel=5
					-13, -18, -11, -4, -19, -19, -11, -12, -17,
					-- layer=2 filter=69 channel=6
					-5, 5, 0, -25, 9, 2, 5, -3, 0,
					-- layer=2 filter=69 channel=7
					12, 0, -7, -9, -2, 1, -9, -13, 4,
					-- layer=2 filter=69 channel=8
					7, 4, -5, -1, 0, -7, 9, -1, -10,
					-- layer=2 filter=69 channel=9
					-17, -17, -14, 6, -9, 2, -12, 5, 1,
					-- layer=2 filter=69 channel=10
					-13, -3, -10, -12, -8, -10, -9, -7, -12,
					-- layer=2 filter=69 channel=11
					-14, -2, -10, -6, -9, -19, -23, -20, -12,
					-- layer=2 filter=69 channel=12
					-9, -4, -15, -12, -19, -10, 0, -6, 5,
					-- layer=2 filter=69 channel=13
					0, 8, -1, -10, -1, 0, 7, -1, 8,
					-- layer=2 filter=69 channel=14
					-8, -16, 1, -6, -7, -5, 7, -4, 8,
					-- layer=2 filter=69 channel=15
					-9, -8, -4, -9, -2, 6, -9, 0, -9,
					-- layer=2 filter=69 channel=16
					2, 9, 2, 5, 10, 0, -10, -6, -10,
					-- layer=2 filter=69 channel=17
					2, -8, 3, 7, -5, 0, -4, -9, 6,
					-- layer=2 filter=69 channel=18
					17, 5, -10, 0, -22, -2, 7, -11, -7,
					-- layer=2 filter=69 channel=19
					-3, -14, -9, -19, -9, -13, -4, 3, -1,
					-- layer=2 filter=69 channel=20
					1, 1, 1, -4, -3, 4, -4, 5, 0,
					-- layer=2 filter=69 channel=21
					3, 4, 5, 7, -2, -9, 6, 0, -6,
					-- layer=2 filter=69 channel=22
					2, -1, 3, -1, -2, -1, -3, 4, -7,
					-- layer=2 filter=69 channel=23
					-16, 5, -3, -6, -7, -7, -8, 5, 2,
					-- layer=2 filter=69 channel=24
					-16, -9, -5, 4, 10, 2, 0, -6, -2,
					-- layer=2 filter=69 channel=25
					-10, -3, -13, -17, -8, -3, -14, -15, 0,
					-- layer=2 filter=69 channel=26
					-7, 4, -4, -6, 9, -7, 1, -9, 0,
					-- layer=2 filter=69 channel=27
					-4, -16, -4, -11, -7, 6, -14, 6, 15,
					-- layer=2 filter=69 channel=28
					8, -6, 0, -1, 10, 2, -3, -11, -16,
					-- layer=2 filter=69 channel=29
					-9, 1, 5, -3, -3, 0, -5, 0, 0,
					-- layer=2 filter=69 channel=30
					1, -8, 0, -4, 6, -2, -5, 6, 0,
					-- layer=2 filter=69 channel=31
					1, 2, -7, 0, -7, -11, -3, -6, -8,
					-- layer=2 filter=69 channel=32
					0, -7, -4, 4, -5, -2, -7, -10, -6,
					-- layer=2 filter=69 channel=33
					-7, -1, 6, -17, -19, 0, 6, -10, 7,
					-- layer=2 filter=69 channel=34
					0, -9, -4, 0, -22, -1, 6, 2, 3,
					-- layer=2 filter=69 channel=35
					12, -7, -9, -1, 12, 5, -2, 0, -13,
					-- layer=2 filter=69 channel=36
					4, 1, -6, -2, -6, -5, -9, -8, -5,
					-- layer=2 filter=69 channel=37
					0, -10, -15, -21, -9, -8, -17, -13, -4,
					-- layer=2 filter=69 channel=38
					-21, -12, -2, -18, -5, -6, -12, -6, -6,
					-- layer=2 filter=69 channel=39
					-12, -11, -7, 1, 7, 4, 0, 4, -1,
					-- layer=2 filter=69 channel=40
					-3, -10, 6, -11, -1, 0, 5, 13, -17,
					-- layer=2 filter=69 channel=41
					-11, -3, -11, -3, -10, -6, -9, -3, 8,
					-- layer=2 filter=69 channel=42
					0, -9, 4, -2, -3, 3, 12, -9, 6,
					-- layer=2 filter=69 channel=43
					7, -2, -9, -4, 0, -17, -11, -19, -13,
					-- layer=2 filter=69 channel=44
					6, -2, 8, -9, 5, 10, 7, -9, -7,
					-- layer=2 filter=69 channel=45
					-3, -3, -13, -1, -8, 11, 14, -8, 6,
					-- layer=2 filter=69 channel=46
					-13, -14, 0, -2, 3, 1, -12, -13, -2,
					-- layer=2 filter=69 channel=47
					10, -11, 5, 0, -2, 8, 0, 3, 1,
					-- layer=2 filter=69 channel=48
					2, 3, 2, 4, 8, 6, 0, 6, 8,
					-- layer=2 filter=69 channel=49
					19, -1, -2, 5, -19, -6, -4, -19, 3,
					-- layer=2 filter=69 channel=50
					11, 2, -8, -3, -2, 5, -2, 3, -6,
					-- layer=2 filter=69 channel=51
					-4, -5, -22, -13, -9, -21, -4, -17, -9,
					-- layer=2 filter=69 channel=52
					3, -15, -2, -15, -14, -18, -2, -19, 0,
					-- layer=2 filter=69 channel=53
					-4, -11, 5, 8, 7, 11, -8, 9, 5,
					-- layer=2 filter=69 channel=54
					0, 8, -2, -1, -6, -9, -10, -14, -8,
					-- layer=2 filter=69 channel=55
					-9, 7, -10, 4, 4, -8, -3, 4, -8,
					-- layer=2 filter=69 channel=56
					-10, -21, -16, 1, -20, -7, -16, -6, -19,
					-- layer=2 filter=69 channel=57
					0, 7, -3, -9, 2, 0, -2, 3, 0,
					-- layer=2 filter=69 channel=58
					-4, 0, 4, -1, -18, -18, -6, 0, 8,
					-- layer=2 filter=69 channel=59
					-8, 5, 0, -16, -5, -10, 2, 4, 8,
					-- layer=2 filter=69 channel=60
					-12, -4, 0, -6, -13, -18, 3, -13, -13,
					-- layer=2 filter=69 channel=61
					-3, 4, -2, -27, 3, -11, 5, 2, 0,
					-- layer=2 filter=69 channel=62
					-5, 2, 0, -11, -21, -25, 2, -15, -5,
					-- layer=2 filter=69 channel=63
					-14, -9, 3, -15, 4, -8, 2, -10, -4,
					-- layer=2 filter=69 channel=64
					-11, 0, -6, -1, 5, 0, 5, -8, -5,
					-- layer=2 filter=69 channel=65
					-2, -9, -17, -4, -2, 0, -5, 3, 0,
					-- layer=2 filter=69 channel=66
					7, 3, 1, -10, 6, 0, -7, -1, 7,
					-- layer=2 filter=69 channel=67
					-7, -7, -9, 5, -6, -13, 0, -4, -10,
					-- layer=2 filter=69 channel=68
					1, -11, 5, -4, -4, 1, -8, -7, -3,
					-- layer=2 filter=69 channel=69
					-1, -6, -2, -12, 0, -8, 14, 3, 0,
					-- layer=2 filter=69 channel=70
					0, -6, 5, -3, -1, -7, -1, -5, 0,
					-- layer=2 filter=69 channel=71
					-10, -4, -13, -2, -12, 11, -19, -7, -6,
					-- layer=2 filter=69 channel=72
					5, -4, 4, -9, -13, 5, 1, 0, 3,
					-- layer=2 filter=69 channel=73
					5, -10, -1, -6, 13, 1, -4, 0, 14,
					-- layer=2 filter=69 channel=74
					-11, -1, -11, -3, 6, -3, -5, -2, -8,
					-- layer=2 filter=69 channel=75
					-3, -6, 7, 5, 0, -5, 2, 2, 6,
					-- layer=2 filter=69 channel=76
					0, 5, -1, -5, -12, 0, -10, 6, 7,
					-- layer=2 filter=69 channel=77
					-8, 1, 0, 7, 2, -3, -1, -7, -1,
					-- layer=2 filter=69 channel=78
					-9, -16, -5, 1, -17, -10, -22, -12, -7,
					-- layer=2 filter=69 channel=79
					7, -6, -9, 0, 7, -3, 2, 8, 2,
					-- layer=2 filter=69 channel=80
					-5, 0, 6, -1, -3, -6, -4, -2, 5,
					-- layer=2 filter=69 channel=81
					-1, 0, -10, 2, 6, 0, 0, -7, -7,
					-- layer=2 filter=69 channel=82
					0, -3, -7, -7, 4, 7, -9, 10, 1,
					-- layer=2 filter=69 channel=83
					-6, 0, -5, -7, 11, 6, -1, -3, -2,
					-- layer=2 filter=69 channel=84
					-7, -7, -5, 3, -8, 8, 7, -2, -5,
					-- layer=2 filter=69 channel=85
					-7, -1, 0, -1, -3, 7, -9, 10, 0,
					-- layer=2 filter=69 channel=86
					5, 4, 5, 0, -7, -3, -7, -8, 3,
					-- layer=2 filter=69 channel=87
					9, -1, -19, 4, -6, -22, -12, -7, -19,
					-- layer=2 filter=69 channel=88
					-16, -14, 2, -2, -9, 9, 5, -3, -11,
					-- layer=2 filter=69 channel=89
					-5, -5, -2, 3, -16, -13, -7, 0, 4,
					-- layer=2 filter=69 channel=90
					6, 4, -6, 7, 9, 9, -8, 1, 2,
					-- layer=2 filter=69 channel=91
					0, 4, 2, -13, -3, 0, -6, 6, 0,
					-- layer=2 filter=69 channel=92
					-5, 4, -3, -5, -5, -13, 0, 7, 8,
					-- layer=2 filter=69 channel=93
					-5, -10, 3, 10, 4, 4, 8, 0, 5,
					-- layer=2 filter=69 channel=94
					-14, 0, 4, -21, -10, -5, -10, -6, 0,
					-- layer=2 filter=69 channel=95
					-2, 4, 12, -7, 9, 1, -12, -3, 5,
					-- layer=2 filter=69 channel=96
					0, 10, -18, -3, 8, -6, -14, -15, -11,
					-- layer=2 filter=69 channel=97
					-4, 0, -14, -13, -7, -9, 3, 2, 7,
					-- layer=2 filter=69 channel=98
					15, -1, -2, -4, 15, 0, -4, -7, -8,
					-- layer=2 filter=69 channel=99
					-14, -5, -2, -17, -15, -7, -20, 16, 0,
					-- layer=2 filter=69 channel=100
					-11, -15, -9, -8, 0, 0, -13, -4, -13,
					-- layer=2 filter=69 channel=101
					-10, -13, -13, -9, -7, 0, -2, 1, -4,
					-- layer=2 filter=69 channel=102
					20, 5, -2, 15, -18, -14, 6, -10, -9,
					-- layer=2 filter=69 channel=103
					7, -2, 8, -5, 4, 2, 5, 9, -14,
					-- layer=2 filter=69 channel=104
					11, 9, -14, -2, -21, -1, 3, -9, -4,
					-- layer=2 filter=69 channel=105
					5, 4, -7, 8, 1, 0, 0, 7, 0,
					-- layer=2 filter=69 channel=106
					0, -10, -5, -7, 1, -4, -6, 1, -2,
					-- layer=2 filter=69 channel=107
					8, -1, -10, -1, 8, 10, 3, 0, 2,
					-- layer=2 filter=69 channel=108
					-15, -15, 1, -12, -22, -3, -7, -4, 1,
					-- layer=2 filter=69 channel=109
					-7, -11, 6, -2, 0, 7, 0, -7, 5,
					-- layer=2 filter=69 channel=110
					-11, 0, 11, -16, -7, 8, -1, 10, -1,
					-- layer=2 filter=69 channel=111
					10, 8, 3, -9, -3, 2, 6, 8, -5,
					-- layer=2 filter=69 channel=112
					-14, -13, -14, -18, -4, 4, -15, -7, -20,
					-- layer=2 filter=69 channel=113
					-6, -4, -4, 2, -2, 5, 2, 0, 6,
					-- layer=2 filter=69 channel=114
					0, -4, -3, -4, -4, -7, 8, -3, -1,
					-- layer=2 filter=69 channel=115
					3, -9, 10, -2, -10, -4, 4, -5, -7,
					-- layer=2 filter=69 channel=116
					9, 9, -18, 0, -13, -7, 2, -9, -8,
					-- layer=2 filter=69 channel=117
					5, -1, -10, -15, -5, -6, -8, -6, 9,
					-- layer=2 filter=69 channel=118
					-8, -1, -15, -11, -7, -8, -9, -15, -4,
					-- layer=2 filter=69 channel=119
					0, -8, -17, 8, -26, -2, -9, -14, -9,
					-- layer=2 filter=69 channel=120
					-5, -8, 2, 10, 2, -7, -3, 4, -2,
					-- layer=2 filter=69 channel=121
					-5, -9, 2, 9, 3, -1, 7, -7, 0,
					-- layer=2 filter=69 channel=122
					-1, 7, -9, -5, -5, 5, -9, -7, 0,
					-- layer=2 filter=69 channel=123
					6, -1, 0, -11, -20, -1, -5, -9, 0,
					-- layer=2 filter=69 channel=124
					-2, -6, -6, -11, -17, -2, -5, -1, -11,
					-- layer=2 filter=69 channel=125
					2, 1, 5, 4, -5, -10, 2, -9, -7,
					-- layer=2 filter=69 channel=126
					-3, 0, 9, -2, 0, 0, -4, -8, 2,
					-- layer=2 filter=69 channel=127
					-6, -12, -18, -7, -5, -16, -2, -12, -13,
					-- layer=2 filter=70 channel=0
					17, 7, 15, 16, 7, 22, 1, 10, -10,
					-- layer=2 filter=70 channel=1
					-24, -27, -16, -39, -63, -55, -9, 12, 22,
					-- layer=2 filter=70 channel=2
					-4, -2, 7, 4, 2, 5, 8, 3, -5,
					-- layer=2 filter=70 channel=3
					19, -12, 0, 9, 4, 3, -12, -15, 6,
					-- layer=2 filter=70 channel=4
					-8, -1, -1, -2, 4, -6, -10, -40, -18,
					-- layer=2 filter=70 channel=5
					7, -6, 12, 3, -4, 2, 20, 6, 8,
					-- layer=2 filter=70 channel=6
					10, 45, 16, 12, 37, 10, 0, 14, 29,
					-- layer=2 filter=70 channel=7
					-57, -110, -37, -82, -112, -98, -19, -11, -8,
					-- layer=2 filter=70 channel=8
					0, -2, 7, 8, 0, 5, -4, -3, -2,
					-- layer=2 filter=70 channel=9
					21, 19, 21, 15, 6, -3, -10, -39, 0,
					-- layer=2 filter=70 channel=10
					28, 17, 9, 21, 5, 3, -6, 4, 12,
					-- layer=2 filter=70 channel=11
					-4, -5, 1, -4, 0, 2, 0, -14, -8,
					-- layer=2 filter=70 channel=12
					-49, -47, -43, -39, -71, -53, -5, 9, 29,
					-- layer=2 filter=70 channel=13
					8, -7, -5, -5, -1, 2, -3, 6, -10,
					-- layer=2 filter=70 channel=14
					-32, -50, -29, -37, -67, -46, -3, -3, -2,
					-- layer=2 filter=70 channel=15
					45, -9, -3, 51, 12, 26, 3, 59, 12,
					-- layer=2 filter=70 channel=16
					0, -34, -42, 11, 8, -15, 15, -12, 21,
					-- layer=2 filter=70 channel=17
					-3, -6, 5, 11, -4, 7, 0, 0, 5,
					-- layer=2 filter=70 channel=18
					23, 6, 0, 15, 15, 21, 9, -1, -14,
					-- layer=2 filter=70 channel=19
					-23, 17, 37, -66, -22, 9, 1, 41, 54,
					-- layer=2 filter=70 channel=20
					2, -4, -1, 8, -3, -6, -7, 12, 8,
					-- layer=2 filter=70 channel=21
					0, -4, 10, -11, 2, 1, 1, -1, -4,
					-- layer=2 filter=70 channel=22
					-7, -4, 6, 0, 10, 7, 7, 5, -4,
					-- layer=2 filter=70 channel=23
					38, 12, 6, 12, 12, -16, -16, -6, -18,
					-- layer=2 filter=70 channel=24
					-5, 14, -13, 14, 9, -19, 5, 0, -6,
					-- layer=2 filter=70 channel=25
					-9, -2, 0, 12, 7, 14, 16, -8, -4,
					-- layer=2 filter=70 channel=26
					-6, 4, 6, 8, 6, 2, 10, -8, -2,
					-- layer=2 filter=70 channel=27
					-17, -29, 14, -15, -22, 18, 6, -16, 6,
					-- layer=2 filter=70 channel=28
					-42, -115, -61, -95, -85, -27, -56, -58, -46,
					-- layer=2 filter=70 channel=29
					-1, 4, 9, 4, 10, 1, -4, -9, -4,
					-- layer=2 filter=70 channel=30
					-1, 28, 15, 6, 27, 3, 21, -27, -4,
					-- layer=2 filter=70 channel=31
					-22, 14, -69, -22, -27, -29, -36, 49, 16,
					-- layer=2 filter=70 channel=32
					5, 9, 4, -5, 0, 0, 10, 2, 1,
					-- layer=2 filter=70 channel=33
					-30, -21, -3, -92, -66, -31, -7, 4, 33,
					-- layer=2 filter=70 channel=34
					-27, -12, 20, -44, -9, 54, 10, 23, 37,
					-- layer=2 filter=70 channel=35
					-77, -81, -18, -74, -51, -17, -57, -52, -40,
					-- layer=2 filter=70 channel=36
					2, 6, 1, -7, 8, -6, -7, -7, -8,
					-- layer=2 filter=70 channel=37
					3, -14, 6, 2, 4, 13, 11, 12, 7,
					-- layer=2 filter=70 channel=38
					-4, -8, 13, 0, -1, 10, 9, -23, -5,
					-- layer=2 filter=70 channel=39
					40, 1, -1, 5, -19, -21, -39, -34, -24,
					-- layer=2 filter=70 channel=40
					26, -1, -6, 20, -44, -1, 3, -31, 11,
					-- layer=2 filter=70 channel=41
					-8, -1, 4, 2, 6, -2, 10, 8, -3,
					-- layer=2 filter=70 channel=42
					14, 23, -13, 4, -23, -20, 2, 14, 0,
					-- layer=2 filter=70 channel=43
					15, -15, 25, -12, 2, 17, -20, -50, 9,
					-- layer=2 filter=70 channel=44
					-6, -1, 4, -4, -6, -8, -5, -3, -2,
					-- layer=2 filter=70 channel=45
					17, 6, 12, 8, 5, 27, 23, -18, 30,
					-- layer=2 filter=70 channel=46
					0, 12, 6, -3, -7, -32, -14, 22, -9,
					-- layer=2 filter=70 channel=47
					-23, -91, -16, -10, -58, -2, 24, -22, 28,
					-- layer=2 filter=70 channel=48
					2, 5, -1, -7, 2, -5, 0, 0, 1,
					-- layer=2 filter=70 channel=49
					49, 40, -15, 33, 29, -2, -9, 44, -1,
					-- layer=2 filter=70 channel=50
					-3, 3, -2, 0, 1, 2, -15, 2, 10,
					-- layer=2 filter=70 channel=51
					10, -7, 18, 13, 3, 4, 12, -8, 8,
					-- layer=2 filter=70 channel=52
					-11, 28, 4, -2, 6, 8, -16, -10, 2,
					-- layer=2 filter=70 channel=53
					27, 51, 12, 25, 34, -9, 11, 60, -9,
					-- layer=2 filter=70 channel=54
					-27, -57, -37, -37, -43, -40, -9, 13, -10,
					-- layer=2 filter=70 channel=55
					10, 16, 6, 15, 8, 6, 8, -8, 2,
					-- layer=2 filter=70 channel=56
					5, -28, 4, -5, -23, 14, 3, -19, -7,
					-- layer=2 filter=70 channel=57
					-8, 7, -9, 5, -6, -6, -1, -13, 7,
					-- layer=2 filter=70 channel=58
					-65, -72, -33, -56, -77, -38, -7, -4, 14,
					-- layer=2 filter=70 channel=59
					-79, -58, 29, -12, -32, 13, 15, 55, 39,
					-- layer=2 filter=70 channel=60
					-2, -6, -6, -19, -32, -25, 50, -16, 10,
					-- layer=2 filter=70 channel=61
					9, 2, 25, 46, 1, 1, 33, -39, -7,
					-- layer=2 filter=70 channel=62
					22, 35, 18, 19, 33, 20, 28, 52, 19,
					-- layer=2 filter=70 channel=63
					-1, 7, -14, 19, -13, -2, 12, -2, -26,
					-- layer=2 filter=70 channel=64
					5, 1, -21, 2, 0, -25, -9, -22, -22,
					-- layer=2 filter=70 channel=65
					4, 46, 24, 32, -2, -14, 7, -1, -7,
					-- layer=2 filter=70 channel=66
					17, 8, 41, 34, -21, 12, 11, -5, 33,
					-- layer=2 filter=70 channel=67
					7, 27, 20, 9, 11, 4, -23, -6, 3,
					-- layer=2 filter=70 channel=68
					0, -2, 9, -6, -2, 9, -5, 5, -4,
					-- layer=2 filter=70 channel=69
					14, -6, -4, 15, 11, -15, -9, -4, 0,
					-- layer=2 filter=70 channel=70
					-44, -69, 1, -67, -77, 4, -25, -33, -15,
					-- layer=2 filter=70 channel=71
					5, -3, 27, 0, -20, 9, 5, -33, 11,
					-- layer=2 filter=70 channel=72
					-42, -92, -61, -115, -136, -39, -35, -7, -57,
					-- layer=2 filter=70 channel=73
					-14, -4, -33, 13, 36, 29, 43, 38, 32,
					-- layer=2 filter=70 channel=74
					18, 19, 14, 4, 1, 5, -2, -8, -16,
					-- layer=2 filter=70 channel=75
					-65, -95, 36, 5, -18, 0, 28, 3, 22,
					-- layer=2 filter=70 channel=76
					34, 2, 23, 33, 50, 1, -11, 19, 6,
					-- layer=2 filter=70 channel=77
					6, -11, -8, 8, -7, 8, -3, 5, 8,
					-- layer=2 filter=70 channel=78
					12, 9, -9, 14, 3, 4, 1, 7, -5,
					-- layer=2 filter=70 channel=79
					-7, -6, 10, 6, -6, -7, -5, 6, -8,
					-- layer=2 filter=70 channel=80
					28, 0, 10, 13, 9, -6, -4, -10, -13,
					-- layer=2 filter=70 channel=81
					10, 6, 5, 2, 9, 3, 5, 8, 7,
					-- layer=2 filter=70 channel=82
					7, 2, -6, -8, -9, 11, -9, -8, 6,
					-- layer=2 filter=70 channel=83
					2, -2, 6, -5, -1, 19, 1, -30, 0,
					-- layer=2 filter=70 channel=84
					-1, -5, 5, -1, -3, -9, 1, 2, -7,
					-- layer=2 filter=70 channel=85
					8, 9, -9, 4, -4, 4, 9, -4, 4,
					-- layer=2 filter=70 channel=86
					-6, 0, -11, -4, -4, -13, -1, -8, 2,
					-- layer=2 filter=70 channel=87
					-40, -12, -1, 0, 47, 12, -81, -11, 14,
					-- layer=2 filter=70 channel=88
					-15, 6, 4, 16, 18, 0, 12, 10, 1,
					-- layer=2 filter=70 channel=89
					-55, -39, -5, -48, -40, -38, -4, 35, 15,
					-- layer=2 filter=70 channel=90
					0, -7, -5, -6, -10, 3, 8, 8, -11,
					-- layer=2 filter=70 channel=91
					-22, -52, -2, 1, -23, 5, 39, 11, 58,
					-- layer=2 filter=70 channel=92
					-30, -51, -23, -44, -71, -40, -14, 9, -9,
					-- layer=2 filter=70 channel=93
					-10, 41, -23, -12, -20, 16, -6, -26, 14,
					-- layer=2 filter=70 channel=94
					42, 13, 27, 43, 7, 58, 48, 33, -28,
					-- layer=2 filter=70 channel=95
					-1, -10, -15, -7, 0, -7, 1, -3, 3,
					-- layer=2 filter=70 channel=96
					23, 67, 51, 52, 79, 12, 25, 53, 29,
					-- layer=2 filter=70 channel=97
					-15, 11, -15, 5, 8, -12, -7, -24, -1,
					-- layer=2 filter=70 channel=98
					-27, -137, -51, -55, -65, -42, -15, -66, -39,
					-- layer=2 filter=70 channel=99
					2, 15, 3, 38, 6, -9, 29, 25, 10,
					-- layer=2 filter=70 channel=100
					-8, 20, 6, 5, 9, 26, -12, -9, 8,
					-- layer=2 filter=70 channel=101
					-2, -12, 6, 3, -7, -4, -1, -10, 16,
					-- layer=2 filter=70 channel=102
					-11, 34, 27, 34, 45, 19, 27, 42, 38,
					-- layer=2 filter=70 channel=103
					-22, 21, 4, 41, 16, -11, -22, -44, 39,
					-- layer=2 filter=70 channel=104
					48, 4, -3, 38, 43, 32, 0, 55, -3,
					-- layer=2 filter=70 channel=105
					9, -50, 68, -40, 5, -11, -26, -16, -31,
					-- layer=2 filter=70 channel=106
					-1, -16, 0, -4, -19, 6, 19, -19, 19,
					-- layer=2 filter=70 channel=107
					22, 52, -36, 23, -7, -9, 14, 46, -5,
					-- layer=2 filter=70 channel=108
					5, 10, 23, 10, -6, 19, 34, -10, 20,
					-- layer=2 filter=70 channel=109
					2, 11, 9, -2, 1, 6, 6, 10, 5,
					-- layer=2 filter=70 channel=110
					-47, -20, -35, -24, -9, -33, 4, -15, 18,
					-- layer=2 filter=70 channel=111
					11, 0, -2, -12, 10, 1, 2, 7, -4,
					-- layer=2 filter=70 channel=112
					0, 8, 21, 22, -10, -25, 5, 14, -6,
					-- layer=2 filter=70 channel=113
					-1, 17, -4, -9, 0, -14, 6, -20, 2,
					-- layer=2 filter=70 channel=114
					11, 0, 19, -12, -9, 14, -3, -2, 0,
					-- layer=2 filter=70 channel=115
					7, 5, -1, -12, -8, -9, -8, -3, -6,
					-- layer=2 filter=70 channel=116
					-49, 30, 0, 4, 26, 22, -31, -17, 32,
					-- layer=2 filter=70 channel=117
					-29, -61, -53, -85, -63, -82, -11, -15, 1,
					-- layer=2 filter=70 channel=118
					19, 0, 14, 22, 32, 22, -6, -10, 25,
					-- layer=2 filter=70 channel=119
					-12, -34, -19, 20, -7, -23, 8, 26, 19,
					-- layer=2 filter=70 channel=120
					0, -2, 0, 0, 3, 2, 1, 10, 0,
					-- layer=2 filter=70 channel=121
					0, 9, 0, -6, 0, 1, 0, -10, 0,
					-- layer=2 filter=70 channel=122
					9, 15, -7, -14, 1, 2, -6, 21, 15,
					-- layer=2 filter=70 channel=123
					-92, -91, -56, -75, -77, -63, -66, -8, -25,
					-- layer=2 filter=70 channel=124
					33, -27, -43, 14, -11, -11, 14, 52, -5,
					-- layer=2 filter=70 channel=125
					0, 11, 9, 8, 5, 4, -3, 8, 0,
					-- layer=2 filter=70 channel=126
					-56, 33, 6, 7, 25, 2, 41, 22, 24,
					-- layer=2 filter=70 channel=127
					-1, -6, 11, 0, -13, -11, -3, 2, 18,
					-- layer=2 filter=71 channel=0
					-16, -21, -8, -22, -30, -4, 21, 16, 38,
					-- layer=2 filter=71 channel=1
					16, -1, 31, 0, 8, -29, 9, -8, -16,
					-- layer=2 filter=71 channel=2
					7, -8, 3, 1, 1, 4, 9, 3, 2,
					-- layer=2 filter=71 channel=3
					1, 2, -33, 13, -37, -19, 15, 17, 3,
					-- layer=2 filter=71 channel=4
					26, 15, 11, 14, -15, -6, 28, 4, 7,
					-- layer=2 filter=71 channel=5
					-70, -57, 12, -61, -67, 42, -44, -23, 44,
					-- layer=2 filter=71 channel=6
					-12, 64, 3, -1, 22, 24, -8, -10, 23,
					-- layer=2 filter=71 channel=7
					9, -11, 40, 12, -27, 14, 29, -23, 8,
					-- layer=2 filter=71 channel=8
					0, 3, 3, -3, -5, -5, 7, 5, -9,
					-- layer=2 filter=71 channel=9
					25, 15, 11, -5, 5, -37, -25, 5, 20,
					-- layer=2 filter=71 channel=10
					8, -14, -44, -27, -46, -9, 12, -25, 3,
					-- layer=2 filter=71 channel=11
					-32, -32, 28, -39, -22, 45, -23, -13, 32,
					-- layer=2 filter=71 channel=12
					28, 23, -2, -2, 0, -14, 11, -26, 39,
					-- layer=2 filter=71 channel=13
					7, -8, -6, -1, 0, 6, -2, -7, -4,
					-- layer=2 filter=71 channel=14
					6, 7, 33, 31, 19, 16, -12, -33, 9,
					-- layer=2 filter=71 channel=15
					-31, -47, -23, 1, -57, 13, -18, -6, -44,
					-- layer=2 filter=71 channel=16
					2, -10, -30, 11, 4, 11, 0, -17, -69,
					-- layer=2 filter=71 channel=17
					3, 6, -7, 4, -8, 5, 2, 9, 9,
					-- layer=2 filter=71 channel=18
					-11, -16, 0, -12, -16, 5, -59, -26, 56,
					-- layer=2 filter=71 channel=19
					-39, -14, 3, -48, 9, -28, -20, -4, -62,
					-- layer=2 filter=71 channel=20
					-1, -8, 7, -7, -1, 2, 9, 0, 8,
					-- layer=2 filter=71 channel=21
					8, 3, 20, 16, -6, 14, 11, 5, -2,
					-- layer=2 filter=71 channel=22
					2, 11, 5, 6, 2, -8, 3, -4, 7,
					-- layer=2 filter=71 channel=23
					35, -7, -6, 32, 6, -5, 52, 4, -28,
					-- layer=2 filter=71 channel=24
					27, 12, 0, 35, -5, 6, 12, -8, -1,
					-- layer=2 filter=71 channel=25
					9, 13, 3, 60, 25, 32, 37, 26, 22,
					-- layer=2 filter=71 channel=26
					8, -8, -5, -5, 2, -5, -5, -9, 0,
					-- layer=2 filter=71 channel=27
					-100, -84, -2, -82, -69, 18, -72, -41, 29,
					-- layer=2 filter=71 channel=28
					9, -6, -9, 24, 17, 38, 32, 9, -6,
					-- layer=2 filter=71 channel=29
					9, 6, 3, -7, 1, 7, -8, 4, -7,
					-- layer=2 filter=71 channel=30
					-17, 21, 7, -11, -1, 33, 18, -8, -41,
					-- layer=2 filter=71 channel=31
					-26, -27, -28, -22, -5, -2, -7, 27, 16,
					-- layer=2 filter=71 channel=32
					-9, -8, 4, 2, 6, 12, 3, 7, 4,
					-- layer=2 filter=71 channel=33
					6, 6, 42, -7, -46, 34, 39, 3, 17,
					-- layer=2 filter=71 channel=34
					-41, -21, -2, -50, 67, -18, -21, -6, 0,
					-- layer=2 filter=71 channel=35
					-12, -32, -75, 6, 0, -4, 36, 5, -7,
					-- layer=2 filter=71 channel=36
					-1, -7, 11, -7, 1, -4, -8, -8, -4,
					-- layer=2 filter=71 channel=37
					-47, -30, 23, -66, -48, 46, -83, -22, 21,
					-- layer=2 filter=71 channel=38
					-76, -61, 40, -25, -44, 19, -21, -15, 2,
					-- layer=2 filter=71 channel=39
					37, -3, -27, 2, -60, -24, -7, -36, -48,
					-- layer=2 filter=71 channel=40
					-14, -28, -57, -46, -28, -17, -26, -27, 0,
					-- layer=2 filter=71 channel=41
					3, -4, 5, 2, -8, 9, 10, 4, 3,
					-- layer=2 filter=71 channel=42
					50, 10, -11, 14, 14, -19, 54, 17, -23,
					-- layer=2 filter=71 channel=43
					-40, -33, -8, -57, -56, -13, -48, -47, 7,
					-- layer=2 filter=71 channel=44
					-10, 0, -7, -6, -3, 1, -7, 3, 5,
					-- layer=2 filter=71 channel=45
					-28, 4, -66, -37, -41, -12, 17, -31, -47,
					-- layer=2 filter=71 channel=46
					25, 5, 4, 2, -23, 0, 8, -32, -55,
					-- layer=2 filter=71 channel=47
					24, 24, 13, 35, 18, 29, 28, -6, -18,
					-- layer=2 filter=71 channel=48
					3, -2, 8, -4, 3, 5, -6, -7, 11,
					-- layer=2 filter=71 channel=49
					16, 52, -37, 12, 1, -30, -57, -44, -2,
					-- layer=2 filter=71 channel=50
					18, -7, 11, 6, -19, 5, -28, -16, -25,
					-- layer=2 filter=71 channel=51
					-45, -30, 49, -29, -18, 34, -16, 0, 15,
					-- layer=2 filter=71 channel=52
					-22, -21, 28, -47, -18, -6, -51, 3, 7,
					-- layer=2 filter=71 channel=53
					13, 72, 49, 8, 55, -24, -25, -25, -19,
					-- layer=2 filter=71 channel=54
					-2, -7, -16, 11, 4, 9, 38, -13, -10,
					-- layer=2 filter=71 channel=55
					5, -10, 9, 0, 6, -6, -6, -8, -10,
					-- layer=2 filter=71 channel=56
					-44, -47, 24, -53, -47, 14, -57, -17, 31,
					-- layer=2 filter=71 channel=57
					0, 21, -9, 3, -1, -16, 0, 5, -7,
					-- layer=2 filter=71 channel=58
					0, 14, -33, -7, -30, 0, 10, -16, 2,
					-- layer=2 filter=71 channel=59
					-70, 9, 28, -35, -42, -32, -17, -13, -23,
					-- layer=2 filter=71 channel=60
					-14, 21, 10, -40, -13, -27, -26, -36, -38,
					-- layer=2 filter=71 channel=61
					-25, 27, 9, 7, 42, 0, -15, -6, 4,
					-- layer=2 filter=71 channel=62
					-20, 29, -12, -48, 21, 15, -32, -40, -34,
					-- layer=2 filter=71 channel=63
					11, 1, -17, 15, -16, -19, 16, 4, -19,
					-- layer=2 filter=71 channel=64
					-1, -7, -14, 16, 6, -44, 23, -7, -53,
					-- layer=2 filter=71 channel=65
					-7, 35, 37, 2, 23, 1, -12, -4, -29,
					-- layer=2 filter=71 channel=66
					-3, -9, -7, 52, -13, -25, -39, -1, 22,
					-- layer=2 filter=71 channel=67
					-13, -12, 11, -42, -7, 17, -33, -26, -23,
					-- layer=2 filter=71 channel=68
					3, 2, -8, 10, 8, -4, -8, 0, 0,
					-- layer=2 filter=71 channel=69
					23, 17, -15, 17, 1, -17, 15, -9, -47,
					-- layer=2 filter=71 channel=70
					-2, -22, -56, 0, -11, 18, 34, -10, -7,
					-- layer=2 filter=71 channel=71
					-80, -73, 0, -17, 2, 55, -19, -4, 64,
					-- layer=2 filter=71 channel=72
					3, -31, 50, 4, -16, 7, 36, 50, 0,
					-- layer=2 filter=71 channel=73
					-31, 25, 37, -13, 7, 44, -11, -30, 6,
					-- layer=2 filter=71 channel=74
					0, 3, 7, 12, -9, 5, 23, -10, -9,
					-- layer=2 filter=71 channel=75
					12, 32, -17, 30, 18, -46, -7, -14, 43,
					-- layer=2 filter=71 channel=76
					-9, 17, 7, -39, 35, 10, 14, -9, -6,
					-- layer=2 filter=71 channel=77
					-3, -9, 8, -6, 5, -1, 8, 2, 1,
					-- layer=2 filter=71 channel=78
					-4, 7, -3, -10, 1, 35, 1, 2, 21,
					-- layer=2 filter=71 channel=79
					3, -10, 1, 10, 3, 4, 3, 2, -7,
					-- layer=2 filter=71 channel=80
					30, 1, -31, 32, 0, -7, 27, -34, -33,
					-- layer=2 filter=71 channel=81
					-16, -5, -10, -15, -18, -15, -12, -10, 1,
					-- layer=2 filter=71 channel=82
					-7, 1, 5, 2, 4, 6, 5, 12, 5,
					-- layer=2 filter=71 channel=83
					32, 18, -3, 13, -13, -8, 27, 23, -39,
					-- layer=2 filter=71 channel=84
					-2, -2, 4, -3, 7, -7, -5, -8, 3,
					-- layer=2 filter=71 channel=85
					-2, -13, -9, -1, -6, -11, 0, 3, -4,
					-- layer=2 filter=71 channel=86
					-12, -9, 3, -3, -7, 5, 2, -19, -14,
					-- layer=2 filter=71 channel=87
					28, 26, 30, -4, 39, 35, 31, -3, 1,
					-- layer=2 filter=71 channel=88
					-1, 17, 9, -17, 5, -19, 3, -31, -7,
					-- layer=2 filter=71 channel=89
					3, 8, 21, 33, -4, -18, 20, 13, -10,
					-- layer=2 filter=71 channel=90
					-4, 6, -4, 6, 1, -3, 1, 5, 6,
					-- layer=2 filter=71 channel=91
					20, 11, -2, 15, -14, -58, 46, -1, 13,
					-- layer=2 filter=71 channel=92
					10, -14, 7, 2, 9, -45, 31, 1, -4,
					-- layer=2 filter=71 channel=93
					32, 55, -14, 40, -23, 19, 27, 25, -2,
					-- layer=2 filter=71 channel=94
					-20, 40, -12, 1, 20, 3, -7, 14, 30,
					-- layer=2 filter=71 channel=95
					0, 8, 13, 1, 0, -9, -1, 4, -9,
					-- layer=2 filter=71 channel=96
					-22, 10, 7, 31, 33, 0, 24, 22, -12,
					-- layer=2 filter=71 channel=97
					2, 30, -29, 37, -4, 9, 16, 22, 17,
					-- layer=2 filter=71 channel=98
					26, -13, -23, 21, 16, 17, 28, 7, -21,
					-- layer=2 filter=71 channel=99
					1, 3, -28, -23, 23, 20, -67, -31, -18,
					-- layer=2 filter=71 channel=100
					17, -2, 17, -44, 7, 18, -16, -3, 29,
					-- layer=2 filter=71 channel=101
					-2, -31, 12, 18, 1, 29, 20, 4, 14,
					-- layer=2 filter=71 channel=102
					-31, 12, 44, 18, 15, -5, -33, -32, -30,
					-- layer=2 filter=71 channel=103
					-20, -31, -12, -9, -20, -23, -15, -7, 24,
					-- layer=2 filter=71 channel=104
					-1, 60, -9, -17, 3, -24, -75, -13, -6,
					-- layer=2 filter=71 channel=105
					19, -2, -2, -34, 2, 12, -9, -20, 51,
					-- layer=2 filter=71 channel=106
					6, 2, 9, 49, -11, 22, 30, 20, 1,
					-- layer=2 filter=71 channel=107
					-15, 3, 8, -4, -21, 49, 43, 35, 21,
					-- layer=2 filter=71 channel=108
					-91, -39, 15, -41, -9, 14, -57, -89, -8,
					-- layer=2 filter=71 channel=109
					16, -7, 6, 11, 0, 0, 10, 12, 13,
					-- layer=2 filter=71 channel=110
					11, -10, -1, 17, 29, -35, 12, -4, -11,
					-- layer=2 filter=71 channel=111
					9, 3, 7, -5, -7, -4, 1, 8, -1,
					-- layer=2 filter=71 channel=112
					-12, 26, -6, -13, -4, 16, 2, 7, 26,
					-- layer=2 filter=71 channel=113
					10, -3, -21, -8, 0, 0, 20, 28, -62,
					-- layer=2 filter=71 channel=114
					-8, -14, -5, -11, 1, 7, -7, -5, 16,
					-- layer=2 filter=71 channel=115
					-9, -5, -11, -6, -3, -3, 6, 2, -4,
					-- layer=2 filter=71 channel=116
					0, -4, 23, -9, 10, 11, -26, -11, -3,
					-- layer=2 filter=71 channel=117
					1, -14, 35, 30, -5, 30, 2, -49, -49,
					-- layer=2 filter=71 channel=118
					-27, -22, -31, -23, -31, -36, 7, -19, -15,
					-- layer=2 filter=71 channel=119
					-28, 0, -29, -8, -2, 0, 19, 0, 34,
					-- layer=2 filter=71 channel=120
					7, -7, 0, -10, 9, 8, -7, 4, -10,
					-- layer=2 filter=71 channel=121
					2, 6, 0, 10, 4, -2, 0, 8, -4,
					-- layer=2 filter=71 channel=122
					0, 9, 5, -4, 5, 0, -4, 13, 1,
					-- layer=2 filter=71 channel=123
					19, 0, 47, 9, 14, 35, -5, 0, -33,
					-- layer=2 filter=71 channel=124
					18, -3, 3, 19, -15, 9, 62, 22, -44,
					-- layer=2 filter=71 channel=125
					4, -2, -6, 6, 1, 9, 5, 6, 10,
					-- layer=2 filter=71 channel=126
					23, 3, 33, 20, -4, -22, 36, 24, 17,
					-- layer=2 filter=71 channel=127
					-22, -34, 0, -32, 5, 13, 54, 41, -19,
					-- layer=2 filter=72 channel=0
					7, 2, 5, -10, -3, 4, -3, 0, 3,
					-- layer=2 filter=72 channel=1
					3, 4, 6, 12, -10, -7, -2, -4, -10,
					-- layer=2 filter=72 channel=2
					-2, -2, -2, -1, -6, -3, -4, -3, 1,
					-- layer=2 filter=72 channel=3
					-5, -1, -9, -6, -6, -10, 2, 3, 1,
					-- layer=2 filter=72 channel=4
					7, -5, -17, -5, -2, -4, 5, 2, -1,
					-- layer=2 filter=72 channel=5
					-6, -8, -10, -14, -17, 0, -8, -9, -1,
					-- layer=2 filter=72 channel=6
					-5, 3, 2, 6, 5, -10, 0, -10, -1,
					-- layer=2 filter=72 channel=7
					-4, 7, -2, -3, -1, 0, -13, 0, 9,
					-- layer=2 filter=72 channel=8
					-3, -6, 3, 11, 10, 7, 0, 8, -5,
					-- layer=2 filter=72 channel=9
					-9, -2, 2, -5, -10, 2, -10, -7, -9,
					-- layer=2 filter=72 channel=10
					-6, 6, 0, 0, 0, -10, -13, 0, 3,
					-- layer=2 filter=72 channel=11
					-18, -11, -7, -3, -8, -3, -11, -9, 3,
					-- layer=2 filter=72 channel=12
					-9, -3, -1, -7, -12, -10, 6, 0, -5,
					-- layer=2 filter=72 channel=13
					-6, -5, -9, -7, 0, -8, 3, -3, 7,
					-- layer=2 filter=72 channel=14
					5, 3, -7, 6, -11, -3, -4, -12, -8,
					-- layer=2 filter=72 channel=15
					3, -12, 5, -9, 8, 3, -9, 1, -4,
					-- layer=2 filter=72 channel=16
					-9, -4, 6, -12, 0, 4, -3, -10, -2,
					-- layer=2 filter=72 channel=17
					0, -9, 0, 0, 1, 6, 4, -10, -11,
					-- layer=2 filter=72 channel=18
					-8, -5, -9, 5, 3, -5, -3, 5, -7,
					-- layer=2 filter=72 channel=19
					-11, -4, -8, -2, -2, -8, 8, 8, -7,
					-- layer=2 filter=72 channel=20
					-7, 5, -5, -6, 6, 4, 0, -12, -3,
					-- layer=2 filter=72 channel=21
					-7, -2, 5, -10, -2, 1, 2, 8, -8,
					-- layer=2 filter=72 channel=22
					5, 2, 1, 11, 7, 0, 4, -2, 10,
					-- layer=2 filter=72 channel=23
					-2, -13, 2, 1, -7, 5, -6, 0, -10,
					-- layer=2 filter=72 channel=24
					0, 3, -8, -10, -3, -10, -4, -11, -7,
					-- layer=2 filter=72 channel=25
					-16, -4, 0, -4, -14, -13, -13, -20, -7,
					-- layer=2 filter=72 channel=26
					-6, -8, 6, -10, 0, 9, -8, -8, 2,
					-- layer=2 filter=72 channel=27
					-16, -11, 0, 2, 6, -4, 5, -14, 1,
					-- layer=2 filter=72 channel=28
					-10, 3, -4, -6, -6, 5, -3, -12, 1,
					-- layer=2 filter=72 channel=29
					7, -11, 1, 0, 0, 0, 7, 3, 8,
					-- layer=2 filter=72 channel=30
					1, -2, -16, -9, -11, -4, -10, -2, -5,
					-- layer=2 filter=72 channel=31
					0, -4, 1, -12, -5, 5, 0, 10, -1,
					-- layer=2 filter=72 channel=32
					6, 0, -1, -2, -2, 4, -7, -11, -7,
					-- layer=2 filter=72 channel=33
					2, 3, 3, -8, 6, -9, -11, -1, 8,
					-- layer=2 filter=72 channel=34
					2, -4, -8, -8, -5, 0, 1, -8, 4,
					-- layer=2 filter=72 channel=35
					-2, -6, -12, 6, 4, -3, -17, 2, -9,
					-- layer=2 filter=72 channel=36
					-8, -7, -1, -5, 2, 4, -4, -1, 7,
					-- layer=2 filter=72 channel=37
					-10, -6, -8, 1, -7, -3, 3, -4, 4,
					-- layer=2 filter=72 channel=38
					-7, 2, 7, -7, -3, -2, -11, -7, 1,
					-- layer=2 filter=72 channel=39
					1, -4, -5, 0, -3, -2, 0, -8, 3,
					-- layer=2 filter=72 channel=40
					-8, 5, -1, -5, 0, 11, -10, 9, -10,
					-- layer=2 filter=72 channel=41
					5, 1, -1, 5, -1, 8, -4, -4, 7,
					-- layer=2 filter=72 channel=42
					-14, -7, -15, -12, -14, -10, -1, 4, -8,
					-- layer=2 filter=72 channel=43
					0, -10, -8, 0, 5, -10, 5, -8, 3,
					-- layer=2 filter=72 channel=44
					-7, 1, -8, -5, 6, 8, -4, 6, -4,
					-- layer=2 filter=72 channel=45
					2, -7, 3, -10, 6, -3, -5, -5, 10,
					-- layer=2 filter=72 channel=46
					-4, -1, 4, 2, 0, -6, -1, -2, 5,
					-- layer=2 filter=72 channel=47
					-6, -3, 0, 5, -1, 8, -7, -7, 0,
					-- layer=2 filter=72 channel=48
					6, -3, 8, 2, 7, 9, -4, 8, 8,
					-- layer=2 filter=72 channel=49
					-10, -11, 2, 2, -3, -15, -12, -6, -17,
					-- layer=2 filter=72 channel=50
					3, 0, -7, 0, -4, 8, 0, -2, -8,
					-- layer=2 filter=72 channel=51
					-14, -8, -10, -9, 2, -3, 0, -7, 2,
					-- layer=2 filter=72 channel=52
					-16, -19, -11, 0, -4, 5, -2, -5, 1,
					-- layer=2 filter=72 channel=53
					-9, 0, -10, 4, -1, -6, -3, 2, -9,
					-- layer=2 filter=72 channel=54
					-10, -12, 1, -11, -5, -3, -13, -6, 5,
					-- layer=2 filter=72 channel=55
					7, 8, 6, -8, -10, 10, -7, 1, -1,
					-- layer=2 filter=72 channel=56
					-13, -3, -3, -12, -8, -2, -5, -1, 1,
					-- layer=2 filter=72 channel=57
					1, 3, -3, -3, -8, -11, -10, 3, -3,
					-- layer=2 filter=72 channel=58
					-10, 5, -9, 3, -13, -5, -11, 4, 0,
					-- layer=2 filter=72 channel=59
					-9, 2, -1, 9, -2, -15, 4, -3, 6,
					-- layer=2 filter=72 channel=60
					-2, 0, 0, 1, -1, 4, 3, -4, -14,
					-- layer=2 filter=72 channel=61
					-8, -7, -2, -12, 1, -11, 5, -14, 5,
					-- layer=2 filter=72 channel=62
					-10, -7, -6, -9, 7, -8, 1, 2, -3,
					-- layer=2 filter=72 channel=63
					-6, 5, -2, -2, -12, -15, 0, -12, 3,
					-- layer=2 filter=72 channel=64
					0, -3, -11, 6, 5, 5, -1, 0, -5,
					-- layer=2 filter=72 channel=65
					-9, -7, 4, -6, -3, -1, 2, 8, -3,
					-- layer=2 filter=72 channel=66
					-1, -6, -4, 6, -7, -2, 9, 0, -1,
					-- layer=2 filter=72 channel=67
					2, -8, -10, -2, 4, -7, -4, -7, -3,
					-- layer=2 filter=72 channel=68
					-3, 2, -7, 8, 8, -2, 4, -12, -10,
					-- layer=2 filter=72 channel=69
					3, -8, 4, -3, -4, -14, -10, -14, -1,
					-- layer=2 filter=72 channel=70
					-7, 5, -18, 5, -7, -7, -4, -11, 2,
					-- layer=2 filter=72 channel=71
					-8, 0, 7, -1, -6, 1, -3, 1, -4,
					-- layer=2 filter=72 channel=72
					-11, 1, -13, 11, 5, -10, -2, -13, -4,
					-- layer=2 filter=72 channel=73
					-7, -5, -11, -2, -4, 5, 11, 1, -6,
					-- layer=2 filter=72 channel=74
					5, -2, -8, -4, 2, -6, -3, -1, 2,
					-- layer=2 filter=72 channel=75
					-10, -3, 8, -7, -4, 7, 11, -9, 0,
					-- layer=2 filter=72 channel=76
					-3, -11, 7, -3, -12, 8, -8, 9, -2,
					-- layer=2 filter=72 channel=77
					0, -3, -2, -2, -4, -9, 8, 6, -1,
					-- layer=2 filter=72 channel=78
					0, 3, -6, -9, -6, -1, -1, -9, 2,
					-- layer=2 filter=72 channel=79
					7, -2, 7, -9, -11, 0, -3, 8, 2,
					-- layer=2 filter=72 channel=80
					-7, -11, 2, 0, -6, -2, 2, -8, 5,
					-- layer=2 filter=72 channel=81
					7, 2, 5, -10, 1, -1, 0, -2, 9,
					-- layer=2 filter=72 channel=82
					-8, -7, -4, 8, 4, 2, -6, -6, 3,
					-- layer=2 filter=72 channel=83
					-7, 0, -6, -11, 1, -9, 6, 7, -4,
					-- layer=2 filter=72 channel=84
					-2, 4, 7, -3, 3, 5, 1, 10, -2,
					-- layer=2 filter=72 channel=85
					-15, 6, 4, 3, -4, 1, -8, 5, -7,
					-- layer=2 filter=72 channel=86
					1, 2, 4, 1, 7, 6, -7, 5, 7,
					-- layer=2 filter=72 channel=87
					4, 0, 2, -9, -6, -7, 1, -13, 2,
					-- layer=2 filter=72 channel=88
					-3, -12, -16, -9, 4, 4, -2, -4, -7,
					-- layer=2 filter=72 channel=89
					3, 1, 1, 10, 0, -15, -10, -7, 0,
					-- layer=2 filter=72 channel=90
					-5, -4, 7, 9, 5, -10, 4, 1, -9,
					-- layer=2 filter=72 channel=91
					4, -2, 1, -4, 2, -9, 4, -15, -4,
					-- layer=2 filter=72 channel=92
					1, 5, 0, 12, 5, 0, -11, -3, -2,
					-- layer=2 filter=72 channel=93
					5, 11, 3, 4, 0, -11, 1, -6, 3,
					-- layer=2 filter=72 channel=94
					-6, -5, -10, 0, -10, 2, 10, -13, -9,
					-- layer=2 filter=72 channel=95
					-2, 0, -9, -1, 0, -4, -9, 8, 4,
					-- layer=2 filter=72 channel=96
					-8, -10, 5, -1, 1, -8, -1, -15, 2,
					-- layer=2 filter=72 channel=97
					0, 3, -1, -6, -3, -2, 0, -12, -9,
					-- layer=2 filter=72 channel=98
					9, 0, -17, -10, 0, 9, 6, -3, -4,
					-- layer=2 filter=72 channel=99
					-3, -3, -1, 1, -2, -4, -3, 0, 4,
					-- layer=2 filter=72 channel=100
					-2, -10, 0, -6, -2, 1, 7, 5, -6,
					-- layer=2 filter=72 channel=101
					5, -15, 2, 6, -12, -12, -2, -13, 6,
					-- layer=2 filter=72 channel=102
					-8, -5, -7, -1, -14, -1, 0, -4, 0,
					-- layer=2 filter=72 channel=103
					7, -9, 2, 3, 5, 5, -6, 0, -8,
					-- layer=2 filter=72 channel=104
					3, 0, 8, 9, 5, 10, 5, 7, -8,
					-- layer=2 filter=72 channel=105
					0, -6, -8, 0, -10, -8, -5, 1, -1,
					-- layer=2 filter=72 channel=106
					-4, -1, -1, -18, 0, -12, 0, -18, -15,
					-- layer=2 filter=72 channel=107
					0, 11, 2, 9, 2, 9, -2, -4, 10,
					-- layer=2 filter=72 channel=108
					-2, -8, -7, 6, -1, 5, 0, -3, -8,
					-- layer=2 filter=72 channel=109
					7, -11, -10, 0, 1, 8, 4, 7, 4,
					-- layer=2 filter=72 channel=110
					4, 1, -1, 1, 1, -10, -4, -10, -16,
					-- layer=2 filter=72 channel=111
					-5, -11, 7, -6, 3, 11, -10, 8, 1,
					-- layer=2 filter=72 channel=112
					-3, 0, -4, -5, -7, -10, -11, 8, 0,
					-- layer=2 filter=72 channel=113
					6, -4, -5, 8, -8, -4, -1, -5, -11,
					-- layer=2 filter=72 channel=114
					2, -9, 5, 1, 7, -1, -8, -2, 9,
					-- layer=2 filter=72 channel=115
					10, 9, -7, 5, -10, -7, 0, 10, -10,
					-- layer=2 filter=72 channel=116
					-14, -10, 8, 0, -5, 1, -11, -3, -6,
					-- layer=2 filter=72 channel=117
					-12, 3, 0, 2, -10, 0, 0, -8, 14,
					-- layer=2 filter=72 channel=118
					-3, -9, -8, 8, -3, 7, 7, 0, -10,
					-- layer=2 filter=72 channel=119
					-9, -3, 3, -2, -9, 1, 7, -2, -1,
					-- layer=2 filter=72 channel=120
					8, -1, -2, -7, 9, -4, -1, 8, -1,
					-- layer=2 filter=72 channel=121
					1, -10, -2, -5, 7, 7, -4, 4, 5,
					-- layer=2 filter=72 channel=122
					4, 3, -2, 10, 0, -11, 5, -4, -7,
					-- layer=2 filter=72 channel=123
					-11, -12, -2, 0, 0, -9, 4, -5, 0,
					-- layer=2 filter=72 channel=124
					2, -14, 3, -1, 1, -8, -1, 18, -4,
					-- layer=2 filter=72 channel=125
					9, -5, 5, 0, 6, 6, 8, 7, 7,
					-- layer=2 filter=72 channel=126
					-8, 7, 0, 4, -4, -2, -9, 8, 1,
					-- layer=2 filter=72 channel=127
					3, -9, -7, 0, -2, -11, -11, 4, 6,
					-- layer=2 filter=73 channel=0
					-9, -9, -8, -3, -1, -11, 8, -8, 0,
					-- layer=2 filter=73 channel=1
					0, 6, 0, -4, -2, -3, 5, -3, -11,
					-- layer=2 filter=73 channel=2
					7, 2, -4, -2, -8, 7, -4, 0, -1,
					-- layer=2 filter=73 channel=3
					5, -11, -5, 8, 0, 4, -6, 6, 4,
					-- layer=2 filter=73 channel=4
					-2, -5, -6, -2, -9, 5, 6, -2, -1,
					-- layer=2 filter=73 channel=5
					9, 0, -8, -7, 6, 0, -6, 0, 5,
					-- layer=2 filter=73 channel=6
					-2, 3, -12, -6, -2, 2, 0, 0, -5,
					-- layer=2 filter=73 channel=7
					-6, -15, 9, -10, -6, -3, 3, 6, 0,
					-- layer=2 filter=73 channel=8
					7, 6, 6, -7, -1, -10, -7, 1, -7,
					-- layer=2 filter=73 channel=9
					-3, -11, -12, 6, -11, 1, -3, -2, 2,
					-- layer=2 filter=73 channel=10
					5, -5, -8, 7, -4, 0, 4, -10, -3,
					-- layer=2 filter=73 channel=11
					-12, 5, 1, 3, -6, 8, -11, -5, -6,
					-- layer=2 filter=73 channel=12
					-13, -6, -7, 3, 0, 0, -7, 5, -12,
					-- layer=2 filter=73 channel=13
					7, -6, -10, -1, -1, 7, 4, -5, -4,
					-- layer=2 filter=73 channel=14
					-8, -7, 5, 0, 0, -1, 5, 5, 7,
					-- layer=2 filter=73 channel=15
					1, 0, -2, -10, -3, -9, -9, 5, -9,
					-- layer=2 filter=73 channel=16
					7, -10, 8, 0, -12, 6, 1, 0, -1,
					-- layer=2 filter=73 channel=17
					7, -5, 4, -9, -1, 8, 3, -6, 3,
					-- layer=2 filter=73 channel=18
					-8, -10, -11, 0, -3, 4, -15, 10, -12,
					-- layer=2 filter=73 channel=19
					-11, -10, -15, -11, -7, -4, 0, 2, -12,
					-- layer=2 filter=73 channel=20
					2, -4, 0, -1, -8, -7, 9, -9, -2,
					-- layer=2 filter=73 channel=21
					10, -2, -4, -6, -3, 4, -1, -9, 6,
					-- layer=2 filter=73 channel=22
					5, 9, 1, -9, 6, 10, 2, 1, 3,
					-- layer=2 filter=73 channel=23
					-1, 7, -11, -3, -3, -10, 3, -6, -9,
					-- layer=2 filter=73 channel=24
					-1, -6, 2, 0, 8, 0, -2, 5, -5,
					-- layer=2 filter=73 channel=25
					0, -8, 2, -5, -2, 4, -5, -8, 3,
					-- layer=2 filter=73 channel=26
					8, 8, 8, -5, 9, 6, 0, 4, -9,
					-- layer=2 filter=73 channel=27
					0, 4, 1, 0, -3, 0, -6, -10, 2,
					-- layer=2 filter=73 channel=28
					5, 5, 4, 1, -7, -2, 4, -11, -1,
					-- layer=2 filter=73 channel=29
					-1, -5, -4, -5, -10, 1, -5, -10, -10,
					-- layer=2 filter=73 channel=30
					-7, 6, -2, 7, 3, 0, 6, -9, 7,
					-- layer=2 filter=73 channel=31
					-8, 6, 2, 6, 6, -7, 9, 3, -8,
					-- layer=2 filter=73 channel=32
					2, -8, 0, -7, 7, -9, -2, -11, -7,
					-- layer=2 filter=73 channel=33
					-16, -5, -7, -4, -4, -8, 1, 7, 3,
					-- layer=2 filter=73 channel=34
					-2, -11, 3, 3, 2, -7, -3, 1, -4,
					-- layer=2 filter=73 channel=35
					-5, -14, -2, 3, -7, -4, -7, 1, 3,
					-- layer=2 filter=73 channel=36
					0, 5, -9, -4, -3, 1, -1, 0, 1,
					-- layer=2 filter=73 channel=37
					-5, 0, 6, 0, 4, 2, -3, 0, -9,
					-- layer=2 filter=73 channel=38
					-5, 3, -12, 0, 0, 0, 4, -4, 0,
					-- layer=2 filter=73 channel=39
					4, -7, 0, -3, -3, 3, -3, -7, -9,
					-- layer=2 filter=73 channel=40
					-1, 0, 0, -9, 2, 3, 7, 3, 0,
					-- layer=2 filter=73 channel=41
					-8, -4, -4, 6, -7, 4, 7, 8, -8,
					-- layer=2 filter=73 channel=42
					-3, 4, -6, 6, -3, -11, 0, -9, 0,
					-- layer=2 filter=73 channel=43
					-5, -8, -3, 2, -12, -1, 0, 6, -1,
					-- layer=2 filter=73 channel=44
					-4, 5, -4, -9, 3, 3, -8, -4, 4,
					-- layer=2 filter=73 channel=45
					-4, 8, -5, 8, -11, 0, 2, -7, 2,
					-- layer=2 filter=73 channel=46
					-3, 7, 5, 0, -11, -12, -8, 5, -6,
					-- layer=2 filter=73 channel=47
					-4, -2, 9, -8, -3, 1, 4, -5, -8,
					-- layer=2 filter=73 channel=48
					2, -6, 2, 2, 0, 8, -5, 10, 7,
					-- layer=2 filter=73 channel=49
					-11, 0, -9, -3, -9, -4, -4, 5, -9,
					-- layer=2 filter=73 channel=50
					-10, -5, -7, 4, -1, 5, -8, -7, 7,
					-- layer=2 filter=73 channel=51
					-2, -1, -13, -9, 5, -3, -9, -10, -9,
					-- layer=2 filter=73 channel=52
					1, -3, 3, -12, -11, 5, 0, 4, 6,
					-- layer=2 filter=73 channel=53
					-6, -4, 5, 0, -8, -5, 1, -5, 5,
					-- layer=2 filter=73 channel=54
					-9, 5, 2, 2, 3, -4, -10, -1, -7,
					-- layer=2 filter=73 channel=55
					9, -1, 2, 3, 0, -9, -2, 0, 2,
					-- layer=2 filter=73 channel=56
					5, -4, 0, -3, -11, 7, 0, 5, -9,
					-- layer=2 filter=73 channel=57
					-3, 0, 5, 3, -6, 1, -4, -7, 5,
					-- layer=2 filter=73 channel=58
					-4, -6, -8, -6, -6, 0, 0, 0, 4,
					-- layer=2 filter=73 channel=59
					-15, -9, -3, -6, 6, -9, -6, 3, 0,
					-- layer=2 filter=73 channel=60
					3, -11, 3, -2, -2, 5, 2, -8, -12,
					-- layer=2 filter=73 channel=61
					-14, -10, 10, -4, -13, 2, 6, -9, 2,
					-- layer=2 filter=73 channel=62
					-16, 1, -8, -2, 4, -11, -7, 3, -16,
					-- layer=2 filter=73 channel=63
					0, -1, 0, 8, 1, 0, -4, -2, -5,
					-- layer=2 filter=73 channel=64
					-3, -1, 2, 7, -2, 0, 1, -6, 0,
					-- layer=2 filter=73 channel=65
					-8, -7, 8, 0, -9, -2, 0, -8, -12,
					-- layer=2 filter=73 channel=66
					-8, -2, -7, -9, 7, 5, -1, -7, -10,
					-- layer=2 filter=73 channel=67
					4, -11, -6, -8, -6, -12, -12, -6, 1,
					-- layer=2 filter=73 channel=68
					3, -3, -7, 0, -9, -6, 4, -4, 0,
					-- layer=2 filter=73 channel=69
					0, 0, 0, 4, 0, -5, 6, 6, 6,
					-- layer=2 filter=73 channel=70
					0, 3, 10, -5, 6, 9, -3, -6, 7,
					-- layer=2 filter=73 channel=71
					-2, -7, -10, -4, 6, 1, 1, -3, -10,
					-- layer=2 filter=73 channel=72
					0, 1, -12, 4, -16, -14, -14, -1, -2,
					-- layer=2 filter=73 channel=73
					5, -8, -13, -4, 9, 6, 0, 3, 0,
					-- layer=2 filter=73 channel=74
					7, -8, 0, -10, -1, 6, -10, -5, 8,
					-- layer=2 filter=73 channel=75
					-7, -2, 6, -10, -8, -2, -8, 0, 9,
					-- layer=2 filter=73 channel=76
					-5, -5, 6, 3, -5, -10, 4, -10, 7,
					-- layer=2 filter=73 channel=77
					-4, -1, -9, -6, 0, -6, 1, -2, 4,
					-- layer=2 filter=73 channel=78
					2, -11, -11, -3, 3, -9, 0, -8, -8,
					-- layer=2 filter=73 channel=79
					7, -5, 2, 0, -2, 3, 4, 2, -10,
					-- layer=2 filter=73 channel=80
					-10, 0, -9, 7, -1, 2, -3, -5, 6,
					-- layer=2 filter=73 channel=81
					-8, 2, 8, -9, 0, -3, -10, -4, -6,
					-- layer=2 filter=73 channel=82
					-3, 4, -1, 2, 9, 7, -8, -9, -3,
					-- layer=2 filter=73 channel=83
					1, 0, -8, -13, 0, 0, 4, -1, -7,
					-- layer=2 filter=73 channel=84
					4, 7, -7, -3, -6, -7, 0, -1, 7,
					-- layer=2 filter=73 channel=85
					3, -7, -3, -7, 0, 8, -5, 3, -5,
					-- layer=2 filter=73 channel=86
					0, 8, 7, 1, 9, 6, 5, 9, 0,
					-- layer=2 filter=73 channel=87
					0, -13, -7, 2, -4, 2, 0, -4, -2,
					-- layer=2 filter=73 channel=88
					-4, 3, 0, 5, 0, -4, 3, 2, -2,
					-- layer=2 filter=73 channel=89
					-7, -3, -6, -8, 0, -6, -3, -5, 0,
					-- layer=2 filter=73 channel=90
					-1, 5, 7, 4, 2, -9, 1, 0, 9,
					-- layer=2 filter=73 channel=91
					-3, 5, -3, -2, -2, -5, -7, -10, -1,
					-- layer=2 filter=73 channel=92
					6, -1, -3, -11, -13, -2, -8, -3, 1,
					-- layer=2 filter=73 channel=93
					8, 6, 4, -2, -8, 8, 5, 0, 2,
					-- layer=2 filter=73 channel=94
					3, -10, 5, 3, -4, -4, 9, 1, -2,
					-- layer=2 filter=73 channel=95
					0, -8, 3, 1, 2, -7, 6, -5, -11,
					-- layer=2 filter=73 channel=96
					-4, -1, 2, 0, -9, -7, -11, 2, -1,
					-- layer=2 filter=73 channel=97
					-7, 2, -6, 5, -11, 5, -5, -3, -5,
					-- layer=2 filter=73 channel=98
					-5, 8, 1, -11, -5, 9, -17, 4, -2,
					-- layer=2 filter=73 channel=99
					-7, 6, -5, -6, -6, -10, 1, -9, 7,
					-- layer=2 filter=73 channel=100
					-3, -6, 2, 2, -5, -14, -2, -6, 0,
					-- layer=2 filter=73 channel=101
					5, 5, 8, -5, 4, 0, -3, 0, 2,
					-- layer=2 filter=73 channel=102
					-12, -8, 1, 1, 5, -8, 2, 3, -9,
					-- layer=2 filter=73 channel=103
					0, -5, -1, 8, -8, 7, -6, 4, -8,
					-- layer=2 filter=73 channel=104
					-8, 7, 8, -9, -11, 1, 1, 2, 0,
					-- layer=2 filter=73 channel=105
					7, -1, 7, 3, -5, -3, -3, -5, -10,
					-- layer=2 filter=73 channel=106
					-6, 4, 2, -8, -6, 0, 0, -6, -3,
					-- layer=2 filter=73 channel=107
					-6, 7, 9, -8, 6, -10, 5, 9, 5,
					-- layer=2 filter=73 channel=108
					-1, -8, -2, -7, 0, -10, -2, -3, -7,
					-- layer=2 filter=73 channel=109
					4, -5, 0, 4, 3, 6, 0, 0, -1,
					-- layer=2 filter=73 channel=110
					5, 8, 6, 2, 6, 2, -2, -1, -6,
					-- layer=2 filter=73 channel=111
					1, -10, 0, 4, 10, -7, -9, -8, -3,
					-- layer=2 filter=73 channel=112
					-3, -10, -5, 1, -10, -6, 3, 1, -4,
					-- layer=2 filter=73 channel=113
					-3, 2, -10, 7, -1, -10, 3, 1, -3,
					-- layer=2 filter=73 channel=114
					7, 6, 8, 8, 5, 8, -10, -7, 3,
					-- layer=2 filter=73 channel=115
					-2, -1, 5, -10, -9, 0, 6, 9, -6,
					-- layer=2 filter=73 channel=116
					-8, -5, -5, -2, -3, 4, -11, -2, 2,
					-- layer=2 filter=73 channel=117
					3, -2, -8, -2, -4, -7, -8, -1, 2,
					-- layer=2 filter=73 channel=118
					-11, 0, 3, 4, 1, 1, -7, -7, -5,
					-- layer=2 filter=73 channel=119
					-3, -11, -9, 2, -11, 5, -6, -11, 5,
					-- layer=2 filter=73 channel=120
					-6, -8, 2, 6, 0, 7, 5, 5, 10,
					-- layer=2 filter=73 channel=121
					-5, -10, -2, 4, 0, 6, 5, -6, -10,
					-- layer=2 filter=73 channel=122
					3, 0, 1, 4, 7, -5, -9, 7, 3,
					-- layer=2 filter=73 channel=123
					1, -10, 4, 5, -1, -8, 2, 9, -4,
					-- layer=2 filter=73 channel=124
					-11, -6, 1, -11, 2, 3, -1, -1, -7,
					-- layer=2 filter=73 channel=125
					0, -7, -9, -9, 2, 10, 8, -10, -2,
					-- layer=2 filter=73 channel=126
					0, -8, 3, -1, -1, 8, 6, 8, 3,
					-- layer=2 filter=73 channel=127
					-5, -10, -9, 4, -6, -12, -3, 7, 3,
					-- layer=2 filter=74 channel=0
					-14, -22, 2, 0, -25, -11, -1, -1, 33,
					-- layer=2 filter=74 channel=1
					-4, -10, 37, 20, 32, 51, -24, 18, -11,
					-- layer=2 filter=74 channel=2
					-11, -3, -9, 8, -5, -1, 3, 6, 10,
					-- layer=2 filter=74 channel=3
					24, 27, -15, 32, -7, 3, -44, -12, 36,
					-- layer=2 filter=74 channel=4
					1, 0, -6, -3, 21, 4, 0, 27, -18,
					-- layer=2 filter=74 channel=5
					-19, -38, -18, -15, -4, 10, -14, 21, 17,
					-- layer=2 filter=74 channel=6
					-10, -19, -24, -34, -1, -27, 19, -30, 34,
					-- layer=2 filter=74 channel=7
					-34, 11, -20, -4, 22, 16, 43, 46, 57,
					-- layer=2 filter=74 channel=8
					-4, -8, 2, -1, -4, 3, -9, 8, -2,
					-- layer=2 filter=74 channel=9
					20, 8, -6, 23, -15, -30, -3, -48, -11,
					-- layer=2 filter=74 channel=10
					-1, -4, -25, 13, -6, -29, -4, 20, 27,
					-- layer=2 filter=74 channel=11
					-28, -32, -15, 5, 3, -6, 10, 5, 16,
					-- layer=2 filter=74 channel=12
					-28, -5, -3, 3, 22, 76, -13, -6, -4,
					-- layer=2 filter=74 channel=13
					0, -5, 3, 0, 7, 4, 3, -8, 0,
					-- layer=2 filter=74 channel=14
					-14, 21, 28, 3, 29, 54, -12, -9, 1,
					-- layer=2 filter=74 channel=15
					-47, -80, 6, -77, 67, 20, -59, 26, -19,
					-- layer=2 filter=74 channel=16
					10, -1, 6, -14, -6, -17, -5, 2, 4,
					-- layer=2 filter=74 channel=17
					-4, -10, 4, 4, 1, 0, 4, 8, 2,
					-- layer=2 filter=74 channel=18
					-34, -48, -42, 0, -12, 0, 20, 7, -35,
					-- layer=2 filter=74 channel=19
					-10, -23, -31, -2, 6, -45, -15, -38, -8,
					-- layer=2 filter=74 channel=20
					-5, -1, 6, 3, 9, 9, 7, -6, 3,
					-- layer=2 filter=74 channel=21
					10, 5, 26, 7, -7, 11, 2, -9, -10,
					-- layer=2 filter=74 channel=22
					-9, -8, -2, -3, 0, -8, -8, 5, -10,
					-- layer=2 filter=74 channel=23
					0, -16, 38, -8, -13, 6, 10, 7, 8,
					-- layer=2 filter=74 channel=24
					7, -13, -10, 17, 14, 20, -4, 1, 10,
					-- layer=2 filter=74 channel=25
					-32, -39, -24, 21, 16, 30, -17, 1, 28,
					-- layer=2 filter=74 channel=26
					-5, -4, -3, 0, -3, -4, 5, 10, 8,
					-- layer=2 filter=74 channel=27
					-10, -27, 18, 2, 2, 11, -2, -7, 21,
					-- layer=2 filter=74 channel=28
					-23, -18, -46, -39, 8, 22, -1, -21, 17,
					-- layer=2 filter=74 channel=29
					7, 10, -7, 1, -7, -9, 4, 1, -8,
					-- layer=2 filter=74 channel=30
					3, 4, 12, -10, -30, -14, 8, -14, 1,
					-- layer=2 filter=74 channel=31
					-72, -61, -61, -43, 0, -35, -57, -17, 46,
					-- layer=2 filter=74 channel=32
					-4, 6, 2, 8, 0, 4, -1, 2, 3,
					-- layer=2 filter=74 channel=33
					-23, 0, 14, -22, -7, 20, -5, 7, 25,
					-- layer=2 filter=74 channel=34
					-34, -68, -44, -2, -9, 15, 29, -8, -2,
					-- layer=2 filter=74 channel=35
					-70, -24, -61, -51, 13, -2, 2, -3, 26,
					-- layer=2 filter=74 channel=36
					-7, -9, -3, 19, 4, -5, 5, 7, -1,
					-- layer=2 filter=74 channel=37
					-10, -19, 0, 17, 3, -8, 1, 2, 3,
					-- layer=2 filter=74 channel=38
					6, -18, -12, -7, 13, -25, 20, 38, 12,
					-- layer=2 filter=74 channel=39
					0, -4, 3, -7, -14, -24, -63, -24, 12,
					-- layer=2 filter=74 channel=40
					-24, -26, 0, -42, 31, 27, -14, -68, 11,
					-- layer=2 filter=74 channel=41
					-12, -8, 0, -5, -7, 8, 6, 7, 10,
					-- layer=2 filter=74 channel=42
					-1, 26, 8, -7, -11, -5, -13, 0, 1,
					-- layer=2 filter=74 channel=43
					-45, -43, -13, -11, 17, -3, -27, 11, 34,
					-- layer=2 filter=74 channel=44
					6, 2, 5, -2, 10, -3, -5, -4, 9,
					-- layer=2 filter=74 channel=45
					-84, -6, -8, -47, -22, -23, -22, 0, 58,
					-- layer=2 filter=74 channel=46
					26, 4, 19, 16, 2, -11, 15, 13, 10,
					-- layer=2 filter=74 channel=47
					15, -14, -13, -12, 15, 45, 9, -7, 29,
					-- layer=2 filter=74 channel=48
					-5, 2, 0, -4, -10, -3, -1, -8, 7,
					-- layer=2 filter=74 channel=49
					-14, 10, -14, 33, -20, 20, 0, -15, -16,
					-- layer=2 filter=74 channel=50
					16, -9, 9, 13, -13, 1, -17, -4, -6,
					-- layer=2 filter=74 channel=51
					-10, -15, 4, 6, -11, -2, -1, 6, 10,
					-- layer=2 filter=74 channel=52
					-47, -2, 26, 12, 29, -11, 11, 17, -16,
					-- layer=2 filter=74 channel=53
					-5, 8, -15, 19, 8, 22, -38, -39, -23,
					-- layer=2 filter=74 channel=54
					-29, -10, 10, -16, 13, 39, 14, 6, 5,
					-- layer=2 filter=74 channel=55
					5, -3, 5, 4, 5, 11, 1, 3, 6,
					-- layer=2 filter=74 channel=56
					-10, -32, -13, -2, -13, -15, 24, -5, 0,
					-- layer=2 filter=74 channel=57
					12, 8, -2, -5, -1, -8, 7, -4, -2,
					-- layer=2 filter=74 channel=58
					-28, -25, -33, -30, 20, 59, 28, 14, 30,
					-- layer=2 filter=74 channel=59
					0, -8, 8, 15, -21, -33, -13, 12, 34,
					-- layer=2 filter=74 channel=60
					-9, -6, 2, -4, 48, 27, -20, 13, -4,
					-- layer=2 filter=74 channel=61
					0, 23, 4, -22, 37, 4, -16, -25, 32,
					-- layer=2 filter=74 channel=62
					-2, -30, -23, 15, -19, -41, 21, -23, -3,
					-- layer=2 filter=74 channel=63
					16, -2, 4, 9, 8, 22, -23, -5, -7,
					-- layer=2 filter=74 channel=64
					36, 40, 30, 7, 26, -12, -18, -2, -11,
					-- layer=2 filter=74 channel=65
					7, 8, -22, -6, 46, -31, -14, 21, 2,
					-- layer=2 filter=74 channel=66
					-9, 10, 4, -23, 6, -13, 0, -12, 56,
					-- layer=2 filter=74 channel=67
					45, 19, -15, 20, -7, -38, 38, 0, -34,
					-- layer=2 filter=74 channel=68
					-1, 3, -6, 8, 0, -1, 12, 1, -1,
					-- layer=2 filter=74 channel=69
					17, 22, 32, 4, -4, 2, -7, -10, -18,
					-- layer=2 filter=74 channel=70
					-48, -40, -11, -40, 12, 33, -7, 7, 15,
					-- layer=2 filter=74 channel=71
					-15, 15, 26, 0, -14, 20, -18, -33, 5,
					-- layer=2 filter=74 channel=72
					-18, 37, 17, -4, 17, 26, 7, 0, 16,
					-- layer=2 filter=74 channel=73
					16, 13, -42, 25, 27, -18, 40, -4, 43,
					-- layer=2 filter=74 channel=74
					13, 12, -15, -21, -32, -34, 10, 32, -11,
					-- layer=2 filter=74 channel=75
					-1, 2, -38, -16, 38, 34, -23, -23, -3,
					-- layer=2 filter=74 channel=76
					-5, 6, -9, 40, 13, -35, 8, -11, 44,
					-- layer=2 filter=74 channel=77
					1, 5, -9, -8, 3, 4, -5, 1, 2,
					-- layer=2 filter=74 channel=78
					-27, -24, -67, 35, 8, -17, 24, 10, 0,
					-- layer=2 filter=74 channel=79
					6, -3, 11, 6, 10, -2, 2, -7, 1,
					-- layer=2 filter=74 channel=80
					22, 17, 12, 0, -3, -13, 3, -24, -11,
					-- layer=2 filter=74 channel=81
					-1, -1, 10, -3, -11, 4, 3, -1, 3,
					-- layer=2 filter=74 channel=82
					3, -12, 0, -3, -7, 8, 5, -6, 4,
					-- layer=2 filter=74 channel=83
					26, 14, 2, -22, 1, 15, -4, 40, -27,
					-- layer=2 filter=74 channel=84
					4, -8, 10, -4, 3, -5, 1, 6, 9,
					-- layer=2 filter=74 channel=85
					6, -5, -7, 3, -11, 4, -14, -5, 12,
					-- layer=2 filter=74 channel=86
					8, 17, 2, 1, 6, 6, 1, -5, -4,
					-- layer=2 filter=74 channel=87
					-83, -34, 1, 0, 12, -21, 23, 15, 3,
					-- layer=2 filter=74 channel=88
					11, 17, 3, -32, 6, -19, -26, 11, -6,
					-- layer=2 filter=74 channel=89
					-22, 5, -6, 15, -17, 16, -9, -3, -5,
					-- layer=2 filter=74 channel=90
					-7, -2, -3, 8, 2, -6, 0, -7, 0,
					-- layer=2 filter=74 channel=91
					-33, -23, -18, -9, 3, 26, -3, -16, -22,
					-- layer=2 filter=74 channel=92
					-44, -22, 0, 16, 17, 34, -32, 16, -8,
					-- layer=2 filter=74 channel=93
					-25, 11, -36, -76, -24, 12, -41, -48, -23,
					-- layer=2 filter=74 channel=94
					55, 42, 21, 34, 41, 48, 33, -29, 46,
					-- layer=2 filter=74 channel=95
					-2, -10, -1, 0, 6, 4, 1, 0, -13,
					-- layer=2 filter=74 channel=96
					3, -5, 24, 7, -32, 41, -15, -32, -31,
					-- layer=2 filter=74 channel=97
					-3, 30, -10, 14, 19, 6, -24, 1, -13,
					-- layer=2 filter=74 channel=98
					-2, 5, -13, -11, 47, 20, 25, 17, 29,
					-- layer=2 filter=74 channel=99
					-25, 1, 10, 19, 0, -43, -35, -6, -9,
					-- layer=2 filter=74 channel=100
					-10, -3, -11, -7, -4, -13, 0, 17, 13,
					-- layer=2 filter=74 channel=101
					-47, -29, 17, -14, -19, 30, -17, -27, 24,
					-- layer=2 filter=74 channel=102
					20, -41, -7, 36, -18, 38, 13, -70, -46,
					-- layer=2 filter=74 channel=103
					-52, 0, -36, -3, 16, -1, 0, 26, 20,
					-- layer=2 filter=74 channel=104
					-2, -3, -18, 23, -29, 40, -1, -35, -35,
					-- layer=2 filter=74 channel=105
					0, 35, -26, -29, -28, -58, 40, 10, 15,
					-- layer=2 filter=74 channel=106
					-13, -29, -16, -1, 6, 40, -22, -3, 10,
					-- layer=2 filter=74 channel=107
					6, -20, -30, 13, 17, -5, -41, 7, -56,
					-- layer=2 filter=74 channel=108
					3, -6, 4, 47, -30, 11, 6, -39, 17,
					-- layer=2 filter=74 channel=109
					18, 0, -10, 7, 8, -11, 12, 8, 3,
					-- layer=2 filter=74 channel=110
					24, 21, 48, -22, 5, 10, -23, 2, 14,
					-- layer=2 filter=74 channel=111
					-8, 3, 8, 7, -5, 2, -9, -11, 4,
					-- layer=2 filter=74 channel=112
					0, -26, 1, 17, 36, -13, -15, 0, 33,
					-- layer=2 filter=74 channel=113
					16, -1, 0, -4, 4, 16, 3, 19, 0,
					-- layer=2 filter=74 channel=114
					-9, -19, -10, -10, -13, -17, -18, -6, -1,
					-- layer=2 filter=74 channel=115
					0, -5, -1, 5, -4, 0, -4, 9, -6,
					-- layer=2 filter=74 channel=116
					-49, -45, -7, -7, 21, 2, 12, -18, 7,
					-- layer=2 filter=74 channel=117
					8, 30, 9, -52, 5, 24, -3, 19, -11,
					-- layer=2 filter=74 channel=118
					-12, -33, -43, 25, -14, -17, 2, -9, 2,
					-- layer=2 filter=74 channel=119
					6, -16, -45, -14, -5, -17, 9, 25, -30,
					-- layer=2 filter=74 channel=120
					1, 1, -4, 8, -10, 4, -8, -5, 1,
					-- layer=2 filter=74 channel=121
					-10, -7, -10, 0, 6, -5, -12, 4, 8,
					-- layer=2 filter=74 channel=122
					-12, -9, -15, -8, 11, 3, -3, -14, 0,
					-- layer=2 filter=74 channel=123
					-26, 4, 19, 1, 24, 45, 38, 8, 3,
					-- layer=2 filter=74 channel=124
					-29, -70, -5, -33, 39, -5, 0, 28, 37,
					-- layer=2 filter=74 channel=125
					6, -1, 4, -8, 8, -2, -5, 3, 2,
					-- layer=2 filter=74 channel=126
					-6, -1, 37, -9, -20, -25, -22, -24, -28,
					-- layer=2 filter=74 channel=127
					3, -25, 21, 5, 30, 28, -12, 24, 3,
					-- layer=2 filter=75 channel=0
					13, 15, -21, 26, 13, 0, 20, 21, -6,
					-- layer=2 filter=75 channel=1
					-20, 19, -5, -49, 0, 18, -42, -23, -17,
					-- layer=2 filter=75 channel=2
					-5, -7, 7, 2, 0, 8, -5, 6, 0,
					-- layer=2 filter=75 channel=3
					-6, 37, 13, -8, 34, 15, -58, 2, 38,
					-- layer=2 filter=75 channel=4
					-8, 12, 7, -11, -12, 31, 2, -11, 10,
					-- layer=2 filter=75 channel=5
					0, 9, -3, 11, 14, -6, 2, -25, 5,
					-- layer=2 filter=75 channel=6
					-47, -61, -60, -16, -50, -29, 38, -44, -17,
					-- layer=2 filter=75 channel=7
					12, 28, -25, -1, 36, 22, 49, 48, 13,
					-- layer=2 filter=75 channel=8
					-7, -3, -4, 10, 11, -6, 0, -7, 4,
					-- layer=2 filter=75 channel=9
					-29, -23, 10, -30, 2, 30, -7, -5, 10,
					-- layer=2 filter=75 channel=10
					15, 21, -9, 2, 9, -10, -10, 11, 43,
					-- layer=2 filter=75 channel=11
					1, -18, -15, 8, -7, 3, 9, -6, -6,
					-- layer=2 filter=75 channel=12
					-22, 12, 11, -36, -2, 35, 10, 16, -1,
					-- layer=2 filter=75 channel=13
					0, -5, 0, -2, 8, -6, -5, -8, 3,
					-- layer=2 filter=75 channel=14
					-43, -8, -9, -43, -17, 0, -8, -7, -37,
					-- layer=2 filter=75 channel=15
					30, -5, -16, -40, -10, 46, 16, -76, 93,
					-- layer=2 filter=75 channel=16
					-9, 21, 21, -38, -19, 49, -40, -38, 21,
					-- layer=2 filter=75 channel=17
					-7, 9, -5, 3, -5, -4, 3, -4, 0,
					-- layer=2 filter=75 channel=18
					39, 39, 27, 28, -32, 52, -7, -26, -6,
					-- layer=2 filter=75 channel=19
					-2, -12, 0, -20, 48, 43, -51, 13, -9,
					-- layer=2 filter=75 channel=20
					-5, 3, -3, 3, 8, -3, 0, -7, -5,
					-- layer=2 filter=75 channel=21
					22, 18, 7, -5, 4, 12, 11, -13, -5,
					-- layer=2 filter=75 channel=22
					-2, 0, -6, 7, 4, 2, 10, 7, 7,
					-- layer=2 filter=75 channel=23
					-54, 10, 16, -20, -6, 41, -33, -28, -21,
					-- layer=2 filter=75 channel=24
					6, 16, 5, -4, 16, 17, -30, 15, 18,
					-- layer=2 filter=75 channel=25
					7, -4, -8, 19, 1, 6, -2, -9, 1,
					-- layer=2 filter=75 channel=26
					3, -2, -6, -9, 9, -2, 10, 2, -1,
					-- layer=2 filter=75 channel=27
					-3, 3, -4, -11, 39, 31, -38, -18, -36,
					-- layer=2 filter=75 channel=28
					12, 12, -16, 21, 72, 27, -10, 36, 20,
					-- layer=2 filter=75 channel=29
					2, 7, -4, 8, 3, 8, 10, 2, -6,
					-- layer=2 filter=75 channel=30
					-15, 3, 18, 14, -14, 4, -3, -5, 0,
					-- layer=2 filter=75 channel=31
					-17, -44, -25, -23, 12, -10, -58, -42, -17,
					-- layer=2 filter=75 channel=32
					9, -3, 2, -3, 4, -7, -4, 0, 5,
					-- layer=2 filter=75 channel=33
					15, 14, -20, -34, -34, -4, -54, -28, -41,
					-- layer=2 filter=75 channel=34
					31, -11, -48, 17, -44, 8, -11, 17, -42,
					-- layer=2 filter=75 channel=35
					3, 13, -23, 14, 1, 17, -37, 18, 20,
					-- layer=2 filter=75 channel=36
					-4, 4, 8, -10, 3, -5, -5, -4, -6,
					-- layer=2 filter=75 channel=37
					7, -2, -7, 23, -14, 7, 5, -17, -3,
					-- layer=2 filter=75 channel=38
					-15, -8, -2, -2, 18, 11, 11, -20, -20,
					-- layer=2 filter=75 channel=39
					-43, 16, 20, -31, -18, 33, -2, 0, 31,
					-- layer=2 filter=75 channel=40
					58, 17, -21, -44, -40, 35, -19, -22, 9,
					-- layer=2 filter=75 channel=41
					-2, 7, 10, 7, 5, 8, 1, 0, -6,
					-- layer=2 filter=75 channel=42
					-53, 33, 14, -39, 29, 14, -36, -2, 1,
					-- layer=2 filter=75 channel=43
					0, 13, 2, -18, 23, 23, -71, -19, 22,
					-- layer=2 filter=75 channel=44
					-6, 9, 3, -6, 11, -5, -2, -1, 11,
					-- layer=2 filter=75 channel=45
					-6, 40, 9, -87, 29, 64, -58, 5, -6,
					-- layer=2 filter=75 channel=46
					-35, -5, 6, 20, -13, 6, 0, 11, 14,
					-- layer=2 filter=75 channel=47
					57, 45, 25, 9, 12, 42, -2, 38, -8,
					-- layer=2 filter=75 channel=48
					1, -4, 4, 3, 0, -8, 4, 2, -5,
					-- layer=2 filter=75 channel=49
					25, 16, 30, -18, -11, 45, -19, -21, 29,
					-- layer=2 filter=75 channel=50
					21, 6, 22, -9, 5, -3, 10, 3, -6,
					-- layer=2 filter=75 channel=51
					5, -14, 6, 29, 8, -14, 29, -13, -13,
					-- layer=2 filter=75 channel=52
					13, 2, -31, 14, -31, -14, -16, -8, 19,
					-- layer=2 filter=75 channel=53
					25, -38, 21, -43, 55, 16, -21, -35, 29,
					-- layer=2 filter=75 channel=54
					31, 15, 6, -6, 6, 27, 10, -17, 9,
					-- layer=2 filter=75 channel=55
					2, 0, -6, 0, 7, -1, -5, 8, -2,
					-- layer=2 filter=75 channel=56
					-3, 3, -20, 1, -5, 17, 8, -15, 12,
					-- layer=2 filter=75 channel=57
					13, -6, 0, 13, 9, -4, 17, 4, -5,
					-- layer=2 filter=75 channel=58
					3, -17, -1, -22, 4, 45, 18, 10, 1,
					-- layer=2 filter=75 channel=59
					-7, -19, 6, -48, 22, 9, -13, -48, -26,
					-- layer=2 filter=75 channel=60
					32, -3, -33, 18, 18, -62, -19, 27, -36,
					-- layer=2 filter=75 channel=61
					41, 10, 6, 49, 23, -13, 37, 17, -44,
					-- layer=2 filter=75 channel=62
					-13, -56, -28, -27, -60, 8, -10, -22, -23,
					-- layer=2 filter=75 channel=63
					5, 13, -14, -31, 16, 9, 3, 10, 4,
					-- layer=2 filter=75 channel=64
					-33, -6, 8, -37, -31, 0, -44, -18, -5,
					-- layer=2 filter=75 channel=65
					18, -36, -2, 29, -29, -69, 1, -36, -12,
					-- layer=2 filter=75 channel=66
					37, 36, 15, -22, 5, 25, -39, 10, 49,
					-- layer=2 filter=75 channel=67
					-10, -6, 4, 14, 34, 42, -18, 5, 13,
					-- layer=2 filter=75 channel=68
					-2, -8, 10, 8, -9, 7, 3, 2, 9,
					-- layer=2 filter=75 channel=69
					-36, 4, 20, -57, 0, 10, -44, -26, 6,
					-- layer=2 filter=75 channel=70
					13, 5, -54, -6, 4, 0, -14, 26, 14,
					-- layer=2 filter=75 channel=71
					-26, 9, -9, -7, 39, 19, -53, -23, -13,
					-- layer=2 filter=75 channel=72
					28, 6, -25, -29, 4, -8, -24, 19, 2,
					-- layer=2 filter=75 channel=73
					47, 9, -24, 0, 62, 16, 1, 75, 38,
					-- layer=2 filter=75 channel=74
					-6, -4, -11, -10, 14, 19, 11, 11, 11,
					-- layer=2 filter=75 channel=75
					-60, -30, -70, -51, 12, 14, 5, 53, -11,
					-- layer=2 filter=75 channel=76
					18, -58, 49, -58, 12, 27, -8, -6, 53,
					-- layer=2 filter=75 channel=77
					9, -5, 3, 3, 3, 10, 1, 1, 2,
					-- layer=2 filter=75 channel=78
					27, 4, -12, 12, -14, 2, 10, -15, 20,
					-- layer=2 filter=75 channel=79
					-6, -3, -3, -1, -3, 0, -2, 0, 0,
					-- layer=2 filter=75 channel=80
					-51, -5, 15, -41, -36, 27, -40, 26, 46,
					-- layer=2 filter=75 channel=81
					-3, 7, 0, -2, 0, 3, -1, -1, 0,
					-- layer=2 filter=75 channel=82
					0, 3, 8, 1, 5, -4, 6, -6, 6,
					-- layer=2 filter=75 channel=83
					-34, -1, 9, -40, 14, 31, -20, -30, -19,
					-- layer=2 filter=75 channel=84
					4, -7, -6, -2, -7, 8, 5, -5, -8,
					-- layer=2 filter=75 channel=85
					-4, -15, 3, -9, 12, 14, -8, -7, -1,
					-- layer=2 filter=75 channel=86
					-5, 8, 4, -1, 4, 10, 1, -12, 9,
					-- layer=2 filter=75 channel=87
					5, 26, 1, 20, -77, 32, -22, 0, 42,
					-- layer=2 filter=75 channel=88
					-7, -27, -9, -7, -21, 17, 6, -25, -2,
					-- layer=2 filter=75 channel=89
					-60, -38, -36, -44, -18, -11, -2, -8, 6,
					-- layer=2 filter=75 channel=90
					-5, -11, 3, 4, -10, 1, -3, -5, -7,
					-- layer=2 filter=75 channel=91
					-42, -29, -26, -62, -10, -14, -21, 31, 21,
					-- layer=2 filter=75 channel=92
					-31, 0, -4, -31, -5, 22, -2, -7, -5,
					-- layer=2 filter=75 channel=93
					-1, -59, -36, 24, -91, -43, 34, -13, 9,
					-- layer=2 filter=75 channel=94
					23, 12, -25, -26, 5, -11, 15, -6, 12,
					-- layer=2 filter=75 channel=95
					6, -5, -9, -7, 1, 3, -11, 2, 0,
					-- layer=2 filter=75 channel=96
					7, -60, -17, 12, -30, -62, 45, 18, 13,
					-- layer=2 filter=75 channel=97
					-13, 21, 17, -15, 23, 44, -51, 20, 17,
					-- layer=2 filter=75 channel=98
					31, 25, -25, 8, 11, 25, -8, 50, -17,
					-- layer=2 filter=75 channel=99
					-13, -15, -7, 29, 20, -32, -8, -14, -10,
					-- layer=2 filter=75 channel=100
					-11, -16, -17, -28, 4, 12, -33, -29, 21,
					-- layer=2 filter=75 channel=101
					8, 4, -24, 15, 42, 8, -49, 19, -10,
					-- layer=2 filter=75 channel=102
					13, -18, -4, 28, -10, -2, -17, -34, 2,
					-- layer=2 filter=75 channel=103
					-38, -25, 32, -2, 10, -50, 0, 14, -59,
					-- layer=2 filter=75 channel=104
					0, 2, -1, -21, -46, 27, 5, -24, 27,
					-- layer=2 filter=75 channel=105
					-8, 6, 34, -14, 22, 25, -26, -21, 6,
					-- layer=2 filter=75 channel=106
					3, 11, -18, 8, 15, -1, 0, 8, 6,
					-- layer=2 filter=75 channel=107
					-16, 19, 33, -7, 9, 30, 21, -20, -17,
					-- layer=2 filter=75 channel=108
					-51, 20, -8, 5, 30, 13, -17, -72, -21,
					-- layer=2 filter=75 channel=109
					17, -8, 5, 9, 14, 0, 5, -10, 7,
					-- layer=2 filter=75 channel=110
					-23, -5, -5, -8, -40, -24, -20, -12, -3,
					-- layer=2 filter=75 channel=111
					-2, 7, -1, 10, -11, 3, -6, 11, 6,
					-- layer=2 filter=75 channel=112
					15, 26, 15, 27, 14, -31, 10, -16, -29,
					-- layer=2 filter=75 channel=113
					20, -16, 12, 4, 21, -20, -19, 1, 11,
					-- layer=2 filter=75 channel=114
					-13, -5, -6, 12, -4, -10, -24, -11, -8,
					-- layer=2 filter=75 channel=115
					8, 4, -4, -3, 1, 10, 11, -7, 5,
					-- layer=2 filter=75 channel=116
					29, 8, -19, -34, -79, 23, -35, -33, 14,
					-- layer=2 filter=75 channel=117
					32, 25, -56, -21, 20, 48, 51, 18, -21,
					-- layer=2 filter=75 channel=118
					-12, -10, 37, -47, -1, 20, -26, 16, 58,
					-- layer=2 filter=75 channel=119
					-11, 62, 50, 16, 13, 72, -28, 2, 16,
					-- layer=2 filter=75 channel=120
					2, 8, 3, -8, 7, -6, 9, -5, -10,
					-- layer=2 filter=75 channel=121
					0, 11, 5, 0, -2, -3, 4, 5, 1,
					-- layer=2 filter=75 channel=122
					-5, 2, -11, -3, 4, 10, -2, 7, -3,
					-- layer=2 filter=75 channel=123
					11, 14, 6, -13, 32, 7, 35, 35, 3,
					-- layer=2 filter=75 channel=124
					-12, -3, 13, -37, 37, 13, 15, 7, 43,
					-- layer=2 filter=75 channel=125
					-1, -5, 7, 10, 9, 6, 5, 5, 9,
					-- layer=2 filter=75 channel=126
					18, -5, 21, -26, 43, 18, -11, 59, 38,
					-- layer=2 filter=75 channel=127
					-1, 21, -1, -9, 20, -13, -20, -44, 8,
					-- layer=2 filter=76 channel=0
					-11, 7, -9, 4, -2, -13, 3, -3, 7,
					-- layer=2 filter=76 channel=1
					-7, -17, -17, -6, -10, 5, 3, -7, -13,
					-- layer=2 filter=76 channel=2
					-4, -8, -8, 7, -2, -6, 11, -8, 7,
					-- layer=2 filter=76 channel=3
					-12, -2, -4, 6, 0, 0, 0, -2, -8,
					-- layer=2 filter=76 channel=4
					6, -2, -12, 5, -6, -3, 0, 2, -12,
					-- layer=2 filter=76 channel=5
					-1, -5, -12, -2, -11, -8, 0, 1, 3,
					-- layer=2 filter=76 channel=6
					-9, -9, 0, -7, -10, 1, -10, 7, -2,
					-- layer=2 filter=76 channel=7
					-5, 7, 5, 5, -5, 4, 16, 10, 3,
					-- layer=2 filter=76 channel=8
					-9, -9, 5, -3, 0, 5, -5, 6, 3,
					-- layer=2 filter=76 channel=9
					-10, -7, -4, 7, -11, 7, 3, -10, -8,
					-- layer=2 filter=76 channel=10
					-7, -1, 11, 9, -3, -14, 0, -7, 1,
					-- layer=2 filter=76 channel=11
					-7, -9, -12, -5, 4, -2, 0, -7, 2,
					-- layer=2 filter=76 channel=12
					-18, -22, -9, -12, 0, -4, 12, 12, 8,
					-- layer=2 filter=76 channel=13
					0, 0, 4, -6, 3, -8, 5, -3, 6,
					-- layer=2 filter=76 channel=14
					-4, -18, -18, -13, -4, 8, -1, -6, -2,
					-- layer=2 filter=76 channel=15
					-8, -6, -2, 6, 2, -3, 0, -5, -5,
					-- layer=2 filter=76 channel=16
					-5, -2, -8, 2, 1, 4, -4, 0, -4,
					-- layer=2 filter=76 channel=17
					7, 0, 6, 8, -6, -1, -7, 1, -1,
					-- layer=2 filter=76 channel=18
					-11, -13, -3, -6, 6, -15, -8, 4, -18,
					-- layer=2 filter=76 channel=19
					-16, -1, -14, -7, -2, 6, 4, 6, -9,
					-- layer=2 filter=76 channel=20
					7, 3, 7, 6, 12, 2, 9, 11, 7,
					-- layer=2 filter=76 channel=21
					5, 2, -7, 7, 5, 5, 2, 8, -6,
					-- layer=2 filter=76 channel=22
					0, -4, -4, 4, -2, 9, 5, -10, 10,
					-- layer=2 filter=76 channel=23
					-3, 3, -12, 3, -13, -14, 6, 0, 1,
					-- layer=2 filter=76 channel=24
					-11, -11, -14, 6, 3, 0, -3, -11, -4,
					-- layer=2 filter=76 channel=25
					4, -9, -17, -7, 4, 0, 1, 4, 14,
					-- layer=2 filter=76 channel=26
					-3, 2, 7, -6, -4, 0, 6, -1, 9,
					-- layer=2 filter=76 channel=27
					-15, -4, -6, -6, -3, -4, -8, -9, -2,
					-- layer=2 filter=76 channel=28
					-11, -2, 14, -6, -12, -11, -7, 8, -8,
					-- layer=2 filter=76 channel=29
					4, -7, 6, -7, -7, 7, -3, 8, -10,
					-- layer=2 filter=76 channel=30
					-3, -7, -4, 0, -4, -2, -13, -3, -7,
					-- layer=2 filter=76 channel=31
					-6, 5, -7, -6, 2, -7, 2, -5, -8,
					-- layer=2 filter=76 channel=32
					-5, 11, 1, -1, 4, -2, 0, 9, -11,
					-- layer=2 filter=76 channel=33
					-13, 5, -13, -2, 13, 8, 2, -4, -10,
					-- layer=2 filter=76 channel=34
					-9, -13, -5, -3, -13, -10, 1, -1, -6,
					-- layer=2 filter=76 channel=35
					-6, -7, 5, 0, 1, -14, -2, 0, -4,
					-- layer=2 filter=76 channel=36
					-4, -3, 7, 2, -11, 9, -1, -9, -8,
					-- layer=2 filter=76 channel=37
					-5, 0, 0, -6, 0, -3, -11, -8, 4,
					-- layer=2 filter=76 channel=38
					-9, -8, 0, -4, -2, -3, -2, -10, -7,
					-- layer=2 filter=76 channel=39
					-8, -4, -10, -7, -7, -6, 2, 5, 4,
					-- layer=2 filter=76 channel=40
					8, -8, -2, -3, 5, 1, -7, -1, -7,
					-- layer=2 filter=76 channel=41
					8, -7, -11, -9, -1, -5, 2, 7, 8,
					-- layer=2 filter=76 channel=42
					-2, -10, -7, -3, -4, 0, -12, 6, 4,
					-- layer=2 filter=76 channel=43
					-5, -2, 5, 2, -6, 2, 3, 0, -9,
					-- layer=2 filter=76 channel=44
					-4, -5, -7, -10, 7, 3, 4, 8, 1,
					-- layer=2 filter=76 channel=45
					-9, -4, 1, -7, 0, 0, 1, -2, 2,
					-- layer=2 filter=76 channel=46
					7, -5, -10, 2, 2, -9, 8, -7, -6,
					-- layer=2 filter=76 channel=47
					-17, -8, -3, -4, -16, -17, -1, -10, -16,
					-- layer=2 filter=76 channel=48
					-9, 2, -2, -1, -1, -5, -5, -4, 0,
					-- layer=2 filter=76 channel=49
					-13, -11, 3, 3, -12, 4, -16, -12, -1,
					-- layer=2 filter=76 channel=50
					7, 1, -5, 0, -7, -10, 3, -10, -6,
					-- layer=2 filter=76 channel=51
					6, -5, -8, -2, 1, -9, -15, -10, 0,
					-- layer=2 filter=76 channel=52
					-2, 2, -3, 1, 4, -11, -11, -6, -5,
					-- layer=2 filter=76 channel=53
					8, -4, -2, 5, 7, 6, -13, -4, -9,
					-- layer=2 filter=76 channel=54
					-3, 1, 4, -6, 0, 2, -3, 15, 1,
					-- layer=2 filter=76 channel=55
					9, 5, 1, 3, 5, 4, 6, -9, -2,
					-- layer=2 filter=76 channel=56
					-1, 0, -8, 0, -5, -8, -11, 0, 6,
					-- layer=2 filter=76 channel=57
					7, 4, -8, -10, -8, 2, -5, -1, -9,
					-- layer=2 filter=76 channel=58
					-12, -24, -11, -6, -1, -1, 3, 8, 4,
					-- layer=2 filter=76 channel=59
					-5, -8, -15, -17, 2, 3, 1, -11, 6,
					-- layer=2 filter=76 channel=60
					4, -3, 3, 4, -1, 0, 4, 2, -9,
					-- layer=2 filter=76 channel=61
					1, 2, -10, 0, -11, -5, -7, 6, -11,
					-- layer=2 filter=76 channel=62
					-1, -8, 6, -2, -10, -4, -6, 5, -6,
					-- layer=2 filter=76 channel=63
					-9, -8, 0, -3, -6, 1, -11, -5, -9,
					-- layer=2 filter=76 channel=64
					0, 0, 0, -5, -1, 0, 1, 0, -7,
					-- layer=2 filter=76 channel=65
					-9, 4, 5, -6, -3, -11, -11, -1, -13,
					-- layer=2 filter=76 channel=66
					-5, -3, 9, 3, -6, 1, 9, -1, 3,
					-- layer=2 filter=76 channel=67
					-7, 8, 5, 9, -5, -1, 4, -10, -10,
					-- layer=2 filter=76 channel=68
					4, 0, -5, -2, 4, -2, 8, -1, -11,
					-- layer=2 filter=76 channel=69
					-11, 4, 2, -3, 5, -11, -10, 2, 7,
					-- layer=2 filter=76 channel=70
					-12, -5, -4, -7, 2, -7, -14, -10, -13,
					-- layer=2 filter=76 channel=71
					-3, -11, -15, -16, -3, -6, -8, 0, -9,
					-- layer=2 filter=76 channel=72
					-1, -4, 5, -6, 12, -4, -10, 0, -6,
					-- layer=2 filter=76 channel=73
					2, 6, -4, -4, -8, 0, 14, -10, -13,
					-- layer=2 filter=76 channel=74
					6, -6, 4, 3, 3, 0, -11, 0, -8,
					-- layer=2 filter=76 channel=75
					0, 8, -8, 0, 9, 0, 7, -6, -9,
					-- layer=2 filter=76 channel=76
					-3, 4, -9, -2, -7, -18, -4, 0, 0,
					-- layer=2 filter=76 channel=77
					10, 5, -4, 0, 7, 1, 6, 0, 4,
					-- layer=2 filter=76 channel=78
					-9, -9, -2, 0, -2, -14, 5, -13, 4,
					-- layer=2 filter=76 channel=79
					-2, 0, 4, -5, 0, -6, -7, -5, 10,
					-- layer=2 filter=76 channel=80
					-5, -4, 6, 2, 1, 4, -3, -6, 2,
					-- layer=2 filter=76 channel=81
					5, 5, -9, -2, 6, 10, 4, 2, 3,
					-- layer=2 filter=76 channel=82
					2, -4, 9, 0, 8, 8, -3, 4, 5,
					-- layer=2 filter=76 channel=83
					0, -6, -2, 0, 5, -6, -10, -11, -9,
					-- layer=2 filter=76 channel=84
					4, -7, 4, 0, 8, -6, 3, 2, -3,
					-- layer=2 filter=76 channel=85
					-3, -10, -6, 7, -6, -1, 3, 5, 11,
					-- layer=2 filter=76 channel=86
					-15, -13, -15, 2, -14, 4, -14, 0, -2,
					-- layer=2 filter=76 channel=87
					5, -2, 1, 0, -7, -16, -6, -10, 3,
					-- layer=2 filter=76 channel=88
					-6, -6, 0, 4, -14, -12, -7, 0, 0,
					-- layer=2 filter=76 channel=89
					-15, -5, -20, -6, 3, -10, 2, -6, 2,
					-- layer=2 filter=76 channel=90
					-5, 6, 4, -9, 0, -1, 0, 2, -7,
					-- layer=2 filter=76 channel=91
					-8, -4, -20, 0, 2, -5, 0, -6, 4,
					-- layer=2 filter=76 channel=92
					0, -18, -12, 1, -10, 0, 7, 7, 5,
					-- layer=2 filter=76 channel=93
					-8, 0, -9, -4, 3, -6, -6, 3, -3,
					-- layer=2 filter=76 channel=94
					-2, 0, 1, -2, -10, 3, -12, 0, 6,
					-- layer=2 filter=76 channel=95
					4, -2, -8, -9, 0, -3, -1, 0, -5,
					-- layer=2 filter=76 channel=96
					7, -2, 1, -5, -15, -4, -18, -14, -15,
					-- layer=2 filter=76 channel=97
					5, -6, 5, 8, -16, -13, -12, -11, -11,
					-- layer=2 filter=76 channel=98
					-12, 8, 0, -4, 1, -5, -7, -14, -18,
					-- layer=2 filter=76 channel=99
					-13, -5, -6, -6, -14, -6, 2, -2, -9,
					-- layer=2 filter=76 channel=100
					-8, 0, -12, -8, 3, -9, -6, 4, -7,
					-- layer=2 filter=76 channel=101
					-9, -15, -3, -18, -4, -6, -10, -14, -18,
					-- layer=2 filter=76 channel=102
					-2, -4, 4, -10, -12, 5, -10, -7, -11,
					-- layer=2 filter=76 channel=103
					0, 9, -10, -8, 6, 6, 8, -5, 1,
					-- layer=2 filter=76 channel=104
					-9, 3, -12, -3, -6, -3, -12, 0, 6,
					-- layer=2 filter=76 channel=105
					5, -6, -2, -3, -4, -11, -10, 4, 5,
					-- layer=2 filter=76 channel=106
					2, -13, -10, -5, -11, -14, -5, -5, 3,
					-- layer=2 filter=76 channel=107
					2, -1, -6, -5, 6, -7, -8, -3, 4,
					-- layer=2 filter=76 channel=108
					-7, 0, 1, -2, -10, -4, -6, 1, 4,
					-- layer=2 filter=76 channel=109
					9, 10, 10, 4, -4, -9, 8, 5, -9,
					-- layer=2 filter=76 channel=110
					-1, -5, 8, -3, 0, -13, -11, -8, 2,
					-- layer=2 filter=76 channel=111
					-7, 1, -1, 6, 0, 6, -5, -4, -2,
					-- layer=2 filter=76 channel=112
					-15, -11, -8, -7, -10, -2, -5, -3, -9,
					-- layer=2 filter=76 channel=113
					-11, -8, 0, -9, 2, 2, -13, 0, -5,
					-- layer=2 filter=76 channel=114
					-2, 0, -6, 8, 0, -6, 9, -9, -7,
					-- layer=2 filter=76 channel=115
					6, 1, -1, 6, -5, -4, -2, 4, -1,
					-- layer=2 filter=76 channel=116
					-1, -11, -6, 2, -7, -8, -10, 3, 2,
					-- layer=2 filter=76 channel=117
					-14, 5, 2, -2, -1, 4, 2, 0, -7,
					-- layer=2 filter=76 channel=118
					6, 7, -9, 5, 3, -16, 1, -11, 3,
					-- layer=2 filter=76 channel=119
					4, -9, -9, -10, -10, -11, 0, -2, 0,
					-- layer=2 filter=76 channel=120
					9, 8, -1, 9, 10, -2, 0, 5, 1,
					-- layer=2 filter=76 channel=121
					-1, -3, -6, -1, -8, -6, -11, -2, 0,
					-- layer=2 filter=76 channel=122
					6, 3, -4, 0, 2, 2, 6, 3, 5,
					-- layer=2 filter=76 channel=123
					-18, -6, -8, 0, 8, 0, 9, 6, -7,
					-- layer=2 filter=76 channel=124
					-1, 2, -10, -7, 2, -9, -6, 4, -1,
					-- layer=2 filter=76 channel=125
					0, 6, -5, -5, -1, -1, -10, 1, -5,
					-- layer=2 filter=76 channel=126
					-1, -3, 5, -3, 8, -6, 4, 9, -10,
					-- layer=2 filter=76 channel=127
					-9, -1, 2, -1, -11, 4, -7, -7, 2,
					-- layer=2 filter=77 channel=0
					12, 18, 35, -7, -31, -2, 19, -3, 4,
					-- layer=2 filter=77 channel=1
					19, -21, -2, -43, -23, -14, 2, -9, -20,
					-- layer=2 filter=77 channel=2
					-2, 10, 7, 10, 7, -5, 10, -5, -9,
					-- layer=2 filter=77 channel=3
					-26, -3, 0, 10, -3, -25, 6, 2, -29,
					-- layer=2 filter=77 channel=4
					3, 52, 48, -29, 27, 0, -27, -24, -45,
					-- layer=2 filter=77 channel=5
					55, 26, 34, 16, -19, -9, -50, -31, -13,
					-- layer=2 filter=77 channel=6
					5, -5, 6, -10, -56, 26, 0, -24, 15,
					-- layer=2 filter=77 channel=7
					-4, 3, 18, 15, 29, 30, 22, 27, 15,
					-- layer=2 filter=77 channel=8
					-5, -6, -4, 2, 4, -4, 8, 8, -8,
					-- layer=2 filter=77 channel=9
					21, 30, -13, -44, -13, 16, -39, -17, -41,
					-- layer=2 filter=77 channel=10
					-11, 8, 32, 15, 10, 28, 21, -38, -5,
					-- layer=2 filter=77 channel=11
					-12, 21, 3, -21, 6, -10, -24, 14, 3,
					-- layer=2 filter=77 channel=12
					15, 9, 26, -11, -14, -19, 8, 10, -19,
					-- layer=2 filter=77 channel=13
					-1, 9, -9, -8, 8, -8, -3, -11, -1,
					-- layer=2 filter=77 channel=14
					-7, -3, -19, -21, -4, -14, 1, 35, 29,
					-- layer=2 filter=77 channel=15
					55, -3, 23, -21, 44, -24, 0, 0, -46,
					-- layer=2 filter=77 channel=16
					36, 12, 0, 13, -1, -29, -10, -43, -18,
					-- layer=2 filter=77 channel=17
					-10, -3, -3, -2, -6, 9, 2, -8, -1,
					-- layer=2 filter=77 channel=18
					18, 46, 35, -51, 17, -27, -7, 8, -9,
					-- layer=2 filter=77 channel=19
					-37, -62, -22, -10, 22, -6, -20, -27, -29,
					-- layer=2 filter=77 channel=20
					0, -4, 9, -3, 4, -6, -4, 6, -4,
					-- layer=2 filter=77 channel=21
					9, -4, -3, -6, -4, 8, -3, 5, 17,
					-- layer=2 filter=77 channel=22
					-5, -9, 4, -7, 7, -2, 8, -2, 0,
					-- layer=2 filter=77 channel=23
					9, -15, 4, 4, 2, 8, 35, 40, 32,
					-- layer=2 filter=77 channel=24
					-39, -19, -31, 3, 19, 14, 40, 35, 34,
					-- layer=2 filter=77 channel=25
					-92, -35, -36, -20, 0, 23, 36, 53, 40,
					-- layer=2 filter=77 channel=26
					3, -10, -5, 0, 4, -6, 2, -4, 10,
					-- layer=2 filter=77 channel=27
					9, 16, 39, 26, 24, 26, -39, -66, -64,
					-- layer=2 filter=77 channel=28
					1, 31, 13, 25, 12, 15, 40, -11, 5,
					-- layer=2 filter=77 channel=29
					4, 10, -8, 6, 8, -9, 7, -6, -2,
					-- layer=2 filter=77 channel=30
					1, 11, 32, -4, 15, 0, -3, -16, 12,
					-- layer=2 filter=77 channel=31
					-34, 0, 14, -9, -17, 63, -32, -53, -71,
					-- layer=2 filter=77 channel=32
					2, -3, 8, -5, 3, 6, 0, 0, 1,
					-- layer=2 filter=77 channel=33
					-22, 7, 1, -39, 0, -32, 3, 9, -20,
					-- layer=2 filter=77 channel=34
					2, -45, -31, -20, -2, -22, 2, -4, 0,
					-- layer=2 filter=77 channel=35
					-50, 10, -18, -29, 8, -9, 12, 23, 9,
					-- layer=2 filter=77 channel=36
					14, 2, 14, -3, 3, 6, -1, -3, 8,
					-- layer=2 filter=77 channel=37
					21, 10, 14, -3, 20, 0, -47, -22, 2,
					-- layer=2 filter=77 channel=38
					1, 27, 20, 0, -26, 7, -73, -40, -11,
					-- layer=2 filter=77 channel=39
					-2, -28, 9, -17, -3, 5, -20, 41, 22,
					-- layer=2 filter=77 channel=40
					-42, 9, -29, -42, 33, -10, 2, 21, 4,
					-- layer=2 filter=77 channel=41
					-1, 2, 1, 3, -3, 0, 0, 0, 8,
					-- layer=2 filter=77 channel=42
					9, -32, 10, 24, -15, 7, 35, 59, 21,
					-- layer=2 filter=77 channel=43
					20, 33, 43, 8, 35, -14, -52, -39, -40,
					-- layer=2 filter=77 channel=44
					0, 1, 9, -10, 3, -5, -3, 2, 1,
					-- layer=2 filter=77 channel=45
					-23, -4, -16, 15, 31, 19, -18, -4, 9,
					-- layer=2 filter=77 channel=46
					-6, 16, 18, -20, 1, 18, 3, -7, 11,
					-- layer=2 filter=77 channel=47
					51, 87, 38, 25, -17, 17, 2, -17, -3,
					-- layer=2 filter=77 channel=48
					-5, 0, 2, 7, -7, 11, -3, 0, 5,
					-- layer=2 filter=77 channel=49
					36, 43, 37, 5, 52, 41, 0, 71, 22,
					-- layer=2 filter=77 channel=50
					18, 4, 11, 21, 0, 10, 1, 10, 11,
					-- layer=2 filter=77 channel=51
					36, 37, 6, -10, -9, -8, -21, -17, 6,
					-- layer=2 filter=77 channel=52
					40, 22, 1, -41, -45, -38, -41, -20, -27,
					-- layer=2 filter=77 channel=53
					40, -28, -3, -42, -29, 3, -12, 28, -17,
					-- layer=2 filter=77 channel=54
					-40, -36, 26, -10, -33, -37, 20, 22, -5,
					-- layer=2 filter=77 channel=55
					-15, 9, -2, 5, 12, 13, -8, 4, -4,
					-- layer=2 filter=77 channel=56
					17, 29, 43, -1, 0, 17, -36, -9, 10,
					-- layer=2 filter=77 channel=57
					0, 7, -7, -13, -8, 0, 2, 1, 9,
					-- layer=2 filter=77 channel=58
					-18, -12, 35, -16, 12, -12, -14, 9, 14,
					-- layer=2 filter=77 channel=59
					18, -16, -10, 22, 0, -3, -34, -55, -81,
					-- layer=2 filter=77 channel=60
					-18, -15, 38, -7, -22, 1, 43, 17, 4,
					-- layer=2 filter=77 channel=61
					31, 14, 0, 7, -29, 22, 29, -4, 33,
					-- layer=2 filter=77 channel=62
					-14, -29, 28, -3, -18, 11, 37, -1, 0,
					-- layer=2 filter=77 channel=63
					19, -6, -5, 14, 20, 0, 21, 22, -12,
					-- layer=2 filter=77 channel=64
					6, -19, -4, 7, 7, -5, 43, 36, 16,
					-- layer=2 filter=77 channel=65
					20, 10, 10, -9, -39, 8, 1, -52, -5,
					-- layer=2 filter=77 channel=66
					42, 6, 24, -13, 7, -36, 40, 0, 17,
					-- layer=2 filter=77 channel=67
					20, 10, 23, -16, 2, -15, 3, -25, -8,
					-- layer=2 filter=77 channel=68
					6, -2, -7, -5, -5, -3, -10, -7, -10,
					-- layer=2 filter=77 channel=69
					15, -22, -8, -3, 11, 20, 15, 23, 25,
					-- layer=2 filter=77 channel=70
					-64, 11, 11, -23, -11, 5, 0, -9, 1,
					-- layer=2 filter=77 channel=71
					-16, -32, -18, 17, 58, 21, -26, -20, -6,
					-- layer=2 filter=77 channel=72
					-2, -2, -22, -1, 2, 6, 21, 11, 27,
					-- layer=2 filter=77 channel=73
					69, 16, 11, 69, 60, 90, 51, 57, 30,
					-- layer=2 filter=77 channel=74
					-13, -5, 9, -7, -8, 2, 32, -6, 4,
					-- layer=2 filter=77 channel=75
					-18, -21, -36, -42, -31, 3, 0, 18, 23,
					-- layer=2 filter=77 channel=76
					28, 0, -7, -68, -41, 12, -27, -38, -10,
					-- layer=2 filter=77 channel=77
					-1, 3, 9, 3, 0, 0, -10, 5, 5,
					-- layer=2 filter=77 channel=78
					2, -21, -8, 12, -18, -6, 9, 42, 2,
					-- layer=2 filter=77 channel=79
					-6, -3, -3, 3, 7, 8, -3, 0, -8,
					-- layer=2 filter=77 channel=80
					33, 6, 23, 3, -2, -2, -21, -20, -40,
					-- layer=2 filter=77 channel=81
					0, 8, -9, 2, -8, 0, 10, -4, -3,
					-- layer=2 filter=77 channel=82
					-7, 8, 8, 7, -10, 8, -6, 11, -4,
					-- layer=2 filter=77 channel=83
					-8, -13, 9, -13, -2, -1, 10, -1, -22,
					-- layer=2 filter=77 channel=84
					-2, 9, -6, -5, -2, 3, -9, 3, -7,
					-- layer=2 filter=77 channel=85
					-8, 10, 8, 11, -11, -14, 10, 6, -6,
					-- layer=2 filter=77 channel=86
					-17, -5, -14, -12, -12, -24, -1, 6, -2,
					-- layer=2 filter=77 channel=87
					-23, -1, 14, -13, -22, -12, -28, 15, 29,
					-- layer=2 filter=77 channel=88
					3, -11, -8, -6, -15, -2, 17, 1, 3,
					-- layer=2 filter=77 channel=89
					-5, -4, -24, -12, -2, -36, 37, 36, 4,
					-- layer=2 filter=77 channel=90
					-2, 1, -8, 1, -1, -3, -3, 5, 7,
					-- layer=2 filter=77 channel=91
					0, -19, 24, 0, -32, -9, 40, 18, -9,
					-- layer=2 filter=77 channel=92
					18, -3, 3, -46, -31, -11, -10, 13, 3,
					-- layer=2 filter=77 channel=93
					-14, -51, 52, -15, -44, 18, -15, -103, -46,
					-- layer=2 filter=77 channel=94
					39, -9, 34, -6, -66, 13, 10, 0, -37,
					-- layer=2 filter=77 channel=95
					9, -5, 0, 12, -1, 0, 9, -10, -1,
					-- layer=2 filter=77 channel=96
					38, -25, -12, 0, -80, -73, 31, -13, -58,
					-- layer=2 filter=77 channel=97
					7, 18, -26, -12, 8, 5, -17, 21, -23,
					-- layer=2 filter=77 channel=98
					5, 33, 33, 13, 21, 11, 6, 10, 17,
					-- layer=2 filter=77 channel=99
					19, -10, -1, 1, 5, -5, -31, -34, 6,
					-- layer=2 filter=77 channel=100
					-24, 18, 23, -5, -19, 9, 8, -21, -54,
					-- layer=2 filter=77 channel=101
					-54, -47, -66, -16, 48, 25, -49, -15, -21,
					-- layer=2 filter=77 channel=102
					32, 4, 32, -61, -7, 0, -11, -9, -22,
					-- layer=2 filter=77 channel=103
					0, 11, 26, -55, -53, 33, -24, -35, -51,
					-- layer=2 filter=77 channel=104
					40, 5, 56, -19, 20, -15, -6, 13, 15,
					-- layer=2 filter=77 channel=105
					8, -5, -45, 19, 24, -25, 19, -5, 30,
					-- layer=2 filter=77 channel=106
					-57, -31, -23, -21, 5, 0, 7, -1, 4,
					-- layer=2 filter=77 channel=107
					-43, 13, 7, -29, -23, 24, -48, -17, 26,
					-- layer=2 filter=77 channel=108
					1, 17, -5, 6, 4, -9, -33, -57, -63,
					-- layer=2 filter=77 channel=109
					5, 8, 12, 10, -11, -1, 0, -5, 11,
					-- layer=2 filter=77 channel=110
					-28, -22, -34, -8, -17, -10, 66, 78, 64,
					-- layer=2 filter=77 channel=111
					7, -5, 5, 7, -9, -5, -6, 6, 11,
					-- layer=2 filter=77 channel=112
					-4, 20, 32, -2, 6, 2, 16, 1, 22,
					-- layer=2 filter=77 channel=113
					4, -7, 42, -22, 36, -11, 0, 12, 7,
					-- layer=2 filter=77 channel=114
					3, -1, 7, -3, -15, -4, -20, 2, 6,
					-- layer=2 filter=77 channel=115
					-1, 5, 0, -2, 9, -4, -8, -5, -5,
					-- layer=2 filter=77 channel=116
					6, 0, 18, -59, -13, -40, -26, -15, -11,
					-- layer=2 filter=77 channel=117
					-23, -22, 8, -5, 23, 17, -5, -17, -25,
					-- layer=2 filter=77 channel=118
					37, 54, 29, 27, 20, 4, -11, -13, -11,
					-- layer=2 filter=77 channel=119
					0, 32, 5, -19, 1, 16, 26, -4, -31,
					-- layer=2 filter=77 channel=120
					-5, 4, -4, 5, -4, 5, 0, 0, -7,
					-- layer=2 filter=77 channel=121
					-8, 0, 6, 3, -5, -4, 3, 7, 1,
					-- layer=2 filter=77 channel=122
					0, -1, -8, -6, -6, -18, 9, -8, 0,
					-- layer=2 filter=77 channel=123
					0, 22, 8, -4, 14, 15, -4, 7, -8,
					-- layer=2 filter=77 channel=124
					-24, -42, -13, 1, -28, -12, -7, -27, -1,
					-- layer=2 filter=77 channel=125
					4, -4, 7, -4, -6, -11, 2, -5, -1,
					-- layer=2 filter=77 channel=126
					42, 28, -15, -1, -35, 13, 21, -33, -5,
					-- layer=2 filter=77 channel=127
					8, -23, -31, -53, -1, -17, 3, -33, 4,
					-- layer=2 filter=78 channel=0
					-1, -3, 0, 3, -8, -5, 3, 9, -8,
					-- layer=2 filter=78 channel=1
					-11, -10, 2, -1, 1, -2, -13, -11, -19,
					-- layer=2 filter=78 channel=2
					-3, 4, 0, 8, -3, 5, -2, 5, 6,
					-- layer=2 filter=78 channel=3
					-9, 5, 1, -4, -9, -8, -17, -13, -3,
					-- layer=2 filter=78 channel=4
					0, -8, -14, -2, 0, 1, -2, -11, -7,
					-- layer=2 filter=78 channel=5
					-8, 1, -5, -3, -6, -5, -17, -2, -6,
					-- layer=2 filter=78 channel=6
					0, -10, -10, -12, 9, 10, -16, 4, -6,
					-- layer=2 filter=78 channel=7
					-7, -4, -4, -5, -11, 6, -23, -8, 4,
					-- layer=2 filter=78 channel=8
					11, 2, -4, -2, -10, -6, -7, 7, -7,
					-- layer=2 filter=78 channel=9
					-4, 1, 0, 7, -5, -2, -6, -10, 3,
					-- layer=2 filter=78 channel=10
					-4, -1, -1, 0, -9, 1, -3, -5, 4,
					-- layer=2 filter=78 channel=11
					-11, -4, -5, -5, -5, 5, -10, -5, -6,
					-- layer=2 filter=78 channel=12
					-6, -9, -15, -14, -13, -7, -18, -17, -1,
					-- layer=2 filter=78 channel=13
					10, -1, 2, -6, 1, 0, 11, 10, -7,
					-- layer=2 filter=78 channel=14
					-2, 5, -5, -5, 4, 5, -8, 7, -3,
					-- layer=2 filter=78 channel=15
					0, -10, -6, 3, -8, -9, 7, -3, 5,
					-- layer=2 filter=78 channel=16
					-2, 5, -7, -6, 1, -1, 2, 3, -2,
					-- layer=2 filter=78 channel=17
					0, 1, 10, -1, 6, -8, -11, 5, -3,
					-- layer=2 filter=78 channel=18
					-4, -3, -12, 5, -20, -3, -17, -15, 0,
					-- layer=2 filter=78 channel=19
					-4, -4, -16, -7, -2, 1, -6, -10, -11,
					-- layer=2 filter=78 channel=20
					-10, 4, 9, 6, -4, 0, 3, 9, 2,
					-- layer=2 filter=78 channel=21
					-8, -8, 6, -3, 0, -5, -8, 2, 2,
					-- layer=2 filter=78 channel=22
					2, 3, -2, 5, -2, -4, -3, 8, 7,
					-- layer=2 filter=78 channel=23
					-14, 0, -18, -17, -2, -6, -9, 6, 1,
					-- layer=2 filter=78 channel=24
					0, -5, 8, 3, 0, -13, -10, 2, -3,
					-- layer=2 filter=78 channel=25
					-7, -13, -15, -7, -5, 1, -5, 2, 8,
					-- layer=2 filter=78 channel=26
					6, -7, 3, 3, -1, 6, 9, 8, 6,
					-- layer=2 filter=78 channel=27
					-10, -6, -6, -13, -11, 1, 0, -11, -9,
					-- layer=2 filter=78 channel=28
					-9, -10, -4, -24, -16, -2, -4, -12, 9,
					-- layer=2 filter=78 channel=29
					-1, -7, -6, 4, 1, -1, 3, -5, 4,
					-- layer=2 filter=78 channel=30
					-1, 5, -6, -7, -11, -7, -10, 0, 3,
					-- layer=2 filter=78 channel=31
					9, 2, -7, -9, -2, 10, -2, 3, 10,
					-- layer=2 filter=78 channel=32
					-12, -7, 5, 1, -5, 7, -9, -5, -1,
					-- layer=2 filter=78 channel=33
					3, -16, 6, 0, 5, -14, -12, 1, 0,
					-- layer=2 filter=78 channel=34
					-6, -4, -5, -2, -13, 9, 4, -12, 5,
					-- layer=2 filter=78 channel=35
					0, 9, -14, -4, -12, -5, -8, -9, -10,
					-- layer=2 filter=78 channel=36
					-1, 1, -2, -2, 4, -9, -8, -2, -11,
					-- layer=2 filter=78 channel=37
					-10, -4, -11, 1, -2, 6, 1, 3, -11,
					-- layer=2 filter=78 channel=38
					1, -5, 7, 1, -2, -7, -1, 0, 1,
					-- layer=2 filter=78 channel=39
					3, 2, -12, 2, -5, 5, -3, -2, -4,
					-- layer=2 filter=78 channel=40
					-9, -5, -9, 5, 1, 0, 7, -7, -8,
					-- layer=2 filter=78 channel=41
					5, 1, 0, 8, 3, -8, 8, 10, 11,
					-- layer=2 filter=78 channel=42
					0, 4, -7, 4, -6, 3, 8, -3, -1,
					-- layer=2 filter=78 channel=43
					-2, 2, 2, -11, 0, 0, 0, -9, 3,
					-- layer=2 filter=78 channel=44
					7, -3, 7, 6, -1, -1, 7, -6, 0,
					-- layer=2 filter=78 channel=45
					-2, 4, -5, -2, 4, 2, -9, 6, 5,
					-- layer=2 filter=78 channel=46
					6, -9, -7, 9, -6, 1, -8, 7, -7,
					-- layer=2 filter=78 channel=47
					12, -8, 0, 0, 14, -15, -4, 9, 5,
					-- layer=2 filter=78 channel=48
					7, -4, 1, -7, 5, -6, -3, 7, -5,
					-- layer=2 filter=78 channel=49
					-2, -15, -3, -10, -13, -8, 0, -18, -20,
					-- layer=2 filter=78 channel=50
					0, 5, 2, -8, -2, 8, -9, 10, -2,
					-- layer=2 filter=78 channel=51
					-2, -6, 2, -14, -14, -10, 0, 3, -2,
					-- layer=2 filter=78 channel=52
					0, -5, -12, -2, 0, -13, -11, -2, 0,
					-- layer=2 filter=78 channel=53
					-8, -9, 8, -3, -3, 1, -8, -5, 7,
					-- layer=2 filter=78 channel=54
					-7, -1, 0, 1, 0, -4, -24, -4, -3,
					-- layer=2 filter=78 channel=55
					-6, 1, -5, -3, 8, -7, 3, -8, 2,
					-- layer=2 filter=78 channel=56
					7, 3, -3, 5, -1, 4, -1, -1, 5,
					-- layer=2 filter=78 channel=57
					0, -4, 3, -3, -7, 3, -3, -1, 5,
					-- layer=2 filter=78 channel=58
					4, -3, 0, -10, -12, 4, -7, 0, -20,
					-- layer=2 filter=78 channel=59
					-8, -12, 7, -7, -9, 0, -5, 4, -9,
					-- layer=2 filter=78 channel=60
					-5, 4, 9, -8, 6, 1, -6, -1, 6,
					-- layer=2 filter=78 channel=61
					-1, 12, -8, -11, -13, 0, -6, 3, 8,
					-- layer=2 filter=78 channel=62
					3, 7, 0, -8, -10, 0, -22, -3, 5,
					-- layer=2 filter=78 channel=63
					-4, -2, -3, -3, -1, 0, 0, -4, -5,
					-- layer=2 filter=78 channel=64
					4, 0, -2, 1, -8, 3, 8, 4, 7,
					-- layer=2 filter=78 channel=65
					-5, -2, 4, -11, 5, 5, -2, -10, 5,
					-- layer=2 filter=78 channel=66
					-6, 1, 0, -3, -4, -2, 1, -5, -7,
					-- layer=2 filter=78 channel=67
					-3, -1, 2, 1, -9, -1, 1, -3, -12,
					-- layer=2 filter=78 channel=68
					7, 11, 4, 3, 11, -6, -6, 7, 2,
					-- layer=2 filter=78 channel=69
					2, -8, -14, -4, -15, -10, -11, -3, -3,
					-- layer=2 filter=78 channel=70
					-7, 0, -16, -7, -12, -1, -10, -8, -12,
					-- layer=2 filter=78 channel=71
					3, 8, -6, 7, -8, 5, 8, 4, 0,
					-- layer=2 filter=78 channel=72
					-16, -5, 1, 0, -2, -13, -18, -24, -5,
					-- layer=2 filter=78 channel=73
					-11, -13, -4, -17, 0, -13, -9, -13, 0,
					-- layer=2 filter=78 channel=74
					4, -4, 5, 3, 8, -2, -3, -5, -2,
					-- layer=2 filter=78 channel=75
					0, 5, 0, 6, 10, 0, -7, -3, -6,
					-- layer=2 filter=78 channel=76
					0, 7, -5, 10, -3, 3, 7, -1, 6,
					-- layer=2 filter=78 channel=77
					-3, -4, 2, -3, -10, 10, 0, 2, -9,
					-- layer=2 filter=78 channel=78
					8, 0, -5, -3, 1, -2, -9, -11, -8,
					-- layer=2 filter=78 channel=79
					-6, 5, -2, -7, 4, 7, 8, -6, -3,
					-- layer=2 filter=78 channel=80
					-9, 5, -6, -9, -8, -4, -6, 8, 0,
					-- layer=2 filter=78 channel=81
					0, 9, 10, 2, 8, -5, 3, 6, 5,
					-- layer=2 filter=78 channel=82
					-5, 0, 7, 2, 6, 0, 7, 9, 0,
					-- layer=2 filter=78 channel=83
					-2, 2, -10, 8, -1, 4, -5, 3, 5,
					-- layer=2 filter=78 channel=84
					6, -8, 11, -7, -2, 4, 2, 8, -4,
					-- layer=2 filter=78 channel=85
					-9, -3, 0, 0, 8, -8, -4, -6, -6,
					-- layer=2 filter=78 channel=86
					4, 4, 5, 5, 7, -3, 10, 0, 4,
					-- layer=2 filter=78 channel=87
					-3, -6, 0, 2, -11, 2, 7, -2, -4,
					-- layer=2 filter=78 channel=88
					-12, -6, 3, -7, -12, -2, -8, -8, -7,
					-- layer=2 filter=78 channel=89
					-5, -11, 4, -15, -13, 1, -7, -2, -9,
					-- layer=2 filter=78 channel=90
					-8, -5, -5, 6, 4, 3, -8, 7, -4,
					-- layer=2 filter=78 channel=91
					-12, -7, -26, -18, -1, 1, -11, 0, -8,
					-- layer=2 filter=78 channel=92
					-8, -12, -14, -18, -1, -14, -12, -13, -11,
					-- layer=2 filter=78 channel=93
					-9, -3, 2, -4, -10, 5, -3, -8, -9,
					-- layer=2 filter=78 channel=94
					-23, 0, -5, -3, 3, 2, -16, -16, -1,
					-- layer=2 filter=78 channel=95
					-8, -5, -3, -4, -5, -2, -2, -1, -8,
					-- layer=2 filter=78 channel=96
					-6, 1, 14, -10, -16, -12, -13, -11, 11,
					-- layer=2 filter=78 channel=97
					0, 0, 4, 3, 0, -3, 2, -9, 0,
					-- layer=2 filter=78 channel=98
					-16, -10, -10, -4, 7, 0, 0, -4, -4,
					-- layer=2 filter=78 channel=99
					-11, -5, -12, -9, 0, -5, 0, -8, -8,
					-- layer=2 filter=78 channel=100
					-15, -14, -4, 4, -8, 0, -11, 7, -5,
					-- layer=2 filter=78 channel=101
					-8, 2, -7, -5, 0, 0, 3, 2, -1,
					-- layer=2 filter=78 channel=102
					-9, -15, 4, 6, -5, -20, 2, 2, -16,
					-- layer=2 filter=78 channel=103
					10, 6, -1, -3, 1, 3, -9, -7, -5,
					-- layer=2 filter=78 channel=104
					-2, -6, -3, -12, -1, -9, -1, -13, 0,
					-- layer=2 filter=78 channel=105
					-2, -4, -9, 5, 7, -6, 8, 0, -1,
					-- layer=2 filter=78 channel=106
					-14, -7, -3, -10, -13, -5, 0, 11, 10,
					-- layer=2 filter=78 channel=107
					0, -4, -1, -4, 6, 9, 7, 2, 1,
					-- layer=2 filter=78 channel=108
					-4, 0, 9, 5, -6, 0, -10, -7, -9,
					-- layer=2 filter=78 channel=109
					6, -2, -6, 8, -3, -4, 9, 11, -8,
					-- layer=2 filter=78 channel=110
					-15, -9, 2, -5, 4, -10, -2, -1, -9,
					-- layer=2 filter=78 channel=111
					5, -4, -1, 4, 7, -2, 10, 8, -6,
					-- layer=2 filter=78 channel=112
					-6, 4, -6, -8, 0, -3, -5, -1, 5,
					-- layer=2 filter=78 channel=113
					-1, 0, -9, 1, -2, -12, -5, -10, -5,
					-- layer=2 filter=78 channel=114
					4, -5, 2, 1, 0, -9, -7, 1, 4,
					-- layer=2 filter=78 channel=115
					-1, 6, 0, -8, 0, -3, 1, 3, 1,
					-- layer=2 filter=78 channel=116
					-15, 0, -11, -1, 6, -9, -16, -13, 2,
					-- layer=2 filter=78 channel=117
					-6, -5, -6, -9, -4, -16, -15, 1, 13,
					-- layer=2 filter=78 channel=118
					-6, 6, 1, 8, -4, -2, -3, 1, -6,
					-- layer=2 filter=78 channel=119
					0, -3, -8, -3, -8, -4, -13, -11, -6,
					-- layer=2 filter=78 channel=120
					-5, -1, -1, 5, 9, -9, 8, -1, -6,
					-- layer=2 filter=78 channel=121
					0, -1, 3, 7, 2, 0, 9, 8, -8,
					-- layer=2 filter=78 channel=122
					-7, 4, 6, 9, 10, -10, 2, 4, 3,
					-- layer=2 filter=78 channel=123
					-15, 1, 5, 0, -17, 0, -11, -8, 0,
					-- layer=2 filter=78 channel=124
					3, -4, -5, -10, 0, -7, 0, -8, 1,
					-- layer=2 filter=78 channel=125
					10, -2, 0, 2, 9, -3, -5, 5, -8,
					-- layer=2 filter=78 channel=126
					-9, 9, -7, 8, 8, -4, -6, 5, -9,
					-- layer=2 filter=78 channel=127
					1, -7, -12, 0, -12, -11, 6, 2, 4,
					-- layer=2 filter=79 channel=0
					-8, -5, -9, -6, -12, -1, -7, -5, -4,
					-- layer=2 filter=79 channel=1
					-14, -2, -13, -3, -14, -11, 1, 2, -4,
					-- layer=2 filter=79 channel=2
					5, -8, 6, 5, 5, 8, -2, 9, -4,
					-- layer=2 filter=79 channel=3
					8, -8, 8, -5, 5, 7, 7, 2, -13,
					-- layer=2 filter=79 channel=4
					7, 2, 0, -6, 2, 0, 5, -6, -2,
					-- layer=2 filter=79 channel=5
					-10, -15, 4, -2, -1, -1, 2, 3, -9,
					-- layer=2 filter=79 channel=6
					2, -7, 8, 5, -10, -4, 3, 6, 3,
					-- layer=2 filter=79 channel=7
					-10, -3, 6, 1, 0, 2, 7, 12, -4,
					-- layer=2 filter=79 channel=8
					7, 0, 3, 8, 0, 7, -4, -4, 9,
					-- layer=2 filter=79 channel=9
					-4, 5, 3, 6, 0, -11, 4, -8, -3,
					-- layer=2 filter=79 channel=10
					-3, -10, -3, 8, 6, 5, -4, -11, -8,
					-- layer=2 filter=79 channel=11
					1, -12, 0, 2, -3, -13, 2, -10, 5,
					-- layer=2 filter=79 channel=12
					-1, 7, -2, -9, 4, 0, -10, -10, -7,
					-- layer=2 filter=79 channel=13
					-1, 0, 2, -7, 0, -6, 7, -11, -10,
					-- layer=2 filter=79 channel=14
					-7, 3, 5, 6, -5, -14, -1, 3, 1,
					-- layer=2 filter=79 channel=15
					-7, 5, 3, 0, 0, -5, 3, -2, 1,
					-- layer=2 filter=79 channel=16
					-10, 7, 6, -9, 3, -3, 1, 0, -2,
					-- layer=2 filter=79 channel=17
					-1, 5, 6, -4, -5, 1, -4, -6, 8,
					-- layer=2 filter=79 channel=18
					-1, -1, -15, 2, 4, -7, 3, -3, -9,
					-- layer=2 filter=79 channel=19
					-2, 4, 5, -5, 0, -8, -2, -5, -8,
					-- layer=2 filter=79 channel=20
					-10, 5, 6, 8, 5, -6, 5, 1, 1,
					-- layer=2 filter=79 channel=21
					11, -9, 0, 0, 1, 0, 4, 5, 7,
					-- layer=2 filter=79 channel=22
					-5, 9, -1, 7, 1, -9, 3, 0, -3,
					-- layer=2 filter=79 channel=23
					-12, -12, -9, 1, -6, -10, -7, -3, -2,
					-- layer=2 filter=79 channel=24
					-4, -4, 4, -9, 6, 8, -5, 8, 0,
					-- layer=2 filter=79 channel=25
					-13, -5, 4, 5, -5, 0, -1, -9, -5,
					-- layer=2 filter=79 channel=26
					1, -8, -10, -8, 1, -2, 3, 0, -6,
					-- layer=2 filter=79 channel=27
					1, 3, -13, 0, 6, -10, -5, -3, -7,
					-- layer=2 filter=79 channel=28
					5, -13, -5, -9, -10, -4, 2, 1, -15,
					-- layer=2 filter=79 channel=29
					5, 7, 3, -12, -11, -10, -12, 1, 3,
					-- layer=2 filter=79 channel=30
					-10, 1, 3, -11, 0, -4, 6, 2, -2,
					-- layer=2 filter=79 channel=31
					-6, 4, -5, 5, -5, -7, -9, -9, -3,
					-- layer=2 filter=79 channel=32
					-11, 8, -12, 0, 0, -4, -7, 0, -2,
					-- layer=2 filter=79 channel=33
					5, 2, -1, 3, 3, -11, 6, 2, -6,
					-- layer=2 filter=79 channel=34
					-3, -6, 3, -1, 7, -5, 2, -9, 6,
					-- layer=2 filter=79 channel=35
					-2, 0, -7, -12, -1, 0, -7, -10, 1,
					-- layer=2 filter=79 channel=36
					-8, -11, 4, -8, 6, 4, -8, -10, -6,
					-- layer=2 filter=79 channel=37
					3, -8, -12, -10, 0, 6, -3, 0, 3,
					-- layer=2 filter=79 channel=38
					-5, -11, 5, -5, -7, 3, -3, -12, -7,
					-- layer=2 filter=79 channel=39
					-3, -10, 9, -7, -9, -3, -1, -6, 3,
					-- layer=2 filter=79 channel=40
					-7, 2, -2, -9, -3, -8, -6, -13, 11,
					-- layer=2 filter=79 channel=41
					5, 0, -6, 9, 11, -1, -6, -6, -8,
					-- layer=2 filter=79 channel=42
					2, -9, 7, 8, 4, 0, 7, 7, -13,
					-- layer=2 filter=79 channel=43
					6, 7, 3, -11, 3, 1, -10, -9, -1,
					-- layer=2 filter=79 channel=44
					1, -10, -5, 0, -2, 8, -6, -9, 9,
					-- layer=2 filter=79 channel=45
					-8, 7, 4, 2, 4, -9, 3, -10, 1,
					-- layer=2 filter=79 channel=46
					-3, -7, -6, 2, -9, -5, -9, 1, 9,
					-- layer=2 filter=79 channel=47
					-10, 0, 6, -13, 7, -5, -8, -2, 7,
					-- layer=2 filter=79 channel=48
					2, 10, 3, 6, -4, -7, 5, -4, 10,
					-- layer=2 filter=79 channel=49
					2, -6, -4, -11, -8, -6, -1, 2, -1,
					-- layer=2 filter=79 channel=50
					-9, 5, 10, -3, -7, -1, -6, 6, -10,
					-- layer=2 filter=79 channel=51
					-2, -7, 0, -2, -10, -1, 7, -4, -10,
					-- layer=2 filter=79 channel=52
					-12, -5, 4, 2, -11, -2, -6, -9, -11,
					-- layer=2 filter=79 channel=53
					3, 2, 8, -7, 1, -6, 2, -6, 9,
					-- layer=2 filter=79 channel=54
					-7, 3, -12, 4, -9, -7, 1, -11, -2,
					-- layer=2 filter=79 channel=55
					0, -2, 7, -6, 3, -9, -11, -9, -6,
					-- layer=2 filter=79 channel=56
					-3, 5, 3, -3, -5, -11, -5, 4, 1,
					-- layer=2 filter=79 channel=57
					9, 2, -6, 6, -1, -4, -6, -2, -12,
					-- layer=2 filter=79 channel=58
					-2, 6, 0, 0, 4, 1, -10, -7, -10,
					-- layer=2 filter=79 channel=59
					-10, -5, -8, -7, -10, -6, -6, 4, 0,
					-- layer=2 filter=79 channel=60
					-9, 8, -4, 7, -14, 1, 4, 0, -10,
					-- layer=2 filter=79 channel=61
					1, 5, -5, 0, 0, 3, -10, -4, -6,
					-- layer=2 filter=79 channel=62
					-8, -6, 4, -17, 0, -8, -8, 5, -14,
					-- layer=2 filter=79 channel=63
					-12, 2, 1, 1, 7, -7, -6, 6, -4,
					-- layer=2 filter=79 channel=64
					8, -5, -5, 5, -11, 7, -5, 7, -5,
					-- layer=2 filter=79 channel=65
					-9, -9, -9, -8, 2, -4, 3, -11, 3,
					-- layer=2 filter=79 channel=66
					-8, -11, 11, 8, -10, -2, -9, -2, -2,
					-- layer=2 filter=79 channel=67
					3, 0, 0, -1, 2, 3, -6, -12, -1,
					-- layer=2 filter=79 channel=68
					-7, 5, -7, 2, 2, 0, 1, -11, 4,
					-- layer=2 filter=79 channel=69
					6, 3, 7, -3, 0, -6, -9, 0, -9,
					-- layer=2 filter=79 channel=70
					8, -14, -4, -12, 2, -10, -4, -10, -9,
					-- layer=2 filter=79 channel=71
					-12, -9, -1, -7, 3, -8, 5, 0, 5,
					-- layer=2 filter=79 channel=72
					-10, -14, -1, 1, -5, -10, 2, 0, 0,
					-- layer=2 filter=79 channel=73
					0, -7, 8, 2, -11, 6, -10, 0, 1,
					-- layer=2 filter=79 channel=74
					2, -4, -8, 5, -8, -10, 6, -11, -4,
					-- layer=2 filter=79 channel=75
					-5, 9, -1, -4, -4, -9, -9, -10, 4,
					-- layer=2 filter=79 channel=76
					0, -2, -9, -10, 5, 3, 2, 3, -6,
					-- layer=2 filter=79 channel=77
					-8, 6, -6, 8, 0, 0, -11, 0, 5,
					-- layer=2 filter=79 channel=78
					4, 3, 2, 4, -9, -3, 3, -11, -11,
					-- layer=2 filter=79 channel=79
					-8, 8, -2, -7, 8, -2, -11, -11, -8,
					-- layer=2 filter=79 channel=80
					4, -4, 8, -4, 4, 0, 6, 1, 8,
					-- layer=2 filter=79 channel=81
					-7, -7, 7, 0, -7, -10, -4, -9, 4,
					-- layer=2 filter=79 channel=82
					9, 3, -10, 3, -5, 8, 4, -10, -9,
					-- layer=2 filter=79 channel=83
					0, -1, -8, 5, -8, -2, -7, -4, -1,
					-- layer=2 filter=79 channel=84
					-8, 11, -7, 0, -6, 3, -8, -4, 4,
					-- layer=2 filter=79 channel=85
					-2, 0, 0, 5, -12, -3, -9, -5, 0,
					-- layer=2 filter=79 channel=86
					-11, 0, -2, -1, 6, 2, -6, -2, -4,
					-- layer=2 filter=79 channel=87
					5, -7, -4, -11, -9, 0, 3, 0, 4,
					-- layer=2 filter=79 channel=88
					-3, -8, -5, -10, -1, -7, -8, 4, -7,
					-- layer=2 filter=79 channel=89
					-3, -4, -12, 2, 0, 3, 4, -8, -1,
					-- layer=2 filter=79 channel=90
					2, -1, -4, 7, 2, -9, -4, -1, -6,
					-- layer=2 filter=79 channel=91
					-4, 4, -3, -4, 1, 3, 1, -2, 5,
					-- layer=2 filter=79 channel=92
					-8, -16, 5, -2, -2, 3, -5, 0, 3,
					-- layer=2 filter=79 channel=93
					-5, 3, 0, -16, 6, 0, 0, 3, 3,
					-- layer=2 filter=79 channel=94
					0, -12, 5, -10, 1, -11, -2, -3, 4,
					-- layer=2 filter=79 channel=95
					1, 6, 8, 8, -4, 3, 6, 3, -10,
					-- layer=2 filter=79 channel=96
					-8, -20, -2, -11, -5, -9, 1, 4, 3,
					-- layer=2 filter=79 channel=97
					-1, -5, -11, -9, 0, -11, -1, -8, -9,
					-- layer=2 filter=79 channel=98
					-7, 6, -4, -6, -12, -7, -3, -17, 5,
					-- layer=2 filter=79 channel=99
					0, 7, 6, -13, -5, -10, -16, -4, -1,
					-- layer=2 filter=79 channel=100
					2, 8, 6, 0, -12, 0, 5, -2, -2,
					-- layer=2 filter=79 channel=101
					-6, -14, 5, 4, -1, 2, -7, -5, 5,
					-- layer=2 filter=79 channel=102
					-4, 5, -2, 4, -2, 3, -7, -4, -12,
					-- layer=2 filter=79 channel=103
					0, -3, 2, 1, -7, -4, 5, -9, 0,
					-- layer=2 filter=79 channel=104
					-4, -2, 9, 1, 6, 6, 5, 3, 5,
					-- layer=2 filter=79 channel=105
					-12, 5, -1, 0, 7, -7, 3, -5, 6,
					-- layer=2 filter=79 channel=106
					-7, -3, 3, -6, -7, -14, 1, 2, -8,
					-- layer=2 filter=79 channel=107
					-9, -4, 6, -2, 0, 5, -5, 0, 10,
					-- layer=2 filter=79 channel=108
					-13, -2, -10, -10, -8, 1, 5, 4, -10,
					-- layer=2 filter=79 channel=109
					3, 6, -1, 7, -5, 0, -1, 8, 7,
					-- layer=2 filter=79 channel=110
					-7, -1, 4, 2, 1, -3, 1, 0, 5,
					-- layer=2 filter=79 channel=111
					8, 1, -7, -4, -2, 7, 0, 0, 5,
					-- layer=2 filter=79 channel=112
					2, -2, -7, -7, 2, 3, -10, 4, -1,
					-- layer=2 filter=79 channel=113
					1, -6, -3, -3, -3, -6, 6, -8, -2,
					-- layer=2 filter=79 channel=114
					-5, -4, 3, -2, 3, 6, 8, -8, 0,
					-- layer=2 filter=79 channel=115
					0, -8, 9, 4, -7, 7, -10, -2, 0,
					-- layer=2 filter=79 channel=116
					-11, 7, -11, -10, -7, 3, -6, -2, -12,
					-- layer=2 filter=79 channel=117
					-8, -7, 3, -1, -6, 1, -8, 5, 3,
					-- layer=2 filter=79 channel=118
					-9, 0, 0, 0, 0, -11, -6, -3, 2,
					-- layer=2 filter=79 channel=119
					2, -4, -6, -8, -9, 2, 0, 0, -13,
					-- layer=2 filter=79 channel=120
					-10, -4, 6, -1, -2, -4, 4, -8, 8,
					-- layer=2 filter=79 channel=121
					-10, 0, 6, -11, -9, 6, 1, -6, 0,
					-- layer=2 filter=79 channel=122
					-1, 0, 0, -3, 3, -11, -7, -6, 8,
					-- layer=2 filter=79 channel=123
					-6, -7, 7, -3, 0, -4, 2, -1, -10,
					-- layer=2 filter=79 channel=124
					-10, -8, 3, -7, 4, 2, -1, 3, -9,
					-- layer=2 filter=79 channel=125
					-5, 5, 1, -7, -6, 5, 7, -1, -5,
					-- layer=2 filter=79 channel=126
					-7, -9, -1, -1, 0, -11, 7, -2, -3,
					-- layer=2 filter=79 channel=127
					-2, -10, -12, 0, 8, -9, -11, 0, -1,
					-- layer=2 filter=80 channel=0
					-32, -25, 19, -29, -13, -56, 35, 23, -39,
					-- layer=2 filter=80 channel=1
					-31, -18, -18, -7, 20, 13, -55, -32, -19,
					-- layer=2 filter=80 channel=2
					-10, -3, 2, 6, -9, 8, -3, -2, -1,
					-- layer=2 filter=80 channel=3
					-53, -11, 4, -22, -38, 8, 26, 2, 13,
					-- layer=2 filter=80 channel=4
					-18, -75, 0, 53, -15, -32, 12, 8, 35,
					-- layer=2 filter=80 channel=5
					-5, -35, -12, 1, -10, -37, -4, -71, -80,
					-- layer=2 filter=80 channel=6
					-2, 3, -14, -28, 2, 23, -4, 50, 14,
					-- layer=2 filter=80 channel=7
					-11, -49, -47, -1, -1, -44, 14, -6, 43,
					-- layer=2 filter=80 channel=8
					-6, -10, -8, -10, 4, 2, 3, -6, -7,
					-- layer=2 filter=80 channel=9
					-19, 32, -29, -68, -3, -11, -33, -55, -35,
					-- layer=2 filter=80 channel=10
					-47, -13, -3, -34, -33, -23, 8, -44, -16,
					-- layer=2 filter=80 channel=11
					13, -21, -8, 7, -47, -11, -19, -20, -15,
					-- layer=2 filter=80 channel=12
					-15, -56, -45, -17, 53, 0, -38, -38, -28,
					-- layer=2 filter=80 channel=13
					-8, 6, 0, 6, -5, 4, 5, 3, 9,
					-- layer=2 filter=80 channel=14
					-22, -19, -62, -50, -6, -6, -53, -34, -18,
					-- layer=2 filter=80 channel=15
					5, 47, -29, 16, -24, 2, -54, -43, 25,
					-- layer=2 filter=80 channel=16
					-45, -54, -29, 8, -25, -61, -39, -46, 12,
					-- layer=2 filter=80 channel=17
					-7, -9, 1, 7, -9, -8, 0, 4, 0,
					-- layer=2 filter=80 channel=18
					-12, -34, -20, 21, 2, -31, -8, -38, 18,
					-- layer=2 filter=80 channel=19
					1, -15, -9, 36, 35, 11, -34, -9, 22,
					-- layer=2 filter=80 channel=20
					-7, 8, -7, 3, -9, -2, 4, 10, 0,
					-- layer=2 filter=80 channel=21
					-15, -11, 2, -19, -9, -6, 6, -10, 5,
					-- layer=2 filter=80 channel=22
					-5, -3, -8, -10, 10, 3, 10, -7, -2,
					-- layer=2 filter=80 channel=23
					-50, -28, -1, 0, -33, -16, -5, 10, 17,
					-- layer=2 filter=80 channel=24
					-80, -25, -15, -43, -29, -26, -28, 5, -44,
					-- layer=2 filter=80 channel=25
					-43, -57, -16, -16, -3, -27, -20, 5, -43,
					-- layer=2 filter=80 channel=26
					-6, 7, -7, -4, -9, -5, 0, -8, -7,
					-- layer=2 filter=80 channel=27
					18, 12, -4, -25, 6, -38, -68, -52, -45,
					-- layer=2 filter=80 channel=28
					-61, -89, 11, 19, -2, -44, 12, 9, 51,
					-- layer=2 filter=80 channel=29
					-1, 3, -9, -11, -8, 4, 4, -1, -2,
					-- layer=2 filter=80 channel=30
					11, -12, -1, 16, -62, 12, 19, -24, -22,
					-- layer=2 filter=80 channel=31
					43, 71, 70, 65, 22, 8, -4, 27, 17,
					-- layer=2 filter=80 channel=32
					2, 8, 0, 2, 5, 2, -5, -2, 7,
					-- layer=2 filter=80 channel=33
					-37, -34, -45, 16, -12, -48, -9, 28, -2,
					-- layer=2 filter=80 channel=34
					11, -40, -3, 11, -3, -20, 43, -59, 36,
					-- layer=2 filter=80 channel=35
					-3, -25, 6, 37, -34, -32, 26, 16, 39,
					-- layer=2 filter=80 channel=36
					-2, 9, -3, -1, 0, -5, 0, 0, 2,
					-- layer=2 filter=80 channel=37
					24, 3, -11, -26, -28, -18, -29, -67, -29,
					-- layer=2 filter=80 channel=38
					0, 16, -4, 6, -22, -13, 0, -30, -58,
					-- layer=2 filter=80 channel=39
					-85, -30, -65, -62, -96, 11, -14, -17, -17,
					-- layer=2 filter=80 channel=40
					31, -9, 16, 40, 21, -29, 45, -90, 8,
					-- layer=2 filter=80 channel=41
					-7, 2, 6, -4, 10, 10, -1, 3, 2,
					-- layer=2 filter=80 channel=42
					6, -99, -39, -68, -1, -24, -78, -41, -73,
					-- layer=2 filter=80 channel=43
					-39, 11, 22, -6, -63, -30, -22, -17, -17,
					-- layer=2 filter=80 channel=44
					2, 8, -2, 0, 6, 9, 0, 4, -5,
					-- layer=2 filter=80 channel=45
					0, 17, 4, 44, 1, -14, -14, 1, -2,
					-- layer=2 filter=80 channel=46
					25, -21, -34, 39, -53, -21, 29, -38, -36,
					-- layer=2 filter=80 channel=47
					-35, -49, 19, -5, -33, -34, -1, 8, 53,
					-- layer=2 filter=80 channel=48
					10, -9, 8, 4, 9, 8, 0, 5, -5,
					-- layer=2 filter=80 channel=49
					16, -26, -16, -25, 30, 6, -7, -39, -11,
					-- layer=2 filter=80 channel=50
					-7, -1, -1, -7, 22, 2, -5, 8, 11,
					-- layer=2 filter=80 channel=51
					3, 1, -2, 1, -40, -13, 8, -37, -29,
					-- layer=2 filter=80 channel=52
					56, 23, 11, 1, -56, -31, -35, -15, 11,
					-- layer=2 filter=80 channel=53
					-22, -22, -12, -81, 25, 18, -39, 7, -56,
					-- layer=2 filter=80 channel=54
					1, -49, -8, 17, -5, -29, 27, 7, 6,
					-- layer=2 filter=80 channel=55
					4, 0, 0, -2, -3, 0, 2, -15, 8,
					-- layer=2 filter=80 channel=56
					-9, -8, 8, -10, -21, -13, -20, -66, -21,
					-- layer=2 filter=80 channel=57
					-2, 2, -10, 2, 4, 1, -13, -5, 6,
					-- layer=2 filter=80 channel=58
					-50, -14, -39, -11, -10, -16, -23, -3, -54,
					-- layer=2 filter=80 channel=59
					-46, -4, -59, 24, -32, -8, -53, 42, -11,
					-- layer=2 filter=80 channel=60
					-2, -35, 9, 46, 42, -5, 21, 18, 4,
					-- layer=2 filter=80 channel=61
					-2, 3, -4, 40, 25, 9, 28, 44, 0,
					-- layer=2 filter=80 channel=62
					18, -9, -17, 7, -3, 27, -20, 3, 8,
					-- layer=2 filter=80 channel=63
					-46, -22, -16, -6, -8, 21, 36, 12, -33,
					-- layer=2 filter=80 channel=64
					-21, -37, -35, -33, -45, -10, -12, -42, -16,
					-- layer=2 filter=80 channel=65
					-18, -22, -7, 42, -18, 5, 21, 34, 17,
					-- layer=2 filter=80 channel=66
					28, 15, -14, -2, 24, 76, -37, -4, 8,
					-- layer=2 filter=80 channel=67
					-4, -42, -8, -17, -76, 0, 18, 16, -28,
					-- layer=2 filter=80 channel=68
					6, 9, -4, -1, -2, 2, -1, -7, 0,
					-- layer=2 filter=80 channel=69
					-50, -42, -105, -55, -49, -16, -73, -49, -19,
					-- layer=2 filter=80 channel=70
					-14, -19, 27, 14, -6, -46, 26, 4, 15,
					-- layer=2 filter=80 channel=71
					16, 5, -23, 9, 17, 2, -103, -46, -35,
					-- layer=2 filter=80 channel=72
					-51, -84, -53, 4, 9, -74, -14, 1, 8,
					-- layer=2 filter=80 channel=73
					64, 47, 57, 16, 40, 18, -12, 8, -4,
					-- layer=2 filter=80 channel=74
					-27, -35, -17, 20, -80, -56, 19, -2, -60,
					-- layer=2 filter=80 channel=75
					-37, -51, -30, -29, -3, 60, -21, -50, 22,
					-- layer=2 filter=80 channel=76
					45, 27, 32, 35, -5, 60, -29, 47, 49,
					-- layer=2 filter=80 channel=77
					-10, -3, -8, -10, 1, -8, -8, -5, 8,
					-- layer=2 filter=80 channel=78
					25, -47, -2, 0, -34, -8, -48, -40, 23,
					-- layer=2 filter=80 channel=79
					-2, -10, -8, 8, 5, 2, 7, -9, 0,
					-- layer=2 filter=80 channel=80
					-41, -10, -9, -13, -45, 5, -2, -53, -8,
					-- layer=2 filter=80 channel=81
					4, 4, 8, -6, -1, 0, 10, -11, -11,
					-- layer=2 filter=80 channel=82
					0, 1, -5, 0, 1, -6, -7, 0, 3,
					-- layer=2 filter=80 channel=83
					-30, -7, -7, 15, 30, -8, 16, -11, 15,
					-- layer=2 filter=80 channel=84
					2, 3, 5, 5, -2, -8, -9, -2, -6,
					-- layer=2 filter=80 channel=85
					11, -8, 16, -6, 13, 0, 0, 1, 14,
					-- layer=2 filter=80 channel=86
					-16, -2, 0, -9, -4, -8, 5, -11, 8,
					-- layer=2 filter=80 channel=87
					16, 4, 12, 59, -40, 8, -1, 37, 43,
					-- layer=2 filter=80 channel=88
					-40, -9, -71, 25, -19, 23, 28, 9, -20,
					-- layer=2 filter=80 channel=89
					-56, -51, -37, 18, 4, -7, -106, -34, -19,
					-- layer=2 filter=80 channel=90
					-2, 8, -6, 7, 6, 1, -8, -8, -8,
					-- layer=2 filter=80 channel=91
					-46, -78, -6, 22, 28, -12, -40, -54, -21,
					-- layer=2 filter=80 channel=92
					-2, -35, -11, -5, 46, -22, -69, -41, -26,
					-- layer=2 filter=80 channel=93
					44, -5, 61, 42, 32, 53, 26, 16, 54,
					-- layer=2 filter=80 channel=94
					12, -19, 5, -8, 31, 14, 21, 65, -1,
					-- layer=2 filter=80 channel=95
					-6, 1, -1, -14, 14, -12, 7, -1, -5,
					-- layer=2 filter=80 channel=96
					-21, 2, 2, -7, 52, 39, -21, 28, -17,
					-- layer=2 filter=80 channel=97
					-47, -25, -50, 10, -39, -31, 0, -43, 0,
					-- layer=2 filter=80 channel=98
					-2, -47, -16, -5, -28, -46, 14, 1, 39,
					-- layer=2 filter=80 channel=99
					33, 19, 0, 30, -3, 11, -51, -3, 25,
					-- layer=2 filter=80 channel=100
					-9, -34, -25, 32, -7, -40, -21, -43, 10,
					-- layer=2 filter=80 channel=101
					30, -25, -6, 6, 12, -37, -27, 14, -33,
					-- layer=2 filter=80 channel=102
					28, -24, -1, 21, 10, 12, -29, -11, -6,
					-- layer=2 filter=80 channel=103
					8, -22, 31, 20, 116, 33, 51, 3, 20,
					-- layer=2 filter=80 channel=104
					-19, -28, -4, -49, 4, 1, -22, -28, -12,
					-- layer=2 filter=80 channel=105
					55, 29, -13, 109, -76, -7, -23, 35, 111,
					-- layer=2 filter=80 channel=106
					-77, -61, -32, -35, -4, 12, -19, 40, -12,
					-- layer=2 filter=80 channel=107
					-20, -50, 23, -58, 43, -27, 14, -7, -9,
					-- layer=2 filter=80 channel=108
					-10, 2, -17, -52, -8, -20, -100, -35, -2,
					-- layer=2 filter=80 channel=109
					17, -11, -4, 1, -12, -11, -5, -3, -12,
					-- layer=2 filter=80 channel=110
					-47, -38, -40, -18, 9, -17, -74, -15, -2,
					-- layer=2 filter=80 channel=111
					9, 7, 7, -1, -4, -10, 7, -7, 8,
					-- layer=2 filter=80 channel=112
					2, 7, 10, 22, 13, 28, 32, -5, -9,
					-- layer=2 filter=80 channel=113
					-21, -31, -13, 26, -12, 36, 29, -22, 13,
					-- layer=2 filter=80 channel=114
					-6, 17, 11, 1, -14, 5, -6, -2, 4,
					-- layer=2 filter=80 channel=115
					-4, 0, 7, -2, 3, 1, -7, 0, 0,
					-- layer=2 filter=80 channel=116
					-17, 2, -11, 16, -20, -7, 12, 1, 32,
					-- layer=2 filter=80 channel=117
					22, -12, 12, 43, 54, -15, -7, -14, 0,
					-- layer=2 filter=80 channel=118
					-25, 0, -29, -53, -73, -32, -21, -34, -25,
					-- layer=2 filter=80 channel=119
					-9, -13, 5, 31, 17, -17, 29, 19, 37,
					-- layer=2 filter=80 channel=120
					-6, 5, 7, 5, -9, 8, 5, -4, 4,
					-- layer=2 filter=80 channel=121
					-6, -3, -10, -4, -8, 2, 0, 5, 3,
					-- layer=2 filter=80 channel=122
					-10, -6, -12, -14, 7, -3, -2, -2, 6,
					-- layer=2 filter=80 channel=123
					-7, -37, -51, 16, -33, -34, -3, 29, 55,
					-- layer=2 filter=80 channel=124
					-3, 16, -27, 26, -14, -7, -34, 13, 61,
					-- layer=2 filter=80 channel=125
					8, 8, -5, 3, -4, 9, 3, 7, 8,
					-- layer=2 filter=80 channel=126
					-6, 23, -25, -4, 48, -16, -3, 12, -11,
					-- layer=2 filter=80 channel=127
					-67, -12, -26, 17, -36, 5, 33, -24, 32,
					-- layer=2 filter=81 channel=0
					0, -8, -5, -2, -2, 0, -9, 2, 0,
					-- layer=2 filter=81 channel=1
					-20, -19, -7, 7, -25, -24, 13, -7, 35,
					-- layer=2 filter=81 channel=2
					2, 7, -9, -2, 3, 11, 0, 1, 4,
					-- layer=2 filter=81 channel=3
					7, -4, 10, 11, -14, -22, 31, 8, 7,
					-- layer=2 filter=81 channel=4
					5, -31, -25, 23, -21, -39, 26, 26, -6,
					-- layer=2 filter=81 channel=5
					-1, -24, 2, -17, 8, 21, 2, 8, 2,
					-- layer=2 filter=81 channel=6
					-7, 5, 11, 30, 19, 15, 32, 52, 43,
					-- layer=2 filter=81 channel=7
					2, -14, -14, -53, -39, -32, 2, 19, -13,
					-- layer=2 filter=81 channel=8
					-5, 8, 7, 6, -7, 0, 8, -3, -3,
					-- layer=2 filter=81 channel=9
					24, -4, -24, 48, -4, -23, 7, -14, 7,
					-- layer=2 filter=81 channel=10
					25, 0, 0, 36, 4, 2, 3, 7, -32,
					-- layer=2 filter=81 channel=11
					-12, 0, 13, 6, 1, 0, 17, 10, 0,
					-- layer=2 filter=81 channel=12
					-40, -33, -11, -25, -28, -18, -7, -4, 4,
					-- layer=2 filter=81 channel=13
					-7, -1, 7, -8, -4, 2, 7, -8, -10,
					-- layer=2 filter=81 channel=14
					-40, -30, 5, -18, -17, -13, -10, -10, 47,
					-- layer=2 filter=81 channel=15
					-21, 32, 12, 37, -18, 7, -40, -22, -6,
					-- layer=2 filter=81 channel=16
					29, -10, -14, 20, -36, -76, 19, -19, -53,
					-- layer=2 filter=81 channel=17
					-1, -2, -8, 2, -7, 7, 1, 0, 4,
					-- layer=2 filter=81 channel=18
					-35, -34, 8, -10, 10, 25, 0, 9, -4,
					-- layer=2 filter=81 channel=19
					9, 0, 26, 10, 3, -27, 20, 16, 27,
					-- layer=2 filter=81 channel=20
					-7, 11, 7, 7, 5, 0, 5, 3, 3,
					-- layer=2 filter=81 channel=21
					10, -14, -1, 8, -10, 3, 7, -10, 4,
					-- layer=2 filter=81 channel=22
					-3, 1, 8, 5, -1, 1, -3, -6, -1,
					-- layer=2 filter=81 channel=23
					6, 1, -29, 28, 16, -43, 6, 12, -35,
					-- layer=2 filter=81 channel=24
					26, -3, 2, 33, -26, -31, 27, 13, 3,
					-- layer=2 filter=81 channel=25
					4, -14, 3, 31, 0, -9, 16, 9, 0,
					-- layer=2 filter=81 channel=26
					5, -9, -3, 10, 5, -4, 3, 3, 6,
					-- layer=2 filter=81 channel=27
					16, -7, 10, 13, -18, -8, 18, 11, 0,
					-- layer=2 filter=81 channel=28
					3, 9, -5, 2, -26, 12, -41, -34, -45,
					-- layer=2 filter=81 channel=29
					5, -8, 6, -5, -6, 10, -7, -9, -9,
					-- layer=2 filter=81 channel=30
					3, -22, -44, 3, -1, -8, 10, 1, -1,
					-- layer=2 filter=81 channel=31
					-10, 28, 16, 33, -17, -39, -47, -1, -17,
					-- layer=2 filter=81 channel=32
					3, 3, -7, 0, 1, 2, -1, -3, 5,
					-- layer=2 filter=81 channel=33
					-2, -48, 14, -11, -17, -37, 31, 19, 18,
					-- layer=2 filter=81 channel=34
					23, 0, 3, 14, 37, 35, 3, 41, 6,
					-- layer=2 filter=81 channel=35
					11, -33, -15, -12, -7, 23, -33, -17, -65,
					-- layer=2 filter=81 channel=36
					-1, -5, -13, -11, 5, -4, -10, 0, -2,
					-- layer=2 filter=81 channel=37
					-18, -5, 20, -24, -7, 8, 10, -5, -3,
					-- layer=2 filter=81 channel=38
					-7, -20, 6, -2, -8, -3, 3, 1, 15,
					-- layer=2 filter=81 channel=39
					11, -2, -18, 13, 22, -63, 15, -40, -65,
					-- layer=2 filter=81 channel=40
					-11, 9, 38, 27, 27, 79, -9, -2, -37,
					-- layer=2 filter=81 channel=41
					5, -6, 2, 5, -9, 11, 7, -8, 0,
					-- layer=2 filter=81 channel=42
					32, 6, -30, 7, -3, -48, -2, -31, -27,
					-- layer=2 filter=81 channel=43
					2, -43, 7, 26, 18, 13, 7, -29, -56,
					-- layer=2 filter=81 channel=44
					-4, -1, 0, -2, 9, 0, 1, -4, 2,
					-- layer=2 filter=81 channel=45
					-40, 11, -12, -6, -39, -61, 10, -3, -35,
					-- layer=2 filter=81 channel=46
					17, 0, -17, 11, 8, -21, 10, -5, -39,
					-- layer=2 filter=81 channel=47
					24, 11, 25, -17, -18, -40, 10, 5, -59,
					-- layer=2 filter=81 channel=48
					-1, 8, -5, 7, 9, -9, 5, 4, 2,
					-- layer=2 filter=81 channel=49
					-31, -1, -16, -9, 13, -20, -11, -14, 13,
					-- layer=2 filter=81 channel=50
					-12, 9, -10, -1, -3, 15, 2, -4, 1,
					-- layer=2 filter=81 channel=51
					0, -8, -3, -1, 7, 18, -4, 4, 3,
					-- layer=2 filter=81 channel=52
					-20, -24, 0, -6, -28, 13, 23, -13, -9,
					-- layer=2 filter=81 channel=53
					-7, -16, -16, 8, -43, -71, -15, 3, -3,
					-- layer=2 filter=81 channel=54
					-7, -14, 6, 8, 24, 8, 22, 48, 2,
					-- layer=2 filter=81 channel=55
					6, -10, 6, 11, -9, 0, 0, 1, -4,
					-- layer=2 filter=81 channel=56
					-2, -7, 16, 1, -9, 10, 5, 5, 11,
					-- layer=2 filter=81 channel=57
					-14, -4, 11, -17, -8, -4, -20, 0, -4,
					-- layer=2 filter=81 channel=58
					-35, -8, -18, -26, -41, -33, -18, -21, -6,
					-- layer=2 filter=81 channel=59
					-16, -37, -24, -8, -31, -44, 3, 8, 26,
					-- layer=2 filter=81 channel=60
					-34, -27, 0, 1, -26, -21, 2, 11, 29,
					-- layer=2 filter=81 channel=61
					-6, 17, 31, 16, 3, 34, -27, 5, 40,
					-- layer=2 filter=81 channel=62
					13, -17, 1, 9, -13, 0, 29, 29, 23,
					-- layer=2 filter=81 channel=63
					3, 8, -18, 7, 9, -47, 15, 10, 4,
					-- layer=2 filter=81 channel=64
					22, 6, -28, 55, 3, -47, 43, -4, -37,
					-- layer=2 filter=81 channel=65
					-7, 19, 21, 8, 13, 45, 2, 40, 30,
					-- layer=2 filter=81 channel=66
					4, 12, -9, -21, 3, 32, 37, 0, 42,
					-- layer=2 filter=81 channel=67
					30, -1, -25, 17, 6, -36, -2, -17, -22,
					-- layer=2 filter=81 channel=68
					-4, -9, 3, -3, -8, 4, -5, 5, 9,
					-- layer=2 filter=81 channel=69
					17, -15, -28, 13, 4, -36, 31, -19, -10,
					-- layer=2 filter=81 channel=70
					-1, -19, 9, -18, 2, 25, -17, 7, -4,
					-- layer=2 filter=81 channel=71
					9, 15, 48, -2, -31, 3, 9, -21, 0,
					-- layer=2 filter=81 channel=72
					2, -7, 28, -25, 11, 1, -45, -13, 33,
					-- layer=2 filter=81 channel=73
					45, 60, 19, -30, 14, -26, -96, 2, 3,
					-- layer=2 filter=81 channel=74
					0, -1, -22, 12, 18, -37, -11, -2, -22,
					-- layer=2 filter=81 channel=75
					18, 30, -34, -47, -38, -6, -21, 8, 23,
					-- layer=2 filter=81 channel=76
					26, 46, 27, 28, -12, 12, 16, -42, -30,
					-- layer=2 filter=81 channel=77
					10, -5, -8, 8, 6, -3, -7, -1, 3,
					-- layer=2 filter=81 channel=78
					-16, -18, 2, 7, 16, -7, 11, 8, -6,
					-- layer=2 filter=81 channel=79
					10, 5, 2, 4, -2, -8, 10, -4, 7,
					-- layer=2 filter=81 channel=80
					35, 15, 1, 32, 9, -30, 19, -23, -46,
					-- layer=2 filter=81 channel=81
					12, 7, -3, -3, 0, 7, 8, 0, 14,
					-- layer=2 filter=81 channel=82
					0, -5, -5, 7, -3, 2, 1, 4, 8,
					-- layer=2 filter=81 channel=83
					25, -6, -40, 8, 4, -25, 28, 0, -3,
					-- layer=2 filter=81 channel=84
					4, 0, 5, 8, 9, -3, -4, -2, 11,
					-- layer=2 filter=81 channel=85
					-2, 1, -17, -14, 3, -6, -12, 1, 7,
					-- layer=2 filter=81 channel=86
					-2, 9, -2, 4, 19, -10, 17, 3, 3,
					-- layer=2 filter=81 channel=87
					-2, -26, 17, -32, 21, -1, 7, -18, -26,
					-- layer=2 filter=81 channel=88
					-22, -25, -28, -4, 21, -16, 12, 5, 3,
					-- layer=2 filter=81 channel=89
					-6, -13, 2, -32, 0, -13, -32, -18, 3,
					-- layer=2 filter=81 channel=90
					-5, 10, 2, -1, -4, -2, 9, 5, -7,
					-- layer=2 filter=81 channel=91
					6, -30, -10, -13, -80, -13, -48, -50, -28,
					-- layer=2 filter=81 channel=92
					-18, -26, -32, -33, -41, -36, -9, -22, 3,
					-- layer=2 filter=81 channel=93
					-34, -31, -3, 30, -22, -29, 17, 28, -42,
					-- layer=2 filter=81 channel=94
					54, -4, 21, 11, 10, 6, -13, 43, -2,
					-- layer=2 filter=81 channel=95
					2, 0, -22, 1, -15, -21, -10, 3, 3,
					-- layer=2 filter=81 channel=96
					-55, 31, -22, -80, 31, 16, -26, 33, 9,
					-- layer=2 filter=81 channel=97
					-4, -5, -14, 24, -26, -57, 40, 11, 8,
					-- layer=2 filter=81 channel=98
					15, 30, 39, 12, 10, 28, -10, 2, -41,
					-- layer=2 filter=81 channel=99
					-6, -7, 10, 21, -26, -6, 27, 0, -64,
					-- layer=2 filter=81 channel=100
					2, 9, -22, 67, -17, 0, 0, -4, -23,
					-- layer=2 filter=81 channel=101
					3, -19, 26, -8, -39, -32, -10, -36, -16,
					-- layer=2 filter=81 channel=102
					-18, 4, 7, -51, -26, 25, 8, 1, 14,
					-- layer=2 filter=81 channel=103
					-16, -55, -74, 6, 21, -7, -28, -8, 21,
					-- layer=2 filter=81 channel=104
					-26, 3, -6, -25, 20, -11, -17, 12, 7,
					-- layer=2 filter=81 channel=105
					-25, 28, -21, 26, 2, -7, -31, -41, -9,
					-- layer=2 filter=81 channel=106
					14, -11, -4, 16, -41, -30, 0, -13, -11,
					-- layer=2 filter=81 channel=107
					10, -8, -52, -16, 44, -41, -33, 20, 1,
					-- layer=2 filter=81 channel=108
					-21, -21, 16, -19, -50, 4, 1, -13, 34,
					-- layer=2 filter=81 channel=109
					-6, -4, -4, 4, 15, 3, 5, 14, 12,
					-- layer=2 filter=81 channel=110
					23, 23, -16, 51, 33, -29, 23, -7, -19,
					-- layer=2 filter=81 channel=111
					4, -3, 1, 4, 2, -7, -3, -7, -7,
					-- layer=2 filter=81 channel=112
					6, -10, -5, -4, -10, 4, -38, 8, 9,
					-- layer=2 filter=81 channel=113
					17, -1, -31, 10, -6, -8, 0, -11, 11,
					-- layer=2 filter=81 channel=114
					-7, 5, -7, -13, -5, -16, 3, -12, -8,
					-- layer=2 filter=81 channel=115
					-2, 2, 8, 7, 4, -4, 2, 1, -4,
					-- layer=2 filter=81 channel=116
					-14, 0, 23, -34, -4, 35, -4, -4, -11,
					-- layer=2 filter=81 channel=117
					25, -5, 0, -10, -10, -64, -22, 52, 1,
					-- layer=2 filter=81 channel=118
					25, 3, 4, 10, 16, 0, 16, 4, -16,
					-- layer=2 filter=81 channel=119
					4, -73, -56, 26, -5, -14, 26, -2, -11,
					-- layer=2 filter=81 channel=120
					-1, -4, -7, 1, 7, 2, -9, -10, 7,
					-- layer=2 filter=81 channel=121
					-4, -5, -1, 1, -6, -8, -9, 0, 4,
					-- layer=2 filter=81 channel=122
					-5, 5, 0, -1, 9, 4, 0, 16, 0,
					-- layer=2 filter=81 channel=123
					22, 15, 30, -4, -15, -26, 12, 0, -6,
					-- layer=2 filter=81 channel=124
					27, 0, -1, 77, 14, -22, 20, -2, 17,
					-- layer=2 filter=81 channel=125
					-3, 4, -4, 6, 0, 2, -5, -3, 7,
					-- layer=2 filter=81 channel=126
					-24, -34, -84, -5, 12, -39, -41, 8, -28,
					-- layer=2 filter=81 channel=127
					-20, -44, -4, 0, 17, -36, -6, -8, 24,
					-- layer=2 filter=82 channel=0
					-2, -1, 4, 0, 6, 2, -12, -2, -13,
					-- layer=2 filter=82 channel=1
					-2, -10, -7, 6, -9, -3, -9, -5, -5,
					-- layer=2 filter=82 channel=2
					-3, 6, -5, 0, -2, 6, 0, -2, -2,
					-- layer=2 filter=82 channel=3
					-1, -6, 11, 7, -3, 2, 10, 4, 0,
					-- layer=2 filter=82 channel=4
					6, -4, -7, -7, -3, -1, 0, -9, -3,
					-- layer=2 filter=82 channel=5
					3, -7, -11, -3, -6, 5, -6, -1, -5,
					-- layer=2 filter=82 channel=6
					-9, 8, -10, -12, 4, -4, -2, -11, 6,
					-- layer=2 filter=82 channel=7
					-5, -6, -1, -2, 2, -13, 4, 3, -1,
					-- layer=2 filter=82 channel=8
					8, 2, 0, -3, -3, 5, -7, 4, 7,
					-- layer=2 filter=82 channel=9
					5, 5, -10, -12, -12, -10, -1, 1, 6,
					-- layer=2 filter=82 channel=10
					-9, -7, -1, 5, -8, 1, -1, 6, 7,
					-- layer=2 filter=82 channel=11
					0, -7, -2, 2, 3, -1, 0, -8, 4,
					-- layer=2 filter=82 channel=12
					0, 0, 0, -9, -5, -13, 5, 0, -3,
					-- layer=2 filter=82 channel=13
					-6, 0, 0, -10, -7, 5, 1, -7, -1,
					-- layer=2 filter=82 channel=14
					-11, 2, -5, 0, -4, -2, 7, -8, -1,
					-- layer=2 filter=82 channel=15
					4, -2, 0, -3, 4, -5, -5, -11, -12,
					-- layer=2 filter=82 channel=16
					3, 0, 2, 3, 8, -2, 2, -9, 0,
					-- layer=2 filter=82 channel=17
					2, 10, 3, 8, 1, -5, 5, 9, -8,
					-- layer=2 filter=82 channel=18
					4, 0, 2, 3, 1, 0, 0, 6, -1,
					-- layer=2 filter=82 channel=19
					-5, -3, 0, -8, 0, -11, -6, -14, 4,
					-- layer=2 filter=82 channel=20
					-3, 8, -2, 0, 2, -4, 2, -3, -6,
					-- layer=2 filter=82 channel=21
					-9, -11, 8, -8, 0, -6, 8, 2, -10,
					-- layer=2 filter=82 channel=22
					0, 2, 0, 2, 6, -1, -9, -5, 6,
					-- layer=2 filter=82 channel=23
					-8, 7, 8, 7, 0, -5, 0, -2, 6,
					-- layer=2 filter=82 channel=24
					-9, -9, 0, 3, -6, -1, -8, 0, -8,
					-- layer=2 filter=82 channel=25
					8, -5, -6, -7, -11, -7, 3, -6, -3,
					-- layer=2 filter=82 channel=26
					2, 9, 0, -8, -8, 3, -7, 0, 8,
					-- layer=2 filter=82 channel=27
					-6, 4, -8, 0, -3, -1, 4, 3, 1,
					-- layer=2 filter=82 channel=28
					8, 3, 3, -7, 10, -10, -10, -10, -8,
					-- layer=2 filter=82 channel=29
					8, -5, 4, -1, -12, -3, -7, 7, -10,
					-- layer=2 filter=82 channel=30
					-2, -12, 5, 3, -11, -6, -4, -1, 4,
					-- layer=2 filter=82 channel=31
					3, -9, 2, -3, -8, -9, 2, 3, -2,
					-- layer=2 filter=82 channel=32
					-4, 6, 8, -9, 5, 3, -11, -9, -6,
					-- layer=2 filter=82 channel=33
					-3, -11, -9, -4, -3, -9, 0, 8, -3,
					-- layer=2 filter=82 channel=34
					-13, -10, -6, -10, 2, 0, 0, 7, -6,
					-- layer=2 filter=82 channel=35
					-6, 6, -11, 9, 2, -9, -6, 0, -12,
					-- layer=2 filter=82 channel=36
					5, 0, -11, -5, 6, 1, 3, 0, -4,
					-- layer=2 filter=82 channel=37
					-1, -9, -9, 7, -1, -8, -10, -11, -2,
					-- layer=2 filter=82 channel=38
					-2, 4, -11, 3, 2, -12, 8, -5, -1,
					-- layer=2 filter=82 channel=39
					6, -5, -4, 0, 0, -8, 0, 8, -12,
					-- layer=2 filter=82 channel=40
					-10, -13, 7, 5, -10, -10, 2, 4, -10,
					-- layer=2 filter=82 channel=41
					0, -7, 6, -6, -2, 6, -7, -2, -1,
					-- layer=2 filter=82 channel=42
					-3, -5, 10, 4, -4, -14, -7, 0, -10,
					-- layer=2 filter=82 channel=43
					-9, -10, -1, -6, 6, -7, -4, -8, 1,
					-- layer=2 filter=82 channel=44
					9, 0, 1, 5, 1, -9, 0, -7, -4,
					-- layer=2 filter=82 channel=45
					-9, -7, 4, 6, -9, -5, 7, -9, 1,
					-- layer=2 filter=82 channel=46
					-4, 3, -8, -4, -7, -2, -2, 5, -10,
					-- layer=2 filter=82 channel=47
					3, 0, 0, -9, -1, -10, -7, 0, -2,
					-- layer=2 filter=82 channel=48
					-5, 2, -2, -8, 8, -6, 2, 1, -6,
					-- layer=2 filter=82 channel=49
					-2, -2, -2, 0, 0, -6, -12, 1, 0,
					-- layer=2 filter=82 channel=50
					-4, -1, -1, -8, 4, -8, -4, -3, 6,
					-- layer=2 filter=82 channel=51
					-10, -7, -13, -1, -2, -2, 6, 2, -5,
					-- layer=2 filter=82 channel=52
					0, 4, 4, 2, -12, -13, -3, -4, -6,
					-- layer=2 filter=82 channel=53
					-1, 6, 2, 0, 3, -7, -2, -8, 3,
					-- layer=2 filter=82 channel=54
					3, -1, 10, 2, 6, -5, 6, -4, 7,
					-- layer=2 filter=82 channel=55
					4, -8, 3, -10, 1, -2, 6, 0, -5,
					-- layer=2 filter=82 channel=56
					2, -1, 4, -3, 2, -9, -8, -1, -1,
					-- layer=2 filter=82 channel=57
					1, -2, -2, 7, -8, 8, -3, 1, 0,
					-- layer=2 filter=82 channel=58
					2, 4, -11, 3, -1, -2, 4, 5, -9,
					-- layer=2 filter=82 channel=59
					7, -6, 1, 2, -8, -4, 1, 3, -8,
					-- layer=2 filter=82 channel=60
					5, -3, -9, 3, -11, -1, -1, -13, -3,
					-- layer=2 filter=82 channel=61
					-2, -15, 3, -2, -9, -9, 3, 4, 0,
					-- layer=2 filter=82 channel=62
					2, -10, -4, -11, 6, -4, -12, 7, -14,
					-- layer=2 filter=82 channel=63
					-8, -6, -7, -6, -8, -10, -9, -11, -11,
					-- layer=2 filter=82 channel=64
					0, 0, -7, 0, -9, -11, 0, 0, 5,
					-- layer=2 filter=82 channel=65
					-3, -2, 1, -7, -5, -4, -5, -9, 0,
					-- layer=2 filter=82 channel=66
					0, -6, -8, -6, -1, 8, -3, 9, -8,
					-- layer=2 filter=82 channel=67
					5, -2, 1, -10, -5, 8, 8, -11, -4,
					-- layer=2 filter=82 channel=68
					-6, -12, 7, 8, 2, -8, 2, -12, -5,
					-- layer=2 filter=82 channel=69
					9, 11, -1, 9, -9, -9, -7, -8, -7,
					-- layer=2 filter=82 channel=70
					-11, 9, 2, -7, 9, -7, 5, -4, -6,
					-- layer=2 filter=82 channel=71
					-2, 1, -2, -1, -2, 2, 5, 0, 0,
					-- layer=2 filter=82 channel=72
					-4, -10, 7, -9, 0, -3, -6, -13, -7,
					-- layer=2 filter=82 channel=73
					2, 6, 5, 4, 0, 1, -6, 6, -5,
					-- layer=2 filter=82 channel=74
					10, -9, 5, 3, -3, -4, -11, 8, -10,
					-- layer=2 filter=82 channel=75
					-8, 3, 2, 5, -3, -3, -1, -9, 3,
					-- layer=2 filter=82 channel=76
					1, -2, -4, 8, 5, -2, -7, 6, 4,
					-- layer=2 filter=82 channel=77
					-10, 4, 7, -10, 7, 10, 7, 5, -5,
					-- layer=2 filter=82 channel=78
					0, -11, -4, 5, 1, -5, 2, -2, -6,
					-- layer=2 filter=82 channel=79
					0, -1, -6, -1, -7, -8, 0, 2, 1,
					-- layer=2 filter=82 channel=80
					2, 4, 9, -7, 1, 4, 4, -11, 5,
					-- layer=2 filter=82 channel=81
					-6, -8, -9, -11, -5, -1, -6, 4, 8,
					-- layer=2 filter=82 channel=82
					10, 10, -1, 4, 3, 7, 6, 3, 11,
					-- layer=2 filter=82 channel=83
					-11, 2, -2, -8, -1, -8, -9, 0, -2,
					-- layer=2 filter=82 channel=84
					-5, -7, -5, -9, -1, 1, 4, 0, 9,
					-- layer=2 filter=82 channel=85
					-4, 8, 1, -4, -1, 0, -9, -4, -7,
					-- layer=2 filter=82 channel=86
					-4, 0, -4, 3, -11, 1, 6, -5, -6,
					-- layer=2 filter=82 channel=87
					-8, 2, -4, -2, -1, -8, -6, 2, -8,
					-- layer=2 filter=82 channel=88
					-9, 0, -1, 1, -2, -3, -3, 0, -10,
					-- layer=2 filter=82 channel=89
					-8, 5, 4, -5, -1, 1, -7, -4, 0,
					-- layer=2 filter=82 channel=90
					-9, -3, 0, -1, 5, -2, 2, 7, 0,
					-- layer=2 filter=82 channel=91
					-9, 0, -12, -7, 1, 5, -11, -6, -7,
					-- layer=2 filter=82 channel=92
					-7, -6, 6, -12, -8, -4, -2, -4, -9,
					-- layer=2 filter=82 channel=93
					-1, -4, -6, -4, 0, -1, -6, -11, 3,
					-- layer=2 filter=82 channel=94
					-5, -3, 1, 8, 6, -7, -11, -9, -11,
					-- layer=2 filter=82 channel=95
					9, -9, -6, -3, -7, -9, 5, -10, 7,
					-- layer=2 filter=82 channel=96
					-12, 10, -4, -5, -8, 0, 2, 3, -14,
					-- layer=2 filter=82 channel=97
					-4, 5, -9, -4, -11, -4, 1, -6, 6,
					-- layer=2 filter=82 channel=98
					-1, -8, 3, -11, 7, 4, -5, -8, 6,
					-- layer=2 filter=82 channel=99
					3, -8, -4, 6, 3, -11, -9, -7, 0,
					-- layer=2 filter=82 channel=100
					8, 0, -6, 7, 8, -10, -2, 5, 1,
					-- layer=2 filter=82 channel=101
					2, -11, 0, -13, 2, -6, 0, -12, -13,
					-- layer=2 filter=82 channel=102
					5, -4, 4, -3, -3, 2, 0, -5, -7,
					-- layer=2 filter=82 channel=103
					-5, -7, -4, -7, -2, 0, 4, -3, 0,
					-- layer=2 filter=82 channel=104
					-6, -2, -8, -5, -10, 0, -8, 5, 6,
					-- layer=2 filter=82 channel=105
					-7, 3, 0, 9, -1, 7, 5, 0, -8,
					-- layer=2 filter=82 channel=106
					-8, -8, -14, 0, -1, 0, -9, -1, -14,
					-- layer=2 filter=82 channel=107
					2, 5, 9, -7, -1, 2, 8, -5, -6,
					-- layer=2 filter=82 channel=108
					-7, -6, -8, -9, 5, 3, -12, -8, -2,
					-- layer=2 filter=82 channel=109
					7, 1, 3, -2, 0, -8, 7, -5, -4,
					-- layer=2 filter=82 channel=110
					-4, 8, 6, 4, -8, -2, 0, -2, -3,
					-- layer=2 filter=82 channel=111
					-5, 4, -8, 10, 4, 3, -8, -9, -7,
					-- layer=2 filter=82 channel=112
					-4, -2, -3, 7, -5, -4, 2, -13, -8,
					-- layer=2 filter=82 channel=113
					-2, 3, -2, 0, -11, 2, 2, 8, 0,
					-- layer=2 filter=82 channel=114
					-5, 6, -8, 5, 4, 5, 4, 0, -6,
					-- layer=2 filter=82 channel=115
					9, -2, 2, 3, -7, 0, 0, -7, -3,
					-- layer=2 filter=82 channel=116
					-2, -2, 7, -1, -5, -3, -9, -4, -13,
					-- layer=2 filter=82 channel=117
					3, 7, -10, -6, -3, -13, -2, 6, 6,
					-- layer=2 filter=82 channel=118
					5, 0, -1, 4, 8, -10, -9, 2, -6,
					-- layer=2 filter=82 channel=119
					-15, -8, -7, -10, -5, 8, 4, 7, 4,
					-- layer=2 filter=82 channel=120
					9, 10, -5, -6, -3, -8, -9, -7, 3,
					-- layer=2 filter=82 channel=121
					-9, 2, 1, -9, -10, -6, 0, -6, 0,
					-- layer=2 filter=82 channel=122
					0, 4, 0, -8, 5, -7, -5, 2, -8,
					-- layer=2 filter=82 channel=123
					2, -13, -10, -3, -10, -6, 2, 1, -11,
					-- layer=2 filter=82 channel=124
					0, 4, 2, -10, 6, -5, 5, -1, 8,
					-- layer=2 filter=82 channel=125
					0, 10, 4, -10, 0, 2, -7, -3, -4,
					-- layer=2 filter=82 channel=126
					-2, 2, 2, 5, 6, -6, 0, 1, -8,
					-- layer=2 filter=82 channel=127
					3, -4, -10, 3, 1, -8, -8, 6, 9,
					-- layer=2 filter=83 channel=0
					23, -7, -3, -19, -6, -8, 6, -11, -1,
					-- layer=2 filter=83 channel=1
					-12, -21, -11, -7, -11, 14, -11, -8, 11,
					-- layer=2 filter=83 channel=2
					-2, 3, -2, 9, 6, 3, -2, -7, 8,
					-- layer=2 filter=83 channel=3
					-12, -9, -18, -39, -36, -38, 0, 22, 26,
					-- layer=2 filter=83 channel=4
					39, 32, 11, -39, -14, -15, -16, -28, 5,
					-- layer=2 filter=83 channel=5
					12, -9, 1, 5, 0, 0, -3, -7, -23,
					-- layer=2 filter=83 channel=6
					16, 6, 7, 32, 58, 17, -13, 54, 36,
					-- layer=2 filter=83 channel=7
					35, 12, 39, -25, 44, 45, -14, 3, 11,
					-- layer=2 filter=83 channel=8
					-4, 0, -11, 5, 6, -5, 0, 2, 0,
					-- layer=2 filter=83 channel=9
					25, 9, -47, 37, -8, -23, 4, 12, -35,
					-- layer=2 filter=83 channel=10
					0, 5, -16, -1, -35, -33, -2, -13, -24,
					-- layer=2 filter=83 channel=11
					-10, -27, -22, 5, 5, -18, 10, 8, 10,
					-- layer=2 filter=83 channel=12
					-15, -16, -4, -23, 12, 14, -26, 25, 21,
					-- layer=2 filter=83 channel=13
					2, 9, -5, 8, 10, -3, 10, -7, -5,
					-- layer=2 filter=83 channel=14
					-1, -16, 21, -1, 6, 22, -6, -8, 8,
					-- layer=2 filter=83 channel=15
					-10, 22, 11, 38, -1, -47, -27, -13, -30,
					-- layer=2 filter=83 channel=16
					47, 58, 8, 9, 3, -24, 2, 35, 9,
					-- layer=2 filter=83 channel=17
					-5, 7, 0, -1, 5, 7, -8, 5, -1,
					-- layer=2 filter=83 channel=18
					43, 10, 52, 0, 19, 15, -1, -16, -6,
					-- layer=2 filter=83 channel=19
					-25, 7, 17, 3, -9, 20, 6, 15, 8,
					-- layer=2 filter=83 channel=20
					0, -5, 3, 9, -1, 2, 0, 3, -3,
					-- layer=2 filter=83 channel=21
					-9, -4, -24, -3, -3, -11, -4, 1, -20,
					-- layer=2 filter=83 channel=22
					5, 9, -9, -1, 9, -5, -5, 2, 0,
					-- layer=2 filter=83 channel=23
					-9, 1, -8, -28, 1, 9, -11, 6, 17,
					-- layer=2 filter=83 channel=24
					23, 17, -20, -56, -37, -62, 18, 5, -24,
					-- layer=2 filter=83 channel=25
					-9, -26, -6, -45, -36, -45, 36, 32, 1,
					-- layer=2 filter=83 channel=26
					-3, 0, 1, 9, 1, 2, 0, -9, 8,
					-- layer=2 filter=83 channel=27
					9, 15, 13, 36, 22, 2, -19, -18, -41,
					-- layer=2 filter=83 channel=28
					4, 14, 8, -5, -21, 30, -32, -29, 18,
					-- layer=2 filter=83 channel=29
					1, 8, 4, 2, 9, 10, -3, 5, -4,
					-- layer=2 filter=83 channel=30
					13, 12, 5, 36, 0, -1, 3, -17, -19,
					-- layer=2 filter=83 channel=31
					47, 13, 37, -14, -62, 6, 61, -13, 43,
					-- layer=2 filter=83 channel=32
					-1, 8, -2, -1, 3, 4, 0, 5, -9,
					-- layer=2 filter=83 channel=33
					-4, 13, 57, 6, -29, 0, -33, -15, 26,
					-- layer=2 filter=83 channel=34
					-6, 7, -41, 53, 15, 5, -1, -10, -25,
					-- layer=2 filter=83 channel=35
					9, 8, 7, 0, 24, 2, 0, -9, 22,
					-- layer=2 filter=83 channel=36
					2, 3, -10, 1, 0, 4, -6, -12, -3,
					-- layer=2 filter=83 channel=37
					-5, 0, -4, 28, 3, 13, 0, -8, 7,
					-- layer=2 filter=83 channel=38
					1, 15, 2, 49, 4, -1, -14, -28, -32,
					-- layer=2 filter=83 channel=39
					48, -15, -16, -27, -12, -13, 13, 1, -22,
					-- layer=2 filter=83 channel=40
					27, 0, 3, -10, 9, 46, -6, 58, -19,
					-- layer=2 filter=83 channel=41
					-7, 11, 4, -6, -5, 4, 3, 10, 10,
					-- layer=2 filter=83 channel=42
					-17, -13, 11, 5, 16, 13, -55, -2, 15,
					-- layer=2 filter=83 channel=43
					38, 31, -4, -27, 10, -21, -27, -18, -35,
					-- layer=2 filter=83 channel=44
					1, -10, 3, 6, -5, 1, -11, 6, 2,
					-- layer=2 filter=83 channel=45
					22, 6, 27, -12, -82, -13, 9, -14, -18,
					-- layer=2 filter=83 channel=46
					11, 13, -25, 7, -15, -37, -20, -21, -27,
					-- layer=2 filter=83 channel=47
					35, 36, 18, 55, 14, 35, -5, 18, 6,
					-- layer=2 filter=83 channel=48
					6, -10, 2, 6, 0, -7, -1, 5, -11,
					-- layer=2 filter=83 channel=49
					-6, 9, 14, -2, 25, 17, -16, -12, -28,
					-- layer=2 filter=83 channel=50
					-17, 5, 5, -9, -2, -2, -13, -30, -5,
					-- layer=2 filter=83 channel=51
					-23, -24, 2, -3, -1, 2, 19, -2, 1,
					-- layer=2 filter=83 channel=52
					-36, -30, -19, -7, 3, 3, -2, 0, 19,
					-- layer=2 filter=83 channel=53
					0, 3, -16, 5, 17, 4, -19, -2, -14,
					-- layer=2 filter=83 channel=54
					-47, -14, -16, -39, 3, -21, 12, 17, 32,
					-- layer=2 filter=83 channel=55
					-5, 2, -8, 2, 7, 0, 8, 3, -2,
					-- layer=2 filter=83 channel=56
					4, -12, -22, -1, -14, -1, -16, 11, 3,
					-- layer=2 filter=83 channel=57
					-3, 0, 2, -3, 4, 4, -10, -7, -8,
					-- layer=2 filter=83 channel=58
					-11, 36, -7, 22, 14, 16, -23, 18, 0,
					-- layer=2 filter=83 channel=59
					28, 35, -8, 6, 32, 1, -12, -4, -20,
					-- layer=2 filter=83 channel=60
					-3, -22, 12, 27, 8, -36, -25, -34, -71,
					-- layer=2 filter=83 channel=61
					-7, 0, -12, -20, 19, -25, -36, 5, -73,
					-- layer=2 filter=83 channel=62
					-31, -11, -3, 35, 14, 27, -21, 31, 23,
					-- layer=2 filter=83 channel=63
					29, -26, -1, -23, 1, -4, -34, -4, -39,
					-- layer=2 filter=83 channel=64
					2, 0, -24, -13, 0, 17, -9, -20, -1,
					-- layer=2 filter=83 channel=65
					6, -6, 9, 19, 11, 15, -10, 3, -14,
					-- layer=2 filter=83 channel=66
					-38, -11, -33, -2, 35, -36, -21, 48, 30,
					-- layer=2 filter=83 channel=67
					16, 49, -16, 19, 10, -51, 17, -42, -66,
					-- layer=2 filter=83 channel=68
					8, -8, -3, 4, 3, 11, 8, -6, -2,
					-- layer=2 filter=83 channel=69
					13, -2, -39, 19, 28, -7, -28, -5, -12,
					-- layer=2 filter=83 channel=70
					0, 26, 6, 15, -20, 17, -34, -43, -1,
					-- layer=2 filter=83 channel=71
					-11, 2, -6, -9, 9, 3, -5, 9, -5,
					-- layer=2 filter=83 channel=72
					-59, -15, 39, -3, -17, 0, -16, -19, 9,
					-- layer=2 filter=83 channel=73
					37, 21, 10, -3, 3, -23, -26, -30, -42,
					-- layer=2 filter=83 channel=74
					2, 1, -16, 7, 15, -29, -9, -35, -24,
					-- layer=2 filter=83 channel=75
					-5, -27, 19, 0, 6, -4, 8, -13, 55,
					-- layer=2 filter=83 channel=76
					22, -29, -44, 26, 15, -27, 1, -7, 0,
					-- layer=2 filter=83 channel=77
					2, 8, -7, 8, -3, 5, 0, 6, 6,
					-- layer=2 filter=83 channel=78
					-24, -33, -6, -24, -17, 1, 9, 12, 28,
					-- layer=2 filter=83 channel=79
					5, 5, 8, -8, -7, -8, -8, 0, -3,
					-- layer=2 filter=83 channel=80
					22, 30, -20, -32, -28, -59, -62, -68, -26,
					-- layer=2 filter=83 channel=81
					-6, -5, 0, -5, -11, -18, -9, -1, -2,
					-- layer=2 filter=83 channel=82
					8, -4, 12, -7, -6, 3, -2, 4, 11,
					-- layer=2 filter=83 channel=83
					8, -16, -10, -10, -21, -23, -36, -28, -21,
					-- layer=2 filter=83 channel=84
					1, -7, -1, 0, -2, 2, 6, 1, 0,
					-- layer=2 filter=83 channel=85
					-14, 4, 12, -1, -8, 2, -11, 7, -16,
					-- layer=2 filter=83 channel=86
					-4, -3, -8, -9, 9, -4, -10, 7, 12,
					-- layer=2 filter=83 channel=87
					36, 43, -31, -15, -7, -40, -3, -10, -42,
					-- layer=2 filter=83 channel=88
					33, 9, -1, 32, 4, 17, 2, 1, -19,
					-- layer=2 filter=83 channel=89
					-22, -10, -10, 3, 17, 11, 0, 2, 25,
					-- layer=2 filter=83 channel=90
					-1, 7, 10, 2, 8, -11, 5, 4, 9,
					-- layer=2 filter=83 channel=91
					-19, 9, -3, 33, 18, -5, 12, 11, 5,
					-- layer=2 filter=83 channel=92
					-17, -14, 10, 6, 15, 17, -9, -24, 7,
					-- layer=2 filter=83 channel=93
					6, -5, 35, 14, 2, 33, -1, 23, 37,
					-- layer=2 filter=83 channel=94
					-26, 2, 4, -28, 12, 0, 6, 34, 20,
					-- layer=2 filter=83 channel=95
					2, -3, 8, -3, -9, -10, 1, 8, -2,
					-- layer=2 filter=83 channel=96
					47, -21, -13, 25, 77, 36, 51, 90, 24,
					-- layer=2 filter=83 channel=97
					31, 43, 14, 1, -27, 11, -51, -44, 8,
					-- layer=2 filter=83 channel=98
					-9, 6, 5, 8, -12, 21, -16, -18, 6,
					-- layer=2 filter=83 channel=99
					-44, -25, 4, 38, 39, 14, 28, 12, 19,
					-- layer=2 filter=83 channel=100
					28, -13, -16, 23, 8, -37, -45, -56, -54,
					-- layer=2 filter=83 channel=101
					-18, -13, 3, -17, -11, 8, -26, 11, 11,
					-- layer=2 filter=83 channel=102
					6, -18, -16, 8, 35, -14, 19, 34, 33,
					-- layer=2 filter=83 channel=103
					-19, -31, -9, -17, -23, 12, 23, -33, -9,
					-- layer=2 filter=83 channel=104
					6, 19, -23, -30, 37, 9, -10, -15, 0,
					-- layer=2 filter=83 channel=105
					-13, -16, -6, 63, -7, 2, -1, 31, 18,
					-- layer=2 filter=83 channel=106
					-29, 25, 2, -22, -24, -1, -4, -8, -13,
					-- layer=2 filter=83 channel=107
					-12, 0, 27, -9, -16, -20, -6, 39, -36,
					-- layer=2 filter=83 channel=108
					-26, -12, 5, -9, 20, 5, -5, -1, 2,
					-- layer=2 filter=83 channel=109
					4, 5, 3, -2, -3, -8, -14, 3, -8,
					-- layer=2 filter=83 channel=110
					21, 11, 5, -11, 24, 16, 37, 13, 7,
					-- layer=2 filter=83 channel=111
					11, 11, 12, -2, -4, 6, -6, 9, 2,
					-- layer=2 filter=83 channel=112
					23, 29, 14, 14, 31, 10, 30, -13, -25,
					-- layer=2 filter=83 channel=113
					-2, 7, 0, 28, -20, 20, -46, -31, -40,
					-- layer=2 filter=83 channel=114
					7, 5, 10, 5, -1, 0, 5, 0, -4,
					-- layer=2 filter=83 channel=115
					6, 4, -3, 3, 1, -3, -1, 7, -11,
					-- layer=2 filter=83 channel=116
					7, 13, -24, 3, 32, -50, 15, 20, -21,
					-- layer=2 filter=83 channel=117
					-46, 2, 9, -4, 31, 0, 3, -12, 31,
					-- layer=2 filter=83 channel=118
					22, 17, -10, -12, -13, -15, -17, 0, 1,
					-- layer=2 filter=83 channel=119
					43, 18, 12, 10, 23, 5, 9, -7, -5,
					-- layer=2 filter=83 channel=120
					-6, -2, 0, 8, -2, 10, -10, 5, -5,
					-- layer=2 filter=83 channel=121
					-8, -7, -8, 8, -6, 3, 6, -6, 5,
					-- layer=2 filter=83 channel=122
					-5, -3, 7, 16, 0, 4, 1, -1, 5,
					-- layer=2 filter=83 channel=123
					-9, -9, 45, 4, -25, 25, 3, 21, 22,
					-- layer=2 filter=83 channel=124
					6, 8, -45, 38, -14, -3, -22, -1, 13,
					-- layer=2 filter=83 channel=125
					0, -3, 8, 6, -3, 0, -8, 5, 1,
					-- layer=2 filter=83 channel=126
					19, -1, 1, -19, 17, -55, -43, -7, -29,
					-- layer=2 filter=83 channel=127
					-7, -19, -4, 11, -3, 14, -31, -17, -21,
					-- layer=2 filter=84 channel=0
					11, -3, -1, -10, -2, 0, 3, 6, -6,
					-- layer=2 filter=84 channel=1
					-11, -22, -19, -21, -12, -8, -2, -9, -7,
					-- layer=2 filter=84 channel=2
					7, -4, -1, -5, -5, -6, -3, 2, 6,
					-- layer=2 filter=84 channel=3
					-6, -22, 1, -12, 6, 12, -22, -12, -14,
					-- layer=2 filter=84 channel=4
					-7, -11, -24, -11, -10, 0, -9, 5, -14,
					-- layer=2 filter=84 channel=5
					10, -12, -2, 5, -25, -16, -8, -13, -6,
					-- layer=2 filter=84 channel=6
					-13, 4, 15, -4, 4, -6, 4, -1, -2,
					-- layer=2 filter=84 channel=7
					1, -4, -7, -2, 6, -15, 7, 6, -17,
					-- layer=2 filter=84 channel=8
					-1, -5, 9, -8, -4, -3, -11, 4, -1,
					-- layer=2 filter=84 channel=9
					0, 10, 3, -6, 1, 8, 0, -2, -8,
					-- layer=2 filter=84 channel=10
					-11, -14, -1, -4, -24, -6, 5, -20, 15,
					-- layer=2 filter=84 channel=11
					-11, -4, -13, -23, -11, 0, -7, -5, -8,
					-- layer=2 filter=84 channel=12
					1, -13, -23, -9, -9, 6, -2, -17, -9,
					-- layer=2 filter=84 channel=13
					0, -3, 1, 1, 3, 1, -9, -9, -1,
					-- layer=2 filter=84 channel=14
					0, 4, -24, -6, 1, -11, -8, -8, -16,
					-- layer=2 filter=84 channel=15
					0, -4, 2, -19, 11, -8, -7, -9, -7,
					-- layer=2 filter=84 channel=16
					-3, -12, -9, 1, -8, -7, 0, 1, -8,
					-- layer=2 filter=84 channel=17
					1, 4, -7, 9, -7, -2, 6, 2, -8,
					-- layer=2 filter=84 channel=18
					0, -4, -10, 0, 2, 3, -16, 6, -2,
					-- layer=2 filter=84 channel=19
					-8, -11, -17, -6, -22, -19, 14, -5, -3,
					-- layer=2 filter=84 channel=20
					6, -5, -1, -6, 4, -4, 1, -7, 3,
					-- layer=2 filter=84 channel=21
					-5, -6, 5, -5, 4, -7, -3, 7, -6,
					-- layer=2 filter=84 channel=22
					0, 10, 4, 9, 6, 3, -9, 0, -1,
					-- layer=2 filter=84 channel=23
					-3, -13, -10, -3, -11, -15, 3, -4, -18,
					-- layer=2 filter=84 channel=24
					-8, -9, -2, -10, -6, -4, -11, 0, 9,
					-- layer=2 filter=84 channel=25
					-5, 3, 6, -13, -2, 2, -6, 1, 16,
					-- layer=2 filter=84 channel=26
					3, -3, 0, -8, 9, 10, -7, 1, -2,
					-- layer=2 filter=84 channel=27
					-10, -10, -14, 10, 5, 0, -5, 1, -6,
					-- layer=2 filter=84 channel=28
					-1, -11, 15, -12, -2, -1, -21, -8, -3,
					-- layer=2 filter=84 channel=29
					-3, -2, -1, -2, -11, -1, 6, 2, -8,
					-- layer=2 filter=84 channel=30
					0, -5, -1, -5, -2, -14, 2, 0, -7,
					-- layer=2 filter=84 channel=31
					-9, 11, 3, -5, 2, -11, -17, -5, -3,
					-- layer=2 filter=84 channel=32
					0, -8, 3, 0, -11, 6, -5, -8, 0,
					-- layer=2 filter=84 channel=33
					-8, -10, -3, -6, 1, -7, -2, 1, 0,
					-- layer=2 filter=84 channel=34
					0, 6, -7, 0, -17, -8, 11, -13, -15,
					-- layer=2 filter=84 channel=35
					-15, -5, 3, -8, 2, 1, 8, 9, -17,
					-- layer=2 filter=84 channel=36
					-11, -3, -10, 0, -10, -10, -1, 0, -3,
					-- layer=2 filter=84 channel=37
					-5, -9, 0, -1, -14, -12, -12, -12, -17,
					-- layer=2 filter=84 channel=38
					-4, -9, -16, 0, -14, 7, 3, -16, 1,
					-- layer=2 filter=84 channel=39
					-22, 0, -3, 1, -3, -12, 14, -8, -22,
					-- layer=2 filter=84 channel=40
					-1, -7, 8, 0, -9, -8, -2, -17, 2,
					-- layer=2 filter=84 channel=41
					-6, -4, -7, 9, -4, -6, 3, 0, 6,
					-- layer=2 filter=84 channel=42
					-15, -13, -9, -8, 10, 7, -18, 0, -21,
					-- layer=2 filter=84 channel=43
					-9, -3, -12, -6, -14, 8, -22, 2, -16,
					-- layer=2 filter=84 channel=44
					8, -5, 5, 5, -8, -6, 6, 4, 3,
					-- layer=2 filter=84 channel=45
					-5, 1, 6, 1, 12, -8, 5, 4, 8,
					-- layer=2 filter=84 channel=46
					0, 2, -1, -2, -15, 16, -3, 2, 11,
					-- layer=2 filter=84 channel=47
					-22, -7, -2, -1, -18, -9, -3, -10, -8,
					-- layer=2 filter=84 channel=48
					2, -11, 4, -8, 10, 7, 1, 7, 8,
					-- layer=2 filter=84 channel=49
					-6, -10, 3, -14, -28, -1, -22, -18, -16,
					-- layer=2 filter=84 channel=50
					-2, -9, -1, 7, -5, 0, -4, -6, 8,
					-- layer=2 filter=84 channel=51
					-2, -8, -10, -14, -6, -3, -6, -17, -10,
					-- layer=2 filter=84 channel=52
					-8, -25, -10, -15, -1, -5, -8, -6, -12,
					-- layer=2 filter=84 channel=53
					-7, 4, -3, 1, 5, 6, -1, -4, -2,
					-- layer=2 filter=84 channel=54
					-15, -13, 0, -18, -12, -10, -18, -5, -5,
					-- layer=2 filter=84 channel=55
					-6, 1, 5, -11, -7, 5, -4, 4, -1,
					-- layer=2 filter=84 channel=56
					-1, -17, -18, -8, -12, -3, -10, -6, -11,
					-- layer=2 filter=84 channel=57
					-8, -11, -1, -8, 4, -2, 1, 5, -10,
					-- layer=2 filter=84 channel=58
					13, 0, -11, 6, -3, -7, 4, -8, 3,
					-- layer=2 filter=84 channel=59
					-3, 1, -1, 18, -1, 0, -8, -11, -9,
					-- layer=2 filter=84 channel=60
					-6, 0, -8, 1, -2, -2, -22, -15, -13,
					-- layer=2 filter=84 channel=61
					-5, 0, 2, 18, -17, -14, -1, -19, -3,
					-- layer=2 filter=84 channel=62
					-8, 5, -22, -11, 4, -26, -7, -12, -12,
					-- layer=2 filter=84 channel=63
					-8, 3, 2, 3, -19, -1, -4, -4, -13,
					-- layer=2 filter=84 channel=64
					-9, -3, -6, -2, -11, 1, 10, 12, -4,
					-- layer=2 filter=84 channel=65
					-4, -13, -7, -13, -12, 2, -13, -12, -18,
					-- layer=2 filter=84 channel=66
					-1, -6, -7, -6, 7, 0, 1, 0, -5,
					-- layer=2 filter=84 channel=67
					-9, -5, 4, -10, 2, -15, -7, -9, 4,
					-- layer=2 filter=84 channel=68
					0, -6, -11, -4, 5, -4, 2, -4, -6,
					-- layer=2 filter=84 channel=69
					8, 6, -20, 9, 7, -7, -19, -18, -2,
					-- layer=2 filter=84 channel=70
					-15, -14, -15, -16, -2, -12, -3, -4, -9,
					-- layer=2 filter=84 channel=71
					20, -11, 6, 2, 0, 2, -1, -1, -20,
					-- layer=2 filter=84 channel=72
					-6, -19, 4, 14, 13, -25, -4, 5, -17,
					-- layer=2 filter=84 channel=73
					-10, 6, 15, -17, -21, -5, -13, 1, -6,
					-- layer=2 filter=84 channel=74
					-4, -5, 5, -7, -7, -1, 5, -4, 2,
					-- layer=2 filter=84 channel=75
					2, 1, -8, -18, -4, 0, -3, -8, -13,
					-- layer=2 filter=84 channel=76
					-18, -4, 10, -14, 1, 2, -6, -22, -6,
					-- layer=2 filter=84 channel=77
					9, 0, -10, 7, 6, -3, 8, 8, 5,
					-- layer=2 filter=84 channel=78
					-13, -6, 0, -15, -6, 5, -5, -17, -11,
					-- layer=2 filter=84 channel=79
					8, 0, -10, 0, 4, 0, 4, -7, -7,
					-- layer=2 filter=84 channel=80
					-6, -7, -1, -4, -2, -6, -1, 3, -5,
					-- layer=2 filter=84 channel=81
					-9, -1, -10, 6, -8, 1, 9, -4, -1,
					-- layer=2 filter=84 channel=82
					-12, 0, -10, 8, -8, -11, -11, 2, 5,
					-- layer=2 filter=84 channel=83
					-13, 5, -6, -9, -4, -6, -12, 2, -4,
					-- layer=2 filter=84 channel=84
					5, -8, 9, 5, -8, 1, -1, 1, 8,
					-- layer=2 filter=84 channel=85
					0, -11, -7, -3, -9, 7, -5, 8, 4,
					-- layer=2 filter=84 channel=86
					-11, -7, 3, 5, -5, 8, 10, 9, -1,
					-- layer=2 filter=84 channel=87
					0, -5, 0, -9, 7, 2, -9, 8, 7,
					-- layer=2 filter=84 channel=88
					8, -2, 4, -10, -7, -5, -15, -17, -1,
					-- layer=2 filter=84 channel=89
					-11, -2, -5, 5, -1, 8, -3, -22, 0,
					-- layer=2 filter=84 channel=90
					8, -4, 9, -4, 7, 2, -10, -6, 8,
					-- layer=2 filter=84 channel=91
					14, -6, -8, -10, 11, -14, -12, -12, -28,
					-- layer=2 filter=84 channel=92
					0, -10, -15, -1, 4, -1, 7, -14, 2,
					-- layer=2 filter=84 channel=93
					-11, -3, 16, -20, 6, -17, -8, -18, -5,
					-- layer=2 filter=84 channel=94
					-21, -8, -3, 16, -12, 1, -21, -13, -10,
					-- layer=2 filter=84 channel=95
					-1, 5, 4, -3, -9, -2, -1, 8, -8,
					-- layer=2 filter=84 channel=96
					17, 6, -5, 1, 0, -11, -21, -7, -17,
					-- layer=2 filter=84 channel=97
					-7, -12, -3, -19, -8, -5, -10, 4, -6,
					-- layer=2 filter=84 channel=98
					-24, 0, -12, -4, -4, -17, -9, -6, -14,
					-- layer=2 filter=84 channel=99
					-8, 9, -24, -12, -7, -24, -4, 0, 10,
					-- layer=2 filter=84 channel=100
					-2, -12, -24, 6, -11, 3, -7, 3, -13,
					-- layer=2 filter=84 channel=101
					-13, -28, 5, -10, 5, -6, -4, -7, 0,
					-- layer=2 filter=84 channel=102
					12, 4, -21, -1, 1, -6, -5, 2, -13,
					-- layer=2 filter=84 channel=103
					3, -4, 0, 6, 4, 2, 9, -10, 6,
					-- layer=2 filter=84 channel=104
					-6, -11, -8, 7, -1, -3, -10, 3, -20,
					-- layer=2 filter=84 channel=105
					-7, -7, 7, 1, -3, -7, 1, -3, -15,
					-- layer=2 filter=84 channel=106
					-3, -16, -4, 2, -17, 5, 9, -2, 13,
					-- layer=2 filter=84 channel=107
					0, 9, 0, -18, 8, 1, 0, 5, -9,
					-- layer=2 filter=84 channel=108
					2, 11, -16, 17, 8, -1, -2, -3, -13,
					-- layer=2 filter=84 channel=109
					-4, 4, -2, -6, 4, -9, 7, 4, -4,
					-- layer=2 filter=84 channel=110
					-7, -8, -14, -1, -16, -10, 2, 4, -17,
					-- layer=2 filter=84 channel=111
					-1, 10, -4, -5, 0, -4, -8, 0, 8,
					-- layer=2 filter=84 channel=112
					-5, 2, 3, -14, -8, -1, 1, -6, 10,
					-- layer=2 filter=84 channel=113
					0, 5, 0, -14, -12, -12, 8, -5, 0,
					-- layer=2 filter=84 channel=114
					9, -8, 7, 0, 4, -11, 4, -6, -3,
					-- layer=2 filter=84 channel=115
					3, 5, -2, 5, 4, -7, -3, -5, 0,
					-- layer=2 filter=84 channel=116
					-1, -15, -6, -13, 2, -4, -8, -5, -7,
					-- layer=2 filter=84 channel=117
					-4, -3, -10, -3, -12, -6, -7, -5, -6,
					-- layer=2 filter=84 channel=118
					-6, -3, -13, -7, -12, 5, -6, -13, -7,
					-- layer=2 filter=84 channel=119
					-7, -13, -16, 1, -3, -18, -11, 3, -8,
					-- layer=2 filter=84 channel=120
					2, 0, 2, -7, -3, 9, 6, 9, 2,
					-- layer=2 filter=84 channel=121
					8, -6, -3, 6, 0, -9, -7, -1, -1,
					-- layer=2 filter=84 channel=122
					-8, -7, 0, 10, 3, 1, 0, 5, 5,
					-- layer=2 filter=84 channel=123
					-8, 6, -2, 1, 1, -3, 10, -16, -29,
					-- layer=2 filter=84 channel=124
					4, -13, 6, -1, 11, 14, -12, -14, 2,
					-- layer=2 filter=84 channel=125
					-1, -12, 0, 6, 0, -2, -3, 9, -6,
					-- layer=2 filter=84 channel=126
					5, 14, 8, 2, 7, -9, -10, -4, -8,
					-- layer=2 filter=84 channel=127
					3, 1, -7, 1, 1, -21, 0, -13, -19,
					-- layer=2 filter=85 channel=0
					10, 15, 7, 12, 26, 26, 0, 10, 0,
					-- layer=2 filter=85 channel=1
					24, 14, -37, 5, -2, -4, 0, -22, -15,
					-- layer=2 filter=85 channel=2
					-7, -11, -9, 6, -9, 0, -5, -3, 4,
					-- layer=2 filter=85 channel=3
					-27, -7, -9, -35, 16, -4, 7, 3, -2,
					-- layer=2 filter=85 channel=4
					19, 21, -5, 11, 18, 23, -32, -12, -19,
					-- layer=2 filter=85 channel=5
					-14, -25, -14, -11, 13, -7, 18, 42, -14,
					-- layer=2 filter=85 channel=6
					27, -42, -19, -2, -58, -30, 23, -25, -69,
					-- layer=2 filter=85 channel=7
					-60, -38, -13, -11, -14, -19, -5, 14, 38,
					-- layer=2 filter=85 channel=8
					7, -11, 6, 7, -8, 2, 9, -3, -4,
					-- layer=2 filter=85 channel=9
					0, 3, -4, -8, 16, -19, 2, 13, 15,
					-- layer=2 filter=85 channel=10
					22, 9, 3, 0, 23, 16, 15, 10, -13,
					-- layer=2 filter=85 channel=11
					-16, -27, -18, 8, 0, -12, 25, 14, -7,
					-- layer=2 filter=85 channel=12
					29, 22, -37, 12, 11, 29, -5, -7, 0,
					-- layer=2 filter=85 channel=13
					-11, -5, -7, 3, -11, -6, 5, 5, -11,
					-- layer=2 filter=85 channel=14
					16, 8, -24, 14, -23, -20, 13, -20, -17,
					-- layer=2 filter=85 channel=15
					-4, -1, 55, -48, -54, -25, -21, -17, -131,
					-- layer=2 filter=85 channel=16
					-4, -7, -17, -28, -17, -22, -18, 0, 23,
					-- layer=2 filter=85 channel=17
					7, 4, -7, -1, -9, -6, 2, 8, -6,
					-- layer=2 filter=85 channel=18
					4, -73, -54, -5, -65, 20, 0, -38, -49,
					-- layer=2 filter=85 channel=19
					-18, -12, 20, 21, 10, -8, -22, -45, -40,
					-- layer=2 filter=85 channel=20
					10, 0, -5, -3, 3, -7, 6, 7, -11,
					-- layer=2 filter=85 channel=21
					-23, -12, -12, 0, -4, -7, -31, -23, 0,
					-- layer=2 filter=85 channel=22
					4, -5, 4, 5, -3, 1, 10, -11, 0,
					-- layer=2 filter=85 channel=23
					23, 3, -27, 14, -3, -3, 7, 8, 30,
					-- layer=2 filter=85 channel=24
					8, 7, -5, -2, 16, -12, 18, 17, 21,
					-- layer=2 filter=85 channel=25
					-9, -9, 6, 6, 6, 9, 25, 12, 14,
					-- layer=2 filter=85 channel=26
					3, 6, -7, -6, 2, 0, -6, -3, -1,
					-- layer=2 filter=85 channel=27
					20, 18, 35, 21, 17, 17, -21, -26, -1,
					-- layer=2 filter=85 channel=28
					26, 15, 6, -18, -13, 28, -54, -28, 32,
					-- layer=2 filter=85 channel=29
					4, 0, -3, -8, 6, 10, 7, 7, 10,
					-- layer=2 filter=85 channel=30
					14, 3, 19, 14, 10, -22, 0, 0, 2,
					-- layer=2 filter=85 channel=31
					-24, 41, 78, -34, -1, -51, 36, 30, -67,
					-- layer=2 filter=85 channel=32
					-3, -7, -6, 4, 0, -3, 2, 0, 6,
					-- layer=2 filter=85 channel=33
					-43, 7, -2, 30, 0, -24, 11, 22, 16,
					-- layer=2 filter=85 channel=34
					6, -78, -32, -7, 31, -17, 70, 23, 33,
					-- layer=2 filter=85 channel=35
					3, 23, 20, -38, -11, 8, -23, -34, 37,
					-- layer=2 filter=85 channel=36
					-3, 1, -3, -2, 1, 5, 2, 9, -13,
					-- layer=2 filter=85 channel=37
					-6, -25, -11, 8, -1, -21, 21, 27, -28,
					-- layer=2 filter=85 channel=38
					1, 27, 15, 5, 22, -8, 1, 0, -9,
					-- layer=2 filter=85 channel=39
					6, -2, 13, 3, 1, -29, -2, -12, 21,
					-- layer=2 filter=85 channel=40
					-76, -23, 37, -53, -37, -15, 12, -42, -3,
					-- layer=2 filter=85 channel=41
					3, -2, 6, 7, 9, -8, 6, 8, 6,
					-- layer=2 filter=85 channel=42
					-4, -6, -10, 5, 0, 10, -10, 35, 36,
					-- layer=2 filter=85 channel=43
					-11, -21, -14, -32, 17, -22, -11, 20, -9,
					-- layer=2 filter=85 channel=44
					6, -8, -2, 8, -6, -3, -5, -4, 3,
					-- layer=2 filter=85 channel=45
					-3, 25, 3, -15, 14, 8, -69, -74, 20,
					-- layer=2 filter=85 channel=46
					17, 2, 9, 21, 15, -8, 18, -7, -27,
					-- layer=2 filter=85 channel=47
					9, 43, 35, 10, 23, 30, -31, -37, 44,
					-- layer=2 filter=85 channel=48
					0, -1, 4, 10, -9, 10, -5, 0, 3,
					-- layer=2 filter=85 channel=49
					40, -49, -7, -3, -42, 35, 3, -45, 15,
					-- layer=2 filter=85 channel=50
					-2, -7, 0, 4, -26, -35, -2, -12, 2,
					-- layer=2 filter=85 channel=51
					-3, -4, 18, 6, 12, -20, 16, 42, -10,
					-- layer=2 filter=85 channel=52
					-23, -40, 6, -2, -35, -23, -35, -36, -32,
					-- layer=2 filter=85 channel=53
					39, -60, 26, -19, -51, 15, -30, -36, -52,
					-- layer=2 filter=85 channel=54
					-21, -18, -27, 3, -9, -8, 12, -27, 3,
					-- layer=2 filter=85 channel=55
					6, 0, 11, -4, 8, 4, -8, 1, -3,
					-- layer=2 filter=85 channel=56
					-5, -25, -33, 19, -8, -8, 23, 34, -6,
					-- layer=2 filter=85 channel=57
					-12, 0, -6, -9, -10, -7, 11, -4, 9,
					-- layer=2 filter=85 channel=58
					-12, 48, -36, -9, 20, 32, 5, -21, 21,
					-- layer=2 filter=85 channel=59
					-5, 22, -1, 10, -3, 13, -33, -58, 15,
					-- layer=2 filter=85 channel=60
					10, 5, 20, -11, 7, 19, -1, -23, -31,
					-- layer=2 filter=85 channel=61
					4, 4, 43, -17, 8, 3, -51, -18, -6,
					-- layer=2 filter=85 channel=62
					7, -95, 25, 36, -33, -60, 41, -26, -41,
					-- layer=2 filter=85 channel=63
					39, 14, 9, -2, 14, 15, -8, -14, 31,
					-- layer=2 filter=85 channel=64
					26, 3, 4, 9, -1, 2, 17, 20, 20,
					-- layer=2 filter=85 channel=65
					-5, 11, 15, 7, -6, 1, 12, -1, -58,
					-- layer=2 filter=85 channel=66
					17, -13, 3, 8, 30, -32, 1, -12, -33,
					-- layer=2 filter=85 channel=67
					-1, -23, -11, -3, 15, -12, 9, 18, -20,
					-- layer=2 filter=85 channel=68
					-3, 0, -6, -5, 8, -2, -4, 7, 10,
					-- layer=2 filter=85 channel=69
					26, 10, 0, -8, -11, -9, 7, 0, 33,
					-- layer=2 filter=85 channel=70
					8, 17, 25, -4, -13, 11, -43, -6, 18,
					-- layer=2 filter=85 channel=71
					8, 44, 61, 23, 22, 28, -20, -22, 11,
					-- layer=2 filter=85 channel=72
					-8, -19, -3, 16, -11, -16, -1, -13, -13,
					-- layer=2 filter=85 channel=73
					11, -47, 25, -44, 15, 19, 36, -29, 8,
					-- layer=2 filter=85 channel=74
					9, 17, -2, 6, 24, 16, 23, 11, 6,
					-- layer=2 filter=85 channel=75
					-16, 26, -15, -12, 16, 8, -18, -14, 5,
					-- layer=2 filter=85 channel=76
					25, -41, 32, -42, -11, -32, 27, -9, -31,
					-- layer=2 filter=85 channel=77
					-9, 0, 6, -10, 0, 4, 8, 3, 8,
					-- layer=2 filter=85 channel=78
					2, -26, -28, 28, -11, -13, 21, 10, -28,
					-- layer=2 filter=85 channel=79
					1, -2, -3, -4, -1, 0, 4, -7, 3,
					-- layer=2 filter=85 channel=80
					-3, 14, 6, -8, 7, -2, -43, -11, -19,
					-- layer=2 filter=85 channel=81
					-4, 9, -2, -5, -2, 3, -6, -1, 14,
					-- layer=2 filter=85 channel=82
					-4, 9, 11, -8, -3, -5, 6, 5, 9,
					-- layer=2 filter=85 channel=83
					5, 23, 1, 24, 1, 0, -39, -10, -6,
					-- layer=2 filter=85 channel=84
					-2, -6, 0, -5, 11, 2, -7, -5, 4,
					-- layer=2 filter=85 channel=85
					3, 0, -4, -7, -6, -4, -8, -11, 0,
					-- layer=2 filter=85 channel=86
					5, 1, -21, 5, 16, 1, -6, 3, 0,
					-- layer=2 filter=85 channel=87
					-12, -60, 3, -47, -70, -7, -2, 45, 38,
					-- layer=2 filter=85 channel=88
					41, 31, -5, -17, 18, -10, 16, 3, -1,
					-- layer=2 filter=85 channel=89
					-3, 6, -17, 2, -15, 8, 22, -4, 0,
					-- layer=2 filter=85 channel=90
					-7, -11, 2, -3, 11, -3, 7, 7, 7,
					-- layer=2 filter=85 channel=91
					-18, 17, -8, 3, 35, 43, -1, 3, 0,
					-- layer=2 filter=85 channel=92
					-1, 27, -16, -12, -10, 13, 14, -6, -1,
					-- layer=2 filter=85 channel=93
					-19, -63, 59, -2, -44, 22, 53, -36, -88,
					-- layer=2 filter=85 channel=94
					-17, 1, -10, -19, -63, -28, -44, -71, -34,
					-- layer=2 filter=85 channel=95
					0, -6, -4, 4, -12, -15, 1, 3, -12,
					-- layer=2 filter=85 channel=96
					12, -49, -8, 0, -53, 7, 4, -45, 38,
					-- layer=2 filter=85 channel=97
					-17, 37, -12, -2, 32, 17, 10, 11, 30,
					-- layer=2 filter=85 channel=98
					-4, 19, 12, 4, 0, 4, -23, -16, 33,
					-- layer=2 filter=85 channel=99
					-35, 4, 25, -42, -2, -4, -85, -60, -28,
					-- layer=2 filter=85 channel=100
					24, 45, 11, 1, 23, 12, 4, -17, 6,
					-- layer=2 filter=85 channel=101
					-9, 14, 11, -11, -8, 18, -5, -15, -7,
					-- layer=2 filter=85 channel=102
					-9, -104, -28, -10, -51, -12, 7, -73, -33,
					-- layer=2 filter=85 channel=103
					-19, -4, -21, -20, -37, 9, 31, 75, 10,
					-- layer=2 filter=85 channel=104
					15, -40, -11, -1, -74, -2, -6, -79, -5,
					-- layer=2 filter=85 channel=105
					-67, 6, -6, -28, -11, -92, 6, -4, -1,
					-- layer=2 filter=85 channel=106
					1, -13, -12, 7, 13, -3, 7, 20, 6,
					-- layer=2 filter=85 channel=107
					-34, -9, 2, 87, 23, 29, -34, 36, -22,
					-- layer=2 filter=85 channel=108
					25, 17, 36, -7, -9, -5, -36, -37, -6,
					-- layer=2 filter=85 channel=109
					-10, -11, -11, -3, 4, -1, 3, 7, -16,
					-- layer=2 filter=85 channel=110
					10, -17, -1, -58, 7, 2, -19, 9, 26,
					-- layer=2 filter=85 channel=111
					4, -3, 6, 5, 6, 1, 3, 4, -1,
					-- layer=2 filter=85 channel=112
					-5, -6, 52, 8, 18, 4, 12, 20, 5,
					-- layer=2 filter=85 channel=113
					33, 18, 18, 1, 11, 13, 1, 6, 21,
					-- layer=2 filter=85 channel=114
					4, 0, -13, -8, -4, 5, 7, 1, -10,
					-- layer=2 filter=85 channel=115
					-1, 3, -5, 7, -9, -7, 7, -1, 8,
					-- layer=2 filter=85 channel=116
					12, -47, 7, -44, -66, 20, -6, 4, 7,
					-- layer=2 filter=85 channel=117
					-91, -32, -15, -37, -57, -22, -7, -7, -24,
					-- layer=2 filter=85 channel=118
					2, 2, 3, 7, 7, 16, -8, 9, -3,
					-- layer=2 filter=85 channel=119
					27, 0, -34, 9, -19, -13, 26, -40, 21,
					-- layer=2 filter=85 channel=120
					8, 5, -1, -7, 5, -8, 9, 5, 2,
					-- layer=2 filter=85 channel=121
					-8, 7, 0, -5, -6, 0, -2, 6, -5,
					-- layer=2 filter=85 channel=122
					-1, -12, 6, -6, -5, 5, -2, -5, -1,
					-- layer=2 filter=85 channel=123
					-44, -21, 5, 37, -5, -18, -17, -11, -2,
					-- layer=2 filter=85 channel=124
					-62, -60, -22, 8, -40, -28, 6, 21, 10,
					-- layer=2 filter=85 channel=125
					-2, 6, 2, -3, 1, 7, 1, -8, -7,
					-- layer=2 filter=85 channel=126
					-12, 42, 31, -7, 111, 0, 11, 60, 24,
					-- layer=2 filter=85 channel=127
					58, 2, -5, 37, 4, 0, -25, -1, 16,
					-- layer=2 filter=86 channel=0
					4, 3, -3, -3, -2, 2, 0, 3, 5,
					-- layer=2 filter=86 channel=1
					-4, -18, -3, 3, -14, -8, -14, -2, -7,
					-- layer=2 filter=86 channel=2
					8, -7, -1, 3, 0, 0, 1, 2, -2,
					-- layer=2 filter=86 channel=3
					4, -7, -11, -17, 1, -2, 0, -2, 3,
					-- layer=2 filter=86 channel=4
					5, -12, -7, 0, 4, 8, -10, -9, -2,
					-- layer=2 filter=86 channel=5
					3, -8, -9, -7, -19, -3, -3, -10, 4,
					-- layer=2 filter=86 channel=6
					1, -17, 4, 5, 14, -6, -10, -5, -24,
					-- layer=2 filter=86 channel=7
					-9, 10, -13, -2, -10, -10, -13, -13, -4,
					-- layer=2 filter=86 channel=8
					0, -3, -5, 3, 0, -7, 0, -3, -5,
					-- layer=2 filter=86 channel=9
					1, -12, -9, -2, -8, 7, 2, -14, -3,
					-- layer=2 filter=86 channel=10
					0, 4, -1, -8, -8, -4, -1, 2, -1,
					-- layer=2 filter=86 channel=11
					0, 0, 0, -15, -12, -9, 4, -12, -3,
					-- layer=2 filter=86 channel=12
					5, -5, -1, -12, 5, -1, -22, -8, -23,
					-- layer=2 filter=86 channel=13
					5, -2, -3, 5, 8, -6, 0, 4, 4,
					-- layer=2 filter=86 channel=14
					10, -7, -11, 4, -18, -1, -11, -10, -12,
					-- layer=2 filter=86 channel=15
					-6, -2, -12, -7, -3, 4, 4, 0, 6,
					-- layer=2 filter=86 channel=16
					-9, 0, 5, 7, -12, 0, 0, 6, 5,
					-- layer=2 filter=86 channel=17
					11, 8, 1, -3, -7, 6, 8, 5, 8,
					-- layer=2 filter=86 channel=18
					0, 7, -5, -9, -3, -6, -4, -10, 4,
					-- layer=2 filter=86 channel=19
					-11, -25, -7, -2, -10, -17, 0, -4, -6,
					-- layer=2 filter=86 channel=20
					-4, 0, -5, -8, -1, -4, -6, -5, -7,
					-- layer=2 filter=86 channel=21
					-1, -7, 0, -5, -4, 9, -6, 9, 2,
					-- layer=2 filter=86 channel=22
					1, -5, -7, 11, 5, -10, 9, -9, -4,
					-- layer=2 filter=86 channel=23
					-11, -2, 5, 12, -12, 2, 0, 8, 4,
					-- layer=2 filter=86 channel=24
					-12, -9, 2, -6, -1, -12, -3, -8, -12,
					-- layer=2 filter=86 channel=25
					7, -1, -11, 0, 8, 5, -3, -6, -4,
					-- layer=2 filter=86 channel=26
					-3, 7, 6, 0, -9, -4, 0, 1, -5,
					-- layer=2 filter=86 channel=27
					1, 3, -17, -2, -10, -19, -13, -7, -3,
					-- layer=2 filter=86 channel=28
					-8, -27, -10, -6, -4, -11, -15, -3, 4,
					-- layer=2 filter=86 channel=29
					4, 1, 3, 2, -5, -2, -7, 1, -4,
					-- layer=2 filter=86 channel=30
					-4, -6, -3, -12, -2, -8, -1, -9, 2,
					-- layer=2 filter=86 channel=31
					-3, -4, 0, 4, -3, -20, 11, 16, 9,
					-- layer=2 filter=86 channel=32
					2, 10, -9, -6, -8, -1, -4, -4, 4,
					-- layer=2 filter=86 channel=33
					3, 1, -2, 6, 0, -4, -8, -7, -9,
					-- layer=2 filter=86 channel=34
					-7, -10, 2, 4, -12, -11, -3, -6, -7,
					-- layer=2 filter=86 channel=35
					-14, -10, -4, 7, -4, 0, -11, 2, -10,
					-- layer=2 filter=86 channel=36
					8, 0, -1, 5, 0, -6, -4, 3, -3,
					-- layer=2 filter=86 channel=37
					-9, -1, -4, -4, -10, -9, 0, -13, -10,
					-- layer=2 filter=86 channel=38
					5, 9, -7, -18, -13, -6, -17, 6, -22,
					-- layer=2 filter=86 channel=39
					-7, 9, -9, 4, 0, -9, -1, -3, -7,
					-- layer=2 filter=86 channel=40
					8, -9, 2, -3, 12, -14, -13, 0, 7,
					-- layer=2 filter=86 channel=41
					-7, -8, -5, -1, -7, 11, 3, 5, -6,
					-- layer=2 filter=86 channel=42
					0, -10, 7, -10, 0, -1, 3, -6, -11,
					-- layer=2 filter=86 channel=43
					4, -6, -5, -13, -16, 7, -4, 0, -4,
					-- layer=2 filter=86 channel=44
					0, -4, -4, 2, 1, 8, -4, -4, 2,
					-- layer=2 filter=86 channel=45
					8, -9, -14, -1, -12, -8, 1, -7, 9,
					-- layer=2 filter=86 channel=46
					1, -13, 2, -10, 0, 3, 3, 0, -5,
					-- layer=2 filter=86 channel=47
					5, -15, -2, -3, 1, -4, -2, 0, -3,
					-- layer=2 filter=86 channel=48
					-6, 6, -2, 2, 2, 2, 4, 9, 7,
					-- layer=2 filter=86 channel=49
					-6, 3, -19, -11, -29, -22, -8, -3, -21,
					-- layer=2 filter=86 channel=50
					0, -8, -5, -7, 0, 0, 4, -5, -7,
					-- layer=2 filter=86 channel=51
					-6, -4, -12, -7, -8, -8, -13, 0, -6,
					-- layer=2 filter=86 channel=52
					-6, -21, -8, 0, -23, -2, -22, -26, -3,
					-- layer=2 filter=86 channel=53
					-7, -2, 1, 3, 0, -8, 2, 6, -2,
					-- layer=2 filter=86 channel=54
					-3, -14, -21, -10, 0, -12, -2, -16, -14,
					-- layer=2 filter=86 channel=55
					2, 4, 6, -1, 9, 2, -3, 8, 1,
					-- layer=2 filter=86 channel=56
					1, -11, 4, -14, 4, 3, -12, -13, 0,
					-- layer=2 filter=86 channel=57
					6, 0, -9, 0, -7, -4, -8, 0, 6,
					-- layer=2 filter=86 channel=58
					6, -3, 0, 9, -7, -6, -10, -4, -9,
					-- layer=2 filter=86 channel=59
					1, -10, 0, -6, -11, -2, -3, -14, -12,
					-- layer=2 filter=86 channel=60
					-16, -4, -6, -4, 2, -5, -7, -13, -11,
					-- layer=2 filter=86 channel=61
					-23, -5, -5, -14, -3, 3, 0, -12, -17,
					-- layer=2 filter=86 channel=62
					-8, -9, -3, 10, 7, 4, -18, 0, -10,
					-- layer=2 filter=86 channel=63
					0, 2, -5, 7, 2, -1, 4, -11, -10,
					-- layer=2 filter=86 channel=64
					-5, 0, 6, 7, -1, 7, 0, 3, -2,
					-- layer=2 filter=86 channel=65
					3, -20, 4, 0, 5, 1, -10, 1, -1,
					-- layer=2 filter=86 channel=66
					3, 3, 1, -1, 8, 18, -4, -6, 11,
					-- layer=2 filter=86 channel=67
					1, 6, 0, -3, -3, -8, 7, 2, -8,
					-- layer=2 filter=86 channel=68
					-1, 0, 4, 0, 6, -4, -1, 9, 2,
					-- layer=2 filter=86 channel=69
					-1, -8, -10, -18, -13, 6, 0, -10, -9,
					-- layer=2 filter=86 channel=70
					-2, -6, -13, -12, 4, -14, 0, -4, 0,
					-- layer=2 filter=86 channel=71
					4, 0, -3, -13, -11, -2, 6, -10, -10,
					-- layer=2 filter=86 channel=72
					9, 11, -8, -3, -3, -8, 14, 3, 3,
					-- layer=2 filter=86 channel=73
					-7, -10, -16, -16, -26, -8, -1, -8, -1,
					-- layer=2 filter=86 channel=74
					-2, -10, -1, 8, -2, -12, 2, -2, -8,
					-- layer=2 filter=86 channel=75
					-4, -10, 5, 0, 6, 8, -6, -8, 8,
					-- layer=2 filter=86 channel=76
					-1, -7, -7, -4, 3, -12, -14, 0, -9,
					-- layer=2 filter=86 channel=77
					6, -6, 3, 2, -1, 7, 10, 0, 2,
					-- layer=2 filter=86 channel=78
					-15, -3, -14, -16, -9, -8, -12, -2, -6,
					-- layer=2 filter=86 channel=79
					2, 7, 5, -4, -2, 11, 1, 7, -7,
					-- layer=2 filter=86 channel=80
					-10, -3, 7, 4, 8, -3, -5, -5, -5,
					-- layer=2 filter=86 channel=81
					3, -7, 0, 0, -3, -10, 8, 6, -8,
					-- layer=2 filter=86 channel=82
					-3, -5, 10, 1, -7, 4, -4, 11, 7,
					-- layer=2 filter=86 channel=83
					8, -14, -9, 5, 0, -8, 9, 8, -11,
					-- layer=2 filter=86 channel=84
					0, -5, 10, 7, -5, -5, 5, 0, 1,
					-- layer=2 filter=86 channel=85
					9, 1, -8, -4, 7, -7, 0, -3, -9,
					-- layer=2 filter=86 channel=86
					10, -7, 7, -4, -7, 4, 9, -10, -5,
					-- layer=2 filter=86 channel=87
					6, -3, 2, 0, -5, -2, -4, -2, 8,
					-- layer=2 filter=86 channel=88
					2, -9, 7, -10, -12, -10, -6, -11, 5,
					-- layer=2 filter=86 channel=89
					-2, 1, 0, 0, 3, -7, -14, -12, 0,
					-- layer=2 filter=86 channel=90
					-7, 1, 9, -8, -10, 9, 2, -10, -6,
					-- layer=2 filter=86 channel=91
					8, -1, -3, -11, 2, 3, -4, 4, -12,
					-- layer=2 filter=86 channel=92
					1, -5, -12, -2, -4, 0, -3, -3, -13,
					-- layer=2 filter=86 channel=93
					-1, -22, -7, 7, 6, -11, -17, 15, -8,
					-- layer=2 filter=86 channel=94
					-20, -13, 0, -14, -29, -23, -11, -5, -2,
					-- layer=2 filter=86 channel=95
					8, 1, 0, -8, 7, -2, 8, 7, -7,
					-- layer=2 filter=86 channel=96
					-4, 2, 4, -1, -12, -8, -6, -11, -10,
					-- layer=2 filter=86 channel=97
					0, 6, -7, -7, 2, 6, 5, -11, 7,
					-- layer=2 filter=86 channel=98
					1, -23, -11, -6, -8, -25, -19, -11, -10,
					-- layer=2 filter=86 channel=99
					-26, -9, -20, -5, -22, -9, -10, -16, -8,
					-- layer=2 filter=86 channel=100
					13, -10, 6, -11, -10, 7, -4, 0, -2,
					-- layer=2 filter=86 channel=101
					0, -1, -1, 6, -3, 1, -16, -13, -3,
					-- layer=2 filter=86 channel=102
					-7, -1, 4, -4, 4, -5, -18, -3, -7,
					-- layer=2 filter=86 channel=103
					-9, -11, 4, 4, 0, 8, -8, -8, 0,
					-- layer=2 filter=86 channel=104
					-7, -13, 0, 10, 1, -8, 4, -6, 1,
					-- layer=2 filter=86 channel=105
					5, 3, -6, 3, 0, 4, -5, -5, 7,
					-- layer=2 filter=86 channel=106
					-4, 9, -6, -9, 8, 1, 7, 2, -20,
					-- layer=2 filter=86 channel=107
					-2, -2, -4, 1, -3, -14, 3, 5, 11,
					-- layer=2 filter=86 channel=108
					3, -7, 0, -1, 1, -11, -5, -18, -12,
					-- layer=2 filter=86 channel=109
					-9, -8, -8, 11, -1, -6, 7, 2, 3,
					-- layer=2 filter=86 channel=110
					-6, 5, 7, 0, 2, -6, -7, -11, -14,
					-- layer=2 filter=86 channel=111
					0, 7, -5, 6, 0, 0, 3, 10, 8,
					-- layer=2 filter=86 channel=112
					-3, -12, -5, -7, -2, -1, 1, -3, 0,
					-- layer=2 filter=86 channel=113
					4, 1, -9, 1, -13, -10, -12, -4, 1,
					-- layer=2 filter=86 channel=114
					-3, -4, -3, -1, 4, 2, -1, 4, 6,
					-- layer=2 filter=86 channel=115
					-5, 9, 4, -9, -7, 3, 3, -5, 10,
					-- layer=2 filter=86 channel=116
					-13, -2, -3, 0, 0, -4, -10, -18, 9,
					-- layer=2 filter=86 channel=117
					-10, 4, 0, -11, -16, -8, -2, -5, -8,
					-- layer=2 filter=86 channel=118
					3, -2, -2, -7, -6, 0, 0, 0, -12,
					-- layer=2 filter=86 channel=119
					-5, -8, -13, 8, -7, -4, -9, -6, -7,
					-- layer=2 filter=86 channel=120
					-7, -9, 8, -8, -1, 2, 2, 2, 3,
					-- layer=2 filter=86 channel=121
					-3, 3, 1, -8, -7, 7, 5, 4, 10,
					-- layer=2 filter=86 channel=122
					4, -3, 5, 2, 1, 0, -8, -7, 7,
					-- layer=2 filter=86 channel=123
					-8, 7, -8, -8, -5, -15, -19, -23, -23,
					-- layer=2 filter=86 channel=124
					9, 2, -11, -7, -12, -12, -3, -4, 1,
					-- layer=2 filter=86 channel=125
					7, 7, -1, -2, 7, 6, 1, -12, -1,
					-- layer=2 filter=86 channel=126
					8, -7, -7, 0, 5, 3, 6, 7, 9,
					-- layer=2 filter=86 channel=127
					8, 0, 1, -14, -4, -3, -17, -9, -9,
					-- layer=2 filter=87 channel=0
					-15, 2, -19, -3, -10, -13, 0, 6, 16,
					-- layer=2 filter=87 channel=1
					-9, 10, -19, -2, 10, 0, -4, -31, 4,
					-- layer=2 filter=87 channel=2
					4, 0, 3, 0, -5, 2, -1, -7, 9,
					-- layer=2 filter=87 channel=3
					-6, 19, 10, -44, -11, -57, 19, 14, -14,
					-- layer=2 filter=87 channel=4
					15, 11, 37, -33, 20, 16, 29, 11, 29,
					-- layer=2 filter=87 channel=5
					-25, -9, 6, -9, -12, 28, -25, 24, 32,
					-- layer=2 filter=87 channel=6
					-65, -16, -38, -37, 15, 25, -72, -18, -7,
					-- layer=2 filter=87 channel=7
					-14, -20, -52, 25, 0, 0, 63, 33, 27,
					-- layer=2 filter=87 channel=8
					-5, -6, -7, -3, 0, -10, 11, 0, 2,
					-- layer=2 filter=87 channel=9
					22, -2, 3, 0, -2, -34, -31, -18, -21,
					-- layer=2 filter=87 channel=10
					14, 7, 6, 0, 4, -14, 17, 42, 13,
					-- layer=2 filter=87 channel=11
					6, 4, 29, -1, 16, 46, -8, -2, 25,
					-- layer=2 filter=87 channel=12
					-35, 6, -50, -20, -10, -28, -22, -41, 22,
					-- layer=2 filter=87 channel=13
					0, 9, -6, 6, -3, 9, 10, 8, -4,
					-- layer=2 filter=87 channel=14
					10, 4, -1, 10, 0, 10, 15, -34, 5,
					-- layer=2 filter=87 channel=15
					-85, 20, -43, -7, -25, -17, -50, -2, 14,
					-- layer=2 filter=87 channel=16
					-1, 20, -41, -33, -11, -8, -48, -14, -13,
					-- layer=2 filter=87 channel=17
					0, -8, 4, -4, 0, -6, -1, 0, -10,
					-- layer=2 filter=87 channel=18
					8, 3, 34, 37, 54, 52, 4, -12, 35,
					-- layer=2 filter=87 channel=19
					-13, 48, 6, -32, 0, -3, -13, 49, -42,
					-- layer=2 filter=87 channel=20
					0, 4, -5, -10, 2, 4, 1, 2, -11,
					-- layer=2 filter=87 channel=21
					23, 5, 16, 10, 17, -1, -9, -6, -3,
					-- layer=2 filter=87 channel=22
					0, 4, -2, 0, 1, -7, -2, 5, 7,
					-- layer=2 filter=87 channel=23
					-23, 34, 5, -10, 9, 9, 0, 14, 1,
					-- layer=2 filter=87 channel=24
					24, 4, -22, 3, 7, -28, 15, -6, -29,
					-- layer=2 filter=87 channel=25
					8, 15, -4, -12, 5, 22, 14, 4, 10,
					-- layer=2 filter=87 channel=26
					2, -7, 0, 6, -3, 4, 4, -2, 1,
					-- layer=2 filter=87 channel=27
					-12, -6, 18, -27, -20, 14, -7, -20, 26,
					-- layer=2 filter=87 channel=28
					-16, -14, -25, 17, -10, 9, 18, 16, 15,
					-- layer=2 filter=87 channel=29
					0, 5, 1, 8, -3, 10, -9, 11, -2,
					-- layer=2 filter=87 channel=30
					7, 1, 17, -1, -2, 25, 6, -1, 8,
					-- layer=2 filter=87 channel=31
					-19, -7, -65, -72, -89, -12, 24, 25, 6,
					-- layer=2 filter=87 channel=32
					-12, -8, 6, -1, -5, -8, -7, 0, 6,
					-- layer=2 filter=87 channel=33
					-17, 31, 46, -13, -28, -10, -5, -23, 30,
					-- layer=2 filter=87 channel=34
					-47, -18, 67, 29, -20, 11, -29, -20, 3,
					-- layer=2 filter=87 channel=35
					-35, 12, -7, 5, -12, -17, 31, 31, 8,
					-- layer=2 filter=87 channel=36
					1, 0, 0, -8, -3, -4, -11, 2, -7,
					-- layer=2 filter=87 channel=37
					-2, -3, 17, -5, -6, 31, -23, -4, 20,
					-- layer=2 filter=87 channel=38
					-48, -3, 8, -10, -16, 48, -17, -2, 14,
					-- layer=2 filter=87 channel=39
					25, 35, 0, 6, 3, -7, -15, -40, -36,
					-- layer=2 filter=87 channel=40
					-47, -22, -38, 8, -28, -8, -26, -40, 45,
					-- layer=2 filter=87 channel=41
					10, -1, 1, 6, -3, 8, -8, -9, 4,
					-- layer=2 filter=87 channel=42
					19, 44, -10, -18, -18, -42, -31, -2, -25,
					-- layer=2 filter=87 channel=43
					-15, 44, 8, -40, 18, 16, 5, 0, 16,
					-- layer=2 filter=87 channel=44
					-3, -3, -9, -3, -9, -4, 1, 0, -8,
					-- layer=2 filter=87 channel=45
					-34, -41, -18, -36, -30, -17, -12, 13, 1,
					-- layer=2 filter=87 channel=46
					19, 14, -3, 20, -7, 12, 34, 24, 13,
					-- layer=2 filter=87 channel=47
					0, -2, -26, 22, 1, -40, 23, 60, 39,
					-- layer=2 filter=87 channel=48
					2, -2, 6, 6, -7, -4, -6, -11, 10,
					-- layer=2 filter=87 channel=49
					9, -51, -30, 21, 33, 1, -82, -19, -71,
					-- layer=2 filter=87 channel=50
					20, 30, 22, 13, -9, 0, -9, 18, -10,
					-- layer=2 filter=87 channel=51
					-10, 19, 29, -3, 0, 50, -20, 0, -4,
					-- layer=2 filter=87 channel=52
					-84, -37, -29, -27, 21, 37, -7, -30, 9,
					-- layer=2 filter=87 channel=53
					25, -48, -21, 38, 47, -20, 0, 22, -39,
					-- layer=2 filter=87 channel=54
					-51, -48, -51, 5, 21, -1, 33, 36, 48,
					-- layer=2 filter=87 channel=55
					7, -1, 7, 0, -1, 10, -2, -6, 8,
					-- layer=2 filter=87 channel=56
					20, 17, 31, 10, 6, 31, -25, 0, 24,
					-- layer=2 filter=87 channel=57
					-3, 1, -5, 4, -1, -2, -3, 10, -9,
					-- layer=2 filter=87 channel=58
					-64, -20, -54, -31, -49, 5, -21, -44, 28,
					-- layer=2 filter=87 channel=59
					-11, 10, 36, -39, 22, 3, -19, -11, 5,
					-- layer=2 filter=87 channel=60
					-15, 3, -43, 21, -7, 1, 14, -51, -29,
					-- layer=2 filter=87 channel=61
					6, 0, -54, 57, 78, -36, 11, -4, -16,
					-- layer=2 filter=87 channel=62
					-14, 7, 8, 15, 27, 57, -13, -3, -11,
					-- layer=2 filter=87 channel=63
					17, 6, -35, 2, 14, -32, -10, -4, -18,
					-- layer=2 filter=87 channel=64
					7, -5, 2, 0, 24, -21, -15, -12, -6,
					-- layer=2 filter=87 channel=65
					-13, 3, -38, 19, 36, 47, 1, -26, -11,
					-- layer=2 filter=87 channel=66
					-3, 27, -33, -43, -33, -4, 49, -17, 2,
					-- layer=2 filter=87 channel=67
					15, 36, 20, 7, 25, 22, -23, 4, 17,
					-- layer=2 filter=87 channel=68
					1, 11, 6, -9, 4, 3, -6, -4, -5,
					-- layer=2 filter=87 channel=69
					5, 1, -13, 32, 13, -9, 0, -13, -23,
					-- layer=2 filter=87 channel=70
					-53, -48, -7, 0, -28, -14, 12, 25, 19,
					-- layer=2 filter=87 channel=71
					-9, 0, 35, -31, -6, 21, -20, -8, 14,
					-- layer=2 filter=87 channel=72
					13, 35, 20, 8, -56, -25, 31, -3, 11,
					-- layer=2 filter=87 channel=73
					-104, -104, 1, -43, -44, -17, 27, 5, -48,
					-- layer=2 filter=87 channel=74
					5, 21, -1, 16, 3, 13, -10, 13, -18,
					-- layer=2 filter=87 channel=75
					10, 0, -49, 12, -38, 12, -37, -32, 36,
					-- layer=2 filter=87 channel=76
					-29, -49, 15, -63, 2, -38, 18, 0, 25,
					-- layer=2 filter=87 channel=77
					9, 2, 9, 7, 1, 2, 4, 9, -8,
					-- layer=2 filter=87 channel=78
					4, -1, -14, 7, 20, 38, 11, 2, 11,
					-- layer=2 filter=87 channel=79
					2, -1, -8, -12, 5, 4, 0, 7, -10,
					-- layer=2 filter=87 channel=80
					18, 25, 4, -19, 2, 17, 14, 18, -14,
					-- layer=2 filter=87 channel=81
					-3, 18, 0, 6, 1, 1, 5, -10, -1,
					-- layer=2 filter=87 channel=82
					10, -11, 5, -3, -1, 3, -5, 10, 13,
					-- layer=2 filter=87 channel=83
					14, 16, 11, -26, -18, 22, -26, 25, 5,
					-- layer=2 filter=87 channel=84
					0, 11, -3, -11, 7, -5, -11, 10, -10,
					-- layer=2 filter=87 channel=85
					-5, 2, -6, -16, -4, -14, 4, -8, -3,
					-- layer=2 filter=87 channel=86
					15, 0, -15, 9, -5, 3, 10, -4, 0,
					-- layer=2 filter=87 channel=87
					-4, 6, 28, -48, 18, 24, -65, 0, 25,
					-- layer=2 filter=87 channel=88
					8, 33, 11, -15, 18, 7, -28, -23, -13,
					-- layer=2 filter=87 channel=89
					6, 32, -2, 10, 0, 13, 16, -11, 12,
					-- layer=2 filter=87 channel=90
					-2, -3, 4, 0, 11, 0, 1, -2, 4,
					-- layer=2 filter=87 channel=91
					-15, 21, -65, 17, -37, -23, 4, -30, -10,
					-- layer=2 filter=87 channel=92
					-9, 11, -47, -8, -25, -25, 21, -43, 0,
					-- layer=2 filter=87 channel=93
					8, -1, -41, 5, -39, -23, -41, -33, -36,
					-- layer=2 filter=87 channel=94
					48, 19, -29, 35, 62, 19, 36, 57, 19,
					-- layer=2 filter=87 channel=95
					3, 3, 7, -3, 0, -7, -10, 5, 14,
					-- layer=2 filter=87 channel=96
					-1, 19, 28, -42, -12, -5, -18, -34, -15,
					-- layer=2 filter=87 channel=97
					-1, 18, -24, -11, 8, -35, -14, -14, -24,
					-- layer=2 filter=87 channel=98
					-32, -23, -34, 39, 2, -23, 20, 25, 13,
					-- layer=2 filter=87 channel=99
					-45, -22, 1, -13, 13, -35, 1, 8, 4,
					-- layer=2 filter=87 channel=100
					-13, 11, -6, -26, -31, 18, 0, 20, 51,
					-- layer=2 filter=87 channel=101
					13, 18, 22, -58, -2, 21, -26, 6, 28,
					-- layer=2 filter=87 channel=102
					-18, 16, 35, 6, 29, 34, -1, -46, -15,
					-- layer=2 filter=87 channel=103
					32, -5, -3, 2, 1, -9, 27, -20, 38,
					-- layer=2 filter=87 channel=104
					68, 22, -2, 41, 36, 39, 9, 15, -12,
					-- layer=2 filter=87 channel=105
					-22, 28, 9, -51, -15, -27, 14, 7, 96,
					-- layer=2 filter=87 channel=106
					11, 52, 4, -28, -18, 15, -10, 1, -2,
					-- layer=2 filter=87 channel=107
					23, -19, -17, 20, 36, -14, 15, 23, 33,
					-- layer=2 filter=87 channel=108
					18, -40, 0, -38, 1, 0, -18, -57, -19,
					-- layer=2 filter=87 channel=109
					-3, -6, 0, -1, 0, -1, 2, -9, 5,
					-- layer=2 filter=87 channel=110
					-13, 10, -25, -17, 4, -61, 7, -37, -21,
					-- layer=2 filter=87 channel=111
					4, -9, 10, 3, 0, 0, -6, 2, 8,
					-- layer=2 filter=87 channel=112
					10, 6, 4, 15, 1, 4, 8, 18, -12,
					-- layer=2 filter=87 channel=113
					0, -28, -22, 50, -21, -20, 34, 0, -4,
					-- layer=2 filter=87 channel=114
					0, -10, 4, -1, 7, -13, 5, 9, 5,
					-- layer=2 filter=87 channel=115
					6, -2, 6, 7, 0, 4, -6, 1, 2,
					-- layer=2 filter=87 channel=116
					-20, 21, 37, -9, 11, 31, -78, -37, 34,
					-- layer=2 filter=87 channel=117
					-3, -3, -5, 21, -4, 9, 30, -7, -3,
					-- layer=2 filter=87 channel=118
					-24, 8, -8, -35, 9, 5, 1, 6, 21,
					-- layer=2 filter=87 channel=119
					8, 14, 11, 11, 46, 11, 5, 26, 54,
					-- layer=2 filter=87 channel=120
					5, -9, 2, -6, 0, -2, 0, -5, -10,
					-- layer=2 filter=87 channel=121
					2, -1, 2, 3, 0, -9, 8, 7, 1,
					-- layer=2 filter=87 channel=122
					-10, 1, 0, -6, -2, -12, 4, 10, 5,
					-- layer=2 filter=87 channel=123
					-2, 9, 7, -9, 12, -9, 33, 3, -4,
					-- layer=2 filter=87 channel=124
					-12, 53, -14, 7, -18, -27, 56, 42, 80,
					-- layer=2 filter=87 channel=125
					1, -1, 7, -4, -7, 6, 3, -6, 4,
					-- layer=2 filter=87 channel=126
					20, -14, -1, -7, -31, -22, 41, -41, -58,
					-- layer=2 filter=87 channel=127
					-5, -21, 5, -22, -5, -10, 43, 19, 17,
					-- layer=2 filter=88 channel=0
					17, 0, 17, -10, -20, -13, -31, -29, -6,
					-- layer=2 filter=88 channel=1
					-30, -26, -15, 19, -17, -16, 3, 20, 35,
					-- layer=2 filter=88 channel=2
					1, 5, -5, -7, -6, -1, 5, 5, -3,
					-- layer=2 filter=88 channel=3
					9, 46, -2, -29, -26, 39, -9, -34, -30,
					-- layer=2 filter=88 channel=4
					-50, 1, -42, -60, -9, -39, -23, 6, 51,
					-- layer=2 filter=88 channel=5
					27, 14, 21, -29, -27, 11, -50, -57, 15,
					-- layer=2 filter=88 channel=6
					-43, -24, 48, 8, 23, 7, 17, 17, 26,
					-- layer=2 filter=88 channel=7
					64, 17, 19, 31, -28, 41, 15, 56, 0,
					-- layer=2 filter=88 channel=8
					7, -7, -2, -1, -3, -7, 0, -7, 6,
					-- layer=2 filter=88 channel=9
					32, 52, 4, -2, 12, -32, -39, -14, -36,
					-- layer=2 filter=88 channel=10
					15, 13, 9, -27, -39, -5, 12, -39, -12,
					-- layer=2 filter=88 channel=11
					-20, 2, 10, -25, -16, 0, -36, -9, 6,
					-- layer=2 filter=88 channel=12
					-24, -27, 13, 19, 1, -15, 23, 49, 22,
					-- layer=2 filter=88 channel=13
					-2, -6, -4, 0, 8, 8, -4, -4, -4,
					-- layer=2 filter=88 channel=14
					-17, -8, 2, 22, -6, -2, 11, 31, 42,
					-- layer=2 filter=88 channel=15
					12, -2, 50, -38, -9, 65, -42, 26, 69,
					-- layer=2 filter=88 channel=16
					-10, 0, -24, -1, 1, -53, 8, -14, -56,
					-- layer=2 filter=88 channel=17
					-7, -5, -9, 9, -2, -8, -10, -5, -11,
					-- layer=2 filter=88 channel=18
					0, -8, 2, 7, 8, -9, -5, 34, 29,
					-- layer=2 filter=88 channel=19
					15, 10, 20, -4, -6, -17, 14, 47, 19,
					-- layer=2 filter=88 channel=20
					3, 7, 6, -8, 0, 6, 0, 2, 5,
					-- layer=2 filter=88 channel=21
					-20, -2, -1, -6, 13, 8, -1, -3, 14,
					-- layer=2 filter=88 channel=22
					-7, 4, -3, -10, 0, 6, 9, -11, 11,
					-- layer=2 filter=88 channel=23
					-35, -26, -34, -24, -10, -14, 33, 17, 4,
					-- layer=2 filter=88 channel=24
					19, 25, 3, -25, -10, -11, -49, -53, -68,
					-- layer=2 filter=88 channel=25
					-1, 7, 12, -51, -22, -22, -54, -42, -61,
					-- layer=2 filter=88 channel=26
					1, -2, -10, 2, -8, -7, 8, 8, -3,
					-- layer=2 filter=88 channel=27
					33, 35, 10, -19, -5, -13, -74, -68, -59,
					-- layer=2 filter=88 channel=28
					-20, -1, 2, 38, 15, 20, 42, -2, -48,
					-- layer=2 filter=88 channel=29
					0, 8, 4, 7, -3, 0, 4, -2, 9,
					-- layer=2 filter=88 channel=30
					9, 3, 18, -13, -16, 0, -63, -14, 30,
					-- layer=2 filter=88 channel=31
					-68, -40, -40, -57, -55, -41, 2, -17, -52,
					-- layer=2 filter=88 channel=32
					-8, 0, 8, -4, -6, -11, 7, 1, 8,
					-- layer=2 filter=88 channel=33
					27, 36, -5, 13, -43, 23, -5, -15, 27,
					-- layer=2 filter=88 channel=34
					30, -47, -21, -12, 5, -22, -4, 13, -36,
					-- layer=2 filter=88 channel=35
					37, 9, 33, 28, -1, 17, 5, -20, -61,
					-- layer=2 filter=88 channel=36
					-2, 14, -8, -1, -3, 0, 10, -5, 2,
					-- layer=2 filter=88 channel=37
					-19, -17, 11, -14, 8, 8, -46, -18, 14,
					-- layer=2 filter=88 channel=38
					18, 19, 3, -5, -12, 20, -62, -56, 8,
					-- layer=2 filter=88 channel=39
					1, -18, -14, 0, -7, 26, 15, -25, -59,
					-- layer=2 filter=88 channel=40
					30, -56, 65, -11, 24, -31, -42, -4, 19,
					-- layer=2 filter=88 channel=41
					5, 0, -1, 9, 9, -6, 3, -9, -11,
					-- layer=2 filter=88 channel=42
					-15, 3, -18, 16, 18, 0, 19, 36, -67,
					-- layer=2 filter=88 channel=43
					31, 46, 22, -40, 33, 0, -50, -22, 17,
					-- layer=2 filter=88 channel=44
					-8, -5, 9, 1, -4, -7, 5, 4, -6,
					-- layer=2 filter=88 channel=45
					4, -29, -25, -24, -84, -32, -38, -30, -44,
					-- layer=2 filter=88 channel=46
					15, -5, -19, -36, -16, 20, -12, -55, -3,
					-- layer=2 filter=88 channel=47
					-47, -32, -55, -32, -15, -16, 37, 11, -14,
					-- layer=2 filter=88 channel=48
					0, 3, 6, -5, -8, 8, -7, 1, -12,
					-- layer=2 filter=88 channel=49
					-1, -1, -39, 18, 3, 3, -17, 15, 7,
					-- layer=2 filter=88 channel=50
					9, -6, -4, 17, 7, 18, 3, 6, 9,
					-- layer=2 filter=88 channel=51
					-23, -9, 8, -32, -16, 15, -17, -27, 5,
					-- layer=2 filter=88 channel=52
					-35, -42, -4, -37, -10, 38, -38, 18, 28,
					-- layer=2 filter=88 channel=53
					20, 19, 29, 29, 19, 26, -17, 35, 17,
					-- layer=2 filter=88 channel=54
					-48, -47, -33, 3, -8, -19, 19, 23, 8,
					-- layer=2 filter=88 channel=55
					3, 6, -10, -9, -7, 1, 2, 0, 5,
					-- layer=2 filter=88 channel=56
					0, -1, 30, -59, 5, 15, -11, -14, -11,
					-- layer=2 filter=88 channel=57
					-10, 1, 13, 0, -9, 3, -7, -5, -10,
					-- layer=2 filter=88 channel=58
					-11, 5, 20, 57, 8, -27, 8, 7, 24,
					-- layer=2 filter=88 channel=59
					2, -13, -2, 25, -26, 0, -12, -29, -19,
					-- layer=2 filter=88 channel=60
					6, -53, -21, 22, -8, -24, 42, 12, 33,
					-- layer=2 filter=88 channel=61
					14, -55, 28, 20, -17, 12, 34, -8, 33,
					-- layer=2 filter=88 channel=62
					0, -48, -12, 9, 4, 1, 30, 16, 18,
					-- layer=2 filter=88 channel=63
					-26, -53, -47, -23, -10, -7, 9, 3, -12,
					-- layer=2 filter=88 channel=64
					-27, 0, -46, 5, 19, -7, -2, 9, -4,
					-- layer=2 filter=88 channel=65
					0, -31, 45, 7, -3, 16, 41, 17, 45,
					-- layer=2 filter=88 channel=66
					1, 11, 20, -33, -12, -8, -16, 5, -17,
					-- layer=2 filter=88 channel=67
					26, 40, 6, -10, 8, 11, -51, -120, 18,
					-- layer=2 filter=88 channel=68
					5, -3, -5, -1, -8, -7, 3, 5, 3,
					-- layer=2 filter=88 channel=69
					-22, -8, -39, 27, 27, -2, 0, 14, -13,
					-- layer=2 filter=88 channel=70
					9, 6, 8, 41, 9, 0, 5, -44, -43,
					-- layer=2 filter=88 channel=71
					25, 34, 17, -18, -13, -13, -71, -22, -23,
					-- layer=2 filter=88 channel=72
					-38, -4, -1, 12, -4, 12, 41, 34, -15,
					-- layer=2 filter=88 channel=73
					0, -30, -62, 38, -4, 0, -8, 7, -18,
					-- layer=2 filter=88 channel=74
					-29, 2, -3, -13, 0, 21, -62, -65, -14,
					-- layer=2 filter=88 channel=75
					29, 1, 72, 19, 30, -6, 25, 32, 45,
					-- layer=2 filter=88 channel=76
					-62, 28, -39, 39, 23, -21, -44, 24, 43,
					-- layer=2 filter=88 channel=77
					-7, -8, -1, 2, -2, 4, -10, 7, -3,
					-- layer=2 filter=88 channel=78
					-19, -26, 11, -28, -12, 25, -22, 11, 22,
					-- layer=2 filter=88 channel=79
					-8, -2, 7, -8, -1, -2, 0, -7, 8,
					-- layer=2 filter=88 channel=80
					-2, -8, -70, -61, 9, -29, -46, -14, -11,
					-- layer=2 filter=88 channel=81
					3, 19, 17, 7, 10, 16, -1, 13, -1,
					-- layer=2 filter=88 channel=82
					5, -2, -7, 12, 1, -2, -6, -8, -9,
					-- layer=2 filter=88 channel=83
					-5, -28, -4, -11, 1, -3, 11, -10, 1,
					-- layer=2 filter=88 channel=84
					-7, -6, 0, 7, 1, -10, 0, 2, 0,
					-- layer=2 filter=88 channel=85
					20, 4, 0, -4, -4, -2, 3, 1, -2,
					-- layer=2 filter=88 channel=86
					-14, 8, 3, -11, 15, 9, -8, -14, 3,
					-- layer=2 filter=88 channel=87
					-16, -1, -5, -8, 2, -14, -16, -7, 23,
					-- layer=2 filter=88 channel=88
					-17, -30, -3, -8, 16, -1, -33, -24, 12,
					-- layer=2 filter=88 channel=89
					-9, -8, 15, 43, 2, 8, 22, 14, 38,
					-- layer=2 filter=88 channel=90
					-8, -7, 5, 1, 0, 0, -5, -8, -9,
					-- layer=2 filter=88 channel=91
					-12, 31, 30, 43, 0, -10, 13, 11, -36,
					-- layer=2 filter=88 channel=92
					-33, 0, -6, 34, 8, 11, 3, 22, 0,
					-- layer=2 filter=88 channel=93
					9, 9, 26, 7, 21, -8, 19, 31, 41,
					-- layer=2 filter=88 channel=94
					-6, -33, 2, 24, 2, -18, 29, 27, 45,
					-- layer=2 filter=88 channel=95
					5, 5, -2, -3, -6, -10, 0, 17, 0,
					-- layer=2 filter=88 channel=96
					-4, 19, -10, 2, -15, 31, -10, 48, 35,
					-- layer=2 filter=88 channel=97
					37, 55, 2, -21, 8, -38, -35, -52, -25,
					-- layer=2 filter=88 channel=98
					-23, -59, -25, 20, -13, 13, 40, -13, -32,
					-- layer=2 filter=88 channel=99
					-12, -16, 25, -1, -13, -2, 28, 32, 59,
					-- layer=2 filter=88 channel=100
					23, -4, -23, 11, -9, -18, -58, -45, -5,
					-- layer=2 filter=88 channel=101
					9, 41, 39, -15, -22, -27, -90, -24, -32,
					-- layer=2 filter=88 channel=102
					-3, 0, 15, -27, 20, 24, -27, 47, 46,
					-- layer=2 filter=88 channel=103
					-7, 16, -38, 54, 28, 41, 49, 12, 38,
					-- layer=2 filter=88 channel=104
					-16, 0, -11, -15, 22, 20, -33, 0, 27,
					-- layer=2 filter=88 channel=105
					-60, 12, -4, 35, -22, -30, 11, 0, 23,
					-- layer=2 filter=88 channel=106
					0, 64, 26, -1, -7, -23, -39, -53, -63,
					-- layer=2 filter=88 channel=107
					26, 61, -5, -23, 4, 47, 25, 67, 18,
					-- layer=2 filter=88 channel=108
					18, 13, 26, -6, 0, 16, -63, 19, 40,
					-- layer=2 filter=88 channel=109
					-14, 1, -10, 2, -3, -5, -25, -17, 6,
					-- layer=2 filter=88 channel=110
					11, 25, 6, 15, 55, 39, 12, -12, -16,
					-- layer=2 filter=88 channel=111
					-5, -2, -10, 0, 0, 9, 4, 0, 7,
					-- layer=2 filter=88 channel=112
					23, -32, 1, 5, -61, -23, 7, -16, -13,
					-- layer=2 filter=88 channel=113
					0, -2, -20, -6, -1, 19, 3, -1, 5,
					-- layer=2 filter=88 channel=114
					0, 0, -10, -12, -17, -24, 5, -11, -16,
					-- layer=2 filter=88 channel=115
					6, 4, 11, -6, 1, 0, 0, 0, -13,
					-- layer=2 filter=88 channel=116
					2, 18, 22, -9, 19, 25, 7, 34, 25,
					-- layer=2 filter=88 channel=117
					-56, -21, -7, 0, -11, 22, 18, 55, 12,
					-- layer=2 filter=88 channel=118
					-2, 29, 17, -61, 0, -9, -47, -11, -17,
					-- layer=2 filter=88 channel=119
					16, -30, -27, 5, 0, -29, -50, 6, -6,
					-- layer=2 filter=88 channel=120
					0, -2, 8, 1, -2, 9, 1, 0, 1,
					-- layer=2 filter=88 channel=121
					0, 8, 6, -7, -11, 0, 3, -10, -1,
					-- layer=2 filter=88 channel=122
					5, 15, 8, 5, -8, -12, 2, 2, -1,
					-- layer=2 filter=88 channel=123
					-39, -50, -16, -20, -16, -12, 46, 39, 7,
					-- layer=2 filter=88 channel=124
					-5, -2, 13, 8, 2, 7, 11, 36, 56,
					-- layer=2 filter=88 channel=125
					-8, 1, 12, -4, 0, -11, 4, -5, -5,
					-- layer=2 filter=88 channel=126
					32, 28, 13, -23, -36, 18, -20, -39, 27,
					-- layer=2 filter=88 channel=127
					-67, -36, -15, -33, -59, -18, 19, 17, 43,
					-- layer=2 filter=89 channel=0
					-54, -9, -19, 16, 7, 12, 19, 22, 22,
					-- layer=2 filter=89 channel=1
					1, 0, -12, -25, -50, -12, -15, -111, -62,
					-- layer=2 filter=89 channel=2
					-1, 4, -5, 3, -8, 8, 8, -6, 4,
					-- layer=2 filter=89 channel=3
					-32, -7, -34, -19, -3, 13, 29, 62, 51,
					-- layer=2 filter=89 channel=4
					-16, -46, -42, -28, 17, -24, 6, 7, 0,
					-- layer=2 filter=89 channel=5
					-2, -6, -37, -4, -15, -5, -11, 10, 22,
					-- layer=2 filter=89 channel=6
					47, 1, 29, 4, 45, 13, 10, 21, -35,
					-- layer=2 filter=89 channel=7
					5, -17, -9, 58, 7, 57, 35, 29, 34,
					-- layer=2 filter=89 channel=8
					0, 10, 5, -7, 10, 9, -7, -7, 6,
					-- layer=2 filter=89 channel=9
					-15, 10, -37, -60, -1, -47, -5, 8, 2,
					-- layer=2 filter=89 channel=10
					-49, -13, -26, 0, 2, 19, 33, 46, 50,
					-- layer=2 filter=89 channel=11
					-4, -15, -18, -12, 6, 3, 10, 21, 19,
					-- layer=2 filter=89 channel=12
					-6, -27, -16, -33, -65, -63, -15, -58, -36,
					-- layer=2 filter=89 channel=13
					-8, 0, -3, 2, -8, -6, 4, -1, 11,
					-- layer=2 filter=89 channel=14
					-9, -35, -27, -33, -82, -76, -43, -26, -73,
					-- layer=2 filter=89 channel=15
					20, 0, 14, -30, -20, -7, 25, 49, -11,
					-- layer=2 filter=89 channel=16
					-9, 6, 30, -9, 32, 24, -31, -10, -34,
					-- layer=2 filter=89 channel=17
					-9, 6, 8, 6, 0, -9, -8, -4, 1,
					-- layer=2 filter=89 channel=18
					18, -31, 14, -21, -37, -8, -17, -17, 3,
					-- layer=2 filter=89 channel=19
					8, 18, 19, 16, 19, 34, 43, -11, -16,
					-- layer=2 filter=89 channel=20
					-6, 8, 0, 2, 3, 8, 7, 9, -1,
					-- layer=2 filter=89 channel=21
					-14, -10, -10, -5, -21, -2, -6, -5, -22,
					-- layer=2 filter=89 channel=22
					1, 1, 0, -3, -8, 8, 5, -2, 6,
					-- layer=2 filter=89 channel=23
					-22, 0, 12, -32, 33, 8, 65, 43, 16,
					-- layer=2 filter=89 channel=24
					-17, 0, -5, -20, -21, -16, 18, 27, 22,
					-- layer=2 filter=89 channel=25
					-28, -18, -2, -16, -11, -3, 28, 36, 41,
					-- layer=2 filter=89 channel=26
					-3, 5, 0, 6, 9, -9, 0, 1, 5,
					-- layer=2 filter=89 channel=27
					30, 36, 36, -11, -16, 3, -3, -3, 13,
					-- layer=2 filter=89 channel=28
					-24, -52, -28, 28, 4, 34, 60, 41, 28,
					-- layer=2 filter=89 channel=29
					-3, 1, -12, 5, 1, -2, -3, 3, -9,
					-- layer=2 filter=89 channel=30
					10, -26, -15, -82, -33, -58, -17, 0, 28,
					-- layer=2 filter=89 channel=31
					-4, -77, -88, -23, -68, -53, -29, 35, -16,
					-- layer=2 filter=89 channel=32
					-2, -3, 0, 1, 7, 6, -11, 1, 0,
					-- layer=2 filter=89 channel=33
					1, -69, -46, 9, 8, 11, 31, 38, 22,
					-- layer=2 filter=89 channel=34
					0, 47, 7, 28, -19, 40, -33, -12, 6,
					-- layer=2 filter=89 channel=35
					-5, -7, -11, 39, 16, 37, 59, 42, 50,
					-- layer=2 filter=89 channel=36
					1, 2, 1, 0, 9, -2, 15, -5, -11,
					-- layer=2 filter=89 channel=37
					15, -9, 8, -7, -13, 6, 17, 5, 0,
					-- layer=2 filter=89 channel=38
					23, 21, -4, -47, -7, -47, -30, -12, 9,
					-- layer=2 filter=89 channel=39
					-22, 1, -15, 5, -10, -34, -3, 2, 10,
					-- layer=2 filter=89 channel=40
					-2, 9, 10, 38, -66, -21, 55, 9, -12,
					-- layer=2 filter=89 channel=41
					0, 2, 9, 10, 4, 1, 3, -8, -6,
					-- layer=2 filter=89 channel=42
					9, 28, 15, -27, -21, -25, 33, 52, 21,
					-- layer=2 filter=89 channel=43
					-5, 1, -51, -1, 13, -14, 44, 39, 39,
					-- layer=2 filter=89 channel=44
					6, -11, 12, -7, -3, -8, 1, -3, -2,
					-- layer=2 filter=89 channel=45
					48, 20, 25, 0, 36, 67, 34, 17, 0,
					-- layer=2 filter=89 channel=46
					-15, -2, -41, -10, 21, 1, 1, 4, 7,
					-- layer=2 filter=89 channel=47
					-47, -54, -36, 46, 17, 57, 51, 40, 11,
					-- layer=2 filter=89 channel=48
					5, 9, -9, 5, -1, -2, 3, -5, -11,
					-- layer=2 filter=89 channel=49
					11, 8, 16, 38, -11, -1, -66, -35, -10,
					-- layer=2 filter=89 channel=50
					9, 7, -8, 3, 8, 29, -21, -6, -8,
					-- layer=2 filter=89 channel=51
					-14, -4, -15, -2, -4, 8, 14, 24, 10,
					-- layer=2 filter=89 channel=52
					5, -8, -3, -3, 11, 10, 23, -19, 31,
					-- layer=2 filter=89 channel=53
					-36, 0, -28, -52, -21, -28, -17, -29, 3,
					-- layer=2 filter=89 channel=54
					-13, -17, -30, 10, 8, 21, 40, 10, 40,
					-- layer=2 filter=89 channel=55
					13, -6, 1, 6, -5, 4, -7, 7, 2,
					-- layer=2 filter=89 channel=56
					-13, -23, -12, -5, -13, -11, 11, 29, 15,
					-- layer=2 filter=89 channel=57
					0, 1, -1, 0, -7, 10, 2, 3, -1,
					-- layer=2 filter=89 channel=58
					-15, -37, -27, -33, -65, -73, -6, -52, 3,
					-- layer=2 filter=89 channel=59
					3, 18, 20, 11, -30, -2, 9, -78, -30,
					-- layer=2 filter=89 channel=60
					17, -7, -11, -15, -15, -5, -56, -88, -33,
					-- layer=2 filter=89 channel=61
					3, -17, 38, 5, 4, 12, 10, -28, 3,
					-- layer=2 filter=89 channel=62
					6, -16, -6, -19, 10, 10, -33, -8, -25,
					-- layer=2 filter=89 channel=63
					-9, -17, -28, -38, -41, -4, 26, 23, 11,
					-- layer=2 filter=89 channel=64
					-21, 4, 5, -1, 20, 2, 49, 60, 35,
					-- layer=2 filter=89 channel=65
					34, -12, 4, -21, 36, 7, 17, -3, -38,
					-- layer=2 filter=89 channel=66
					27, 21, -17, -18, -26, 32, 11, -26, -16,
					-- layer=2 filter=89 channel=67
					-56, 5, -68, -102, -4, -37, -45, 0, -23,
					-- layer=2 filter=89 channel=68
					2, -7, 0, 8, 6, 0, -8, 0, -9,
					-- layer=2 filter=89 channel=69
					14, -5, 20, -11, -7, -2, 12, 13, 30,
					-- layer=2 filter=89 channel=70
					-20, -26, -17, 27, 11, 15, 50, 16, 32,
					-- layer=2 filter=89 channel=71
					-13, 19, -17, -16, 3, -4, 29, 28, 28,
					-- layer=2 filter=89 channel=72
					0, -18, -48, -21, -60, -52, 13, 1, -33,
					-- layer=2 filter=89 channel=73
					30, 43, 18, 3, 6, 20, -1, -1, 9,
					-- layer=2 filter=89 channel=74
					-40, -62, -83, -85, -5, -11, 13, 29, 9,
					-- layer=2 filter=89 channel=75
					-59, -26, -29, 8, 31, -27, -50, -41, -89,
					-- layer=2 filter=89 channel=76
					18, -23, -15, -24, 11, 14, -14, -29, 12,
					-- layer=2 filter=89 channel=77
					-4, 0, -3, 0, -9, -11, 8, -6, 6,
					-- layer=2 filter=89 channel=78
					23, 0, 4, 11, 23, 7, 13, 20, 7,
					-- layer=2 filter=89 channel=79
					8, 2, 2, 9, 3, 8, -3, 2, 8,
					-- layer=2 filter=89 channel=80
					-44, -32, -41, -19, -21, -17, -7, 20, 11,
					-- layer=2 filter=89 channel=81
					-16, -13, -6, -20, 2, -23, -7, 4, -7,
					-- layer=2 filter=89 channel=82
					-5, 1, 4, -1, 3, 10, 4, -4, 3,
					-- layer=2 filter=89 channel=83
					-9, 13, 4, -44, -25, -14, 15, 18, 13,
					-- layer=2 filter=89 channel=84
					1, -6, 2, -7, -9, -8, 1, -2, 7,
					-- layer=2 filter=89 channel=85
					7, 13, -7, 4, -13, 3, -11, -12, 4,
					-- layer=2 filter=89 channel=86
					5, -1, 14, 4, 10, -1, 9, -22, -13,
					-- layer=2 filter=89 channel=87
					14, -9, -13, -2, 11, -21, -27, -25, -8,
					-- layer=2 filter=89 channel=88
					29, -25, -27, -85, -2, -86, 5, -6, 24,
					-- layer=2 filter=89 channel=89
					-4, -17, 0, -9, -40, -39, -63, -63, -102,
					-- layer=2 filter=89 channel=90
					3, -2, -6, 7, 4, -7, 5, -1, 10,
					-- layer=2 filter=89 channel=91
					16, -7, -13, -12, -52, -48, -12, -61, -112,
					-- layer=2 filter=89 channel=92
					15, 16, -3, -12, -39, -28, -5, -85, -52,
					-- layer=2 filter=89 channel=93
					31, -7, -7, 43, 35, 18, 49, -31, 4,
					-- layer=2 filter=89 channel=94
					-1, -7, 25, 11, 3, -14, 11, -72, -27,
					-- layer=2 filter=89 channel=95
					14, 17, 4, 6, 3, 6, 12, 7, -2,
					-- layer=2 filter=89 channel=96
					20, 24, 27, 20, 42, 16, 21, 7, 1,
					-- layer=2 filter=89 channel=97
					-19, -4, -23, -43, -8, -16, -11, 23, 19,
					-- layer=2 filter=89 channel=98
					-18, -15, 9, 37, 35, 40, 74, 54, 34,
					-- layer=2 filter=89 channel=99
					-6, 26, 0, 0, 22, 42, -14, 10, -4,
					-- layer=2 filter=89 channel=100
					13, 9, -10, -51, -22, -61, -9, -27, 12,
					-- layer=2 filter=89 channel=101
					-23, -14, -32, -7, -1, 8, 10, 22, -4,
					-- layer=2 filter=89 channel=102
					15, 15, 14, 4, 45, 10, 46, 28, -17,
					-- layer=2 filter=89 channel=103
					-6, 25, 33, -32, 26, 18, 37, 8, -17,
					-- layer=2 filter=89 channel=104
					5, 13, 5, 0, 7, -22, -19, -15, 15,
					-- layer=2 filter=89 channel=105
					-7, -58, -24, -27, 0, -9, 21, -7, -40,
					-- layer=2 filter=89 channel=106
					-39, -37, -34, -49, -45, -8, -8, 16, 0,
					-- layer=2 filter=89 channel=107
					-22, 41, 55, -21, -25, 40, 24, -45, 29,
					-- layer=2 filter=89 channel=108
					17, 44, 34, -23, -9, -23, -39, -44, -36,
					-- layer=2 filter=89 channel=109
					0, -5, -3, 0, -4, 12, 18, 0, 7,
					-- layer=2 filter=89 channel=110
					1, -6, 27, 3, -5, -1, 26, 23, 17,
					-- layer=2 filter=89 channel=111
					-5, -6, 5, 8, 5, -6, 4, 1, -7,
					-- layer=2 filter=89 channel=112
					-28, -9, 3, -11, 5, 24, 27, 4, 31,
					-- layer=2 filter=89 channel=113
					6, -12, -19, -51, -53, -36, 29, 6, 7,
					-- layer=2 filter=89 channel=114
					12, 12, 0, 9, 4, 0, 9, -1, 10,
					-- layer=2 filter=89 channel=115
					4, 9, -7, -4, -4, 0, -3, 4, -6,
					-- layer=2 filter=89 channel=116
					3, 35, -12, -35, 6, 0, -5, -36, -4,
					-- layer=2 filter=89 channel=117
					-29, -14, -4, 4, -1, 6, 16, -43, 0,
					-- layer=2 filter=89 channel=118
					31, 31, -12, 13, 38, 27, 22, 46, 17,
					-- layer=2 filter=89 channel=119
					2, -67, -61, -11, -36, -38, 9, -7, 10,
					-- layer=2 filter=89 channel=120
					0, -9, -1, -2, -5, -6, -9, -7, -10,
					-- layer=2 filter=89 channel=121
					10, 1, -4, 11, 9, 8, 7, 0, 10,
					-- layer=2 filter=89 channel=122
					-9, -7, 15, -2, 10, -10, -15, -1, 15,
					-- layer=2 filter=89 channel=123
					18, -24, -24, 37, 13, 51, 33, 51, -13,
					-- layer=2 filter=89 channel=124
					23, 22, 21, -6, 8, 9, 40, 31, -52,
					-- layer=2 filter=89 channel=125
					-7, 7, 0, 6, 4, 2, 5, 2, 9,
					-- layer=2 filter=89 channel=126
					3, -1, 8, -25, 18, 24, -69, -49, -32,
					-- layer=2 filter=89 channel=127
					31, -5, -11, -66, -38, -87, 6, -14, -25,
					-- layer=2 filter=90 channel=0
					-14, -16, -27, -1, -11, -13, 24, -8, -30,
					-- layer=2 filter=90 channel=1
					-48, -21, 5, -7, 8, -15, -5, 14, -8,
					-- layer=2 filter=90 channel=2
					0, -5, 4, 3, 8, -8, -7, -1, 6,
					-- layer=2 filter=90 channel=3
					38, 4, 29, 2, -4, -7, 11, -15, -4,
					-- layer=2 filter=90 channel=4
					9, -14, -42, -8, -31, -22, -39, -16, -28,
					-- layer=2 filter=90 channel=5
					-5, -21, 1, -2, -32, -26, 23, -1, -7,
					-- layer=2 filter=90 channel=6
					13, -75, -58, 9, 10, -46, 20, 6, -18,
					-- layer=2 filter=90 channel=7
					-20, 10, -14, -17, -10, 10, -6, -29, -16,
					-- layer=2 filter=90 channel=8
					-9, 2, 4, 2, -10, -5, 9, 9, -10,
					-- layer=2 filter=90 channel=9
					16, 10, -24, 7, -4, -44, 2, -21, -19,
					-- layer=2 filter=90 channel=10
					22, -4, -8, 12, 4, 5, 31, -3, -19,
					-- layer=2 filter=90 channel=11
					8, -14, -13, -3, -10, 2, -6, -7, 10,
					-- layer=2 filter=90 channel=12
					-33, 12, 1, 11, 18, -23, -34, -23, -33,
					-- layer=2 filter=90 channel=13
					9, 0, -8, -5, 6, 2, 4, 0, -1,
					-- layer=2 filter=90 channel=14
					-56, -26, -13, -11, 11, -30, -13, -23, -22,
					-- layer=2 filter=90 channel=15
					-18, 11, -5, -11, 22, -16, -6, -30, 33,
					-- layer=2 filter=90 channel=16
					-5, -15, -5, -19, 1, -3, -16, 14, 16,
					-- layer=2 filter=90 channel=17
					-3, 4, -6, -3, -10, -2, 7, -4, 4,
					-- layer=2 filter=90 channel=18
					7, -12, -40, 28, 17, -44, -46, 4, 20,
					-- layer=2 filter=90 channel=19
					-4, 0, 12, -29, -8, 28, 8, 2, 6,
					-- layer=2 filter=90 channel=20
					8, -1, -8, -4, 4, -8, 4, -4, 8,
					-- layer=2 filter=90 channel=21
					8, 3, 5, -14, -7, 4, -14, -14, -8,
					-- layer=2 filter=90 channel=22
					-7, 5, 0, 2, 8, -9, -9, -6, 4,
					-- layer=2 filter=90 channel=23
					25, 28, 18, 12, 0, -1, -5, 10, 8,
					-- layer=2 filter=90 channel=24
					16, 2, -4, 10, 32, 15, -3, 12, 10,
					-- layer=2 filter=90 channel=25
					41, 12, 8, -5, 32, 42, -14, 8, 30,
					-- layer=2 filter=90 channel=26
					1, 1, 3, 4, -6, 0, 5, 2, -7,
					-- layer=2 filter=90 channel=27
					7, -24, 3, 1, -19, -8, 28, -2, -32,
					-- layer=2 filter=90 channel=28
					-4, -59, -46, -6, -4, -6, -39, -44, -45,
					-- layer=2 filter=90 channel=29
					4, -7, 6, 0, -3, -9, -2, 4, -7,
					-- layer=2 filter=90 channel=30
					-7, 28, 3, 12, 6, -32, -23, -23, -7,
					-- layer=2 filter=90 channel=31
					-65, 64, 53, -87, 30, 27, -51, 28, 33,
					-- layer=2 filter=90 channel=32
					-2, 0, -10, 11, 0, 5, 5, 3, 5,
					-- layer=2 filter=90 channel=33
					-37, -31, -12, -7, 20, -27, 0, -34, -38,
					-- layer=2 filter=90 channel=34
					-11, -18, -45, -13, -87, -7, -20, -45, -38,
					-- layer=2 filter=90 channel=35
					18, -1, -6, -10, -44, 22, -14, -8, -3,
					-- layer=2 filter=90 channel=36
					-10, 5, -8, 2, -7, -6, 10, 8, -8,
					-- layer=2 filter=90 channel=37
					-6, -30, -7, -13, -31, -9, 18, -1, 1,
					-- layer=2 filter=90 channel=38
					3, 4, 37, 24, 10, 9, 54, 37, -8,
					-- layer=2 filter=90 channel=39
					33, 18, -4, 22, 33, -11, 9, 10, 28,
					-- layer=2 filter=90 channel=40
					-9, -38, -9, -5, 2, -34, -15, -35, -9,
					-- layer=2 filter=90 channel=41
					-4, -10, -7, -2, 0, -8, 1, 9, 2,
					-- layer=2 filter=90 channel=42
					20, 16, -4, 3, -25, -2, -20, 18, 34,
					-- layer=2 filter=90 channel=43
					36, 21, 6, -4, -8, -4, 1, 30, -18,
					-- layer=2 filter=90 channel=44
					-5, -4, -2, 5, 8, 2, 4, 0, 2,
					-- layer=2 filter=90 channel=45
					-40, -2, 17, -35, -44, -13, 19, 41, 11,
					-- layer=2 filter=90 channel=46
					5, 7, -3, 13, -20, -28, -13, -28, -48,
					-- layer=2 filter=90 channel=47
					1, -43, -41, -29, 3, 0, 26, 0, -39,
					-- layer=2 filter=90 channel=48
					0, 4, 6, -6, -1, -9, 0, -5, 10,
					-- layer=2 filter=90 channel=49
					11, -15, -17, 25, 30, -10, -18, 26, 29,
					-- layer=2 filter=90 channel=50
					0, -6, -1, 22, 24, 13, 10, -5, -4,
					-- layer=2 filter=90 channel=51
					-17, -13, 0, -11, -2, -19, -2, -12, -4,
					-- layer=2 filter=90 channel=52
					-6, 21, -42, -9, -37, -14, -49, 0, 33,
					-- layer=2 filter=90 channel=53
					18, -32, 47, -29, 1, -10, -48, 6, 29,
					-- layer=2 filter=90 channel=54
					-2, -4, 4, -4, -16, 10, -36, -2, -18,
					-- layer=2 filter=90 channel=55
					-2, -4, -4, -10, -2, 6, 0, 2, 2,
					-- layer=2 filter=90 channel=56
					8, -34, -9, -10, -28, -10, 0, 7, -26,
					-- layer=2 filter=90 channel=57
					8, -2, 3, 8, -6, -1, 8, 9, 10,
					-- layer=2 filter=90 channel=58
					-46, -11, 18, 14, -3, -16, -37, 10, -41,
					-- layer=2 filter=90 channel=59
					-34, 16, 51, 12, 33, 6, 25, 51, -4,
					-- layer=2 filter=90 channel=60
					13, 51, 20, 45, 25, 36, 42, 21, 55,
					-- layer=2 filter=90 channel=61
					32, 26, 54, 29, 53, 43, 48, 34, 47,
					-- layer=2 filter=90 channel=62
					-4, -44, -72, -49, -17, -26, -31, 28, -2,
					-- layer=2 filter=90 channel=63
					37, 35, -5, 21, 37, -14, 20, -6, -18,
					-- layer=2 filter=90 channel=64
					3, 8, -17, 20, -4, -7, -17, -12, 9,
					-- layer=2 filter=90 channel=65
					7, 9, -11, 42, 29, 8, 25, 35, 12,
					-- layer=2 filter=90 channel=66
					25, -22, 66, 21, -9, 51, -16, 0, 32,
					-- layer=2 filter=90 channel=67
					2, 2, 15, -6, 15, 17, 16, 2, 8,
					-- layer=2 filter=90 channel=68
					-5, 4, -5, 4, -10, -3, 1, 9, -1,
					-- layer=2 filter=90 channel=69
					11, -26, -25, 17, -6, -1, 0, 3, 9,
					-- layer=2 filter=90 channel=70
					11, -25, -10, -7, -64, -1, -13, -48, -43,
					-- layer=2 filter=90 channel=71
					19, -19, 3, -3, -15, 2, -1, 11, -26,
					-- layer=2 filter=90 channel=72
					-43, 14, -11, -17, 10, -24, -21, -17, -48,
					-- layer=2 filter=90 channel=73
					48, 53, 110, -18, 19, 53, 22, 37, 79,
					-- layer=2 filter=90 channel=74
					14, 23, 4, 10, 25, -2, 21, 0, -19,
					-- layer=2 filter=90 channel=75
					3, -22, -29, 22, -32, 66, 13, 22, -1,
					-- layer=2 filter=90 channel=76
					21, -19, 60, -59, 49, -1, -30, -27, 20,
					-- layer=2 filter=90 channel=77
					-3, -8, 3, 7, 0, -11, -9, -4, -10,
					-- layer=2 filter=90 channel=78
					22, 10, -27, -4, -5, 10, -12, 24, 18,
					-- layer=2 filter=90 channel=79
					10, 6, 9, 5, -9, 3, 0, -1, -5,
					-- layer=2 filter=90 channel=80
					30, -21, -24, 5, -30, -28, -16, -5, 0,
					-- layer=2 filter=90 channel=81
					-5, 6, 6, -6, 4, 11, -1, -1, -4,
					-- layer=2 filter=90 channel=82
					3, 2, -9, 0, 6, -2, -9, -5, -11,
					-- layer=2 filter=90 channel=83
					20, 1, -4, 4, -11, -36, -10, -48, -6,
					-- layer=2 filter=90 channel=84
					-1, -11, -4, 10, 3, 2, 5, -9, -2,
					-- layer=2 filter=90 channel=85
					0, -5, -6, -7, 11, -13, -10, -6, -16,
					-- layer=2 filter=90 channel=86
					19, 21, -11, 4, 4, 10, -4, 0, 0,
					-- layer=2 filter=90 channel=87
					-11, -36, -21, -52, -44, -53, -65, -79, -32,
					-- layer=2 filter=90 channel=88
					-24, 27, -3, 28, 37, -30, 40, 12, 0,
					-- layer=2 filter=90 channel=89
					-64, -12, -3, -29, 0, 0, -28, -19, -30,
					-- layer=2 filter=90 channel=90
					-5, 7, -2, 0, 7, 8, -3, -3, -2,
					-- layer=2 filter=90 channel=91
					-20, 19, -13, -13, 0, 1, -8, -1, -8,
					-- layer=2 filter=90 channel=92
					-35, -5, -1, 25, 44, 3, -22, -11, 1,
					-- layer=2 filter=90 channel=93
					-16, -46, -45, -37, 24, 18, -31, 12, 46,
					-- layer=2 filter=90 channel=94
					16, -7, 14, 12, 28, 33, 39, 30, 16,
					-- layer=2 filter=90 channel=95
					-21, -12, -4, -7, -6, -17, -8, -4, -21,
					-- layer=2 filter=90 channel=96
					-25, -61, -18, -5, -8, -26, -29, -20, -41,
					-- layer=2 filter=90 channel=97
					39, 4, -33, -3, 17, -1, -11, -28, -16,
					-- layer=2 filter=90 channel=98
					21, -13, -52, -1, 0, 1, 4, -33, -57,
					-- layer=2 filter=90 channel=99
					38, 0, 2, 0, 0, 38, 18, 33, 48,
					-- layer=2 filter=90 channel=100
					29, 57, 33, 21, 14, -10, -1, -2, -44,
					-- layer=2 filter=90 channel=101
					30, 6, 17, -3, 2, 21, -50, -11, 7,
					-- layer=2 filter=90 channel=102
					-8, -85, -90, 15, -15, -73, -55, -33, -32,
					-- layer=2 filter=90 channel=103
					-60, -17, -24, -23, -5, -4, -22, 43, 28,
					-- layer=2 filter=90 channel=104
					-13, -29, -8, 9, -8, -23, -26, 12, -7,
					-- layer=2 filter=90 channel=105
					-56, -2, -20, -18, 5, -15, -14, -63, -1,
					-- layer=2 filter=90 channel=106
					-17, -9, -9, -1, -2, 15, -34, -6, -3,
					-- layer=2 filter=90 channel=107
					16, 28, -14, 37, 11, 3, -15, 10, 33,
					-- layer=2 filter=90 channel=108
					-16, -34, -24, 8, -8, -29, 22, 4, -1,
					-- layer=2 filter=90 channel=109
					0, 23, 23, 4, 8, 10, -23, 20, -3,
					-- layer=2 filter=90 channel=110
					13, 24, 18, 16, 56, 26, -14, 16, 34,
					-- layer=2 filter=90 channel=111
					-10, -6, -3, 3, 0, -8, -3, -2, -7,
					-- layer=2 filter=90 channel=112
					-5, 0, 10, -10, -3, 7, 24, 26, 15,
					-- layer=2 filter=90 channel=113
					-11, 23, 20, 28, 9, 14, -12, 6, -4,
					-- layer=2 filter=90 channel=114
					7, -6, -2, 3, 0, -5, 1, -8, 4,
					-- layer=2 filter=90 channel=115
					-9, 2, 9, -7, 6, 6, 7, -5, -2,
					-- layer=2 filter=90 channel=116
					4, -81, -23, -33, -23, -61, -58, -51, -34,
					-- layer=2 filter=90 channel=117
					-9, 39, 22, -16, -7, 57, -10, -14, 20,
					-- layer=2 filter=90 channel=118
					41, 1, -23, 0, -16, -31, 15, 0, -25,
					-- layer=2 filter=90 channel=119
					0, -40, -28, -4, 0, -8, -44, 4, 0,
					-- layer=2 filter=90 channel=120
					-4, -5, -8, 6, 0, -5, -9, 6, 4,
					-- layer=2 filter=90 channel=121
					0, 6, 2, 10, -3, -5, -3, 12, 2,
					-- layer=2 filter=90 channel=122
					-8, 0, 4, 0, 4, 0, 1, -4, -10,
					-- layer=2 filter=90 channel=123
					-13, 16, -9, -39, 46, 11, -28, -13, -38,
					-- layer=2 filter=90 channel=124
					-85, -29, 18, -100, 20, 35, -71, -29, 30,
					-- layer=2 filter=90 channel=125
					-10, -8, -3, 4, 11, -8, -2, -1, 10,
					-- layer=2 filter=90 channel=126
					-33, 21, 86, -10, 18, 13, 2, 23, 43,
					-- layer=2 filter=90 channel=127
					0, 17, 1, 25, 1, -40, 20, 7, -20,
					-- layer=2 filter=91 channel=0
					-20, 17, -10, -26, 13, 19, 0, 4, -8,
					-- layer=2 filter=91 channel=1
					-20, -32, -17, 14, 18, 0, -26, -2, 15,
					-- layer=2 filter=91 channel=2
					11, 10, 10, 4, -5, -6, 2, 7, 10,
					-- layer=2 filter=91 channel=3
					2, 21, 21, 6, -2, 23, 42, 23, 24,
					-- layer=2 filter=91 channel=4
					31, 67, -37, -21, -47, -46, -13, -32, -14,
					-- layer=2 filter=91 channel=5
					11, 3, 11, -8, -3, 5, 11, 4, 22,
					-- layer=2 filter=91 channel=6
					-10, -12, -23, 40, 24, -32, 3, 10, -45,
					-- layer=2 filter=91 channel=7
					28, 24, 31, 8, 32, 86, 8, 45, 21,
					-- layer=2 filter=91 channel=8
					4, -10, -6, -3, -3, 2, -7, -7, -2,
					-- layer=2 filter=91 channel=9
					-16, -3, -13, 12, -1, 28, 3, -2, 17,
					-- layer=2 filter=91 channel=10
					10, 27, 3, -20, 3, 15, 13, -3, -8,
					-- layer=2 filter=91 channel=11
					-17, -6, 13, 11, 12, 2, 2, 17, 25,
					-- layer=2 filter=91 channel=12
					4, 28, 20, 36, 18, 27, 1, 25, 34,
					-- layer=2 filter=91 channel=13
					8, 4, 4, -3, 7, 1, 2, -4, 0,
					-- layer=2 filter=91 channel=14
					-6, -3, 8, 13, -18, 2, -32, -12, 33,
					-- layer=2 filter=91 channel=15
					-14, 0, -61, 36, 22, -16, -31, 65, 34,
					-- layer=2 filter=91 channel=16
					20, 41, 24, -26, -25, -34, -25, -21, -114,
					-- layer=2 filter=91 channel=17
					-2, 11, 7, 0, -3, 1, 4, -1, -8,
					-- layer=2 filter=91 channel=18
					-17, 19, -65, 21, -10, -23, 1, -11, -21,
					-- layer=2 filter=91 channel=19
					-3, -53, -34, 19, 11, 0, 22, 2, -5,
					-- layer=2 filter=91 channel=20
					10, 2, 7, -4, 0, 5, -4, 7, 2,
					-- layer=2 filter=91 channel=21
					1, 18, -7, -24, -14, -20, -10, -12, -14,
					-- layer=2 filter=91 channel=22
					8, -1, 3, 3, -7, -1, 0, -5, -3,
					-- layer=2 filter=91 channel=23
					19, 60, 23, 2, 34, -7, 24, 1, -34,
					-- layer=2 filter=91 channel=24
					-8, 5, 0, -6, -3, 0, -15, -6, -25,
					-- layer=2 filter=91 channel=25
					-41, -2, 16, -19, -5, 19, -6, -19, -1,
					-- layer=2 filter=91 channel=26
					-4, 7, 3, -3, -2, 1, 0, -3, -7,
					-- layer=2 filter=91 channel=27
					-25, -24, -7, -11, 27, 42, -5, 2, 12,
					-- layer=2 filter=91 channel=28
					-66, -12, -27, -16, 0, 66, 13, 24, 37,
					-- layer=2 filter=91 channel=29
					7, 1, 8, -3, 11, 0, 4, 7, -1,
					-- layer=2 filter=91 channel=30
					8, 5, 5, -49, -15, -26, -5, -32, -10,
					-- layer=2 filter=91 channel=31
					-32, -75, -10, -54, 6, -11, 28, 0, 11,
					-- layer=2 filter=91 channel=32
					-5, -3, -8, -6, -2, -10, 3, -1, 5,
					-- layer=2 filter=91 channel=33
					28, 11, -8, 37, -9, 46, -52, -48, 50,
					-- layer=2 filter=91 channel=34
					60, 8, -25, 0, -16, -18, -20, 17, -48,
					-- layer=2 filter=91 channel=35
					-57, -40, -42, 11, -14, 29, 24, 22, 6,
					-- layer=2 filter=91 channel=36
					6, 7, 1, -9, 5, 6, 2, 8, -10,
					-- layer=2 filter=91 channel=37
					-6, -23, 3, 5, 31, 5, 11, 2, 32,
					-- layer=2 filter=91 channel=38
					-7, -12, -17, -3, -9, -2, -33, -4, 19,
					-- layer=2 filter=91 channel=39
					37, 30, 37, 25, 0, -57, -27, -1, -81,
					-- layer=2 filter=91 channel=40
					54, 30, 1, -25, 15, 5, 5, 25, 3,
					-- layer=2 filter=91 channel=41
					-6, -3, 11, -1, 3, 5, -1, -2, 0,
					-- layer=2 filter=91 channel=42
					3, 60, 17, -5, 12, -24, -17, 0, -22,
					-- layer=2 filter=91 channel=43
					-16, 30, -9, -31, 15, 3, 27, 0, 16,
					-- layer=2 filter=91 channel=44
					8, 9, -7, 3, -7, 2, 7, 3, -8,
					-- layer=2 filter=91 channel=45
					31, 10, -1, -70, -56, 1, -35, -16, -17,
					-- layer=2 filter=91 channel=46
					1, -24, 0, -46, -21, -7, 30, -2, 2,
					-- layer=2 filter=91 channel=47
					17, 70, 1, -20, 16, 78, 28, 26, 17,
					-- layer=2 filter=91 channel=48
					-5, 7, -9, -8, 0, -4, -1, -8, 1,
					-- layer=2 filter=91 channel=49
					-25, -15, -66, 2, -20, -17, 24, -7, -49,
					-- layer=2 filter=91 channel=50
					-5, -1, -16, -6, 27, 9, -21, -30, -3,
					-- layer=2 filter=91 channel=51
					-3, 8, 21, -7, 2, 23, 0, 12, 24,
					-- layer=2 filter=91 channel=52
					-3, -34, -1, 10, 45, -32, 21, 22, 48,
					-- layer=2 filter=91 channel=53
					-5, -18, -11, 3, 19, -3, 35, -32, 43,
					-- layer=2 filter=91 channel=54
					7, 25, -13, 39, -4, -8, 15, 37, -5,
					-- layer=2 filter=91 channel=55
					-4, 4, -10, -11, 0, -8, -4, -10, -4,
					-- layer=2 filter=91 channel=56
					-40, -6, 11, 13, 14, 8, 0, 15, 23,
					-- layer=2 filter=91 channel=57
					-1, -14, -6, 7, 4, -2, 9, -3, 2,
					-- layer=2 filter=91 channel=58
					-4, 11, 23, 24, 34, 11, -12, 19, 48,
					-- layer=2 filter=91 channel=59
					10, -62, -37, 31, 36, -19, -20, -19, -25,
					-- layer=2 filter=91 channel=60
					14, -40, -2, 17, -10, -26, 10, 5, -8,
					-- layer=2 filter=91 channel=61
					-39, -43, -15, -29, -12, -20, 7, 3, -49,
					-- layer=2 filter=91 channel=62
					1, -20, -50, 39, 3, -33, 10, -10, -46,
					-- layer=2 filter=91 channel=63
					39, 37, 12, -41, -10, 0, -43, -14, -21,
					-- layer=2 filter=91 channel=64
					9, 44, -5, -12, -22, -9, -76, -30, -24,
					-- layer=2 filter=91 channel=65
					-33, -59, 2, 0, -14, 13, 0, -19, -54,
					-- layer=2 filter=91 channel=66
					-6, -36, -22, 3, -16, -18, 15, -7, -15,
					-- layer=2 filter=91 channel=67
					-26, -10, -32, -93, 4, -21, -43, -28, -9,
					-- layer=2 filter=91 channel=68
					9, -7, 11, -2, 0, -3, 3, -9, -6,
					-- layer=2 filter=91 channel=69
					7, 28, 14, -9, 0, 0, -75, 0, -38,
					-- layer=2 filter=91 channel=70
					-26, -12, -24, -20, -14, 15, 18, 5, 32,
					-- layer=2 filter=91 channel=71
					-25, -6, -30, -27, 8, 50, -18, -42, -1,
					-- layer=2 filter=91 channel=72
					4, -7, -26, 29, 22, 57, -19, -12, 4,
					-- layer=2 filter=91 channel=73
					-36, -42, -35, 22, 21, -95, 11, 54, 41,
					-- layer=2 filter=91 channel=74
					16, 4, 0, -39, -23, -18, 0, -16, -28,
					-- layer=2 filter=91 channel=75
					12, -11, -25, -19, 28, -31, 22, -6, 57,
					-- layer=2 filter=91 channel=76
					25, -62, -34, -32, -49, -39, -3, 12, 4,
					-- layer=2 filter=91 channel=77
					4, 11, -1, 9, -7, 1, -5, -5, -5,
					-- layer=2 filter=91 channel=78
					-25, -8, 6, 0, 8, 13, 15, 15, 0,
					-- layer=2 filter=91 channel=79
					-7, -2, -5, 0, -5, -6, 0, 9, -7,
					-- layer=2 filter=91 channel=80
					53, 16, 7, -30, -21, -54, -46, -41, -55,
					-- layer=2 filter=91 channel=81
					-6, 8, -5, -5, -4, 0, -16, 0, -4,
					-- layer=2 filter=91 channel=82
					12, 4, -6, -8, -1, 10, -2, 1, 3,
					-- layer=2 filter=91 channel=83
					10, 19, 19, -36, -5, 29, -1, -34, -12,
					-- layer=2 filter=91 channel=84
					-2, 8, 7, 3, -4, -3, 5, -4, -2,
					-- layer=2 filter=91 channel=85
					0, 12, -4, 10, -3, 0, 11, -4, -4,
					-- layer=2 filter=91 channel=86
					1, 5, 11, -9, 0, 0, 1, -16, 6,
					-- layer=2 filter=91 channel=87
					29, 0, -80, 20, -44, -87, -4, 0, -60,
					-- layer=2 filter=91 channel=88
					0, 19, 23, 0, -40, 6, -34, -6, -1,
					-- layer=2 filter=91 channel=89
					0, -3, -41, 15, -11, -18, -37, 8, 11,
					-- layer=2 filter=91 channel=90
					9, 5, -7, 5, -3, 0, -7, -5, -3,
					-- layer=2 filter=91 channel=91
					-12, -33, -21, -4, -37, 1, -28, 0, 2,
					-- layer=2 filter=91 channel=92
					-46, 10, -2, 37, 15, 10, -5, 9, 0,
					-- layer=2 filter=91 channel=93
					-22, 13, -38, 27, 14, 10, -32, -20, -3,
					-- layer=2 filter=91 channel=94
					-25, -33, 23, -17, -10, -61, 22, 22, -8,
					-- layer=2 filter=91 channel=95
					-4, -16, -23, -7, -12, -4, -4, -9, -3,
					-- layer=2 filter=91 channel=96
					21, 5, -13, 39, 29, -30, -1, -16, 1,
					-- layer=2 filter=91 channel=97
					-1, 20, 25, -21, -10, 8, -29, -38, 18,
					-- layer=2 filter=91 channel=98
					-1, 15, -16, -16, -8, 57, 28, 15, -3,
					-- layer=2 filter=91 channel=99
					-27, -97, -12, 31, 4, -56, 40, -12, 14,
					-- layer=2 filter=91 channel=100
					34, -21, -26, -27, 8, -36, -12, -15, 8,
					-- layer=2 filter=91 channel=101
					-23, 37, 34, -68, -25, 40, -35, -40, 33,
					-- layer=2 filter=91 channel=102
					1, -4, -20, 25, 25, -34, 15, -12, -37,
					-- layer=2 filter=91 channel=103
					-36, -64, -20, -14, -14, 10, -14, -10, 27,
					-- layer=2 filter=91 channel=104
					19, 0, -29, -12, -2, -43, 13, 10, 0,
					-- layer=2 filter=91 channel=105
					15, 45, -43, 24, -18, 37, 11, 40, -70,
					-- layer=2 filter=91 channel=106
					-38, 7, -8, -20, -22, 43, -46, -27, 3,
					-- layer=2 filter=91 channel=107
					-29, 33, -22, 24, -13, -10, -13, 24, 32,
					-- layer=2 filter=91 channel=108
					-1, -45, -8, -1, 36, 19, -15, 2, 34,
					-- layer=2 filter=91 channel=109
					-3, 0, 7, 10, -14, 4, -7, -3, 2,
					-- layer=2 filter=91 channel=110
					-3, 34, -7, -17, 9, 3, -64, -18, -17,
					-- layer=2 filter=91 channel=111
					4, 0, 2, 7, -2, 4, 5, 9, -8,
					-- layer=2 filter=91 channel=112
					-46, -14, 12, -23, 26, 14, 32, 23, -9,
					-- layer=2 filter=91 channel=113
					-22, -8, -20, -27, -33, 27, -23, 4, -2,
					-- layer=2 filter=91 channel=114
					-3, -1, -3, -1, 9, -13, 10, -4, -7,
					-- layer=2 filter=91 channel=115
					6, 6, 6, -9, -8, -6, 5, -3, -5,
					-- layer=2 filter=91 channel=116
					44, 10, -84, 20, -6, -54, -7, 5, 3,
					-- layer=2 filter=91 channel=117
					-12, -1, -16, -24, -22, -5, -27, 43, 10,
					-- layer=2 filter=91 channel=118
					25, 20, -5, 2, 9, -11, 27, 2, -37,
					-- layer=2 filter=91 channel=119
					17, 39, -26, -8, 3, -23, -6, -10, 6,
					-- layer=2 filter=91 channel=120
					-2, 9, -3, -6, -3, 2, -3, -2, 7,
					-- layer=2 filter=91 channel=121
					-6, -1, 7, 5, 11, -2, 4, -4, 0,
					-- layer=2 filter=91 channel=122
					-6, -7, -2, 15, 7, 1, -3, 1, -4,
					-- layer=2 filter=91 channel=123
					38, -10, -7, 21, 24, 55, 13, 9, 0,
					-- layer=2 filter=91 channel=124
					-3, -15, -49, -5, -40, -31, -16, 10, -22,
					-- layer=2 filter=91 channel=125
					3, 4, 6, -6, 1, 7, -8, -4, -1,
					-- layer=2 filter=91 channel=126
					21, 16, 42, 0, 56, -27, -22, 17, -11,
					-- layer=2 filter=91 channel=127
					-3, 5, -16, 22, -28, -39, -47, -17, 0,
					-- layer=2 filter=92 channel=0
					-4, -18, -4, -15, -19, -4, -17, -13, -2,
					-- layer=2 filter=92 channel=1
					-8, 1, -7, -17, -5, 5, -15, -7, -15,
					-- layer=2 filter=92 channel=2
					1, -4, -5, -7, 6, 7, 3, 0, -8,
					-- layer=2 filter=92 channel=3
					-9, -9, -17, 0, -5, 2, -18, -8, 0,
					-- layer=2 filter=92 channel=4
					-9, -7, 0, -7, -4, 3, -18, -7, -2,
					-- layer=2 filter=92 channel=5
					-18, -9, -10, -1, -8, -10, -10, -4, -7,
					-- layer=2 filter=92 channel=6
					-18, -6, -5, -20, -5, -21, 0, -8, -13,
					-- layer=2 filter=92 channel=7
					-7, -15, -11, -4, 0, 0, -3, -9, -15,
					-- layer=2 filter=92 channel=8
					3, -3, -9, 0, 5, -6, 8, -9, -9,
					-- layer=2 filter=92 channel=9
					-17, -15, -10, 8, -4, -22, -16, -12, -12,
					-- layer=2 filter=92 channel=10
					-2, -11, -11, -6, -7, -12, 1, -2, -13,
					-- layer=2 filter=92 channel=11
					-6, 3, 0, -7, 5, 0, -3, 0, -4,
					-- layer=2 filter=92 channel=12
					-14, -8, -14, -13, 1, 0, -10, -4, 1,
					-- layer=2 filter=92 channel=13
					3, 6, 7, 8, 9, -9, -6, -11, 1,
					-- layer=2 filter=92 channel=14
					-4, -13, -12, 0, -2, -16, 0, -4, -10,
					-- layer=2 filter=92 channel=15
					-15, -8, 0, -20, -14, -8, 0, -7, -2,
					-- layer=2 filter=92 channel=16
					-7, -7, -15, -3, -3, -11, -9, -16, -13,
					-- layer=2 filter=92 channel=17
					-4, 3, -3, 0, -10, 6, 9, -8, 6,
					-- layer=2 filter=92 channel=18
					-16, -13, 0, -8, -17, -4, -5, -14, -19,
					-- layer=2 filter=92 channel=19
					-9, -3, -2, -24, -22, -15, -1, -12, -1,
					-- layer=2 filter=92 channel=20
					-8, -8, 0, 1, 6, 1, -11, -8, 1,
					-- layer=2 filter=92 channel=21
					-5, -5, 0, -11, 0, -12, 1, 0, -11,
					-- layer=2 filter=92 channel=22
					8, 11, -8, 7, 3, -9, 4, -7, 0,
					-- layer=2 filter=92 channel=23
					-22, -18, -17, -21, -12, -4, -1, -13, -15,
					-- layer=2 filter=92 channel=24
					-10, -5, -14, 4, -13, -14, -15, -12, -10,
					-- layer=2 filter=92 channel=25
					-17, 0, -2, -12, 7, 7, 0, -3, 9,
					-- layer=2 filter=92 channel=26
					4, 6, -10, -6, -7, 6, -8, -3, -2,
					-- layer=2 filter=92 channel=27
					-2, 12, 11, 8, -6, 4, -12, -11, -8,
					-- layer=2 filter=92 channel=28
					-2, 3, 1, -17, -11, -10, -3, -3, 4,
					-- layer=2 filter=92 channel=29
					0, 6, 0, -11, 5, -7, 3, -1, 2,
					-- layer=2 filter=92 channel=30
					-2, 0, -5, -13, -5, -10, -20, -15, -17,
					-- layer=2 filter=92 channel=31
					3, -5, -9, -3, -1, -4, 1, -7, 0,
					-- layer=2 filter=92 channel=32
					-8, -3, -2, 8, 0, -1, 6, -7, -4,
					-- layer=2 filter=92 channel=33
					-10, -8, 1, -11, -7, -6, -9, -4, -19,
					-- layer=2 filter=92 channel=34
					2, -17, -10, -5, -7, -6, -4, -15, 1,
					-- layer=2 filter=92 channel=35
					-17, -4, -18, -12, -5, -5, -6, 8, -1,
					-- layer=2 filter=92 channel=36
					-1, 0, -5, -5, -1, 2, -5, 3, -2,
					-- layer=2 filter=92 channel=37
					-8, -3, -12, -7, -3, -5, -1, -11, -6,
					-- layer=2 filter=92 channel=38
					-12, -2, -2, 1, -11, -17, -16, 4, 2,
					-- layer=2 filter=92 channel=39
					-9, -16, -13, -16, 0, -13, -1, 1, 0,
					-- layer=2 filter=92 channel=40
					-6, 0, -7, 4, -9, 6, 10, -5, 0,
					-- layer=2 filter=92 channel=41
					3, -7, 6, -6, 5, -11, -8, 1, 3,
					-- layer=2 filter=92 channel=42
					-18, -17, -9, -13, -7, 0, -6, -15, -6,
					-- layer=2 filter=92 channel=43
					19, -5, -16, 1, -13, -8, -7, 0, -4,
					-- layer=2 filter=92 channel=44
					0, -7, -5, 3, -5, 1, 0, 0, -9,
					-- layer=2 filter=92 channel=45
					-12, 4, -5, 1, -2, -5, 2, -9, -4,
					-- layer=2 filter=92 channel=46
					-5, -8, -3, -3, -1, -19, -15, -5, -15,
					-- layer=2 filter=92 channel=47
					6, 2, 1, 0, 0, -9, -6, -9, -5,
					-- layer=2 filter=92 channel=48
					8, 0, -3, 8, 6, -2, 9, -5, -9,
					-- layer=2 filter=92 channel=49
					-12, -13, -14, -9, -11, -19, -6, -3, -12,
					-- layer=2 filter=92 channel=50
					0, -5, 1, -4, 7, -10, 1, -3, -1,
					-- layer=2 filter=92 channel=51
					-4, -1, -19, -2, 0, -3, -4, -16, -16,
					-- layer=2 filter=92 channel=52
					-9, -11, 5, -19, -5, -15, 0, 0, -13,
					-- layer=2 filter=92 channel=53
					-3, -15, -16, -7, -1, -1, -4, -2, -8,
					-- layer=2 filter=92 channel=54
					-19, -8, -5, -10, -7, -1, -1, -8, -18,
					-- layer=2 filter=92 channel=55
					-7, 0, -1, 8, 5, -1, -6, 10, 1,
					-- layer=2 filter=92 channel=56
					4, -5, -12, 0, 7, 7, -2, 2, 7,
					-- layer=2 filter=92 channel=57
					-11, 5, 1, 8, 0, -3, 2, 1, -1,
					-- layer=2 filter=92 channel=58
					-20, -10, -19, -17, 6, -1, -18, -15, -1,
					-- layer=2 filter=92 channel=59
					0, 0, -10, -3, 10, 9, -8, 0, -1,
					-- layer=2 filter=92 channel=60
					-4, -7, 0, -23, -12, -18, -16, -13, -14,
					-- layer=2 filter=92 channel=61
					0, -9, -1, -13, -16, -20, -15, -16, -11,
					-- layer=2 filter=92 channel=62
					-4, -10, -15, -16, -18, -8, -16, -7, -7,
					-- layer=2 filter=92 channel=63
					-14, -15, -2, -12, -16, -2, -11, -11, -11,
					-- layer=2 filter=92 channel=64
					-17, -10, -5, -20, -11, -1, -8, -7, -11,
					-- layer=2 filter=92 channel=65
					4, -1, 6, 0, -12, -4, 0, -8, -1,
					-- layer=2 filter=92 channel=66
					-11, -11, -3, 0, 8, 10, 1, 4, -5,
					-- layer=2 filter=92 channel=67
					-6, -4, 0, -11, -15, 2, 3, -8, -11,
					-- layer=2 filter=92 channel=68
					-5, -10, 0, -8, -8, -11, -3, -9, 7,
					-- layer=2 filter=92 channel=69
					-3, -9, -10, 0, -10, -6, -15, -1, -9,
					-- layer=2 filter=92 channel=70
					-2, -6, -10, -12, -16, -16, -18, 0, -3,
					-- layer=2 filter=92 channel=71
					-8, 0, -2, -4, 2, 0, 1, 7, -9,
					-- layer=2 filter=92 channel=72
					-14, -14, -1, -22, -2, -5, -17, -5, 0,
					-- layer=2 filter=92 channel=73
					1, 0, -6, -16, -8, 0, -15, -13, -2,
					-- layer=2 filter=92 channel=74
					-15, -22, -5, -16, -2, 0, -8, -15, -14,
					-- layer=2 filter=92 channel=75
					-5, -14, -10, 0, -20, -6, 4, -10, -4,
					-- layer=2 filter=92 channel=76
					-16, -9, -2, -9, -9, 0, 4, 0, -6,
					-- layer=2 filter=92 channel=77
					-5, 8, 4, -8, -2, 7, -9, -10, -10,
					-- layer=2 filter=92 channel=78
					-16, 4, -10, 6, -6, -14, 0, 0, 1,
					-- layer=2 filter=92 channel=79
					3, 5, -5, 2, 3, 0, -10, 4, 0,
					-- layer=2 filter=92 channel=80
					-20, -15, -3, -2, 2, -12, -7, -6, -5,
					-- layer=2 filter=92 channel=81
					7, 8, 11, 1, -6, -3, -7, -5, 5,
					-- layer=2 filter=92 channel=82
					7, 8, -4, -3, -3, 3, 0, 8, 2,
					-- layer=2 filter=92 channel=83
					-9, -15, -7, -14, -18, -5, -4, -12, -10,
					-- layer=2 filter=92 channel=84
					0, -6, 3, 0, -9, 4, 3, -1, -5,
					-- layer=2 filter=92 channel=85
					7, -7, -1, 4, 1, 4, -5, 9, -2,
					-- layer=2 filter=92 channel=86
					9, -11, -7, -5, 0, 4, 8, -6, -4,
					-- layer=2 filter=92 channel=87
					0, -22, -7, -20, -8, -12, -1, -17, -10,
					-- layer=2 filter=92 channel=88
					-8, -1, -4, -12, -3, -5, -10, -10, -12,
					-- layer=2 filter=92 channel=89
					-3, -6, -13, 2, 2, -11, 3, -13, -15,
					-- layer=2 filter=92 channel=90
					-8, -2, -3, -3, -2, 5, -2, 4, 0,
					-- layer=2 filter=92 channel=91
					-21, -8, -4, -4, -4, -7, -4, 11, -11,
					-- layer=2 filter=92 channel=92
					-11, -5, -11, -9, -10, 5, -9, -20, -21,
					-- layer=2 filter=92 channel=93
					1, -4, -11, -5, 0, -3, -5, -3, -11,
					-- layer=2 filter=92 channel=94
					-17, -6, 2, -12, -20, -5, -3, -13, -18,
					-- layer=2 filter=92 channel=95
					9, 9, -6, 1, 0, -5, -4, 1, -10,
					-- layer=2 filter=92 channel=96
					-5, -2, -3, -5, -11, -15, -9, -3, -6,
					-- layer=2 filter=92 channel=97
					-19, -19, -2, -5, -1, -5, -4, -9, -3,
					-- layer=2 filter=92 channel=98
					1, -7, -6, -4, -6, -11, -3, -4, 1,
					-- layer=2 filter=92 channel=99
					-6, -10, 15, -2, 5, 5, -11, -1, 11,
					-- layer=2 filter=92 channel=100
					5, -9, -19, 1, -9, -1, -4, -4, -8,
					-- layer=2 filter=92 channel=101
					0, 0, -7, 3, -6, -11, 5, 2, -3,
					-- layer=2 filter=92 channel=102
					-19, 3, -1, -20, -14, -11, 2, -18, -18,
					-- layer=2 filter=92 channel=103
					0, -5, 4, -1, 0, 0, -14, -12, 0,
					-- layer=2 filter=92 channel=104
					-14, -5, 0, -7, -3, -12, 7, -6, -6,
					-- layer=2 filter=92 channel=105
					-13, -8, 2, 7, 1, -1, -15, 4, -3,
					-- layer=2 filter=92 channel=106
					-26, 0, -10, -2, -7, -5, -7, 0, 0,
					-- layer=2 filter=92 channel=107
					-2, 6, -5, -7, -1, 0, -5, -1, -1,
					-- layer=2 filter=92 channel=108
					-9, -9, -7, -4, -2, -8, -10, 0, -14,
					-- layer=2 filter=92 channel=109
					1, -1, -6, 0, -3, 0, 6, 0, -2,
					-- layer=2 filter=92 channel=110
					-8, -18, -11, -1, -5, 6, -9, -4, -19,
					-- layer=2 filter=92 channel=111
					-3, 1, 3, -6, -6, 6, -5, 2, -3,
					-- layer=2 filter=92 channel=112
					3, 3, -10, 0, 5, 1, -15, 3, 7,
					-- layer=2 filter=92 channel=113
					-16, -1, -19, -9, -16, -9, -11, -7, -15,
					-- layer=2 filter=92 channel=114
					6, -7, 2, -4, -1, -11, -5, 3, 5,
					-- layer=2 filter=92 channel=115
					1, 3, 7, 0, 3, -5, 0, -1, -7,
					-- layer=2 filter=92 channel=116
					-11, 0, -19, -14, -11, -20, 3, -23, -15,
					-- layer=2 filter=92 channel=117
					-7, -4, -12, -5, 3, -3, -8, -10, 0,
					-- layer=2 filter=92 channel=118
					-16, -3, -17, -7, -12, -19, -13, -4, 2,
					-- layer=2 filter=92 channel=119
					0, -8, -14, -17, -5, -6, -2, -11, -19,
					-- layer=2 filter=92 channel=120
					-1, 8, 3, -3, -10, -7, 2, 3, -7,
					-- layer=2 filter=92 channel=121
					-6, -7, 5, 4, -4, 6, -8, -4, -11,
					-- layer=2 filter=92 channel=122
					3, 0, 0, 1, -3, 4, -4, -9, -10,
					-- layer=2 filter=92 channel=123
					-7, -5, 8, -9, -9, -17, -9, -9, -10,
					-- layer=2 filter=92 channel=124
					-14, 1, -8, -10, -18, -7, -17, -8, -17,
					-- layer=2 filter=92 channel=125
					5, -1, -5, -7, 7, 1, 7, 8, 8,
					-- layer=2 filter=92 channel=126
					-14, 0, 4, 3, -6, -7, -7, -15, 2,
					-- layer=2 filter=92 channel=127
					0, 4, -11, -12, -2, -9, 3, -17, -9,
					-- layer=2 filter=93 channel=0
					-6, -25, -28, -14, -1, -20, -9, -37, -1,
					-- layer=2 filter=93 channel=1
					-14, -10, 1, 4, -4, -12, 4, -10, -11,
					-- layer=2 filter=93 channel=2
					0, 0, 10, -4, -2, 8, 0, 7, 0,
					-- layer=2 filter=93 channel=3
					-21, -1, -2, -6, -10, 4, -10, -26, -9,
					-- layer=2 filter=93 channel=4
					-61, -13, -20, -22, -30, -23, -34, -2, -6,
					-- layer=2 filter=93 channel=5
					0, -13, -5, -11, 3, -15, -16, 14, -1,
					-- layer=2 filter=93 channel=6
					-24, 0, 14, -28, -29, -6, -24, 6, 9,
					-- layer=2 filter=93 channel=7
					-23, 6, 7, 13, -12, -4, -22, -7, -6,
					-- layer=2 filter=93 channel=8
					-3, -4, 0, -4, 4, -4, 6, 0, 1,
					-- layer=2 filter=93 channel=9
					9, -4, -10, 6, -8, -20, -20, 2, -6,
					-- layer=2 filter=93 channel=10
					-7, -6, -13, -12, -20, -1, 2, -29, -21,
					-- layer=2 filter=93 channel=11
					0, -6, -2, -17, 5, -11, -3, -7, -9,
					-- layer=2 filter=93 channel=12
					-22, -26, -12, 27, -4, -6, -3, -27, -14,
					-- layer=2 filter=93 channel=13
					-9, -8, -8, -2, -8, -2, 6, -8, -5,
					-- layer=2 filter=93 channel=14
					-3, -17, -22, -3, 10, -13, -10, -14, -24,
					-- layer=2 filter=93 channel=15
					-18, -7, -5, -9, -8, 2, 17, 18, 21,
					-- layer=2 filter=93 channel=16
					-21, -13, -12, -4, -4, 2, 5, -9, -18,
					-- layer=2 filter=93 channel=17
					2, -1, -10, 3, -1, 0, -4, 7, 7,
					-- layer=2 filter=93 channel=18
					-36, -10, -17, -11, -17, -7, -17, 22, 1,
					-- layer=2 filter=93 channel=19
					0, 11, 16, 6, -1, 5, -11, 6, -9,
					-- layer=2 filter=93 channel=20
					-5, 3, 7, -9, -12, -11, 1, 6, -4,
					-- layer=2 filter=93 channel=21
					-7, -10, -9, 0, 4, -7, 8, -1, 1,
					-- layer=2 filter=93 channel=22
					-4, 8, 4, -2, 0, -1, 7, -8, -2,
					-- layer=2 filter=93 channel=23
					-17, -9, -26, -38, -31, -5, -43, -22, -12,
					-- layer=2 filter=93 channel=24
					0, -10, 0, -7, -24, 3, 9, -10, -7,
					-- layer=2 filter=93 channel=25
					-6, -2, 2, 9, 0, -8, 11, 0, 18,
					-- layer=2 filter=93 channel=26
					5, 0, 5, 5, 10, 1, -3, -1, 2,
					-- layer=2 filter=93 channel=27
					31, 14, -1, 6, 16, -5, -13, -17, -16,
					-- layer=2 filter=93 channel=28
					6, -10, -19, -16, -20, 9, -19, -37, -4,
					-- layer=2 filter=93 channel=29
					9, -4, -5, 0, 2, 5, -2, -11, 4,
					-- layer=2 filter=93 channel=30
					-3, -38, -25, -48, -10, -10, -39, -18, -30,
					-- layer=2 filter=93 channel=31
					8, 9, 17, -7, -11, 18, 10, 13, -18,
					-- layer=2 filter=93 channel=32
					0, -8, 4, -1, -12, -8, 1, 1, 4,
					-- layer=2 filter=93 channel=33
					-3, -25, -3, -15, -8, 0, -10, 0, -17,
					-- layer=2 filter=93 channel=34
					-19, -31, -14, -29, 11, -18, -9, -30, 4,
					-- layer=2 filter=93 channel=35
					-22, 1, -2, 2, 0, -7, 12, -6, -5,
					-- layer=2 filter=93 channel=36
					-6, -1, 0, -1, 6, -1, 5, -9, 7,
					-- layer=2 filter=93 channel=37
					7, -5, -7, 0, 12, 7, 3, 1, -6,
					-- layer=2 filter=93 channel=38
					17, 0, -11, -1, -7, -21, -23, -26, -30,
					-- layer=2 filter=93 channel=39
					-27, -5, -9, -28, -10, -12, -17, -24, 1,
					-- layer=2 filter=93 channel=40
					-6, -16, 11, -14, 3, 22, 9, 9, 40,
					-- layer=2 filter=93 channel=41
					-8, -2, -2, -9, -6, -3, 0, -8, -8,
					-- layer=2 filter=93 channel=42
					-11, -17, -9, 6, -25, -1, -6, -28, -17,
					-- layer=2 filter=93 channel=43
					-9, 5, -22, -15, -13, -19, 7, -17, -9,
					-- layer=2 filter=93 channel=44
					-5, -2, -1, 6, 5, 0, 2, -5, -8,
					-- layer=2 filter=93 channel=45
					32, 20, -8, 22, 6, -19, -8, -22, -4,
					-- layer=2 filter=93 channel=46
					6, 1, -22, -21, -21, -24, -13, -27, -18,
					-- layer=2 filter=93 channel=47
					-1, 6, -19, -25, -26, -3, -31, -28, -6,
					-- layer=2 filter=93 channel=48
					-1, 0, 7, -5, 4, 11, 10, 6, 0,
					-- layer=2 filter=93 channel=49
					-21, -36, -6, -8, -30, -14, 2, 7, -11,
					-- layer=2 filter=93 channel=50
					-5, 3, -5, 0, -1, -3, 5, 2, -10,
					-- layer=2 filter=93 channel=51
					0, 1, -15, -23, -15, -9, -9, -8, 1,
					-- layer=2 filter=93 channel=52
					-16, -1, 0, -26, 5, 9, -3, 0, -1,
					-- layer=2 filter=93 channel=53
					-36, 0, 4, -6, 0, 3, 13, -18, 13,
					-- layer=2 filter=93 channel=54
					-24, -8, -6, -6, -19, -3, -23, -5, 7,
					-- layer=2 filter=93 channel=55
					2, -8, 3, 7, -4, -3, 1, -6, 8,
					-- layer=2 filter=93 channel=56
					7, -10, -23, 0, 19, -1, -9, 0, 2,
					-- layer=2 filter=93 channel=57
					-9, -10, -3, 0, -2, 7, -4, 7, 5,
					-- layer=2 filter=93 channel=58
					11, 6, -24, 25, 18, 24, 4, -9, -7,
					-- layer=2 filter=93 channel=59
					0, -11, -3, 12, -19, 2, -13, -18, -11,
					-- layer=2 filter=93 channel=60
					-25, -3, -2, -12, -12, 18, -30, -6, -12,
					-- layer=2 filter=93 channel=61
					4, 3, 12, -22, -24, 8, -21, -39, -5,
					-- layer=2 filter=93 channel=62
					-28, 4, -22, -22, -32, -5, 6, -10, 10,
					-- layer=2 filter=93 channel=63
					-30, -28, -30, -38, -31, -14, -25, -23, -15,
					-- layer=2 filter=93 channel=64
					-28, -26, -12, -28, -13, -29, -13, -7, -14,
					-- layer=2 filter=93 channel=65
					-5, 5, 0, -27, -9, -1, -8, -15, -1,
					-- layer=2 filter=93 channel=66
					2, -15, -24, 0, -9, 3, 1, -1, 0,
					-- layer=2 filter=93 channel=67
					11, -12, -16, 6, -11, -16, -8, -27, 19,
					-- layer=2 filter=93 channel=68
					3, 1, 0, 0, -3, 8, 4, -11, 5,
					-- layer=2 filter=93 channel=69
					-25, -19, -30, -26, -13, -15, -20, -31, -29,
					-- layer=2 filter=93 channel=70
					0, 3, 14, -5, 26, 13, -19, -21, -13,
					-- layer=2 filter=93 channel=71
					10, 9, 10, 10, 1, -24, -10, -10, -27,
					-- layer=2 filter=93 channel=72
					-17, -15, -1, -4, -24, -7, -22, 7, -22,
					-- layer=2 filter=93 channel=73
					0, -13, 19, -12, -15, -12, 25, -3, -1,
					-- layer=2 filter=93 channel=74
					-17, -39, -21, -28, -20, -9, -14, -7, 13,
					-- layer=2 filter=93 channel=75
					-7, -12, -8, 27, 0, -4, 13, 11, -10,
					-- layer=2 filter=93 channel=76
					-18, 7, 0, -20, -13, -2, -19, 14, 7,
					-- layer=2 filter=93 channel=77
					-8, -10, -3, -2, -2, -10, 2, -3, -9,
					-- layer=2 filter=93 channel=78
					-15, -19, -12, -17, -20, -11, 0, -10, -19,
					-- layer=2 filter=93 channel=79
					4, 4, -9, -2, -2, 1, 1, 4, 5,
					-- layer=2 filter=93 channel=80
					-35, -20, -27, -34, -39, -11, -7, -19, -27,
					-- layer=2 filter=93 channel=81
					1, 1, 6, -5, 0, -2, -5, -10, 2,
					-- layer=2 filter=93 channel=82
					7, 3, 4, 5, 2, 7, 3, -1, 1,
					-- layer=2 filter=93 channel=83
					5, -3, -13, 11, -10, -11, -33, -10, -29,
					-- layer=2 filter=93 channel=84
					-5, 7, 0, 2, -7, -9, -5, 0, -5,
					-- layer=2 filter=93 channel=85
					-3, 1, 3, 11, 5, -2, -6, -3, 3,
					-- layer=2 filter=93 channel=86
					3, 4, -1, 10, -7, -11, 6, 0, -4,
					-- layer=2 filter=93 channel=87
					-11, 0, -16, -13, 12, -5, -11, -7, 4,
					-- layer=2 filter=93 channel=88
					1, -43, -11, -30, -16, -15, -26, -39, -17,
					-- layer=2 filter=93 channel=89
					-31, -6, -4, 15, 12, 8, 4, 5, 6,
					-- layer=2 filter=93 channel=90
					0, 3, 1, 6, -6, -2, 6, 0, -6,
					-- layer=2 filter=93 channel=91
					-14, 17, -14, 28, 12, 3, 5, 5, -19,
					-- layer=2 filter=93 channel=92
					-15, -18, -15, 32, -12, 0, -8, 1, -10,
					-- layer=2 filter=93 channel=93
					4, 2, 13, -35, 4, 8, -11, -7, 2,
					-- layer=2 filter=93 channel=94
					-15, -5, 1, -4, -19, -7, -14, -16, 11,
					-- layer=2 filter=93 channel=95
					-9, 2, 5, -5, 1, -7, -6, -2, -5,
					-- layer=2 filter=93 channel=96
					-23, -10, -4, -5, -5, 9, -17, 18, 3,
					-- layer=2 filter=93 channel=97
					-7, -7, -18, 3, -27, -12, 8, -14, -7,
					-- layer=2 filter=93 channel=98
					-18, 12, 12, -16, -17, 0, -20, -29, -12,
					-- layer=2 filter=93 channel=99
					4, 18, 14, -2, 4, 16, -8, 4, 13,
					-- layer=2 filter=93 channel=100
					8, 0, -23, -2, -10, 4, -30, -13, -20,
					-- layer=2 filter=93 channel=101
					1, -12, 15, 13, -2, -2, 4, -18, -20,
					-- layer=2 filter=93 channel=102
					-24, -35, -5, -25, -1, 1, -6, 19, 6,
					-- layer=2 filter=93 channel=103
					5, 1, -14, -4, 8, -12, 9, -28, 0,
					-- layer=2 filter=93 channel=104
					-14, -32, -15, 12, -8, -12, -12, -6, -1,
					-- layer=2 filter=93 channel=105
					-18, 19, -18, -20, -10, 4, -8, 0, 6,
					-- layer=2 filter=93 channel=106
					8, -5, 5, 15, -2, -5, -8, -12, 1,
					-- layer=2 filter=93 channel=107
					23, 1, 17, 17, 6, -19, -15, 1, 10,
					-- layer=2 filter=93 channel=108
					20, 7, -15, 19, 18, -19, -16, 6, -19,
					-- layer=2 filter=93 channel=109
					-7, -4, 2, 7, 5, 2, -2, -6, -10,
					-- layer=2 filter=93 channel=110
					-19, -21, -1, 0, -23, -5, 28, -22, -12,
					-- layer=2 filter=93 channel=111
					7, -6, 2, -1, 7, 8, 5, -1, 4,
					-- layer=2 filter=93 channel=112
					12, 23, -5, -8, -6, 17, -5, -14, 13,
					-- layer=2 filter=93 channel=113
					1, -17, -31, -25, -16, 7, -32, -27, -21,
					-- layer=2 filter=93 channel=114
					2, 7, 0, 11, 4, -9, -9, 4, 4,
					-- layer=2 filter=93 channel=115
					0, -7, 8, -10, 2, -5, 3, 8, 8,
					-- layer=2 filter=93 channel=116
					-4, -12, 1, -22, -12, -1, 12, 3, 10,
					-- layer=2 filter=93 channel=117
					-27, 12, 6, 13, -28, -15, -30, -5, -14,
					-- layer=2 filter=93 channel=118
					-17, -2, -13, -35, -3, -2, -23, -28, -33,
					-- layer=2 filter=93 channel=119
					-37, -10, -43, -10, -9, -18, -48, -10, 0,
					-- layer=2 filter=93 channel=120
					-9, -7, 2, -4, 9, 0, -1, 1, 1,
					-- layer=2 filter=93 channel=121
					-1, -6, -8, -10, 0, -5, 8, -8, 4,
					-- layer=2 filter=93 channel=122
					1, -5, -2, 6, -1, 5, 2, -2, -5,
					-- layer=2 filter=93 channel=123
					-13, -7, 2, -27, -31, -5, -20, -10, 3,
					-- layer=2 filter=93 channel=124
					-13, -16, 10, -25, -9, 8, -16, -8, -17,
					-- layer=2 filter=93 channel=125
					2, -7, -1, 4, 1, 2, -10, 1, 3,
					-- layer=2 filter=93 channel=126
					-18, -28, -4, 6, -14, 7, -15, -13, 18,
					-- layer=2 filter=93 channel=127
					2, -18, -19, -19, -35, -8, -52, -18, -12,
					-- layer=2 filter=94 channel=0
					-13, 1, -28, 0, -9, -12, 0, 22, 11,
					-- layer=2 filter=94 channel=1
					-10, -3, 19, -15, -17, -29, -2, -39, -28,
					-- layer=2 filter=94 channel=2
					4, 6, -9, 3, -6, -5, -10, -12, 0,
					-- layer=2 filter=94 channel=3
					0, -18, -40, -7, -2, -7, -11, -1, 11,
					-- layer=2 filter=94 channel=4
					16, -20, -12, 14, -3, -16, -18, 20, 0,
					-- layer=2 filter=94 channel=5
					-31, -10, 29, 1, -8, 11, 7, 21, 11,
					-- layer=2 filter=94 channel=6
					-3, -81, 0, -21, -30, -32, -7, -12, -11,
					-- layer=2 filter=94 channel=7
					14, -12, -53, 38, 6, 8, 7, -15, -22,
					-- layer=2 filter=94 channel=8
					-1, 4, 5, 0, 2, 9, -6, 8, -2,
					-- layer=2 filter=94 channel=9
					14, -12, -39, -16, -38, -16, -11, -32, -9,
					-- layer=2 filter=94 channel=10
					-4, -11, -27, 7, 2, -36, 10, 19, 18,
					-- layer=2 filter=94 channel=11
					-7, -5, 20, 8, 23, 16, -8, 0, 8,
					-- layer=2 filter=94 channel=12
					16, -12, 16, 28, -9, -17, -2, -36, -22,
					-- layer=2 filter=94 channel=13
					-2, 1, 2, -5, 6, -6, 5, 6, -9,
					-- layer=2 filter=94 channel=14
					0, -12, 17, -17, -30, -20, -20, -38, -42,
					-- layer=2 filter=94 channel=15
					-13, 29, 32, -17, 19, 68, 12, 10, 73,
					-- layer=2 filter=94 channel=16
					19, -9, -34, -2, 25, 8, -16, -13, 20,
					-- layer=2 filter=94 channel=17
					5, -5, -3, -8, 9, -9, 0, 7, 8,
					-- layer=2 filter=94 channel=18
					-10, 0, 40, -19, -15, 24, -7, 15, 24,
					-- layer=2 filter=94 channel=19
					-14, -1, 8, -31, -29, -15, -10, -39, -44,
					-- layer=2 filter=94 channel=20
					-9, -1, 2, 1, -6, 4, -3, 2, 0,
					-- layer=2 filter=94 channel=21
					7, 9, 4, 11, 2, 0, 2, 6, 7,
					-- layer=2 filter=94 channel=22
					-6, -3, 7, 2, 7, 0, 8, -6, 4,
					-- layer=2 filter=94 channel=23
					8, 10, -2, -1, 18, -5, -11, -7, -27,
					-- layer=2 filter=94 channel=24
					6, 0, -32, 11, 10, -19, -21, -19, -16,
					-- layer=2 filter=94 channel=25
					15, 3, -18, 3, 37, 22, -22, 4, 2,
					-- layer=2 filter=94 channel=26
					3, -1, -10, -5, 4, -5, 3, 0, -6,
					-- layer=2 filter=94 channel=27
					-8, 15, 38, -32, 1, 0, -16, -10, -5,
					-- layer=2 filter=94 channel=28
					22, 23, -6, 4, -1, 17, -11, -31, -17,
					-- layer=2 filter=94 channel=29
					-5, 0, -2, -3, 6, 5, 6, -7, -1,
					-- layer=2 filter=94 channel=30
					4, -5, -40, -28, -48, -41, 22, -19, -20,
					-- layer=2 filter=94 channel=31
					-15, -83, -69, -76, 19, -30, -10, 13, -4,
					-- layer=2 filter=94 channel=32
					0, -6, 0, 0, -3, 1, 5, 8, -1,
					-- layer=2 filter=94 channel=33
					18, 46, 31, 42, -7, 9, -6, 0, 14,
					-- layer=2 filter=94 channel=34
					13, 35, 29, 57, -3, 58, 15, 51, 58,
					-- layer=2 filter=94 channel=35
					1, 21, 12, 9, 9, 43, -25, 4, -3,
					-- layer=2 filter=94 channel=36
					3, -7, -6, 10, -5, -2, 0, -4, 2,
					-- layer=2 filter=94 channel=37
					-13, -10, 6, 6, 6, 22, -7, 6, 2,
					-- layer=2 filter=94 channel=38
					-6, -37, 25, -36, -21, 0, -1, -15, 8,
					-- layer=2 filter=94 channel=39
					31, 8, -45, 2, 36, 22, 26, 23, 27,
					-- layer=2 filter=94 channel=40
					43, 44, 21, -49, 14, 14, 19, 35, 45,
					-- layer=2 filter=94 channel=41
					0, 0, 9, -6, -6, 0, 8, -12, -10,
					-- layer=2 filter=94 channel=42
					15, 8, -15, -19, 28, -1, -6, -23, -21,
					-- layer=2 filter=94 channel=43
					1, 23, 34, -38, 15, 11, -9, 17, 45,
					-- layer=2 filter=94 channel=44
					-7, -5, -5, 4, -1, -13, -5, -8, -5,
					-- layer=2 filter=94 channel=45
					26, 22, -23, -2, -39, -67, -16, -1, 7,
					-- layer=2 filter=94 channel=46
					-16, -19, -8, -17, -27, -24, 26, -30, 7,
					-- layer=2 filter=94 channel=47
					32, 37, -4, 4, -7, -24, -12, 0, 0,
					-- layer=2 filter=94 channel=48
					8, 3, -4, -7, -8, -11, 10, 4, -5,
					-- layer=2 filter=94 channel=49
					-27, 0, 5, -69, -29, -27, -30, -38, 10,
					-- layer=2 filter=94 channel=50
					7, 5, 10, 26, 3, 9, 8, -1, -8,
					-- layer=2 filter=94 channel=51
					-11, -18, -12, -7, -5, 17, 17, 14, -5,
					-- layer=2 filter=94 channel=52
					5, 43, 48, 17, -40, -2, -9, -1, 12,
					-- layer=2 filter=94 channel=53
					24, -78, 25, -50, -62, -60, 9, -38, -18,
					-- layer=2 filter=94 channel=54
					35, 17, 22, 30, 17, 22, 26, 20, 7,
					-- layer=2 filter=94 channel=55
					0, 0, 0, -7, 7, 11, -2, 1, 7,
					-- layer=2 filter=94 channel=56
					-1, -21, 9, -2, 18, 17, -17, -15, -7,
					-- layer=2 filter=94 channel=57
					9, -13, 0, -6, 4, -3, 2, -12, -17,
					-- layer=2 filter=94 channel=58
					23, -16, -5, 30, 31, 21, 16, 6, 5,
					-- layer=2 filter=94 channel=59
					36, 17, 78, 11, 14, 48, 14, 15, 14,
					-- layer=2 filter=94 channel=60
					20, 20, 9, 23, 20, 33, 29, 1, -7,
					-- layer=2 filter=94 channel=61
					-43, -23, -53, -18, -41, -40, -14, 19, -35,
					-- layer=2 filter=94 channel=62
					4, -4, 17, 13, -10, 34, 25, 0, 38,
					-- layer=2 filter=94 channel=63
					38, 21, -36, 8, -5, -8, 23, -14, 5,
					-- layer=2 filter=94 channel=64
					8, 0, -30, 8, 21, -18, 3, 25, -32,
					-- layer=2 filter=94 channel=65
					-50, -55, -25, -23, -41, -3, -14, -43, 0,
					-- layer=2 filter=94 channel=66
					13, 60, -5, 30, 24, -1, 1, 38, -15,
					-- layer=2 filter=94 channel=67
					-5, -22, 14, -13, -31, -23, 12, -3, 39,
					-- layer=2 filter=94 channel=68
					-8, 9, 7, 0, 6, 1, 7, -3, 6,
					-- layer=2 filter=94 channel=69
					33, 21, -20, -3, 19, -9, 8, -11, -17,
					-- layer=2 filter=94 channel=70
					9, 25, 9, 17, 7, 6, -4, 0, 12,
					-- layer=2 filter=94 channel=71
					-12, 29, 14, 4, 27, 56, -8, -7, 16,
					-- layer=2 filter=94 channel=72
					7, 21, 55, 32, 13, 14, 40, -48, -39,
					-- layer=2 filter=94 channel=73
					-10, -59, -11, -18, -40, -53, 2, 35, -2,
					-- layer=2 filter=94 channel=74
					15, -27, 19, -16, 2, 2, -3, -6, 5,
					-- layer=2 filter=94 channel=75
					-43, -1, -15, -13, -25, 4, -16, -35, -35,
					-- layer=2 filter=94 channel=76
					33, -40, 26, -67, -27, -15, -11, 15, -73,
					-- layer=2 filter=94 channel=77
					1, 0, -4, 6, -11, -4, -3, -5, -8,
					-- layer=2 filter=94 channel=78
					-10, -31, -17, -10, -10, 31, -21, -15, 29,
					-- layer=2 filter=94 channel=79
					-4, -5, -7, 3, 6, 1, -5, -5, -10,
					-- layer=2 filter=94 channel=80
					14, -3, -47, -17, -1, -35, -23, 5, 24,
					-- layer=2 filter=94 channel=81
					15, 12, 8, 11, 11, -2, -5, -7, 6,
					-- layer=2 filter=94 channel=82
					9, 7, -12, -4, -2, -6, 0, 7, -11,
					-- layer=2 filter=94 channel=83
					17, 18, 15, -16, -8, -26, -25, 2, -3,
					-- layer=2 filter=94 channel=84
					4, -9, -3, 8, 7, 9, -5, -11, -5,
					-- layer=2 filter=94 channel=85
					-1, 14, 4, -12, 16, 1, -6, -1, 8,
					-- layer=2 filter=94 channel=86
					10, 5, 2, 21, -9, 10, 2, -3, 5,
					-- layer=2 filter=94 channel=87
					6, -4, 46, 2, 40, 58, 7, 19, 17,
					-- layer=2 filter=94 channel=88
					26, 23, 19, -10, 12, -3, -14, -10, -31,
					-- layer=2 filter=94 channel=89
					19, 8, 58, 16, 4, -1, 5, -37, -17,
					-- layer=2 filter=94 channel=90
					1, 3, -8, 5, 5, 2, 11, 7, -1,
					-- layer=2 filter=94 channel=91
					23, 21, 18, 30, 31, 20, 6, -55, 0,
					-- layer=2 filter=94 channel=92
					-4, -14, 29, -3, -6, 5, 16, -31, 2,
					-- layer=2 filter=94 channel=93
					8, 1, -32, 0, 3, 23, -19, -28, 49,
					-- layer=2 filter=94 channel=94
					-54, -65, -26, -61, -84, -28, -46, -3, -35,
					-- layer=2 filter=94 channel=95
					-1, 0, -10, 7, 4, 0, -6, 2, -9,
					-- layer=2 filter=94 channel=96
					-22, -52, -7, -30, -44, -18, -43, -7, -39,
					-- layer=2 filter=94 channel=97
					-9, -17, -37, -38, 1, -42, -48, -33, -30,
					-- layer=2 filter=94 channel=98
					43, 35, 5, 13, -1, 32, 2, -9, -14,
					-- layer=2 filter=94 channel=99
					-30, -32, -17, -42, -56, -23, 8, 0, -54,
					-- layer=2 filter=94 channel=100
					2, 13, 25, -6, 36, 36, 11, 17, 37,
					-- layer=2 filter=94 channel=101
					-21, 11, -4, -3, 2, 25, -27, 26, 21,
					-- layer=2 filter=94 channel=102
					-59, -65, -9, -30, -68, -32, -42, -16, -28,
					-- layer=2 filter=94 channel=103
					-28, -46, -38, -66, -65, 9, 56, -34, -23,
					-- layer=2 filter=94 channel=104
					-26, -58, 4, -56, -60, -12, -57, -42, -19,
					-- layer=2 filter=94 channel=105
					0, -58, 57, -3, 16, -43, -48, -68, -30,
					-- layer=2 filter=94 channel=106
					15, 19, -4, 25, 30, 13, -3, -23, 1,
					-- layer=2 filter=94 channel=107
					-32, 23, 27, -27, -10, -2, -28, 15, -24,
					-- layer=2 filter=94 channel=108
					-40, -25, -8, -32, -41, -53, -21, -56, -41,
					-- layer=2 filter=94 channel=109
					-4, -5, 7, -6, -2, -1, 3, 1, 2,
					-- layer=2 filter=94 channel=110
					3, 8, 6, -13, 28, 22, -16, -10, -32,
					-- layer=2 filter=94 channel=111
					0, 5, 7, -7, -9, -8, 1, -2, -8,
					-- layer=2 filter=94 channel=112
					-17, -3, -17, -32, -12, -25, 16, 2, 8,
					-- layer=2 filter=94 channel=113
					26, -30, -39, -28, -17, -38, 16, -30, -1,
					-- layer=2 filter=94 channel=114
					-17, -6, -19, 0, -11, 1, 1, 7, -2,
					-- layer=2 filter=94 channel=115
					-10, -6, -5, -3, -8, 4, 2, -8, -3,
					-- layer=2 filter=94 channel=116
					20, 28, 51, 18, 38, 70, 16, 16, 43,
					-- layer=2 filter=94 channel=117
					-14, -36, -20, -32, -40, -26, -4, -29, -50,
					-- layer=2 filter=94 channel=118
					6, -31, -24, -13, 0, -6, -18, 15, 22,
					-- layer=2 filter=94 channel=119
					-12, 5, 4, 3, -8, 0, 10, 14, 5,
					-- layer=2 filter=94 channel=120
					0, 1, -9, -6, -6, -9, 1, -10, -5,
					-- layer=2 filter=94 channel=121
					-1, -4, -3, 2, 3, 0, -10, 0, -1,
					-- layer=2 filter=94 channel=122
					-7, -16, 5, 4, 0, 2, 0, 7, 2,
					-- layer=2 filter=94 channel=123
					20, 11, 5, 32, 5, 14, 28, -27, -2,
					-- layer=2 filter=94 channel=124
					16, 12, 48, -12, 25, 45, -22, 43, 35,
					-- layer=2 filter=94 channel=125
					7, 8, 12, 5, 0, -2, -5, -5, 5,
					-- layer=2 filter=94 channel=126
					-15, 0, 1, -15, -45, -53, 22, 57, 3,
					-- layer=2 filter=94 channel=127
					-2, -10, 11, -17, 2, -6, -16, -9, 0,
					-- layer=2 filter=95 channel=0
					-2, 15, 10, 31, 1, -33, -8, -13, -36,
					-- layer=2 filter=95 channel=1
					-23, -7, 0, -20, -16, -14, 8, -1, 12,
					-- layer=2 filter=95 channel=2
					-5, 2, 9, 2, 9, -1, 7, 11, 5,
					-- layer=2 filter=95 channel=3
					29, 46, -4, 26, 60, -14, 10, 41, -37,
					-- layer=2 filter=95 channel=4
					0, 19, -5, -7, -7, -5, -50, 7, -25,
					-- layer=2 filter=95 channel=5
					16, 1, -10, 5, 9, -21, 5, 0, -19,
					-- layer=2 filter=95 channel=6
					-2, -127, -23, -31, -76, 24, -8, -24, 66,
					-- layer=2 filter=95 channel=7
					20, 20, -8, 6, 9, 11, -24, -2, 28,
					-- layer=2 filter=95 channel=8
					-8, -3, -3, -5, -5, 9, -9, -6, -7,
					-- layer=2 filter=95 channel=9
					-5, 30, 16, -17, 35, -5, -7, -18, -47,
					-- layer=2 filter=95 channel=10
					22, 40, 17, 24, 58, -36, -8, 16, -20,
					-- layer=2 filter=95 channel=11
					-10, -6, -14, -5, 4, -19, 8, -6, -34,
					-- layer=2 filter=95 channel=12
					21, 23, 6, 3, -1, -11, 12, 6, -16,
					-- layer=2 filter=95 channel=13
					-3, 10, 9, -5, 4, 3, 5, 3, 2,
					-- layer=2 filter=95 channel=14
					-18, -5, 3, -19, -16, -25, 18, 7, -17,
					-- layer=2 filter=95 channel=15
					-32, 21, 17, 5, 63, 64, 42, 17, 31,
					-- layer=2 filter=95 channel=16
					13, -34, -24, 6, 15, 9, -18, -21, 1,
					-- layer=2 filter=95 channel=17
					-12, 7, 9, 0, -1, -11, 2, -3, -9,
					-- layer=2 filter=95 channel=18
					-58, -8, 3, -24, -58, 22, -2, -46, 11,
					-- layer=2 filter=95 channel=19
					-21, -31, 23, 9, -8, 43, 15, -19, 48,
					-- layer=2 filter=95 channel=20
					-7, -2, 4, 8, 6, 5, 5, -4, 6,
					-- layer=2 filter=95 channel=21
					-16, -8, -15, -11, -10, 11, -6, -4, 18,
					-- layer=2 filter=95 channel=22
					1, 5, 2, 7, -3, 4, -8, -7, 4,
					-- layer=2 filter=95 channel=23
					-5, -13, -15, 31, 15, 17, 20, -7, 2,
					-- layer=2 filter=95 channel=24
					3, 25, -10, 4, 25, -19, -19, 7, -43,
					-- layer=2 filter=95 channel=25
					-4, 10, -24, -7, -2, -32, -22, 0, -28,
					-- layer=2 filter=95 channel=26
					-6, 7, 1, 9, 9, 3, -2, 2, -4,
					-- layer=2 filter=95 channel=27
					0, 17, 5, -3, 35, 20, 11, 19, -26,
					-- layer=2 filter=95 channel=28
					-10, 10, 10, -21, 19, 28, 13, 27, -50,
					-- layer=2 filter=95 channel=29
					10, -8, -4, -4, 1, 5, 4, -3, 5,
					-- layer=2 filter=95 channel=30
					-9, -11, -1, -22, -18, -22, 10, 9, -13,
					-- layer=2 filter=95 channel=31
					-18, 2, -48, -55, -45, -67, -15, -55, -96,
					-- layer=2 filter=95 channel=32
					2, 1, 10, 7, 10, -1, 11, -1, -7,
					-- layer=2 filter=95 channel=33
					-11, 27, -7, 23, 48, 16, 30, 25, 8,
					-- layer=2 filter=95 channel=34
					-17, -45, 8, 4, 0, 9, 0, 25, 10,
					-- layer=2 filter=95 channel=35
					9, 11, -23, 6, 76, 70, -2, 36, -13,
					-- layer=2 filter=95 channel=36
					8, 4, 6, -1, -2, -11, 10, -5, 8,
					-- layer=2 filter=95 channel=37
					25, 5, 13, 12, 4, 0, 30, 3, -4,
					-- layer=2 filter=95 channel=38
					0, -27, 6, -11, 21, 0, 20, 22, -1,
					-- layer=2 filter=95 channel=39
					4, -14, -16, 35, 31, -6, 34, -3, 0,
					-- layer=2 filter=95 channel=40
					-64, -48, 3, -1, -11, -51, -16, -25, -14,
					-- layer=2 filter=95 channel=41
					5, 5, -11, -7, -2, 9, -2, 3, 2,
					-- layer=2 filter=95 channel=42
					1, -16, -7, 17, 54, 29, 11, 14, 47,
					-- layer=2 filter=95 channel=43
					22, 33, -49, 25, 39, -33, 14, 32, -41,
					-- layer=2 filter=95 channel=44
					-5, 3, 0, -2, 5, 7, 0, 3, -2,
					-- layer=2 filter=95 channel=45
					-16, -13, -55, -49, -4, -6, 6, 5, -53,
					-- layer=2 filter=95 channel=46
					-12, 8, 4, 4, 3, -10, -11, -6, -47,
					-- layer=2 filter=95 channel=47
					-31, 10, -11, 25, -11, -17, 6, 14, -22,
					-- layer=2 filter=95 channel=48
					4, 0, 9, -8, -7, 0, 4, -4, 3,
					-- layer=2 filter=95 channel=49
					-9, -30, 8, -31, -48, 30, 7, -2, 97,
					-- layer=2 filter=95 channel=50
					-10, -1, 13, -6, -11, 0, -4, -8, 36,
					-- layer=2 filter=95 channel=51
					11, -23, -11, -20, -29, -19, 0, 1, -14,
					-- layer=2 filter=95 channel=52
					19, 14, 74, 20, -17, 38, 30, -16, 49,
					-- layer=2 filter=95 channel=53
					24, -32, -11, 22, -30, -20, -22, 16, 46,
					-- layer=2 filter=95 channel=54
					-16, 24, 10, 9, 20, 8, 0, -16, 25,
					-- layer=2 filter=95 channel=55
					0, 2, -10, 2, 0, 5, 8, 6, 4,
					-- layer=2 filter=95 channel=56
					1, -2, -32, -2, -3, -13, 19, -7, -22,
					-- layer=2 filter=95 channel=57
					-6, 6, -2, 7, 7, -8, 2, 4, 2,
					-- layer=2 filter=95 channel=58
					5, 24, 10, 24, 23, 23, 40, 26, -24,
					-- layer=2 filter=95 channel=59
					4, 7, 34, 35, 34, 23, 34, 5, 17,
					-- layer=2 filter=95 channel=60
					0, -21, 3, -11, -42, 23, 11, 2, 62,
					-- layer=2 filter=95 channel=61
					-60, -76, 15, -13, -111, 15, -27, -90, 60,
					-- layer=2 filter=95 channel=62
					-15, -56, 12, -17, -95, 28, 39, -16, 51,
					-- layer=2 filter=95 channel=63
					-3, -4, -22, 36, -9, -27, 31, -7, -6,
					-- layer=2 filter=95 channel=64
					5, 9, -7, 20, 16, 8, 17, 27, 21,
					-- layer=2 filter=95 channel=65
					-17, -87, -23, -54, -143, 16, -45, -69, 67,
					-- layer=2 filter=95 channel=66
					0, 20, 16, 39, -9, 31, 7, -56, -9,
					-- layer=2 filter=95 channel=67
					-19, -10, 0, 3, 12, -17, -8, -5, -63,
					-- layer=2 filter=95 channel=68
					5, 10, 10, 6, 10, 0, 8, 0, 6,
					-- layer=2 filter=95 channel=69
					7, -30, -8, -6, 18, -10, 20, 18, 39,
					-- layer=2 filter=95 channel=70
					3, 16, 2, 11, 44, 27, 0, 12, -22,
					-- layer=2 filter=95 channel=71
					-14, 5, -20, 1, 24, 6, 8, 23, -10,
					-- layer=2 filter=95 channel=72
					8, -8, 9, -18, 4, 25, 21, 9, 35,
					-- layer=2 filter=95 channel=73
					58, 52, 65, 31, 32, 23, 68, -1, -31,
					-- layer=2 filter=95 channel=74
					0, -13, 10, 25, 28, 8, 22, 0, -39,
					-- layer=2 filter=95 channel=75
					-1, -2, -6, -17, -18, 4, 17, 3, -6,
					-- layer=2 filter=95 channel=76
					16, 16, 24, -38, -12, -13, -19, -58, -10,
					-- layer=2 filter=95 channel=77
					1, -4, -5, 2, 2, 6, 2, 8, -11,
					-- layer=2 filter=95 channel=78
					-24, -7, -52, -1, -27, -32, 5, -17, -3,
					-- layer=2 filter=95 channel=79
					5, -7, -7, 7, 5, -6, -3, 8, -3,
					-- layer=2 filter=95 channel=80
					11, 0, 6, 9, 21, -10, 0, 21, -10,
					-- layer=2 filter=95 channel=81
					8, 5, 10, 0, 0, 4, -1, 17, 19,
					-- layer=2 filter=95 channel=82
					-1, 8, 0, 3, -7, 3, 3, -9, 9,
					-- layer=2 filter=95 channel=83
					6, -17, -5, -5, 4, 38, -15, -7, -11,
					-- layer=2 filter=95 channel=84
					-2, -2, 3, 8, -4, 5, -1, -7, 5,
					-- layer=2 filter=95 channel=85
					-4, 5, -1, -9, 14, 8, 17, 3, -7,
					-- layer=2 filter=95 channel=86
					-1, -9, 17, 1, 7, 11, 5, 0, 3,
					-- layer=2 filter=95 channel=87
					-24, -68, 55, -17, -43, 60, -4, 27, 75,
					-- layer=2 filter=95 channel=88
					-15, -19, -3, -5, 2, -5, 0, 0, -3,
					-- layer=2 filter=95 channel=89
					-10, -21, 14, -16, 8, 20, 17, 5, -5,
					-- layer=2 filter=95 channel=90
					-9, -6, -8, 2, 3, -6, -5, 0, 2,
					-- layer=2 filter=95 channel=91
					32, 32, 7, -16, 12, 27, 20, 40, 11,
					-- layer=2 filter=95 channel=92
					0, 17, 5, 0, 4, 17, 3, 19, 22,
					-- layer=2 filter=95 channel=93
					45, 56, -6, -18, -77, 25, 39, -8, 0,
					-- layer=2 filter=95 channel=94
					-64, -134, -14, -20, -133, -39, -8, -78, 46,
					-- layer=2 filter=95 channel=95
					8, 16, 10, -2, 9, -1, 9, 0, 11,
					-- layer=2 filter=95 channel=96
					-41, -84, -59, 37, -180, -55, -13, -43, 29,
					-- layer=2 filter=95 channel=97
					-10, 21, 9, 11, 53, -12, -8, 26, -41,
					-- layer=2 filter=95 channel=98
					-16, 6, 19, 0, -2, 15, 10, 18, -20,
					-- layer=2 filter=95 channel=99
					1, 7, 49, 18, -36, 28, 23, 2, 60,
					-- layer=2 filter=95 channel=100
					27, 29, 3, 4, 58, 18, -8, 35, -35,
					-- layer=2 filter=95 channel=101
					8, 42, 1, 0, 6, -9, -18, 35, 21,
					-- layer=2 filter=95 channel=102
					-47, -77, -17, 16, -103, 2, -3, -65, 55,
					-- layer=2 filter=95 channel=103
					-14, -19, -38, -17, -30, -30, -30, -30, -20,
					-- layer=2 filter=95 channel=104
					11, -42, -2, -31, -93, 17, -16, -72, 40,
					-- layer=2 filter=95 channel=105
					-19, 25, 73, -17, 0, 13, 33, -18, -37,
					-- layer=2 filter=95 channel=106
					-1, 12, -3, 13, 0, 12, 27, 35, -1,
					-- layer=2 filter=95 channel=107
					-32, 1, -12, 39, 17, 9, -10, -16, 33,
					-- layer=2 filter=95 channel=108
					-12, -23, -28, 19, -15, -6, 6, -27, -22,
					-- layer=2 filter=95 channel=109
					3, 10, 5, 12, 4, -6, 18, 8, 13,
					-- layer=2 filter=95 channel=110
					2, 27, -20, -2, 3, 1, -10, 15, 8,
					-- layer=2 filter=95 channel=111
					-1, -5, -5, -7, 1, 4, -6, -11, -2,
					-- layer=2 filter=95 channel=112
					-13, 28, 22, 16, 38, -4, -18, -37, 16,
					-- layer=2 filter=95 channel=113
					-13, -2, -11, -43, -17, -9, -7, 25, -19,
					-- layer=2 filter=95 channel=114
					3, 5, -5, 10, -5, -4, -14, -3, -2,
					-- layer=2 filter=95 channel=115
					2, 8, 2, -5, 13, -11, 1, -3, 4,
					-- layer=2 filter=95 channel=116
					11, -48, 51, 0, -7, 43, -8, 21, 59,
					-- layer=2 filter=95 channel=117
					-32, 26, 3, -78, -35, 4, -7, -60, -2,
					-- layer=2 filter=95 channel=118
					31, 25, 4, 33, 7, -12, -5, 27, -31,
					-- layer=2 filter=95 channel=119
					-43, 3, -3, 5, -1, 25, -5, 14, 3,
					-- layer=2 filter=95 channel=120
					-6, 7, -2, 0, 4, -7, -2, 4, -9,
					-- layer=2 filter=95 channel=121
					2, 5, -4, -8, 10, 2, -9, -4, 7,
					-- layer=2 filter=95 channel=122
					-7, 0, -1, 0, -15, 0, -4, -3, 3,
					-- layer=2 filter=95 channel=123
					1, 16, 0, 14, 1, 5, 3, -18, 10,
					-- layer=2 filter=95 channel=124
					-48, 3, -19, -19, 29, 11, 15, -5, 2,
					-- layer=2 filter=95 channel=125
					11, -3, 3, 10, 7, -1, -3, 5, 9,
					-- layer=2 filter=95 channel=126
					16, 11, -9, 70, -62, -29, 26, 64, 0,
					-- layer=2 filter=95 channel=127
					-3, 8, 2, -19, -22, -20, -14, -20, -23,
					-- layer=2 filter=96 channel=0
					-17, -14, -23, -18, -1, -11, -6, 2, -6,
					-- layer=2 filter=96 channel=1
					-18, -1, 1, -9, -12, -17, -2, -9, -6,
					-- layer=2 filter=96 channel=2
					-1, -7, -9, 0, 6, 3, 3, -6, 5,
					-- layer=2 filter=96 channel=3
					6, -5, 4, 16, 2, 8, -5, 9, 0,
					-- layer=2 filter=96 channel=4
					-8, -27, -25, 0, -19, -9, -2, -17, -8,
					-- layer=2 filter=96 channel=5
					-12, -15, -5, -23, -5, -22, -17, -17, -9,
					-- layer=2 filter=96 channel=6
					-18, 3, 4, -9, -8, -4, -18, -9, -14,
					-- layer=2 filter=96 channel=7
					-8, -14, 7, 2, 0, 1, 3, 4, -10,
					-- layer=2 filter=96 channel=8
					2, 0, -11, 0, -8, -6, 1, -4, -9,
					-- layer=2 filter=96 channel=9
					3, 3, -6, -4, 1, 10, -16, -1, 13,
					-- layer=2 filter=96 channel=10
					-16, -18, -5, -8, -10, -14, -25, 0, 0,
					-- layer=2 filter=96 channel=11
					-20, -13, -11, -22, -15, -4, -2, -10, -5,
					-- layer=2 filter=96 channel=12
					7, -1, -3, 4, 6, -18, -7, -6, -10,
					-- layer=2 filter=96 channel=13
					4, -3, -4, -9, 6, -6, -5, 2, 3,
					-- layer=2 filter=96 channel=14
					3, 2, 7, 3, 0, -19, -13, -12, -13,
					-- layer=2 filter=96 channel=15
					-13, -14, -10, 0, -12, 6, -7, -24, -1,
					-- layer=2 filter=96 channel=16
					-4, -8, 12, -12, 2, 1, -16, -16, -14,
					-- layer=2 filter=96 channel=17
					-3, -4, -10, -4, -7, -1, -9, -8, 2,
					-- layer=2 filter=96 channel=18
					-2, -15, -24, 5, -11, -9, 6, -8, -4,
					-- layer=2 filter=96 channel=19
					-10, -19, -7, -4, -5, -3, -3, -18, -19,
					-- layer=2 filter=96 channel=20
					8, 8, -3, 0, -2, -4, -11, -5, 5,
					-- layer=2 filter=96 channel=21
					-2, 0, -6, -4, 11, 1, 5, 4, -9,
					-- layer=2 filter=96 channel=22
					-4, 6, 2, 9, 0, 7, 4, 0, 12,
					-- layer=2 filter=96 channel=23
					-17, -13, -17, -21, -12, -12, -4, -5, -21,
					-- layer=2 filter=96 channel=24
					-3, 2, 10, 0, 5, 0, 0, 7, 6,
					-- layer=2 filter=96 channel=25
					-9, 3, 5, 8, 7, 6, 0, 10, 0,
					-- layer=2 filter=96 channel=26
					0, 9, 1, -1, -7, 4, 8, 0, -4,
					-- layer=2 filter=96 channel=27
					-13, 1, -8, -13, -10, -3, -2, -13, -5,
					-- layer=2 filter=96 channel=28
					-15, -9, -17, -15, -13, 13, -26, -11, -14,
					-- layer=2 filter=96 channel=29
					-4, 1, -1, 6, -2, -3, -6, 7, 0,
					-- layer=2 filter=96 channel=30
					-6, -2, -30, -15, -30, -16, -16, -13, 11,
					-- layer=2 filter=96 channel=31
					7, -15, 6, -4, -12, -2, -14, -32, -6,
					-- layer=2 filter=96 channel=32
					-2, -8, -2, -5, 2, 11, -1, 7, 6,
					-- layer=2 filter=96 channel=33
					-16, -16, 5, 17, 8, 6, -6, 0, 0,
					-- layer=2 filter=96 channel=34
					-10, -10, -15, 0, -1, 2, -23, 6, -3,
					-- layer=2 filter=96 channel=35
					-10, -18, -33, -9, -10, -3, -13, -15, -13,
					-- layer=2 filter=96 channel=36
					8, 3, -8, -8, 7, -5, -2, -8, -2,
					-- layer=2 filter=96 channel=37
					-23, -19, -8, -10, -12, 4, -4, -13, -8,
					-- layer=2 filter=96 channel=38
					-2, 4, -5, -10, -14, -21, -1, -20, -15,
					-- layer=2 filter=96 channel=39
					-7, -11, 0, -8, 1, 2, -4, 10, -4,
					-- layer=2 filter=96 channel=40
					-16, -20, -18, -2, -15, 15, -11, -1, 3,
					-- layer=2 filter=96 channel=41
					1, -3, 3, 7, 6, 8, 6, -3, 3,
					-- layer=2 filter=96 channel=42
					-12, -25, -7, -2, -10, -23, -16, -5, 2,
					-- layer=2 filter=96 channel=43
					-9, -25, -21, -7, -19, 3, -18, 6, 3,
					-- layer=2 filter=96 channel=44
					-7, 9, -2, 1, -4, -1, 6, 9, -9,
					-- layer=2 filter=96 channel=45
					-28, -17, -14, -11, -1, 5, 2, -4, 4,
					-- layer=2 filter=96 channel=46
					0, -18, -7, -13, -9, -2, -20, -25, -10,
					-- layer=2 filter=96 channel=47
					-22, -8, -10, -7, 3, 0, -8, -1, -12,
					-- layer=2 filter=96 channel=48
					6, -11, 0, -8, -3, -2, -7, -5, 0,
					-- layer=2 filter=96 channel=49
					3, -25, -6, 7, -9, -12, 1, -4, 6,
					-- layer=2 filter=96 channel=50
					-3, -1, 4, -9, 0, 4, 11, 1, -8,
					-- layer=2 filter=96 channel=51
					-6, -7, -6, -10, -20, -1, 0, -9, -16,
					-- layer=2 filter=96 channel=52
					0, 0, -26, -1, -2, -1, -14, -3, -20,
					-- layer=2 filter=96 channel=53
					4, -8, -5, -14, -21, -3, 3, -5, -10,
					-- layer=2 filter=96 channel=54
					-10, -16, -8, -19, -12, 2, 5, -3, 0,
					-- layer=2 filter=96 channel=55
					0, 1, 6, -7, 7, 7, -4, -7, -7,
					-- layer=2 filter=96 channel=56
					-14, -12, -8, -20, -17, -15, 0, -10, -16,
					-- layer=2 filter=96 channel=57
					7, 3, 6, -4, -9, 4, -10, -1, 2,
					-- layer=2 filter=96 channel=58
					-6, -7, -12, -16, -5, -8, 11, 4, -10,
					-- layer=2 filter=96 channel=59
					-20, -3, 10, -13, 8, -11, 6, -3, -8,
					-- layer=2 filter=96 channel=60
					-6, -3, 3, -10, -13, -23, -14, -15, -26,
					-- layer=2 filter=96 channel=61
					-5, 14, -14, -21, -8, -13, -16, 7, -24,
					-- layer=2 filter=96 channel=62
					-7, 0, -17, -21, -12, -17, -17, 6, -16,
					-- layer=2 filter=96 channel=63
					-14, -2, 1, -9, -7, -14, -7, -7, -46,
					-- layer=2 filter=96 channel=64
					-11, -17, -16, -14, -21, -20, 2, -18, -1,
					-- layer=2 filter=96 channel=65
					-11, 3, -1, -22, 7, -14, -4, -14, -24,
					-- layer=2 filter=96 channel=66
					-11, -3, -3, 3, 3, 2, -10, -8, -1,
					-- layer=2 filter=96 channel=67
					-10, 6, -10, -1, -13, -7, -10, -13, 10,
					-- layer=2 filter=96 channel=68
					0, 7, 4, -5, 8, 6, -1, -2, 3,
					-- layer=2 filter=96 channel=69
					-4, 4, -11, 1, -10, -19, -11, -14, -7,
					-- layer=2 filter=96 channel=70
					-4, -20, -23, -13, -14, 7, -17, -24, -25,
					-- layer=2 filter=96 channel=71
					0, -6, -4, -10, -4, 11, 1, 0, -14,
					-- layer=2 filter=96 channel=72
					-3, -4, 0, 5, 7, 5, -8, -3, -20,
					-- layer=2 filter=96 channel=73
					-6, -2, -9, -2, -20, -11, -3, 2, 2,
					-- layer=2 filter=96 channel=74
					-10, 0, -1, -24, -3, -5, -13, -16, -2,
					-- layer=2 filter=96 channel=75
					0, 6, -11, 4, 7, 1, -8, -10, -7,
					-- layer=2 filter=96 channel=76
					7, -12, -2, 2, 8, -6, 4, -11, -3,
					-- layer=2 filter=96 channel=77
					-11, -11, 2, 5, -3, 9, -5, -11, -2,
					-- layer=2 filter=96 channel=78
					-14, -24, -21, -6, -5, -1, 0, 1, -12,
					-- layer=2 filter=96 channel=79
					-1, 7, 5, 4, -8, 6, -11, 0, 0,
					-- layer=2 filter=96 channel=80
					3, -6, 0, -19, -13, -11, -17, -12, 1,
					-- layer=2 filter=96 channel=81
					8, 5, 8, 7, -11, 5, -2, -5, 1,
					-- layer=2 filter=96 channel=82
					0, 0, -9, -3, 0, 3, -6, 8, -5,
					-- layer=2 filter=96 channel=83
					-7, -29, -21, -8, -13, -3, -22, -26, -5,
					-- layer=2 filter=96 channel=84
					-10, 8, 8, -2, 2, 1, -8, -10, -2,
					-- layer=2 filter=96 channel=85
					-7, -6, -5, 11, 9, -3, -10, 6, 7,
					-- layer=2 filter=96 channel=86
					8, 0, 0, -3, 7, 6, 9, 7, 4,
					-- layer=2 filter=96 channel=87
					-6, -5, -37, 3, -8, 0, -5, -1, -6,
					-- layer=2 filter=96 channel=88
					-5, 6, -26, -2, -13, -21, -16, -17, -13,
					-- layer=2 filter=96 channel=89
					-11, -5, 2, -3, 4, -11, 9, -12, -8,
					-- layer=2 filter=96 channel=90
					0, 7, -6, -5, -4, 4, 5, -3, -8,
					-- layer=2 filter=96 channel=91
					-7, 0, 9, 9, 0, -1, -6, -3, -15,
					-- layer=2 filter=96 channel=92
					-14, 0, -1, 3, 7, -9, 5, 2, 1,
					-- layer=2 filter=96 channel=93
					-11, -2, -8, -18, 15, -1, -32, 12, -2,
					-- layer=2 filter=96 channel=94
					-11, 3, -9, -21, -17, -8, -23, 8, -31,
					-- layer=2 filter=96 channel=95
					2, -4, -7, -7, -10, -6, 8, 1, 4,
					-- layer=2 filter=96 channel=96
					-8, 0, -5, -9, -16, -35, 2, -3, -12,
					-- layer=2 filter=96 channel=97
					5, -7, 8, 5, 0, -4, 0, -4, 12,
					-- layer=2 filter=96 channel=98
					-8, -14, -6, -7, 1, 0, -4, -10, -15,
					-- layer=2 filter=96 channel=99
					-5, -10, -8, -17, 1, 4, -13, -2, -11,
					-- layer=2 filter=96 channel=100
					-5, -22, 0, -27, -19, -32, -29, -25, -18,
					-- layer=2 filter=96 channel=101
					9, 3, -2, 4, 1, 6, 10, 6, 1,
					-- layer=2 filter=96 channel=102
					-5, -12, -6, 13, -17, -14, 5, -26, -9,
					-- layer=2 filter=96 channel=103
					1, -10, 3, 1, 0, 0, -8, 5, 1,
					-- layer=2 filter=96 channel=104
					8, -33, -13, -7, -9, 1, 7, 4, -6,
					-- layer=2 filter=96 channel=105
					-17, -17, -19, 3, -3, 12, -7, -4, -7,
					-- layer=2 filter=96 channel=106
					4, 6, 13, 5, 5, -2, 0, 10, 1,
					-- layer=2 filter=96 channel=107
					0, -1, 9, 0, 8, -9, 6, -10, -5,
					-- layer=2 filter=96 channel=108
					4, -5, -9, -2, -16, -6, 9, -4, 1,
					-- layer=2 filter=96 channel=109
					0, 0, -9, 2, 4, 3, 7, -2, -6,
					-- layer=2 filter=96 channel=110
					-10, -3, -15, 0, -1, -13, 4, -11, -3,
					-- layer=2 filter=96 channel=111
					-3, 4, -3, 7, -9, -8, 9, 0, 0,
					-- layer=2 filter=96 channel=112
					-17, -13, -18, -1, -4, -7, 3, -5, -15,
					-- layer=2 filter=96 channel=113
					-8, 0, -17, -10, -12, -11, -1, -39, 0,
					-- layer=2 filter=96 channel=114
					-8, 12, -5, -8, -8, 1, 1, 0, 6,
					-- layer=2 filter=96 channel=115
					-2, -7, 4, -4, 6, 4, -1, -4, 5,
					-- layer=2 filter=96 channel=116
					0, -10, -16, -4, -2, 16, -17, -5, -8,
					-- layer=2 filter=96 channel=117
					-19, -26, -22, -3, -5, -9, -14, 2, -3,
					-- layer=2 filter=96 channel=118
					-8, -18, -6, -22, -26, -14, -23, -19, -5,
					-- layer=2 filter=96 channel=119
					-20, -32, -9, -13, -21, -6, 2, -1, -7,
					-- layer=2 filter=96 channel=120
					-1, -5, 4, -7, 4, -1, -2, 2, -2,
					-- layer=2 filter=96 channel=121
					-4, -1, 5, -1, 0, 3, -6, 7, 5,
					-- layer=2 filter=96 channel=122
					6, -3, -8, 8, -6, -1, 7, 4, 5,
					-- layer=2 filter=96 channel=123
					-20, -18, -5, -2, 9, -1, -10, -1, -12,
					-- layer=2 filter=96 channel=124
					-12, -10, -10, -13, -25, -4, 7, -10, 1,
					-- layer=2 filter=96 channel=125
					-3, 0, 2, 5, -9, -2, -6, 7, 7,
					-- layer=2 filter=96 channel=126
					-6, -4, -17, -14, 9, -5, -6, 7, -21,
					-- layer=2 filter=96 channel=127
					-17, -7, -21, -15, -16, -27, -15, -22, 1,
					-- layer=2 filter=97 channel=0
					-19, -8, -9, 1, 6, -12, -12, -3, -8,
					-- layer=2 filter=97 channel=1
					-15, -20, -8, -12, -8, -11, 2, -9, -11,
					-- layer=2 filter=97 channel=2
					-9, -10, 3, -4, -1, -7, 7, -8, 6,
					-- layer=2 filter=97 channel=3
					-3, 2, -10, 0, -14, 4, -4, 0, 3,
					-- layer=2 filter=97 channel=4
					7, -7, -10, -9, 0, -1, -2, -8, -1,
					-- layer=2 filter=97 channel=5
					1, -7, 4, 7, -9, -10, -6, 2, 4,
					-- layer=2 filter=97 channel=6
					-3, 10, -3, -6, 0, -3, 10, -1, -12,
					-- layer=2 filter=97 channel=7
					2, -4, -1, 2, -5, -10, -11, 12, -7,
					-- layer=2 filter=97 channel=8
					1, -3, -8, -3, -3, -5, -2, 6, -5,
					-- layer=2 filter=97 channel=9
					-10, -17, -13, -6, -5, -1, -15, -10, 2,
					-- layer=2 filter=97 channel=10
					-15, -5, 4, -4, 3, 5, 0, -15, -1,
					-- layer=2 filter=97 channel=11
					-5, -13, 4, -10, -6, -5, 3, 0, -3,
					-- layer=2 filter=97 channel=12
					-9, -22, -7, 0, -1, -6, -12, -10, -19,
					-- layer=2 filter=97 channel=13
					-7, 0, 1, 8, -11, 5, -4, -7, 10,
					-- layer=2 filter=97 channel=14
					-7, -2, -1, 1, 0, -15, -17, 1, 0,
					-- layer=2 filter=97 channel=15
					-2, -7, 4, -13, -11, -13, -2, 6, -8,
					-- layer=2 filter=97 channel=16
					-3, -8, 2, -12, -8, 1, 3, -6, -5,
					-- layer=2 filter=97 channel=17
					10, -5, 9, -1, 8, -9, -9, 10, 9,
					-- layer=2 filter=97 channel=18
					4, -9, -6, 10, -3, -12, 9, 8, -3,
					-- layer=2 filter=97 channel=19
					1, -7, 6, -7, -1, -20, 10, -5, -3,
					-- layer=2 filter=97 channel=20
					-7, 3, 8, 3, 9, 0, -7, -10, -3,
					-- layer=2 filter=97 channel=21
					10, -2, -7, 5, 7, 8, -7, -2, 9,
					-- layer=2 filter=97 channel=22
					0, 0, 5, 8, 3, -1, 4, 7, 11,
					-- layer=2 filter=97 channel=23
					-9, -6, -10, -18, -15, 0, -9, -6, -5,
					-- layer=2 filter=97 channel=24
					-4, -14, -22, -11, -7, 6, 9, -5, 5,
					-- layer=2 filter=97 channel=25
					-8, -7, -4, -5, -3, -4, -7, -11, -9,
					-- layer=2 filter=97 channel=26
					10, -5, -8, 0, 6, -6, -1, 0, -5,
					-- layer=2 filter=97 channel=27
					-5, -1, -16, 0, -5, 2, -14, -6, -14,
					-- layer=2 filter=97 channel=28
					-3, 14, -1, -6, 3, 6, -4, -4, -19,
					-- layer=2 filter=97 channel=29
					2, -4, 6, -9, -2, -4, 8, -2, -11,
					-- layer=2 filter=97 channel=30
					2, 2, -6, -19, -6, -7, -7, -17, 0,
					-- layer=2 filter=97 channel=31
					8, 5, 0, -9, -8, 4, -9, 0, -10,
					-- layer=2 filter=97 channel=32
					-7, 5, -7, -10, -1, -5, 1, 5, -4,
					-- layer=2 filter=97 channel=33
					-8, -3, -4, 0, -1, -7, 2, -2, -12,
					-- layer=2 filter=97 channel=34
					-5, 0, -4, -9, 3, -5, 2, 3, 5,
					-- layer=2 filter=97 channel=35
					-7, 5, -8, -7, 0, -14, -15, -14, -17,
					-- layer=2 filter=97 channel=36
					-3, 3, -8, 8, -10, -11, -10, 7, 1,
					-- layer=2 filter=97 channel=37
					-9, -15, -11, -9, -11, 3, -11, -13, -6,
					-- layer=2 filter=97 channel=38
					-3, -3, -14, -20, 5, -9, -14, 0, 3,
					-- layer=2 filter=97 channel=39
					1, -14, -6, 0, 1, -9, 2, 1, -11,
					-- layer=2 filter=97 channel=40
					6, 6, 10, -6, 8, -6, -8, 3, 12,
					-- layer=2 filter=97 channel=41
					8, -2, -4, 10, 7, -7, 7, -8, 3,
					-- layer=2 filter=97 channel=42
					0, -16, -16, -4, 0, 0, -1, 0, -12,
					-- layer=2 filter=97 channel=43
					2, -13, -16, 10, 6, -6, -17, 4, 0,
					-- layer=2 filter=97 channel=44
					6, 7, -1, 2, -4, 8, -8, 0, 10,
					-- layer=2 filter=97 channel=45
					-4, 6, -5, -9, 4, 8, -6, 3, 6,
					-- layer=2 filter=97 channel=46
					-1, -11, -12, -21, -7, -2, 0, -9, -3,
					-- layer=2 filter=97 channel=47
					1, 6, 1, 3, -12, 6, -18, -12, -13,
					-- layer=2 filter=97 channel=48
					-9, -11, -4, 0, 0, -4, -7, -8, -7,
					-- layer=2 filter=97 channel=49
					8, -4, -3, 11, -14, -11, -1, -6, -5,
					-- layer=2 filter=97 channel=50
					-9, 0, 2, -5, 10, -8, 10, 5, -11,
					-- layer=2 filter=97 channel=51
					6, -8, -4, 2, -4, -11, 5, -13, -17,
					-- layer=2 filter=97 channel=52
					1, -9, 2, 2, -17, -8, 7, -11, -18,
					-- layer=2 filter=97 channel=53
					5, 0, 5, -14, 0, 5, 0, -9, -3,
					-- layer=2 filter=97 channel=54
					-10, 10, -5, 0, 0, -17, -11, -4, -15,
					-- layer=2 filter=97 channel=55
					7, 9, -4, -9, 7, -2, -3, 0, -6,
					-- layer=2 filter=97 channel=56
					3, -3, -14, 7, 0, 0, 2, -10, -3,
					-- layer=2 filter=97 channel=57
					-1, 6, -9, 0, 0, 1, 6, -5, -4,
					-- layer=2 filter=97 channel=58
					-16, -21, -14, -12, -8, -15, -3, -16, -16,
					-- layer=2 filter=97 channel=59
					-4, 3, -6, -6, -12, -15, 3, -12, -5,
					-- layer=2 filter=97 channel=60
					-9, -15, 2, 2, 4, -1, 7, -13, 2,
					-- layer=2 filter=97 channel=61
					0, 0, 8, -4, 10, -13, 0, -5, 0,
					-- layer=2 filter=97 channel=62
					-1, 1, -1, 2, -13, -13, 1, 7, -1,
					-- layer=2 filter=97 channel=63
					-3, -4, -15, -11, -14, 3, -7, -11, -7,
					-- layer=2 filter=97 channel=64
					-13, 4, 0, -1, -1, -2, -2, -1, 1,
					-- layer=2 filter=97 channel=65
					0, -7, -4, 0, -5, 2, 3, 0, -3,
					-- layer=2 filter=97 channel=66
					0, -2, 5, -6, -3, -1, 4, -1, 6,
					-- layer=2 filter=97 channel=67
					-13, -4, -7, -5, -1, -7, -6, -11, -12,
					-- layer=2 filter=97 channel=68
					2, -10, 0, -5, 7, -3, 2, -3, 1,
					-- layer=2 filter=97 channel=69
					-7, -11, -9, -4, -13, -6, -6, -6, -6,
					-- layer=2 filter=97 channel=70
					7, 14, -11, -5, -13, -3, -14, -17, -2,
					-- layer=2 filter=97 channel=71
					0, -10, -11, 9, 3, -10, 2, -2, -11,
					-- layer=2 filter=97 channel=72
					-6, -1, 0, -7, -7, -5, 1, 8, 2,
					-- layer=2 filter=97 channel=73
					11, 1, -2, 7, 3, 7, 4, -4, 9,
					-- layer=2 filter=97 channel=74
					0, -4, -2, -8, 4, 4, 3, -5, -10,
					-- layer=2 filter=97 channel=75
					4, 8, -9, 0, 2, 5, 8, 3, -1,
					-- layer=2 filter=97 channel=76
					10, -1, 3, -1, -8, -9, 13, 2, 5,
					-- layer=2 filter=97 channel=77
					-5, -8, 8, -4, 11, 1, 3, -1, -3,
					-- layer=2 filter=97 channel=78
					-13, -12, 0, -9, 0, -4, 7, -12, -9,
					-- layer=2 filter=97 channel=79
					-9, 5, 10, -2, 8, -10, 0, 2, -1,
					-- layer=2 filter=97 channel=80
					-17, -13, -13, -11, -10, -12, -9, -2, -10,
					-- layer=2 filter=97 channel=81
					-10, -8, -6, -11, 0, -7, 4, 1, -2,
					-- layer=2 filter=97 channel=82
					-7, 7, 11, 0, 6, 0, 0, -6, 7,
					-- layer=2 filter=97 channel=83
					-12, -7, -19, -21, -2, -3, -17, 1, -12,
					-- layer=2 filter=97 channel=84
					-4, 6, -2, 1, -3, 2, -9, 3, 8,
					-- layer=2 filter=97 channel=85
					-8, -10, -3, -5, -10, 0, -1, 1, 7,
					-- layer=2 filter=97 channel=86
					11, 3, 0, 5, 7, 6, -7, -2, 0,
					-- layer=2 filter=97 channel=87
					9, 8, -8, 9, -16, 8, 1, 0, -1,
					-- layer=2 filter=97 channel=88
					-11, -17, -1, -5, -12, -5, -12, -3, -6,
					-- layer=2 filter=97 channel=89
					-8, -2, -13, -15, 5, -15, -2, -14, -9,
					-- layer=2 filter=97 channel=90
					-7, -7, 0, 1, -7, -4, -10, -1, 4,
					-- layer=2 filter=97 channel=91
					-14, -3, -9, -4, -9, -5, -15, 4, -12,
					-- layer=2 filter=97 channel=92
					-9, -4, -5, -9, -3, -13, -3, -9, -10,
					-- layer=2 filter=97 channel=93
					-8, -5, 5, 5, 0, -1, 0, 6, 5,
					-- layer=2 filter=97 channel=94
					-4, -8, -9, -5, -1, -8, -6, 9, -4,
					-- layer=2 filter=97 channel=95
					1, 10, -8, -1, 0, -3, -2, -3, -8,
					-- layer=2 filter=97 channel=96
					2, 9, -3, 8, -2, 6, -5, -8, 4,
					-- layer=2 filter=97 channel=97
					3, -16, -3, -6, 2, -9, -3, -12, -9,
					-- layer=2 filter=97 channel=98
					-11, 10, -4, 2, -11, -9, 0, -3, -13,
					-- layer=2 filter=97 channel=99
					4, 0, 0, -14, 5, -8, -4, 3, -12,
					-- layer=2 filter=97 channel=100
					-16, -14, -7, -12, -1, 2, -14, -20, -9,
					-- layer=2 filter=97 channel=101
					-11, -9, -3, -12, -4, 7, -11, 0, 0,
					-- layer=2 filter=97 channel=102
					-5, -8, -10, 12, -13, -10, 9, -5, -7,
					-- layer=2 filter=97 channel=103
					-10, -3, -7, 7, -2, -7, -9, 4, 1,
					-- layer=2 filter=97 channel=104
					-5, -7, -1, 8, 2, 4, 10, 1, 0,
					-- layer=2 filter=97 channel=105
					-17, 0, 7, -2, -12, 2, -2, 0, 1,
					-- layer=2 filter=97 channel=106
					8, 1, -13, -14, 11, 0, 3, -6, 8,
					-- layer=2 filter=97 channel=107
					-4, 6, -1, 8, 1, 5, 6, -3, -5,
					-- layer=2 filter=97 channel=108
					-3, -9, -11, 4, -17, -5, -2, -4, -10,
					-- layer=2 filter=97 channel=109
					2, -2, 0, 10, -3, -11, -11, -8, 1,
					-- layer=2 filter=97 channel=110
					-10, -7, -8, -7, -13, -10, 4, 8, -7,
					-- layer=2 filter=97 channel=111
					-4, 4, -9, -8, -6, 3, 9, 0, 12,
					-- layer=2 filter=97 channel=112
					-16, -2, -1, -2, 0, -9, 0, -3, -8,
					-- layer=2 filter=97 channel=113
					-2, -17, -9, -16, -13, -2, -14, -11, 5,
					-- layer=2 filter=97 channel=114
					-4, 8, -9, -7, 8, 4, -3, 3, 0,
					-- layer=2 filter=97 channel=115
					10, 7, 9, -9, 8, 0, -3, -5, 8,
					-- layer=2 filter=97 channel=116
					-1, 4, -16, 3, -20, 5, -9, -6, -12,
					-- layer=2 filter=97 channel=117
					-5, -9, 6, 7, -10, -10, -10, 16, 5,
					-- layer=2 filter=97 channel=118
					-3, 2, 1, -9, -2, 0, -14, -9, -3,
					-- layer=2 filter=97 channel=119
					-5, -4, -1, -9, 4, -8, 0, -4, -13,
					-- layer=2 filter=97 channel=120
					-7, -7, 5, -4, 0, 5, 6, -3, 7,
					-- layer=2 filter=97 channel=121
					9, -8, -11, -12, -11, -8, -4, 9, 6,
					-- layer=2 filter=97 channel=122
					-9, 9, -2, -6, -8, 1, -9, -2, 10,
					-- layer=2 filter=97 channel=123
					-13, 6, -11, -5, -16, -2, 0, -3, -12,
					-- layer=2 filter=97 channel=124
					1, 9, 0, 3, -7, -9, 12, 10, 7,
					-- layer=2 filter=97 channel=125
					-2, 3, 3, 1, 2, 0, -1, 5, 9,
					-- layer=2 filter=97 channel=126
					-4, -3, -7, -12, -7, 2, -3, 3, -9,
					-- layer=2 filter=97 channel=127
					5, -1, -2, -1, 0, -3, -2, -7, 8,
					-- layer=2 filter=98 channel=0
					-23, 1, 7, 9, 4, -5, -14, -21, 0,
					-- layer=2 filter=98 channel=1
					1, 2, -25, 5, -39, -17, -6, -19, -65,
					-- layer=2 filter=98 channel=2
					1, -1, 5, 8, -1, 10, -4, 2, 0,
					-- layer=2 filter=98 channel=3
					-22, -12, 36, -21, 24, 12, -8, 21, 6,
					-- layer=2 filter=98 channel=4
					18, -14, -19, -4, 0, -16, -27, -44, -42,
					-- layer=2 filter=98 channel=5
					0, 12, 19, -18, -7, 0, -15, 12, 9,
					-- layer=2 filter=98 channel=6
					-15, -24, -35, 27, -11, 17, 11, 15, 39,
					-- layer=2 filter=98 channel=7
					33, -23, 48, 30, 14, -4, -11, -48, -21,
					-- layer=2 filter=98 channel=8
					4, -6, 1, -9, -8, 4, -7, -5, -2,
					-- layer=2 filter=98 channel=9
					3, -1, -29, 30, 3, -26, 65, 3, -7,
					-- layer=2 filter=98 channel=10
					-7, 4, 5, -4, -16, 3, -15, 0, -7,
					-- layer=2 filter=98 channel=11
					-7, -6, 3, -37, -1, 10, -13, 17, 3,
					-- layer=2 filter=98 channel=12
					12, -11, -25, 0, -49, -38, -10, -33, -16,
					-- layer=2 filter=98 channel=13
					9, 5, 8, 7, 8, -1, 5, 0, 10,
					-- layer=2 filter=98 channel=14
					2, -11, -25, -36, -39, -32, -4, -12, -33,
					-- layer=2 filter=98 channel=15
					-51, 25, 3, 15, -3, 59, 33, 20, -7,
					-- layer=2 filter=98 channel=16
					45, -21, -15, 77, -2, -74, 62, -31, -58,
					-- layer=2 filter=98 channel=17
					-1, -9, -2, 0, 9, -4, 11, 9, 8,
					-- layer=2 filter=98 channel=18
					5, 1, 13, -1, 0, 19, 3, -10, -6,
					-- layer=2 filter=98 channel=19
					19, -8, -22, 39, 12, 18, 8, -15, -66,
					-- layer=2 filter=98 channel=20
					2, 11, -2, 8, 3, -3, 6, 7, 11,
					-- layer=2 filter=98 channel=21
					-6, -7, -17, 4, -6, -21, 0, 4, -3,
					-- layer=2 filter=98 channel=22
					4, 2, -4, 12, 0, -5, 7, -1, 2,
					-- layer=2 filter=98 channel=23
					45, 10, -50, 44, 20, -33, 53, 0, -16,
					-- layer=2 filter=98 channel=24
					-20, -9, -9, -26, -16, 10, 2, -1, 41,
					-- layer=2 filter=98 channel=25
					-37, -23, -14, -37, -27, 27, -17, 7, 61,
					-- layer=2 filter=98 channel=26
					8, -4, 5, 2, 9, 6, -2, 7, 11,
					-- layer=2 filter=98 channel=27
					24, 17, 1, 16, 11, 12, 1, -9, -15,
					-- layer=2 filter=98 channel=28
					7, -1, 5, 50, 6, -2, 9, -27, -55,
					-- layer=2 filter=98 channel=29
					10, 3, -2, 5, 5, -10, 6, -9, -2,
					-- layer=2 filter=98 channel=30
					-6, 3, -52, 54, 12, -11, 34, -3, -41,
					-- layer=2 filter=98 channel=31
					-77, 20, -22, -56, -6, 13, 10, 0, 0,
					-- layer=2 filter=98 channel=32
					7, 5, 0, 0, 2, -4, 1, -5, -6,
					-- layer=2 filter=98 channel=33
					50, 16, 26, 8, 6, -18, 41, 61, -17,
					-- layer=2 filter=98 channel=34
					-26, -20, 5, 36, 27, 40, 45, 9, 1,
					-- layer=2 filter=98 channel=35
					-14, 0, 16, 41, 0, 16, 11, -20, -23,
					-- layer=2 filter=98 channel=36
					5, 6, -7, 6, -7, -3, -13, -10, 2,
					-- layer=2 filter=98 channel=37
					-1, 1, 9, -18, 4, 27, -5, 13, -5,
					-- layer=2 filter=98 channel=38
					19, 7, -13, 22, -29, 0, 0, -27, -5,
					-- layer=2 filter=98 channel=39
					42, 4, -6, 57, -5, -68, 48, -18, -67,
					-- layer=2 filter=98 channel=40
					-35, -30, 12, -26, -13, 69, 0, 8, 3,
					-- layer=2 filter=98 channel=41
					4, -4, -7, 9, -6, 8, -7, 10, -4,
					-- layer=2 filter=98 channel=42
					49, -11, -17, 65, -25, -60, 38, 27, -39,
					-- layer=2 filter=98 channel=43
					-30, -25, 29, -31, -19, 36, -25, 1, -6,
					-- layer=2 filter=98 channel=44
					-6, 2, 7, -4, 3, -3, -4, -9, -5,
					-- layer=2 filter=98 channel=45
					-76, -14, 25, -24, -5, 7, -4, -30, -25,
					-- layer=2 filter=98 channel=46
					-8, -11, -37, -2, -37, -5, -28, -56, -29,
					-- layer=2 filter=98 channel=47
					-17, -70, 23, 34, -1, 19, 20, 1, -45,
					-- layer=2 filter=98 channel=48
					-5, -7, 3, -5, -2, -7, 5, 0, 0,
					-- layer=2 filter=98 channel=49
					-2, -22, 18, -22, 7, 4, 25, 4, -5,
					-- layer=2 filter=98 channel=50
					13, -17, 1, -5, 7, 7, 2, -1, 0,
					-- layer=2 filter=98 channel=51
					-13, -22, -2, -19, 15, 27, -7, 10, 20,
					-- layer=2 filter=98 channel=52
					-44, -28, 0, -13, 9, -8, -2, 15, -40,
					-- layer=2 filter=98 channel=53
					-14, -15, -33, 40, -14, 7, 1, -5, -35,
					-- layer=2 filter=98 channel=54
					-17, -48, -39, 0, 1, 25, -15, 11, -2,
					-- layer=2 filter=98 channel=55
					-4, 10, -4, 4, 14, 7, 1, -10, 5,
					-- layer=2 filter=98 channel=56
					5, 3, 3, -30, 0, 20, -6, 11, 4,
					-- layer=2 filter=98 channel=57
					-4, 0, -1, 0, -2, 13, -13, 0, 0,
					-- layer=2 filter=98 channel=58
					25, -6, -32, 10, -54, -71, -16, -33, -22,
					-- layer=2 filter=98 channel=59
					28, 13, 18, 10, 12, -31, -5, -34, -60,
					-- layer=2 filter=98 channel=60
					20, -3, -23, -7, -36, -4, -51, -39, -29,
					-- layer=2 filter=98 channel=61
					-11, 44, 18, 6, 11, -4, 0, -26, 0,
					-- layer=2 filter=98 channel=62
					-17, -52, -28, 6, -17, 14, 2, 4, 33,
					-- layer=2 filter=98 channel=63
					12, 2, -25, 11, -14, -71, 16, -12, -79,
					-- layer=2 filter=98 channel=64
					38, 2, -49, 40, -4, -22, 67, 7, -6,
					-- layer=2 filter=98 channel=65
					6, 12, -13, 18, 6, 18, 22, -7, 30,
					-- layer=2 filter=98 channel=66
					-28, 19, 62, 4, -24, -9, -15, -10, 4,
					-- layer=2 filter=98 channel=67
					-3, 13, -13, 59, 7, 8, 50, 41, 0,
					-- layer=2 filter=98 channel=68
					5, 5, -3, -5, 7, -4, -5, 3, -7,
					-- layer=2 filter=98 channel=69
					19, -25, -40, 45, -17, -61, 50, 5, -38,
					-- layer=2 filter=98 channel=70
					-6, -7, -4, 21, -9, 11, -8, -20, -20,
					-- layer=2 filter=98 channel=71
					-21, -25, -20, 18, -4, 19, 4, 5, 28,
					-- layer=2 filter=98 channel=72
					71, 23, 8, -8, -15, -15, -30, -42, -88,
					-- layer=2 filter=98 channel=73
					1, -2, 12, -16, -5, 24, -22, -25, -18,
					-- layer=2 filter=98 channel=74
					15, 9, -41, 0, 6, -37, 10, 14, -99,
					-- layer=2 filter=98 channel=75
					18, 3, -46, -28, -42, -42, -14, -50, 1,
					-- layer=2 filter=98 channel=76
					-23, 9, 4, -24, 53, 62, 34, -11, 42,
					-- layer=2 filter=98 channel=77
					1, 0, -10, 4, -7, -2, 1, -3, -6,
					-- layer=2 filter=98 channel=78
					-40, -21, 0, -27, -5, 12, -7, 18, 36,
					-- layer=2 filter=98 channel=79
					-3, 7, 5, 6, -3, 2, 0, 2, -7,
					-- layer=2 filter=98 channel=80
					27, -55, -69, 16, -19, -81, 0, -25, -36,
					-- layer=2 filter=98 channel=81
					-9, 8, 6, 13, 0, 5, 8, 12, -9,
					-- layer=2 filter=98 channel=82
					1, 8, -5, -4, 2, -10, -6, -5, -3,
					-- layer=2 filter=98 channel=83
					48, -13, -58, 47, 8, -60, 44, -2, -24,
					-- layer=2 filter=98 channel=84
					9, -2, 0, -2, 8, -7, 9, -1, 2,
					-- layer=2 filter=98 channel=85
					-4, -15, -8, 3, -4, 14, 5, 8, -9,
					-- layer=2 filter=98 channel=86
					17, 11, 1, -1, 23, -3, -2, -1, 10,
					-- layer=2 filter=98 channel=87
					-7, 11, -15, 39, 23, 19, -54, -5, 3,
					-- layer=2 filter=98 channel=88
					6, 4, -10, 25, -11, -2, 31, 42, -39,
					-- layer=2 filter=98 channel=89
					12, -4, -15, -38, -35, -73, -23, -19, -54,
					-- layer=2 filter=98 channel=90
					-4, -9, 0, -6, -1, 0, 2, -5, 8,
					-- layer=2 filter=98 channel=91
					36, -8, -22, 37, -29, -81, 37, -18, -16,
					-- layer=2 filter=98 channel=92
					39, -17, 4, 10, -27, -18, 16, -41, -35,
					-- layer=2 filter=98 channel=93
					25, 7, 0, 58, 40, 23, 7, 39, 21,
					-- layer=2 filter=98 channel=94
					-5, 32, -19, 39, 10, 17, -13, -7, -17,
					-- layer=2 filter=98 channel=95
					-2, 11, -3, -1, -9, -2, 2, 12, 6,
					-- layer=2 filter=98 channel=96
					-12, -6, -17, 15, 47, 42, 21, 60, 18,
					-- layer=2 filter=98 channel=97
					10, -6, -16, -8, -38, -33, 1, 4, -8,
					-- layer=2 filter=98 channel=98
					-28, -39, 24, 33, 10, 27, -13, -14, -36,
					-- layer=2 filter=98 channel=99
					-22, -7, 11, 24, 16, 11, 30, -8, -15,
					-- layer=2 filter=98 channel=100
					38, 39, -48, 27, -31, -56, 0, -63, -56,
					-- layer=2 filter=98 channel=101
					-29, -48, -40, -50, -47, 14, -47, -20, 38,
					-- layer=2 filter=98 channel=102
					10, -12, -19, -4, -13, 40, 50, 39, 33,
					-- layer=2 filter=98 channel=103
					-27, -21, -24, -25, 29, 49, 48, 39, 22,
					-- layer=2 filter=98 channel=104
					-14, 9, 5, 5, 39, 23, -9, 25, 7,
					-- layer=2 filter=98 channel=105
					-64, -8, -11, 10, -13, 26, -12, -18, 0,
					-- layer=2 filter=98 channel=106
					7, 25, -12, -19, -31, 19, -25, -8, 25,
					-- layer=2 filter=98 channel=107
					-10, 2, 4, 28, 36, 44, 24, 24, -23,
					-- layer=2 filter=98 channel=108
					-5, 24, -6, -10, -5, -7, 37, -6, 7,
					-- layer=2 filter=98 channel=109
					-15, 8, 2, -1, -10, 5, -4, 11, 0,
					-- layer=2 filter=98 channel=110
					38, -18, -45, 39, -5, -23, 25, -3, -29,
					-- layer=2 filter=98 channel=111
					0, 4, -7, 2, -8, -6, 1, 7, 2,
					-- layer=2 filter=98 channel=112
					2, 21, 9, -1, 0, 13, 2, 3, 21,
					-- layer=2 filter=98 channel=113
					-5, -25, -14, 31, -17, -58, -6, -40, -42,
					-- layer=2 filter=98 channel=114
					-19, -5, -4, 7, 5, 0, -6, -15, -18,
					-- layer=2 filter=98 channel=115
					7, 5, -1, -5, 6, 9, 7, 5, 2,
					-- layer=2 filter=98 channel=116
					13, 22, 6, 23, 17, 22, -12, 30, -17,
					-- layer=2 filter=98 channel=117
					-10, -10, -7, 8, 22, 0, -42, -40, -31,
					-- layer=2 filter=98 channel=118
					-21, -33, 9, -31, 14, 37, -31, 24, 0,
					-- layer=2 filter=98 channel=119
					24, -32, -32, 57, -50, -29, 45, -55, -13,
					-- layer=2 filter=98 channel=120
					-1, -4, 4, 1, -6, 3, 0, 2, 1,
					-- layer=2 filter=98 channel=121
					7, 1, -5, -2, -7, -8, -7, 9, -1,
					-- layer=2 filter=98 channel=122
					12, 2, 10, -1, 9, -5, 14, 18, -8,
					-- layer=2 filter=98 channel=123
					20, 10, 45, 41, 3, 34, 1, -43, -55,
					-- layer=2 filter=98 channel=124
					-13, 9, -4, 22, 17, 6, 26, 2, -52,
					-- layer=2 filter=98 channel=125
					10, 7, 0, 0, -10, -4, 6, -12, 0,
					-- layer=2 filter=98 channel=126
					-20, -8, -28, 5, 7, 11, -16, -33, -1,
					-- layer=2 filter=98 channel=127
					4, 18, -49, 24, -24, -39, 0, -25, -44,
					-- layer=2 filter=99 channel=0
					-11, 8, -4, 2, 8, -18, -6, 12, -20,
					-- layer=2 filter=99 channel=1
					-36, -22, -3, -7, -3, 9, 5, -23, -16,
					-- layer=2 filter=99 channel=2
					5, 8, -5, 7, 1, 0, 2, -6, -2,
					-- layer=2 filter=99 channel=3
					-22, -9, -10, 5, -6, -22, 6, 0, -4,
					-- layer=2 filter=99 channel=4
					-7, -18, -1, -19, -27, -18, -15, -32, 0,
					-- layer=2 filter=99 channel=5
					-21, 18, 4, 12, 4, -14, 22, -6, -6,
					-- layer=2 filter=99 channel=6
					-17, 9, -9, -30, 13, -17, 11, 20, -8,
					-- layer=2 filter=99 channel=7
					22, 1, -27, 2, 11, 4, -23, -7, -3,
					-- layer=2 filter=99 channel=8
					9, 3, 6, -2, 0, -5, -3, 7, 2,
					-- layer=2 filter=99 channel=9
					-9, 2, 5, 15, -11, 13, 31, 7, -5,
					-- layer=2 filter=99 channel=10
					14, 3, -6, 10, 19, -10, -7, -5, -7,
					-- layer=2 filter=99 channel=11
					-10, -26, -13, -5, -20, -26, -9, -8, -11,
					-- layer=2 filter=99 channel=12
					-28, -22, -9, -16, -10, 12, 6, -15, -32,
					-- layer=2 filter=99 channel=13
					-1, 5, -3, 3, -7, -4, -12, -6, -6,
					-- layer=2 filter=99 channel=14
					-35, -22, -29, -18, -4, -6, 12, -5, -19,
					-- layer=2 filter=99 channel=15
					-7, -6, -16, -27, -14, 0, -2, -11, 2,
					-- layer=2 filter=99 channel=16
					-8, 5, -7, 9, 5, -35, -20, -15, -3,
					-- layer=2 filter=99 channel=17
					5, 2, -5, -3, -9, 0, -9, -4, -2,
					-- layer=2 filter=99 channel=18
					-18, -6, 6, -14, -33, 0, 0, -42, 6,
					-- layer=2 filter=99 channel=19
					9, -9, 0, -10, -17, 14, -23, -10, 7,
					-- layer=2 filter=99 channel=20
					-5, 8, -5, -10, -6, 9, 5, 0, -7,
					-- layer=2 filter=99 channel=21
					-10, 3, 0, -12, 0, -5, 8, -12, 1,
					-- layer=2 filter=99 channel=22
					-9, 4, -8, 0, 4, -1, 9, 1, -4,
					-- layer=2 filter=99 channel=23
					-6, -39, 5, -2, -20, -1, -21, -1, -21,
					-- layer=2 filter=99 channel=24
					-11, -7, -5, -1, 0, -2, -20, 18, 3,
					-- layer=2 filter=99 channel=25
					4, 0, -7, -12, 1, 7, -17, 3, -9,
					-- layer=2 filter=99 channel=26
					-2, -1, 4, -10, 0, -7, 0, -9, 8,
					-- layer=2 filter=99 channel=27
					-15, -8, 0, -22, 8, 4, -2, -8, -12,
					-- layer=2 filter=99 channel=28
					14, -32, -13, 19, -20, -4, -19, -18, -16,
					-- layer=2 filter=99 channel=29
					-9, 6, 3, -2, -6, 6, 9, 7, -5,
					-- layer=2 filter=99 channel=30
					-13, -18, 9, -7, -10, -5, -7, 5, 3,
					-- layer=2 filter=99 channel=31
					3, 18, 16, -24, 8, -22, -34, -18, 6,
					-- layer=2 filter=99 channel=32
					4, -9, -8, 0, 1, -9, -1, 5, 4,
					-- layer=2 filter=99 channel=33
					11, -6, -36, -25, -17, -13, -20, -15, -7,
					-- layer=2 filter=99 channel=34
					32, -21, 10, 2, -28, -7, 15, 0, 5,
					-- layer=2 filter=99 channel=35
					30, -3, -22, 9, -21, -20, -4, -24, -9,
					-- layer=2 filter=99 channel=36
					-10, 6, 4, -9, 2, -3, -4, -5, 2,
					-- layer=2 filter=99 channel=37
					-6, 0, 0, -13, -3, -5, 2, -2, 5,
					-- layer=2 filter=99 channel=38
					-26, 2, 0, 0, 7, -15, -6, -2, -20,
					-- layer=2 filter=99 channel=39
					-8, -9, -20, -24, 20, -15, -7, -19, 14,
					-- layer=2 filter=99 channel=40
					7, -32, 0, -34, -21, 5, -36, -47, 34,
					-- layer=2 filter=99 channel=41
					8, -5, 0, 4, 7, -11, -2, 10, 3,
					-- layer=2 filter=99 channel=42
					-1, -2, -9, 6, 4, -3, -2, -28, -21,
					-- layer=2 filter=99 channel=43
					0, 8, 0, 5, -17, -3, -9, -7, -2,
					-- layer=2 filter=99 channel=44
					-7, -1, 9, 7, -10, -4, 10, -3, -3,
					-- layer=2 filter=99 channel=45
					3, 17, 16, 7, 3, -21, -10, -12, -10,
					-- layer=2 filter=99 channel=46
					4, 0, -4, -2, -4, -26, -8, 16, -26,
					-- layer=2 filter=99 channel=47
					13, -18, -21, 13, -27, -4, -36, -13, -33,
					-- layer=2 filter=99 channel=48
					3, 0, -6, 5, 4, 8, 2, 7, 1,
					-- layer=2 filter=99 channel=49
					-36, 15, 10, -17, -11, 16, -13, -7, 12,
					-- layer=2 filter=99 channel=50
					6, 0, 0, -10, -6, -6, -9, 1, 9,
					-- layer=2 filter=99 channel=51
					-11, -4, -11, 0, -12, -17, 1, -8, -5,
					-- layer=2 filter=99 channel=52
					9, -2, -11, -3, -13, 11, -5, 4, 2,
					-- layer=2 filter=99 channel=53
					14, -8, -18, -25, 36, -24, 0, -12, 28,
					-- layer=2 filter=99 channel=54
					-1, 9, -4, 5, -9, 3, -9, -12, 2,
					-- layer=2 filter=99 channel=55
					5, -1, 10, -1, 7, -7, 2, 0, 4,
					-- layer=2 filter=99 channel=56
					-27, -8, -3, -21, -20, -19, 12, -22, -23,
					-- layer=2 filter=99 channel=57
					-7, 2, -8, 1, -3, 3, 5, 6, 0,
					-- layer=2 filter=99 channel=58
					-33, -37, -2, -17, -19, 8, 10, -10, -20,
					-- layer=2 filter=99 channel=59
					-35, -10, -1, -17, -19, -15, 4, 13, 16,
					-- layer=2 filter=99 channel=60
					-22, 16, -12, 0, 32, 10, 13, 28, -1,
					-- layer=2 filter=99 channel=61
					-17, 25, 4, 15, 45, -18, 5, 40, 9,
					-- layer=2 filter=99 channel=62
					-25, -5, -20, -32, -2, -10, 4, 20, -13,
					-- layer=2 filter=99 channel=63
					-15, 7, -6, 9, 16, -14, -25, 17, -5,
					-- layer=2 filter=99 channel=64
					-19, -15, 14, -11, -22, 5, 6, -5, 1,
					-- layer=2 filter=99 channel=65
					-39, -5, -24, 1, 15, -20, -2, 23, -27,
					-- layer=2 filter=99 channel=66
					-34, 35, 1, -1, -25, 14, 3, 6, -24,
					-- layer=2 filter=99 channel=67
					-3, 6, 8, -17, -4, 1, -16, 6, -11,
					-- layer=2 filter=99 channel=68
					7, 8, -11, -8, -7, 8, -7, 0, -1,
					-- layer=2 filter=99 channel=69
					-49, -21, 12, -46, -13, 6, -19, -12, -17,
					-- layer=2 filter=99 channel=70
					17, -10, -8, 12, -3, -19, -6, -14, -11,
					-- layer=2 filter=99 channel=71
					-13, -7, 1, -22, 0, -8, -5, -17, -1,
					-- layer=2 filter=99 channel=72
					39, -5, -15, -1, 14, 3, 0, -3, -15,
					-- layer=2 filter=99 channel=73
					27, 11, 24, 3, 50, -11, -18, 31, 21,
					-- layer=2 filter=99 channel=74
					-3, -6, -8, 12, -1, -11, -23, -10, 5,
					-- layer=2 filter=99 channel=75
					-11, -33, -41, -16, -29, -58, 0, -3, 18,
					-- layer=2 filter=99 channel=76
					-4, -27, -10, -3, 22, -17, -19, 23, 11,
					-- layer=2 filter=99 channel=77
					-6, 0, -10, -7, -9, -9, 7, -6, -9,
					-- layer=2 filter=99 channel=78
					-16, 0, -5, 5, -34, 3, -21, -6, -8,
					-- layer=2 filter=99 channel=79
					7, 4, 3, -7, 0, 0, 0, 6, 9,
					-- layer=2 filter=99 channel=80
					-16, -1, -17, -1, 1, -41, 3, -25, -17,
					-- layer=2 filter=99 channel=81
					-9, -10, 5, 9, 2, 7, -5, -2, 0,
					-- layer=2 filter=99 channel=82
					11, -11, -2, -6, -4, -1, 7, 2, -2,
					-- layer=2 filter=99 channel=83
					-24, -26, -6, -11, -49, -16, -4, -17, -15,
					-- layer=2 filter=99 channel=84
					-7, 9, 5, 2, 0, -5, -8, -5, -5,
					-- layer=2 filter=99 channel=85
					1, -9, 0, 3, 8, -4, -7, -6, -2,
					-- layer=2 filter=99 channel=86
					-6, 3, -10, -4, -2, -11, 1, 2, -2,
					-- layer=2 filter=99 channel=87
					1, -2, -17, -34, -7, 5, -20, -25, 9,
					-- layer=2 filter=99 channel=88
					-43, -19, -18, -18, 18, -10, -23, -2, -9,
					-- layer=2 filter=99 channel=89
					-16, -22, -33, -31, -24, 6, 14, -11, -8,
					-- layer=2 filter=99 channel=90
					8, 1, -3, 5, -3, 10, 0, -2, 1,
					-- layer=2 filter=99 channel=91
					-4, -12, -13, 0, -5, 24, -6, -15, 13,
					-- layer=2 filter=99 channel=92
					-33, -10, -17, -12, -31, 15, 14, -21, -30,
					-- layer=2 filter=99 channel=93
					2, 21, -9, -27, -15, -24, -8, 22, 1,
					-- layer=2 filter=99 channel=94
					-14, 9, -21, -2, 23, -2, 3, 44, 2,
					-- layer=2 filter=99 channel=95
					-12, -3, -6, -7, -8, 8, -5, -7, -11,
					-- layer=2 filter=99 channel=96
					5, -38, 8, -4, -8, 16, 11, -10, 14,
					-- layer=2 filter=99 channel=97
					-39, -28, -20, -20, -13, -14, -2, -2, -7,
					-- layer=2 filter=99 channel=98
					41, 0, -9, 23, -9, 1, -37, 5, -12,
					-- layer=2 filter=99 channel=99
					-1, -10, 12, 27, 5, 22, -20, 21, -8,
					-- layer=2 filter=99 channel=100
					-19, 8, -10, -14, -16, -5, -1, -28, -28,
					-- layer=2 filter=99 channel=101
					-20, 3, -4, -25, -3, 7, -8, -3, 2,
					-- layer=2 filter=99 channel=102
					-18, -28, 15, -16, -21, 22, 16, -21, 24,
					-- layer=2 filter=99 channel=103
					-11, 8, -7, -8, 5, 30, -4, -4, 0,
					-- layer=2 filter=99 channel=104
					-24, 9, -8, -5, -16, 11, 2, 7, 19,
					-- layer=2 filter=99 channel=105
					-3, -18, -5, 3, -7, -13, 10, -1, 4,
					-- layer=2 filter=99 channel=106
					-10, -4, -19, -13, -14, -18, -47, -28, -6,
					-- layer=2 filter=99 channel=107
					19, 30, -8, -18, 25, -5, 24, -8, 7,
					-- layer=2 filter=99 channel=108
					-3, -22, -14, -15, -19, 7, 13, -22, 4,
					-- layer=2 filter=99 channel=109
					-7, 0, 6, -8, -7, 9, -8, 2, -9,
					-- layer=2 filter=99 channel=110
					7, 14, 11, 2, -9, 13, 17, 0, -11,
					-- layer=2 filter=99 channel=111
					3, -8, 3, -9, -1, 1, -2, 7, -2,
					-- layer=2 filter=99 channel=112
					-5, 0, -11, 3, 18, -15, 4, 45, 8,
					-- layer=2 filter=99 channel=113
					-27, -3, 14, 12, 10, 0, -16, 16, 0,
					-- layer=2 filter=99 channel=114
					3, 14, 6, -7, 8, 7, -6, 0, -2,
					-- layer=2 filter=99 channel=115
					9, 3, 2, 3, 2, 8, 1, 7, -6,
					-- layer=2 filter=99 channel=116
					9, -21, 7, -16, -39, 3, -20, -26, 7,
					-- layer=2 filter=99 channel=117
					35, 14, -19, 21, 34, 16, -15, 4, -5,
					-- layer=2 filter=99 channel=118
					2, -12, -11, -19, -10, -11, -1, -21, 5,
					-- layer=2 filter=99 channel=119
					-31, -32, 11, -7, -32, -14, -9, -30, -4,
					-- layer=2 filter=99 channel=120
					-1, -4, 7, -9, -10, -7, 4, -2, 6,
					-- layer=2 filter=99 channel=121
					-7, 6, 6, 0, -1, -5, -2, 6, -6,
					-- layer=2 filter=99 channel=122
					0, -8, -4, -4, -8, 0, 10, 1, 10,
					-- layer=2 filter=99 channel=123
					4, -16, -7, 7, -2, 18, -33, -4, 5,
					-- layer=2 filter=99 channel=124
					-2, -2, -29, -46, 1, 27, -30, -39, -16,
					-- layer=2 filter=99 channel=125
					0, 10, -7, -1, 3, 9, -3, -7, 3,
					-- layer=2 filter=99 channel=126
					6, -8, 7, -4, 32, -17, -2, 19, 8,
					-- layer=2 filter=99 channel=127
					-39, -19, 10, 3, -18, 4, -22, -4, 3,
					-- layer=2 filter=100 channel=0
					10, -29, -6, 9, -32, 1, 1, 12, 9,
					-- layer=2 filter=100 channel=1
					23, 25, -9, -17, -1, 7, -10, 0, -13,
					-- layer=2 filter=100 channel=2
					0, -2, 7, 8, -10, -1, -6, 1, 7,
					-- layer=2 filter=100 channel=3
					-43, -48, 33, 21, -10, 12, 22, 39, 36,
					-- layer=2 filter=100 channel=4
					-7, 4, 12, -3, 35, 8, -30, -4, 19,
					-- layer=2 filter=100 channel=5
					5, -1, -4, -3, -31, -15, 19, -13, 39,
					-- layer=2 filter=100 channel=6
					55, 14, -8, 55, 39, 32, 24, 3, -17,
					-- layer=2 filter=100 channel=7
					-7, -59, 2, 38, 23, 4, -30, 7, 18,
					-- layer=2 filter=100 channel=8
					4, 8, 2, 5, -4, -7, -1, -1, -3,
					-- layer=2 filter=100 channel=9
					-27, -19, -27, -13, -71, 20, 46, 8, -14,
					-- layer=2 filter=100 channel=10
					-23, -40, -4, -2, -11, 3, 27, 14, 14,
					-- layer=2 filter=100 channel=11
					27, 16, -2, 0, -13, 2, -1, -11, 5,
					-- layer=2 filter=100 channel=12
					16, 23, 11, -47, 0, 21, -6, -27, -4,
					-- layer=2 filter=100 channel=13
					0, -5, -11, 10, -1, -3, 8, 3, -7,
					-- layer=2 filter=100 channel=14
					48, 27, 10, -52, -14, 20, -20, -41, -6,
					-- layer=2 filter=100 channel=15
					-26, -25, -14, -61, -34, 0, -19, -89, -32,
					-- layer=2 filter=100 channel=16
					-18, 21, 10, 7, 20, -29, -3, -19, -24,
					-- layer=2 filter=100 channel=17
					6, 0, 1, 3, -8, 2, -9, -8, 0,
					-- layer=2 filter=100 channel=18
					18, 42, 26, -43, 3, 6, -5, -49, -8,
					-- layer=2 filter=100 channel=19
					6, -18, -26, 6, 0, -33, -13, -9, -28,
					-- layer=2 filter=100 channel=20
					-6, -5, 0, -8, 5, 8, -9, 6, -5,
					-- layer=2 filter=100 channel=21
					-3, -10, 5, 4, -6, -11, 18, 2, 11,
					-- layer=2 filter=100 channel=22
					-2, 10, 8, -3, 3, -8, 8, -9, 5,
					-- layer=2 filter=100 channel=23
					-41, 12, -9, 23, 29, 1, -23, 20, 8,
					-- layer=2 filter=100 channel=24
					22, 8, 32, 21, -18, 16, 14, -11, 9,
					-- layer=2 filter=100 channel=25
					15, 5, 36, -11, -21, -2, 11, 6, 42,
					-- layer=2 filter=100 channel=26
					0, 2, 8, 1, -5, 5, -11, 0, 6,
					-- layer=2 filter=100 channel=27
					7, -27, -11, 50, 7, 2, 29, 27, 3,
					-- layer=2 filter=100 channel=28
					-2, -31, 10, -10, -3, -32, 5, 34, 38,
					-- layer=2 filter=100 channel=29
					-4, 3, 0, 0, 0, 8, 5, -11, 5,
					-- layer=2 filter=100 channel=30
					-28, -9, -25, -9, 7, -6, 0, -9, -4,
					-- layer=2 filter=100 channel=31
					46, -93, -93, -14, -37, -11, -5, 23, 46,
					-- layer=2 filter=100 channel=32
					9, 5, -7, 1, -4, -3, 7, -5, 10,
					-- layer=2 filter=100 channel=33
					-3, -52, 12, 3, 0, 25, -14, -34, 42,
					-- layer=2 filter=100 channel=34
					7, 4, -26, -26, 5, 14, 40, 0, -43,
					-- layer=2 filter=100 channel=35
					9, -55, -5, 6, -31, -19, -19, -13, 19,
					-- layer=2 filter=100 channel=36
					3, 0, 3, -14, 10, -8, 6, 1, -8,
					-- layer=2 filter=100 channel=37
					22, 19, 11, -5, 0, 4, 15, -1, 9,
					-- layer=2 filter=100 channel=38
					35, -18, 17, -3, -10, -19, 19, 2, 6,
					-- layer=2 filter=100 channel=39
					-23, 5, -17, 24, 14, -27, -7, 0, -23,
					-- layer=2 filter=100 channel=40
					1, -46, -50, 10, 20, 5, 12, -78, -19,
					-- layer=2 filter=100 channel=41
					-1, 7, -2, -7, 6, -4, -6, -4, 9,
					-- layer=2 filter=100 channel=42
					-6, 28, 11, 4, 12, 9, -7, -7, -6,
					-- layer=2 filter=100 channel=43
					-51, -31, -7, 2, -40, 21, 36, 59, 12,
					-- layer=2 filter=100 channel=44
					6, 0, -3, -6, -5, 10, 0, -2, 11,
					-- layer=2 filter=100 channel=45
					32, -37, 2, 24, 29, 17, -31, -13, -31,
					-- layer=2 filter=100 channel=46
					-20, -13, -20, -2, -2, -25, 11, -16, -9,
					-- layer=2 filter=100 channel=47
					-18, -23, 9, -11, 6, 23, 11, 8, 12,
					-- layer=2 filter=100 channel=48
					-10, 11, 4, 0, -1, 3, 5, 7, 9,
					-- layer=2 filter=100 channel=49
					32, 44, 24, -28, -9, 21, 20, -71, -28,
					-- layer=2 filter=100 channel=50
					-19, 0, 0, -24, -14, -31, -4, 1, 0,
					-- layer=2 filter=100 channel=51
					20, -7, -27, -6, -7, -2, 16, 3, 11,
					-- layer=2 filter=100 channel=52
					1, 2, -25, -6, 44, 7, 31, 30, 28,
					-- layer=2 filter=100 channel=53
					10, -3, 39, -10, -18, 54, -28, -84, -28,
					-- layer=2 filter=100 channel=54
					11, 14, -20, 4, 5, 13, -15, 8, 7,
					-- layer=2 filter=100 channel=55
					-5, -7, -4, -7, 1, -5, -8, 4, -16,
					-- layer=2 filter=100 channel=56
					15, 8, 7, 4, -16, -15, 9, 27, -2,
					-- layer=2 filter=100 channel=57
					-2, -12, -3, -1, -9, 20, -13, 4, 7,
					-- layer=2 filter=100 channel=58
					20, 34, 19, -13, -33, 41, 19, -13, -19,
					-- layer=2 filter=100 channel=59
					1, 18, 44, 12, -30, -8, -26, 21, -41,
					-- layer=2 filter=100 channel=60
					14, 18, -33, -19, 21, -39, -14, -22, 20,
					-- layer=2 filter=100 channel=61
					1, 31, -24, 26, 0, -36, -33, -31, -16,
					-- layer=2 filter=100 channel=62
					20, 31, -6, 12, 44, 23, 1, -35, -27,
					-- layer=2 filter=100 channel=63
					-21, -16, -1, -1, -7, -14, -32, 7, -18,
					-- layer=2 filter=100 channel=64
					0, 7, 25, 14, 6, 26, 21, -3, -23,
					-- layer=2 filter=100 channel=65
					37, 38, -18, 49, 58, -24, 15, -3, 44,
					-- layer=2 filter=100 channel=66
					-6, 9, 17, 8, 8, -32, -23, 6, 30,
					-- layer=2 filter=100 channel=67
					-48, -10, -36, 16, -4, -5, 29, 3, -4,
					-- layer=2 filter=100 channel=68
					-2, 0, -9, -4, 0, 1, 2, 0, -10,
					-- layer=2 filter=100 channel=69
					-16, 17, 12, -5, 13, 18, 0, 4, -31,
					-- layer=2 filter=100 channel=70
					-6, -34, -10, -21, -42, -39, 14, 11, 12,
					-- layer=2 filter=100 channel=71
					7, -34, -13, 41, -2, 0, 29, -2, -20,
					-- layer=2 filter=100 channel=72
					15, 3, 39, 12, 10, -35, -41, -6, 2,
					-- layer=2 filter=100 channel=73
					-20, -21, -46, -74, -60, 29, -46, -78, -44,
					-- layer=2 filter=100 channel=74
					-22, -6, -15, 4, -35, -2, 11, 4, -25,
					-- layer=2 filter=100 channel=75
					19, 41, -9, -31, 14, -15, -10, -48, -8,
					-- layer=2 filter=100 channel=76
					-8, -12, -6, -13, -24, -4, -50, -42, -14,
					-- layer=2 filter=100 channel=77
					12, 10, 0, 3, 7, -7, 11, -6, -7,
					-- layer=2 filter=100 channel=78
					6, 44, 29, -14, 15, 19, -24, -26, 2,
					-- layer=2 filter=100 channel=79
					7, 0, -5, 11, -1, -6, -10, 2, 7,
					-- layer=2 filter=100 channel=80
					-28, -14, -29, -1, -20, 1, -12, 10, -18,
					-- layer=2 filter=100 channel=81
					-7, -12, 1, -5, -5, -9, 4, 4, 7,
					-- layer=2 filter=100 channel=82
					2, 5, 7, -5, -1, -3, -2, 6, 1,
					-- layer=2 filter=100 channel=83
					-10, 13, 20, 21, 2, 0, -3, 0, -18,
					-- layer=2 filter=100 channel=84
					-7, 6, -4, 3, 3, -3, -5, -6, -4,
					-- layer=2 filter=100 channel=85
					-5, -13, -16, -12, -6, -3, -14, 8, -5,
					-- layer=2 filter=100 channel=86
					14, 0, 3, -1, -4, -11, -15, -2, -4,
					-- layer=2 filter=100 channel=87
					13, -14, 33, -5, -9, -9, -28, -25, -2,
					-- layer=2 filter=100 channel=88
					-8, -9, 10, -4, -18, 16, 16, -6, -14,
					-- layer=2 filter=100 channel=89
					21, 3, 28, -45, -23, 18, -36, -55, -30,
					-- layer=2 filter=100 channel=90
					0, 3, 5, 8, -2, 0, 0, -6, 2,
					-- layer=2 filter=100 channel=91
					1, -10, -8, -29, -31, -6, -18, -57, 11,
					-- layer=2 filter=100 channel=92
					29, 22, 19, -22, -10, 11, -14, -21, 0,
					-- layer=2 filter=100 channel=93
					-24, 4, 2, -16, 65, 59, -10, 27, -16,
					-- layer=2 filter=100 channel=94
					16, 11, -10, 3, 39, -32, -42, 5, -49,
					-- layer=2 filter=100 channel=95
					5, 8, 4, 4, -2, 7, -5, -2, -4,
					-- layer=2 filter=100 channel=96
					-8, 57, 4, 14, 53, 18, 0, 61, 43,
					-- layer=2 filter=100 channel=97
					-6, -21, 16, -6, -44, 9, -1, -7, -16,
					-- layer=2 filter=100 channel=98
					5, -44, -1, -26, -28, -26, -18, 6, 25,
					-- layer=2 filter=100 channel=99
					-31, 12, -32, 2, 10, -5, -22, 15, -6,
					-- layer=2 filter=100 channel=100
					5, 5, 25, -7, 7, -10, 5, -23, 18,
					-- layer=2 filter=100 channel=101
					34, -55, -13, 8, -24, -32, 12, -12, -10,
					-- layer=2 filter=100 channel=102
					-27, 36, 13, -18, 20, 15, 2, 3, 26,
					-- layer=2 filter=100 channel=103
					-31, 15, -5, -24, 32, 19, 18, -40, 45,
					-- layer=2 filter=100 channel=104
					10, 26, 43, -27, 25, 34, -30, -60, 7,
					-- layer=2 filter=100 channel=105
					-18, 19, -12, 17, -35, -21, -16, 25, -12,
					-- layer=2 filter=100 channel=106
					0, -7, 7, -28, -32, -11, -1, -24, -1,
					-- layer=2 filter=100 channel=107
					-22, -29, -61, -10, -31, 46, 49, 0, 49,
					-- layer=2 filter=100 channel=108
					3, 11, -6, 1, -8, 1, 18, -5, -11,
					-- layer=2 filter=100 channel=109
					-14, -6, -14, -22, -11, -1, -11, 12, -1,
					-- layer=2 filter=100 channel=110
					17, -5, 43, 11, 23, 17, 3, 11, 19,
					-- layer=2 filter=100 channel=111
					0, -3, 7, -7, 10, 4, 12, 10, -6,
					-- layer=2 filter=100 channel=112
					11, 0, -15, 23, -22, -20, 20, -29, 9,
					-- layer=2 filter=100 channel=113
					-27, -3, 44, 6, -3, 3, 5, -18, -8,
					-- layer=2 filter=100 channel=114
					0, 1, 16, 18, 14, 15, 18, 10, 7,
					-- layer=2 filter=100 channel=115
					-7, 7, 0, 2, 6, 6, 6, -5, -1,
					-- layer=2 filter=100 channel=116
					-10, 5, 21, -18, 24, 18, 1, -19, 12,
					-- layer=2 filter=100 channel=117
					20, -51, -101, 12, 4, 1, -50, 13, -4,
					-- layer=2 filter=100 channel=118
					-13, -8, 8, 0, -18, 0, 9, 10, 19,
					-- layer=2 filter=100 channel=119
					3, 18, -7, -12, -8, -7, 8, -7, 0,
					-- layer=2 filter=100 channel=120
					-8, 3, 2, 10, -7, 9, 3, -10, 9,
					-- layer=2 filter=100 channel=121
					11, -8, 2, -6, -3, 5, 8, 9, 5,
					-- layer=2 filter=100 channel=122
					10, 9, 5, -13, 2, -4, 3, 9, 10,
					-- layer=2 filter=100 channel=123
					-3, -25, -1, -15, 36, -11, -16, -5, 27,
					-- layer=2 filter=100 channel=124
					-42, -39, -3, -17, -30, 31, -11, -37, 14,
					-- layer=2 filter=100 channel=125
					-7, -7, -12, 9, 8, 0, -2, -1, -7,
					-- layer=2 filter=100 channel=126
					-24, -34, -27, -95, -44, -5, -89, 0, -27,
					-- layer=2 filter=100 channel=127
					-8, 18, 14, -10, 0, -2, 11, 4, 5,
					-- layer=2 filter=101 channel=0
					-3, -11, 20, -18, 0, 17, -3, 19, 24,
					-- layer=2 filter=101 channel=1
					-10, -8, 16, 9, 9, -34, -2, -16, -6,
					-- layer=2 filter=101 channel=2
					-2, 9, 0, -2, 5, -6, -7, -7, -1,
					-- layer=2 filter=101 channel=3
					7, 32, 21, -18, 3, 60, -19, -41, 17,
					-- layer=2 filter=101 channel=4
					-8, 30, -24, -16, -19, -19, -13, -15, -24,
					-- layer=2 filter=101 channel=5
					-1, -5, -6, -16, -18, 3, 30, 23, 7,
					-- layer=2 filter=101 channel=6
					-49, -65, -11, 3, -5, -58, 32, 36, 21,
					-- layer=2 filter=101 channel=7
					18, -68, -19, -16, -17, -12, 25, 2, 46,
					-- layer=2 filter=101 channel=8
					7, 3, -4, -2, 3, 0, 8, -4, 0,
					-- layer=2 filter=101 channel=9
					3, 0, 14, 2, 1, 10, -33, 1, 17,
					-- layer=2 filter=101 channel=10
					-4, -4, 4, 8, -5, 33, -24, -5, 28,
					-- layer=2 filter=101 channel=11
					-10, -30, -27, -14, -23, -19, 22, 8, 22,
					-- layer=2 filter=101 channel=12
					-21, -36, 0, 22, -10, -44, -42, -46, -9,
					-- layer=2 filter=101 channel=13
					2, -8, 5, 6, 0, 2, -9, 0, 10,
					-- layer=2 filter=101 channel=14
					-18, -15, 0, 12, -5, -30, -4, -14, -1,
					-- layer=2 filter=101 channel=15
					3, -23, -56, 16, -38, 30, 25, 41, -30,
					-- layer=2 filter=101 channel=16
					-2, 1, -30, -1, -9, 9, -5, -18, -10,
					-- layer=2 filter=101 channel=17
					0, 7, 0, -2, 6, 0, 7, 8, -3,
					-- layer=2 filter=101 channel=18
					22, 51, -75, -5, 8, -51, 19, -9, -24,
					-- layer=2 filter=101 channel=19
					-10, -16, -47, 22, 35, -1, 55, -33, -41,
					-- layer=2 filter=101 channel=20
					-7, 1, -4, 0, 3, -8, -9, 3, -8,
					-- layer=2 filter=101 channel=21
					-9, -5, 5, 15, 4, 2, -17, 0, -3,
					-- layer=2 filter=101 channel=22
					-4, 9, -8, 0, -4, -2, -6, -3, -1,
					-- layer=2 filter=101 channel=23
					-10, 4, 2, -17, 6, 8, -44, -12, 0,
					-- layer=2 filter=101 channel=24
					5, -6, 19, -34, 12, 62, -19, 0, 45,
					-- layer=2 filter=101 channel=25
					-37, -24, -11, -40, 3, 16, -31, -12, 31,
					-- layer=2 filter=101 channel=26
					4, -1, -8, 4, -6, -5, 6, -4, -1,
					-- layer=2 filter=101 channel=27
					17, 32, -7, 27, 15, -5, 14, -3, 13,
					-- layer=2 filter=101 channel=28
					-2, -8, -67, 0, -42, -13, -8, -76, -60,
					-- layer=2 filter=101 channel=29
					0, 8, 9, 2, -2, 3, -3, 4, 3,
					-- layer=2 filter=101 channel=30
					22, -7, 16, 13, 13, 23, 11, 24, -7,
					-- layer=2 filter=101 channel=31
					21, -16, -41, 36, -46, -4, 15, -22, -40,
					-- layer=2 filter=101 channel=32
					2, -2, -7, 8, -4, -5, -7, -3, 1,
					-- layer=2 filter=101 channel=33
					3, 3, 38, -20, -53, -1, -56, -23, -43,
					-- layer=2 filter=101 channel=34
					28, 24, 3, 7, 33, -37, 68, 0, -12,
					-- layer=2 filter=101 channel=35
					-26, -47, -73, -17, -9, -16, -24, -40, -13,
					-- layer=2 filter=101 channel=36
					2, -4, -6, -5, 9, 9, -3, 14, 6,
					-- layer=2 filter=101 channel=37
					-4, -5, 0, 9, 0, -9, 40, 3, 17,
					-- layer=2 filter=101 channel=38
					-28, 10, 12, -17, 26, 0, 16, -7, 7,
					-- layer=2 filter=101 channel=39
					2, 10, 28, -8, 11, 22, -11, -24, 6,
					-- layer=2 filter=101 channel=40
					40, 50, 17, -49, -32, -24, -8, -21, 14,
					-- layer=2 filter=101 channel=41
					-2, 7, -5, -3, 9, 8, 3, 2, 6,
					-- layer=2 filter=101 channel=42
					-21, 13, 26, 9, -8, 19, -47, -17, 0,
					-- layer=2 filter=101 channel=43
					29, 14, -17, 2, 14, 24, -17, -22, 25,
					-- layer=2 filter=101 channel=44
					-2, 6, 0, 8, -5, 10, 2, 8, -7,
					-- layer=2 filter=101 channel=45
					0, 11, -1, -40, -41, -38, -8, -38, -47,
					-- layer=2 filter=101 channel=46
					-5, 26, 21, -5, 4, 1, -20, 1, 20,
					-- layer=2 filter=101 channel=47
					39, 21, -21, -4, -12, 13, 28, -21, -4,
					-- layer=2 filter=101 channel=48
					-5, -4, 10, -10, -2, 11, 7, 2, -4,
					-- layer=2 filter=101 channel=49
					18, 3, -93, 11, -15, -70, 35, 8, 22,
					-- layer=2 filter=101 channel=50
					13, 11, 14, 13, 7, 11, 5, -10, 12,
					-- layer=2 filter=101 channel=51
					-29, -26, -10, -26, -11, 19, 27, 22, 12,
					-- layer=2 filter=101 channel=52
					-18, 12, -23, -20, -4, -33, 55, 26, 7,
					-- layer=2 filter=101 channel=53
					-10, -26, -84, 56, -39, 7, 43, 35, -4,
					-- layer=2 filter=101 channel=54
					-33, -17, -45, -6, -21, -19, 20, 9, 23,
					-- layer=2 filter=101 channel=55
					-7, -2, 4, -5, -4, -6, -6, 15, 2,
					-- layer=2 filter=101 channel=56
					-4, -7, -15, -6, -27, 7, 23, 18, 25,
					-- layer=2 filter=101 channel=57
					5, 2, -2, 2, 5, 11, -5, 9, -8,
					-- layer=2 filter=101 channel=58
					-33, -47, -24, 10, 4, -73, -29, -43, -14,
					-- layer=2 filter=101 channel=59
					-16, -6, 15, -3, 25, -38, -30, -38, 14,
					-- layer=2 filter=101 channel=60
					-63, 25, 2, -60, 34, -11, -3, -4, -15,
					-- layer=2 filter=101 channel=61
					27, -15, 11, -17, -25, 24, 19, 25, 35,
					-- layer=2 filter=101 channel=62
					-13, -45, -63, -10, 17, -34, 52, 6, -29,
					-- layer=2 filter=101 channel=63
					23, 11, 16, -25, 4, 9, -29, -5, 28,
					-- layer=2 filter=101 channel=64
					14, 12, 19, -2, 17, 22, -11, -16, -1,
					-- layer=2 filter=101 channel=65
					-15, -14, 33, -13, 10, 6, 55, -19, 21,
					-- layer=2 filter=101 channel=66
					36, 48, 4, 13, -17, -8, 10, 8, 7,
					-- layer=2 filter=101 channel=67
					2, 30, 18, -8, -5, 20, -30, -35, 13,
					-- layer=2 filter=101 channel=68
					3, -3, -2, 11, 4, -4, 0, 7, 8,
					-- layer=2 filter=101 channel=69
					6, 11, 1, 6, 7, 9, -15, -2, 3,
					-- layer=2 filter=101 channel=70
					-19, -34, -81, -8, -33, -35, 5, -14, -26,
					-- layer=2 filter=101 channel=71
					10, 2, 2, 5, -12, 0, -4, -9, 5,
					-- layer=2 filter=101 channel=72
					-13, -8, 1, 4, -38, -38, -30, -65, -66,
					-- layer=2 filter=101 channel=73
					-3, -3, 9, -23, -36, 69, 86, 47, 19,
					-- layer=2 filter=101 channel=74
					-5, 40, 27, -13, -12, -4, -14, -22, 0,
					-- layer=2 filter=101 channel=75
					43, -68, -35, 63, -35, -59, 20, 0, -8,
					-- layer=2 filter=101 channel=76
					34, -16, 6, 37, -23, -15, 79, -10, 73,
					-- layer=2 filter=101 channel=77
					0, 3, 8, -1, 0, 0, 6, 5, 5,
					-- layer=2 filter=101 channel=78
					-5, -33, -41, -1, -14, -10, 12, 14, 25,
					-- layer=2 filter=101 channel=79
					-4, -4, 4, 11, -5, 0, 1, -1, 10,
					-- layer=2 filter=101 channel=80
					24, 26, 6, 14, 6, 16, -17, -32, -20,
					-- layer=2 filter=101 channel=81
					0, 2, -5, 2, -5, -1, 4, -4, 8,
					-- layer=2 filter=101 channel=82
					-2, 1, -8, -3, -7, 7, -2, -2, 10,
					-- layer=2 filter=101 channel=83
					13, -8, -5, -1, -2, -16, -14, -21, -17,
					-- layer=2 filter=101 channel=84
					1, -5, -5, -3, -6, 1, -6, 7, -4,
					-- layer=2 filter=101 channel=85
					6, -4, 0, 7, 1, 10, 10, 19, 14,
					-- layer=2 filter=101 channel=86
					8, 6, -9, 5, -1, 3, 7, 11, 3,
					-- layer=2 filter=101 channel=87
					-14, 8, -92, -44, -8, -35, -10, 5, -35,
					-- layer=2 filter=101 channel=88
					-28, 18, 38, -16, -4, 0, -21, -13, 19,
					-- layer=2 filter=101 channel=89
					-9, -44, 11, 22, 10, -49, -41, -30, -20,
					-- layer=2 filter=101 channel=90
					-8, -7, -2, -8, 6, 0, 0, 1, -11,
					-- layer=2 filter=101 channel=91
					18, -20, 47, 4, 4, -32, -24, -41, -28,
					-- layer=2 filter=101 channel=92
					-21, -3, 13, 34, 18, -30, -26, -51, -31,
					-- layer=2 filter=101 channel=93
					25, -59, 35, 22, 24, 17, 8, -15, 8,
					-- layer=2 filter=101 channel=94
					39, -22, -29, -10, -15, -34, -3, 47, 10,
					-- layer=2 filter=101 channel=95
					8, -2, -6, 1, 4, 9, -6, 7, 5,
					-- layer=2 filter=101 channel=96
					34, 27, -6, -32, 7, 5, 32, 62, 26,
					-- layer=2 filter=101 channel=97
					29, 31, -5, 0, 8, 8, -14, -16, -1,
					-- layer=2 filter=101 channel=98
					21, -3, -61, -4, -23, -9, 22, -15, -10,
					-- layer=2 filter=101 channel=99
					12, 36, -40, -16, -17, -36, 44, 26, -3,
					-- layer=2 filter=101 channel=100
					-5, 5, 10, 14, 3, -28, -41, -37, -25,
					-- layer=2 filter=101 channel=101
					18, -28, -5, -12, 19, 36, -20, 26, 26,
					-- layer=2 filter=101 channel=102
					7, 22, -26, -5, 8, -44, 26, 46, -7,
					-- layer=2 filter=101 channel=103
					-32, -25, 13, -35, 37, 10, -3, -24, -11,
					-- layer=2 filter=101 channel=104
					13, 36, -53, 2, -39, -36, 30, 29, -6,
					-- layer=2 filter=101 channel=105
					-20, -79, -77, 2, -39, -30, -9, -47, 45,
					-- layer=2 filter=101 channel=106
					-29, -16, -7, -11, 4, 9, -21, -34, 1,
					-- layer=2 filter=101 channel=107
					-24, 8, 19, 9, 9, 10, 1, -7, -12,
					-- layer=2 filter=101 channel=108
					29, 27, -3, 48, 13, -14, 66, 47, 3,
					-- layer=2 filter=101 channel=109
					-5, 1, -6, -2, 2, -3, 0, 14, -7,
					-- layer=2 filter=101 channel=110
					-1, -20, 25, 0, -10, 20, -21, -47, 28,
					-- layer=2 filter=101 channel=111
					-10, 1, 4, -4, -1, 0, 2, -8, 8,
					-- layer=2 filter=101 channel=112
					-17, -14, -6, -57, -6, 40, 14, 5, 17,
					-- layer=2 filter=101 channel=113
					3, -34, 15, -17, 18, 21, -22, 16, -17,
					-- layer=2 filter=101 channel=114
					10, 23, 14, -2, 10, 10, -1, -13, -15,
					-- layer=2 filter=101 channel=115
					-7, -10, 0, -5, -2, -7, -3, 10, 2,
					-- layer=2 filter=101 channel=116
					-19, 24, -88, -32, 2, -33, 29, 31, -23,
					-- layer=2 filter=101 channel=117
					-13, -4, 9, -24, -5, -17, 47, -12, 9,
					-- layer=2 filter=101 channel=118
					3, 29, -3, 14, 7, 16, 19, 0, 9,
					-- layer=2 filter=101 channel=119
					7, 30, -32, -3, 9, -34, -4, -10, -20,
					-- layer=2 filter=101 channel=120
					8, -1, -9, 9, 7, -7, -5, 9, -4,
					-- layer=2 filter=101 channel=121
					-6, 5, 0, -9, 5, -2, -6, 9, 0,
					-- layer=2 filter=101 channel=122
					-3, -10, 8, -1, -2, -4, -8, -3, 0,
					-- layer=2 filter=101 channel=123
					23, -39, -13, -50, -49, 3, 1, -3, -6,
					-- layer=2 filter=101 channel=124
					24, -7, -16, 46, 4, -47, -7, 2, -60,
					-- layer=2 filter=101 channel=125
					5, 6, 9, 6, 8, 1, 1, 8, -7,
					-- layer=2 filter=101 channel=126
					35, 46, 58, 12, 12, 14, 41, -8, 3,
					-- layer=2 filter=101 channel=127
					-27, 6, 6, -17, 7, -10, -25, -5, -9,
					-- layer=2 filter=102 channel=0
					14, -47, 5, 0, -12, -10, -22, -38, -32,
					-- layer=2 filter=102 channel=1
					-1, -6, -17, -20, 12, -21, -42, -27, 4,
					-- layer=2 filter=102 channel=2
					0, 1, -4, -7, -4, -9, 2, 3, 5,
					-- layer=2 filter=102 channel=3
					-17, 2, -24, -6, 3, -26, 25, -15, -32,
					-- layer=2 filter=102 channel=4
					-13, 20, 9, -5, -30, 1, -20, -45, 18,
					-- layer=2 filter=102 channel=5
					-13, -12, -22, -5, 37, 10, -35, -4, -19,
					-- layer=2 filter=102 channel=6
					10, -44, -22, -26, -6, -57, -1, 27, -18,
					-- layer=2 filter=102 channel=7
					14, -2, 9, -32, -27, -23, -32, -21, 6,
					-- layer=2 filter=102 channel=8
					0, 5, -5, 1, -6, 10, 1, 8, -7,
					-- layer=2 filter=102 channel=9
					9, -3, -22, -16, -17, -13, 25, 13, -3,
					-- layer=2 filter=102 channel=10
					-18, -27, -16, 3, -13, -38, 0, -29, -56,
					-- layer=2 filter=102 channel=11
					4, 1, -19, -9, -4, -42, 3, -36, 0,
					-- layer=2 filter=102 channel=12
					15, -10, -3, -4, 15, -10, -4, -17, -8,
					-- layer=2 filter=102 channel=13
					-6, -3, -4, -2, 2, -8, -6, 3, 1,
					-- layer=2 filter=102 channel=14
					-22, -6, -14, -21, -23, -8, -13, -35, 0,
					-- layer=2 filter=102 channel=15
					-19, -9, 5, 22, 2, 0, -6, -24, -18,
					-- layer=2 filter=102 channel=16
					-15, -20, -8, -25, -39, -6, 4, -27, -34,
					-- layer=2 filter=102 channel=17
					0, 8, -7, -1, 7, 5, -1, -9, 4,
					-- layer=2 filter=102 channel=18
					-9, 17, -3, -7, -8, 8, 7, -30, 15,
					-- layer=2 filter=102 channel=19
					2, -30, -23, -44, -15, -23, -27, -24, -7,
					-- layer=2 filter=102 channel=20
					-3, 1, 2, -10, -3, 3, 9, 1, -5,
					-- layer=2 filter=102 channel=21
					0, 10, 4, -4, 1, 7, 1, -1, 4,
					-- layer=2 filter=102 channel=22
					0, -3, -5, 2, 2, 6, 0, 1, -8,
					-- layer=2 filter=102 channel=23
					-11, -18, 31, 12, -6, 39, -22, -4, 13,
					-- layer=2 filter=102 channel=24
					-11, -42, -35, 3, -12, -44, 22, -12, -11,
					-- layer=2 filter=102 channel=25
					-47, -37, -49, -16, -53, -48, -16, -57, -49,
					-- layer=2 filter=102 channel=26
					7, -4, 7, -9, 7, 10, -3, -2, 7,
					-- layer=2 filter=102 channel=27
					9, 12, -9, 24, -5, 8, -21, -36, 6,
					-- layer=2 filter=102 channel=28
					-38, -31, -49, 9, 17, 12, 0, 15, 24,
					-- layer=2 filter=102 channel=29
					-8, -9, -3, 0, 3, 4, -6, 3, 2,
					-- layer=2 filter=102 channel=30
					-22, 6, -31, 15, -7, 1, -7, 18, -57,
					-- layer=2 filter=102 channel=31
					-28, 23, 3, -17, -12, -35, -6, -20, -9,
					-- layer=2 filter=102 channel=32
					-1, -10, 6, 1, -2, 0, 4, -9, -8,
					-- layer=2 filter=102 channel=33
					12, -4, -8, -10, -13, 11, -28, -40, -1,
					-- layer=2 filter=102 channel=34
					-5, 8, -32, -23, 11, 16, -13, -2, -7,
					-- layer=2 filter=102 channel=35
					-24, -4, -14, 18, 55, 13, -20, -21, 3,
					-- layer=2 filter=102 channel=36
					0, 5, 0, 3, -9, 6, 3, -9, 1,
					-- layer=2 filter=102 channel=37
					-3, 16, -11, -14, -19, -26, -4, -4, -5,
					-- layer=2 filter=102 channel=38
					5, 0, -4, -1, 10, -49, -49, -19, -38,
					-- layer=2 filter=102 channel=39
					21, -11, 0, -19, -42, -17, 11, -5, -2,
					-- layer=2 filter=102 channel=40
					-9, 16, -3, 32, -20, -8, 30, -30, 21,
					-- layer=2 filter=102 channel=41
					2, -11, 6, -6, 7, -1, -6, -5, 1,
					-- layer=2 filter=102 channel=42
					-10, -28, -11, 9, -7, 11, 0, -16, 22,
					-- layer=2 filter=102 channel=43
					-15, 12, -10, 5, -10, 2, 16, -12, 9,
					-- layer=2 filter=102 channel=44
					-7, 5, 1, 3, -7, -6, 7, -4, 2,
					-- layer=2 filter=102 channel=45
					-26, 2, -13, -6, -31, -18, -19, -10, -24,
					-- layer=2 filter=102 channel=46
					0, 4, -3, -12, -15, -42, -7, -29, -41,
					-- layer=2 filter=102 channel=47
					-22, -3, -14, -13, -35, -3, 14, -4, -23,
					-- layer=2 filter=102 channel=48
					-1, -1, 1, 8, 6, 5, 6, -2, 2,
					-- layer=2 filter=102 channel=49
					-7, -21, -9, 21, -27, 10, 21, -20, 25,
					-- layer=2 filter=102 channel=50
					2, -6, -9, 3, 6, 7, -5, -2, -1,
					-- layer=2 filter=102 channel=51
					-12, -6, -40, -15, -31, -33, -25, -26, -43,
					-- layer=2 filter=102 channel=52
					7, 35, -7, -7, -41, -13, 0, 21, -7,
					-- layer=2 filter=102 channel=53
					-13, 10, -10, 0, -45, -31, 7, -11, 25,
					-- layer=2 filter=102 channel=54
					-22, -8, 2, -16, 23, -14, -79, -23, 4,
					-- layer=2 filter=102 channel=55
					7, -6, -7, -1, -11, 10, -7, -3, 6,
					-- layer=2 filter=102 channel=56
					0, 8, -20, -7, 17, -38, 16, -32, 13,
					-- layer=2 filter=102 channel=57
					1, -1, 9, -3, -4, 9, 0, -9, -4,
					-- layer=2 filter=102 channel=58
					4, 0, 11, -20, 19, 0, -17, -23, -21,
					-- layer=2 filter=102 channel=59
					33, -44, 0, -50, -3, -17, -11, -2, 32,
					-- layer=2 filter=102 channel=60
					10, -26, -6, -52, 35, 0, -74, 24, -10,
					-- layer=2 filter=102 channel=61
					26, -21, -21, -24, -8, -29, -44, 21, 2,
					-- layer=2 filter=102 channel=62
					-12, -24, -19, -41, -3, -8, -13, 0, -8,
					-- layer=2 filter=102 channel=63
					12, -31, 14, -1, -23, 10, -10, 3, -4,
					-- layer=2 filter=102 channel=64
					-16, -16, 0, -7, -12, 13, 10, 14, 8,
					-- layer=2 filter=102 channel=65
					20, -28, -3, 0, 8, -36, -35, 27, -1,
					-- layer=2 filter=102 channel=66
					26, 8, -26, 0, -14, -9, 0, -12, -2,
					-- layer=2 filter=102 channel=67
					-6, -8, -10, 0, -12, -24, 9, -15, -19,
					-- layer=2 filter=102 channel=68
					-11, 5, 2, -5, -1, -5, 2, -11, -7,
					-- layer=2 filter=102 channel=69
					2, -5, -4, 2, -5, 23, 15, 6, 12,
					-- layer=2 filter=102 channel=70
					-41, -16, -36, 19, 8, 2, -38, -13, 0,
					-- layer=2 filter=102 channel=71
					-12, -16, -16, 11, -26, -31, 3, -45, 10,
					-- layer=2 filter=102 channel=72
					3, -7, 1, 6, -38, 18, -13, 0, 45,
					-- layer=2 filter=102 channel=73
					-25, 42, -1, 22, -18, -13, -8, -37, 7,
					-- layer=2 filter=102 channel=74
					5, -6, 12, -10, -14, -14, -5, -34, -24,
					-- layer=2 filter=102 channel=75
					-10, -50, 13, -4, -41, 18, 32, 31, 22,
					-- layer=2 filter=102 channel=76
					-14, -1, 6, -17, -21, -9, -4, 10, 13,
					-- layer=2 filter=102 channel=77
					-2, 6, -7, -5, -7, 0, -10, -5, -3,
					-- layer=2 filter=102 channel=78
					-9, 4, -14, -27, 1, -26, 0, -18, 12,
					-- layer=2 filter=102 channel=79
					-10, -7, 8, -9, 1, -4, 2, -6, 7,
					-- layer=2 filter=102 channel=80
					-2, -14, -9, 0, -23, -33, 11, -26, -19,
					-- layer=2 filter=102 channel=81
					-3, -9, 4, 7, 6, 5, -8, -9, 2,
					-- layer=2 filter=102 channel=82
					8, -11, 0, -10, 7, 6, -4, 5, 2,
					-- layer=2 filter=102 channel=83
					-11, -26, 0, 1, 12, 1, -7, 15, 11,
					-- layer=2 filter=102 channel=84
					-4, 3, -1, 7, -6, 2, -1, -8, -1,
					-- layer=2 filter=102 channel=85
					-4, 3, -11, 7, -2, 1, -1, 1, 4,
					-- layer=2 filter=102 channel=86
					0, -6, 2, -2, 10, 9, -4, -12, -9,
					-- layer=2 filter=102 channel=87
					15, 38, 40, 25, -30, 40, -27, 8, 18,
					-- layer=2 filter=102 channel=88
					-1, -9, -33, 6, -12, -21, 18, 5, -19,
					-- layer=2 filter=102 channel=89
					9, -16, -12, -36, -19, -12, -1, -38, -2,
					-- layer=2 filter=102 channel=90
					-4, 1, -4, -7, 4, 5, 1, -3, 3,
					-- layer=2 filter=102 channel=91
					-2, -33, -26, -16, 19, -12, 9, 26, 28,
					-- layer=2 filter=102 channel=92
					13, -11, -29, -9, 16, -43, -41, -26, 9,
					-- layer=2 filter=102 channel=93
					-6, 4, 1, -27, -13, -43, -19, 10, -3,
					-- layer=2 filter=102 channel=94
					32, -36, 0, -50, 14, -22, -25, 1, 14,
					-- layer=2 filter=102 channel=95
					0, 4, 5, -7, 3, -13, -5, -11, -11,
					-- layer=2 filter=102 channel=96
					-20, 25, 47, 17, -11, 50, -42, -2, 23,
					-- layer=2 filter=102 channel=97
					0, -8, 5, -3, -8, 12, 29, 0, -4,
					-- layer=2 filter=102 channel=98
					-3, -18, -14, 0, -14, -14, 4, -12, -7,
					-- layer=2 filter=102 channel=99
					0, 5, -34, -40, -56, -23, -26, -48, -36,
					-- layer=2 filter=102 channel=100
					20, -32, 6, 4, 21, 7, -8, 4, 1,
					-- layer=2 filter=102 channel=101
					-12, -27, 0, -2, -14, -25, -1, -23, -37,
					-- layer=2 filter=102 channel=102
					-30, 43, 22, 4, -12, 34, -56, -23, 40,
					-- layer=2 filter=102 channel=103
					-26, -16, 10, -6, -1, -9, -14, 2, -4,
					-- layer=2 filter=102 channel=104
					7, -15, 16, 24, -5, 15, 9, -10, 39,
					-- layer=2 filter=102 channel=105
					3, -28, 12, -36, -35, 23, 4, 3, 49,
					-- layer=2 filter=102 channel=106
					-16, -44, -1, -64, -52, -59, -29, -22, -47,
					-- layer=2 filter=102 channel=107
					-34, -13, 16, -26, -23, -22, -27, -31, 15,
					-- layer=2 filter=102 channel=108
					-30, 27, 3, -9, -7, 24, -17, -16, 23,
					-- layer=2 filter=102 channel=109
					6, 7, 4, -5, -8, 6, 1, 4, -4,
					-- layer=2 filter=102 channel=110
					5, -37, -15, -4, -20, -4, 6, 17, 17,
					-- layer=2 filter=102 channel=111
					7, -8, 3, 3, 10, -5, 2, -8, -8,
					-- layer=2 filter=102 channel=112
					-5, -25, -65, -26, -7, -66, -25, 0, -44,
					-- layer=2 filter=102 channel=113
					-16, -8, -45, -12, 0, 1, -9, 13, -33,
					-- layer=2 filter=102 channel=114
					-2, -7, 8, -2, -4, 1, -9, 1, -5,
					-- layer=2 filter=102 channel=115
					-9, 2, -5, -7, -9, 3, 2, -5, 2,
					-- layer=2 filter=102 channel=116
					0, 55, 18, 22, -12, 49, -31, 3, 34,
					-- layer=2 filter=102 channel=117
					7, -13, 11, -36, -32, -68, -37, -32, -7,
					-- layer=2 filter=102 channel=118
					-9, -13, -1, -8, -20, -1, 17, -14, 9,
					-- layer=2 filter=102 channel=119
					-7, -14, -4, -29, -26, 12, -25, -27, 15,
					-- layer=2 filter=102 channel=120
					9, 5, 0, -4, -2, 7, -9, 2, 1,
					-- layer=2 filter=102 channel=121
					-2, -4, 6, 9, 5, 7, -3, 4, -5,
					-- layer=2 filter=102 channel=122
					0, 0, -10, 3, 3, 4, -8, -4, 6,
					-- layer=2 filter=102 channel=123
					29, 8, 16, -31, -53, 3, -3, -2, 30,
					-- layer=2 filter=102 channel=124
					11, -24, 4, -45, 7, -12, -34, -23, -3,
					-- layer=2 filter=102 channel=125
					-8, 1, -7, -6, 8, 5, 6, -9, 3,
					-- layer=2 filter=102 channel=126
					-22, -38, 16, 4, -50, 6, -21, 3, 32,
					-- layer=2 filter=102 channel=127
					1, -7, 8, -28, -4, 34, 0, -2, 5,
					-- layer=2 filter=103 channel=0
					-9, -21, -10, -33, -16, -5, -15, -23, 2,
					-- layer=2 filter=103 channel=1
					-29, -16, -29, -21, -14, -9, -34, -33, -19,
					-- layer=2 filter=103 channel=2
					-6, -7, 5, 5, -4, -12, 4, -5, -12,
					-- layer=2 filter=103 channel=3
					-9, -24, -8, 0, 1, 0, -32, -14, -11,
					-- layer=2 filter=103 channel=4
					5, 14, 29, -5, 15, 5, 1, 8, -21,
					-- layer=2 filter=103 channel=5
					-5, 14, -14, -12, -23, -1, -29, -37, -14,
					-- layer=2 filter=103 channel=6
					15, -3, -28, -7, -5, -25, 9, -21, 15,
					-- layer=2 filter=103 channel=7
					0, -8, -11, 12, 4, -9, -27, -23, -6,
					-- layer=2 filter=103 channel=8
					-1, -5, 7, -5, 5, 1, 8, -4, -2,
					-- layer=2 filter=103 channel=9
					5, -2, 0, -4, -7, -20, -34, -31, -30,
					-- layer=2 filter=103 channel=10
					-27, -11, -11, -32, -12, 0, -8, -13, 6,
					-- layer=2 filter=103 channel=11
					13, -19, 1, -19, -19, 2, -33, -23, -21,
					-- layer=2 filter=103 channel=12
					-27, 8, -9, -22, -7, 1, -36, -24, -24,
					-- layer=2 filter=103 channel=13
					0, 11, -9, -7, 3, 10, 10, -3, -1,
					-- layer=2 filter=103 channel=14
					-15, -26, -7, -34, -11, -26, -12, -13, -40,
					-- layer=2 filter=103 channel=15
					18, -25, -26, -28, -37, -8, -49, 2, -2,
					-- layer=2 filter=103 channel=16
					-26, -11, -15, -23, -31, -37, -10, -26, -20,
					-- layer=2 filter=103 channel=17
					-10, 5, 7, 4, -2, 0, -3, 1, -2,
					-- layer=2 filter=103 channel=18
					15, 1, 1, 4, -28, -22, -13, -19, -5,
					-- layer=2 filter=103 channel=19
					-22, -11, -28, -24, -14, -1, -47, -38, -11,
					-- layer=2 filter=103 channel=20
					0, -3, 0, 8, 4, 2, -4, 4, 8,
					-- layer=2 filter=103 channel=21
					7, -8, -2, 1, -7, 0, 6, -6, -1,
					-- layer=2 filter=103 channel=22
					-7, 2, -1, 2, 4, -4, 4, -4, -5,
					-- layer=2 filter=103 channel=23
					-12, -10, -13, -13, -15, 0, -6, 11, 18,
					-- layer=2 filter=103 channel=24
					-10, -26, -6, -27, -11, -3, -24, -48, -2,
					-- layer=2 filter=103 channel=25
					5, -13, -10, -22, -9, -14, -35, -6, -14,
					-- layer=2 filter=103 channel=26
					-9, -7, 0, -2, 7, 2, -5, 7, -4,
					-- layer=2 filter=103 channel=27
					-7, -14, -7, 0, -5, -14, -7, -29, -14,
					-- layer=2 filter=103 channel=28
					-1, -7, -6, 23, -18, -8, -3, -6, -16,
					-- layer=2 filter=103 channel=29
					2, -10, 8, 0, 6, 0, -10, 7, 3,
					-- layer=2 filter=103 channel=30
					7, -14, -1, -23, 4, -14, -5, 20, -24,
					-- layer=2 filter=103 channel=31
					41, -9, -6, -14, -22, -8, -16, 0, 4,
					-- layer=2 filter=103 channel=32
					1, 6, -10, 2, -10, 3, 5, 5, -4,
					-- layer=2 filter=103 channel=33
					14, -22, 10, -13, -13, -19, -22, -30, -28,
					-- layer=2 filter=103 channel=34
					-21, 38, -2, 18, -30, 12, 1, -15, -27,
					-- layer=2 filter=103 channel=35
					8, 13, -25, 20, 2, 0, 0, 26, -23,
					-- layer=2 filter=103 channel=36
					-6, 8, 4, 8, 7, 0, 0, 6, 4,
					-- layer=2 filter=103 channel=37
					7, -7, -26, -6, 0, -22, -28, -21, -31,
					-- layer=2 filter=103 channel=38
					4, -8, 4, -10, -3, 9, 4, -14, -17,
					-- layer=2 filter=103 channel=39
					-8, -26, -26, -20, -5, -12, -34, -29, 2,
					-- layer=2 filter=103 channel=40
					20, -7, -9, 4, -1, -19, -34, -11, -8,
					-- layer=2 filter=103 channel=41
					-5, -2, -7, 2, 7, 4, -7, 10, -2,
					-- layer=2 filter=103 channel=42
					-14, -6, -40, -25, -21, 2, -33, -7, -1,
					-- layer=2 filter=103 channel=43
					30, 9, -22, 15, -3, -9, -12, -4, -18,
					-- layer=2 filter=103 channel=44
					-1, 3, -2, 9, 1, 1, -5, 0, -9,
					-- layer=2 filter=103 channel=45
					31, -30, -21, -9, -10, -23, -13, -14, -5,
					-- layer=2 filter=103 channel=46
					-7, 7, -11, -15, 1, 2, 12, -2, 0,
					-- layer=2 filter=103 channel=47
					3, -14, -30, -1, -28, -32, -7, -14, -5,
					-- layer=2 filter=103 channel=48
					0, -7, 2, -3, -11, 2, -7, 1, -3,
					-- layer=2 filter=103 channel=49
					-8, 7, -26, 4, -23, 5, -14, -29, -13,
					-- layer=2 filter=103 channel=50
					-1, 5, -8, 0, -2, -4, -9, -10, -5,
					-- layer=2 filter=103 channel=51
					2, 7, -15, -26, 0, -2, -19, -18, -32,
					-- layer=2 filter=103 channel=52
					14, -19, 1, -32, -11, -44, -14, -3, 3,
					-- layer=2 filter=103 channel=53
					16, -15, -4, -51, -22, -22, -40, -9, -18,
					-- layer=2 filter=103 channel=54
					2, -6, -29, -1, -9, -13, -35, -10, -9,
					-- layer=2 filter=103 channel=55
					0, -5, 8, 1, -8, -1, 3, -8, 2,
					-- layer=2 filter=103 channel=56
					6, -7, 5, -8, -12, -5, -15, -30, -19,
					-- layer=2 filter=103 channel=57
					-1, -7, 9, 11, 4, 10, -3, 4, 10,
					-- layer=2 filter=103 channel=58
					1, 18, -11, -5, -9, -7, -16, -5, -9,
					-- layer=2 filter=103 channel=59
					1, -25, 4, -23, 3, 1, -13, -5, -6,
					-- layer=2 filter=103 channel=60
					-47, 10, -23, 16, -22, 12, -17, -19, 34,
					-- layer=2 filter=103 channel=61
					-25, -2, -18, 17, -2, 2, 4, -15, 24,
					-- layer=2 filter=103 channel=62
					24, 16, -12, 2, -50, -28, 0, -38, 1,
					-- layer=2 filter=103 channel=63
					-30, -14, -6, -12, -14, -1, -10, -2, 28,
					-- layer=2 filter=103 channel=64
					-30, -9, -14, -11, 2, -23, 3, 12, -12,
					-- layer=2 filter=103 channel=65
					-30, -4, -27, 8, -8, -6, 5, -23, 8,
					-- layer=2 filter=103 channel=66
					-29, -11, 15, 5, 3, -11, -1, -24, -11,
					-- layer=2 filter=103 channel=67
					-15, -7, -7, -33, -26, 5, -19, -23, 12,
					-- layer=2 filter=103 channel=68
					-5, -5, 3, 1, 2, -8, -12, 7, 6,
					-- layer=2 filter=103 channel=69
					-2, -19, -18, -2, -15, -26, 8, 13, -19,
					-- layer=2 filter=103 channel=70
					9, 8, -36, -7, -22, -20, -2, 8, -27,
					-- layer=2 filter=103 channel=71
					5, 6, 10, 8, -5, 9, -13, 15, -11,
					-- layer=2 filter=103 channel=72
					-22, -22, -5, 0, -21, 8, 5, -12, -9,
					-- layer=2 filter=103 channel=73
					14, -37, -13, -35, -9, 0, -9, 23, -1,
					-- layer=2 filter=103 channel=74
					-18, -2, -2, -28, 4, 14, 0, 10, 24,
					-- layer=2 filter=103 channel=75
					-14, 2, -17, 10, -16, 7, -6, -40, -31,
					-- layer=2 filter=103 channel=76
					33, -40, 4, -18, -24, 0, -21, -16, -4,
					-- layer=2 filter=103 channel=77
					-5, 5, -2, 3, -9, 1, 5, 4, 5,
					-- layer=2 filter=103 channel=78
					11, -16, -16, -21, -14, -14, -20, -29, -25,
					-- layer=2 filter=103 channel=79
					6, 8, 7, -1, 2, 8, -1, 8, -8,
					-- layer=2 filter=103 channel=80
					0, -5, -11, -14, -3, -4, -8, -11, 2,
					-- layer=2 filter=103 channel=81
					-11, -11, -11, -5, -9, 4, 5, 7, -11,
					-- layer=2 filter=103 channel=82
					-7, 0, -7, -5, 8, 1, 2, 5, 10,
					-- layer=2 filter=103 channel=83
					-19, -17, -4, -19, -22, 6, -24, 8, -23,
					-- layer=2 filter=103 channel=84
					-2, 0, 7, 0, -6, -1, 5, 5, 5,
					-- layer=2 filter=103 channel=85
					-3, 8, 8, 3, 5, -7, 2, 7, -6,
					-- layer=2 filter=103 channel=86
					4, -4, 0, -7, -2, -3, 8, -9, -8,
					-- layer=2 filter=103 channel=87
					24, -17, -10, -15, 12, -45, -24, 1, 3,
					-- layer=2 filter=103 channel=88
					0, -17, -21, -29, -2, -9, -19, -24, 10,
					-- layer=2 filter=103 channel=89
					-33, -12, -12, -36, 3, -9, -2, -3, -25,
					-- layer=2 filter=103 channel=90
					5, 8, -5, -9, -1, -8, -2, 9, 4,
					-- layer=2 filter=103 channel=91
					-24, -26, -19, -12, -24, 4, -10, -12, -10,
					-- layer=2 filter=103 channel=92
					-9, -10, -25, -20, -26, -15, -17, -30, -4,
					-- layer=2 filter=103 channel=93
					-7, 4, -18, 11, -24, -21, 32, 7, -9,
					-- layer=2 filter=103 channel=94
					-7, -24, -23, -18, -8, -8, -36, -14, 27,
					-- layer=2 filter=103 channel=95
					-4, -8, 11, 6, 4, -10, 3, 4, 7,
					-- layer=2 filter=103 channel=96
					-41, -32, 9, -24, 24, -8, -15, 22, 10,
					-- layer=2 filter=103 channel=97
					9, -28, -8, -26, -6, -25, -20, -21, -20,
					-- layer=2 filter=103 channel=98
					14, 3, -16, 5, -35, -10, 4, -16, 2,
					-- layer=2 filter=103 channel=99
					7, -22, 5, -61, -16, -37, 0, -11, -16,
					-- layer=2 filter=103 channel=100
					-11, -5, -21, -11, -9, 18, -10, -4, -3,
					-- layer=2 filter=103 channel=101
					21, -18, 30, -8, -22, -5, -12, 6, 17,
					-- layer=2 filter=103 channel=102
					-20, -8, -2, -4, -2, -10, -25, 40, -20,
					-- layer=2 filter=103 channel=103
					-5, 4, -1, -3, 6, -17, -30, -5, -12,
					-- layer=2 filter=103 channel=104
					16, 0, -14, -1, -9, -4, -31, -18, -16,
					-- layer=2 filter=103 channel=105
					11, -27, 1, -9, -5, -20, 27, 2, -5,
					-- layer=2 filter=103 channel=106
					-11, -28, -1, -31, -8, -2, -25, 0, -23,
					-- layer=2 filter=103 channel=107
					-9, -19, 21, 2, 6, 4, -8, 0, 7,
					-- layer=2 filter=103 channel=108
					-27, -21, -16, -2, -15, -22, -28, 17, -23,
					-- layer=2 filter=103 channel=109
					0, -3, -5, -12, -9, 7, -4, -5, -1,
					-- layer=2 filter=103 channel=110
					-40, -19, -33, -18, -12, -15, -25, -8, 11,
					-- layer=2 filter=103 channel=111
					0, 2, 10, -1, -10, -5, 6, -10, 6,
					-- layer=2 filter=103 channel=112
					-26, -4, -13, 14, -8, -16, 16, 3, 12,
					-- layer=2 filter=103 channel=113
					-22, -15, -12, -11, 2, -27, -5, 5, -26,
					-- layer=2 filter=103 channel=114
					-1, -11, 11, 5, 0, 1, -3, 2, 2,
					-- layer=2 filter=103 channel=115
					-5, -10, 2, -1, 8, 7, 4, 0, 2,
					-- layer=2 filter=103 channel=116
					-12, 5, 9, -4, -6, -29, -20, 4, -18,
					-- layer=2 filter=103 channel=117
					-16, 2, -18, -20, -12, 5, -38, -20, 17,
					-- layer=2 filter=103 channel=118
					-5, -11, -24, -17, -9, -30, -12, -6, -3,
					-- layer=2 filter=103 channel=119
					23, 6, -24, 13, -19, -27, -9, 11, -21,
					-- layer=2 filter=103 channel=120
					-9, 7, -3, -10, -5, -5, -6, -4, 3,
					-- layer=2 filter=103 channel=121
					7, 0, 8, 3, -2, -8, 2, 7, 2,
					-- layer=2 filter=103 channel=122
					-5, -1, 5, 6, -5, -4, -6, -6, 2,
					-- layer=2 filter=103 channel=123
					-6, -16, -16, -18, 4, -33, -7, 2, -7,
					-- layer=2 filter=103 channel=124
					11, -1, -34, -31, -2, -24, -25, -6, -3,
					-- layer=2 filter=103 channel=125
					6, -8, 0, -1, 5, 2, -8, 0, -7,
					-- layer=2 filter=103 channel=126
					-1, -25, 23, -14, 14, 0, -7, 0, 46,
					-- layer=2 filter=103 channel=127
					-16, 0, -16, -13, -21, -25, 0, 0, -8,
					-- layer=2 filter=104 channel=0
					-13, -24, -35, -30, -8, -43, -32, 6, 0,
					-- layer=2 filter=104 channel=1
					23, 14, 26, 19, 0, 1, 10, -3, 10,
					-- layer=2 filter=104 channel=2
					-1, 3, -2, 10, 6, -7, -6, 10, 2,
					-- layer=2 filter=104 channel=3
					1, -1, -33, -26, 41, 1, 21, 24, -2,
					-- layer=2 filter=104 channel=4
					22, 10, 16, 15, 23, -3, -16, 12, -1,
					-- layer=2 filter=104 channel=5
					-99, -51, -62, -44, -34, 0, -33, 27, 9,
					-- layer=2 filter=104 channel=6
					-13, -56, 9, 24, 47, 53, -7, 29, 88,
					-- layer=2 filter=104 channel=7
					6, -34, -8, 14, 2, -6, 14, -8, 14,
					-- layer=2 filter=104 channel=8
					-8, 4, 1, 10, -3, -7, -7, -11, -5,
					-- layer=2 filter=104 channel=9
					14, 17, 14, -3, -18, -26, 23, -39, -34,
					-- layer=2 filter=104 channel=10
					18, 18, 5, -22, 21, -21, -10, 20, 16,
					-- layer=2 filter=104 channel=11
					-64, -69, -50, -43, -12, 3, -9, -8, 28,
					-- layer=2 filter=104 channel=12
					7, -18, -6, 31, 10, -4, 38, 9, 22,
					-- layer=2 filter=104 channel=13
					0, 2, -4, 1, 6, -6, -2, 1, -7,
					-- layer=2 filter=104 channel=14
					33, 21, 18, 22, 2, 6, 18, 10, -12,
					-- layer=2 filter=104 channel=15
					23, 42, 13, 48, 18, -22, -30, 12, 3,
					-- layer=2 filter=104 channel=16
					2, 4, 12, -23, -24, -18, 1, -5, -15,
					-- layer=2 filter=104 channel=17
					-3, -5, -5, -4, 0, 9, -4, 2, 0,
					-- layer=2 filter=104 channel=18
					-18, -9, -24, 9, -2, 9, 1, -31, -21,
					-- layer=2 filter=104 channel=19
					-51, -16, -8, 32, -5, -1, 19, 10, 37,
					-- layer=2 filter=104 channel=20
					-4, 6, 3, -1, -3, 8, -8, 5, -7,
					-- layer=2 filter=104 channel=21
					-11, -9, -15, 7, -4, -2, 6, 6, -13,
					-- layer=2 filter=104 channel=22
					5, 7, 1, 3, -8, 5, -8, -2, -7,
					-- layer=2 filter=104 channel=23
					39, 18, 44, -28, -10, -9, 4, 16, 21,
					-- layer=2 filter=104 channel=24
					2, 6, -39, -6, -17, -35, -32, -29, -65,
					-- layer=2 filter=104 channel=25
					7, -19, -18, 40, 23, 18, -23, -16, 11,
					-- layer=2 filter=104 channel=26
					9, -8, 0, 1, -7, -6, 0, 2, 6,
					-- layer=2 filter=104 channel=27
					-19, 5, -42, -42, -40, -71, -66, -45, -34,
					-- layer=2 filter=104 channel=28
					0, -15, -20, -52, -53, -50, 44, 30, 22,
					-- layer=2 filter=104 channel=29
					-4, -8, 1, -1, 6, 11, 2, 0, -4,
					-- layer=2 filter=104 channel=30
					18, 18, -9, 21, -6, 4, 19, -12, -27,
					-- layer=2 filter=104 channel=31
					-29, 25, -20, -36, -40, -1, -17, 71, 33,
					-- layer=2 filter=104 channel=32
					-7, -5, 0, 7, 7, 4, -4, 2, 0,
					-- layer=2 filter=104 channel=33
					-1, -5, 20, 9, -5, -27, 29, 25, 32,
					-- layer=2 filter=104 channel=34
					-18, 1, -33, 37, 38, 8, -2, 26, -7,
					-- layer=2 filter=104 channel=35
					18, 12, -7, -32, 4, -37, 23, 28, -5,
					-- layer=2 filter=104 channel=36
					-9, -9, -7, -8, 10, -5, -3, 8, -5,
					-- layer=2 filter=104 channel=37
					-70, -44, -37, -45, -26, -5, -22, -9, 16,
					-- layer=2 filter=104 channel=38
					7, 17, -7, -12, 0, -21, -17, 18, 16,
					-- layer=2 filter=104 channel=39
					41, 35, 51, -24, 2, -4, 8, -30, -19,
					-- layer=2 filter=104 channel=40
					-19, -32, -4, 27, 16, -26, 21, 8, 6,
					-- layer=2 filter=104 channel=41
					3, -7, 4, -5, -9, 9, -8, 4, -6,
					-- layer=2 filter=104 channel=42
					25, 30, 51, -7, 13, -10, 0, 28, -11,
					-- layer=2 filter=104 channel=43
					-12, 5, -36, -26, 45, -20, 38, 20, 11,
					-- layer=2 filter=104 channel=44
					-2, 6, 2, -6, 7, -3, -3, -4, -11,
					-- layer=2 filter=104 channel=45
					21, 25, 1, 63, -18, -7, -66, -27, 8,
					-- layer=2 filter=104 channel=46
					42, 22, 3, 19, 19, -5, -21, -17, -25,
					-- layer=2 filter=104 channel=47
					21, -10, 11, -28, -46, -46, 4, 29, 0,
					-- layer=2 filter=104 channel=48
					9, 6, 6, 10, -7, -9, 1, 4, 6,
					-- layer=2 filter=104 channel=49
					-7, -31, -27, 20, -19, -3, -7, -37, -55,
					-- layer=2 filter=104 channel=50
					6, 5, 23, -16, 2, -17, -13, 11, -8,
					-- layer=2 filter=104 channel=51
					-81, -86, -76, -37, -17, -3, -18, -11, 13,
					-- layer=2 filter=104 channel=52
					-78, -22, 16, -31, 24, -1, -12, -12, 7,
					-- layer=2 filter=104 channel=53
					-39, -30, -60, -3, 9, 5, 13, 60, 1,
					-- layer=2 filter=104 channel=54
					-4, 25, 12, -6, 2, 29, 17, 21, 41,
					-- layer=2 filter=104 channel=55
					16, 4, 9, 12, 4, 10, 2, 13, -5,
					-- layer=2 filter=104 channel=56
					-24, -33, -78, -16, -44, -21, -15, -3, 9,
					-- layer=2 filter=104 channel=57
					0, 4, 6, 16, -17, 1, 10, 8, 0,
					-- layer=2 filter=104 channel=58
					-8, -29, -18, 27, 7, -5, 13, 35, 30,
					-- layer=2 filter=104 channel=59
					-13, 2, 38, -17, 6, -29, 14, 7, 21,
					-- layer=2 filter=104 channel=60
					-17, 15, -31, -23, -14, -12, -26, -46, 3,
					-- layer=2 filter=104 channel=61
					20, -37, -20, -17, -12, -52, -41, -55, -13,
					-- layer=2 filter=104 channel=62
					-46, -50, -29, 10, 17, 23, -7, -15, 55,
					-- layer=2 filter=104 channel=63
					31, 29, 39, -14, -10, -10, -45, -22, 11,
					-- layer=2 filter=104 channel=64
					13, 43, 9, 1, 2, 5, -34, -34, -45,
					-- layer=2 filter=104 channel=65
					-3, -42, -19, 9, 25, -13, -3, -20, 53,
					-- layer=2 filter=104 channel=66
					23, 7, 33, 27, 8, 6, -14, 9, -19,
					-- layer=2 filter=104 channel=67
					25, 9, 7, -20, -16, -3, -6, -26, -40,
					-- layer=2 filter=104 channel=68
					-6, 10, -5, -7, 3, -8, -5, 7, 1,
					-- layer=2 filter=104 channel=69
					38, 48, 46, 0, 10, 5, -12, -20, -41,
					-- layer=2 filter=104 channel=70
					18, 0, -12, -7, -4, -22, 14, 37, 12,
					-- layer=2 filter=104 channel=71
					-12, 28, -69, 23, 23, -84, 18, 17, 4,
					-- layer=2 filter=104 channel=72
					43, -17, 42, 5, -13, -21, -15, -19, 12,
					-- layer=2 filter=104 channel=73
					-5, -24, -37, 68, -52, 37, 13, 11, 0,
					-- layer=2 filter=104 channel=74
					29, 27, 20, 3, -3, -11, -42, -44, -15,
					-- layer=2 filter=104 channel=75
					4, -26, -13, -20, 3, 2, 29, 4, 24,
					-- layer=2 filter=104 channel=76
					-16, -44, -19, 23, -50, 8, -21, 0, 0,
					-- layer=2 filter=104 channel=77
					6, 8, -1, 0, -7, 7, -1, -4, 0,
					-- layer=2 filter=104 channel=78
					-64, -70, -71, -27, -19, 7, -16, -46, 0,
					-- layer=2 filter=104 channel=79
					-4, 7, -2, -8, 7, -8, 8, 0, -3,
					-- layer=2 filter=104 channel=80
					24, 13, 26, 3, 4, 25, 9, 16, -6,
					-- layer=2 filter=104 channel=81
					7, -6, 7, 8, 8, -2, -6, 4, 4,
					-- layer=2 filter=104 channel=82
					-2, -5, -8, 7, 7, 6, 9, 0, 4,
					-- layer=2 filter=104 channel=83
					13, 22, 11, -6, -33, -10, 6, 8, -1,
					-- layer=2 filter=104 channel=84
					2, -3, -3, -7, -2, 11, -7, 7, 11,
					-- layer=2 filter=104 channel=85
					11, -9, -4, 8, -1, 4, -9, 3, 6,
					-- layer=2 filter=104 channel=86
					6, -11, -9, 14, -12, -19, -12, 12, 1,
					-- layer=2 filter=104 channel=87
					-3, 30, -6, -18, 77, 7, 11, 25, 5,
					-- layer=2 filter=104 channel=88
					43, 46, 15, 21, 13, -20, -12, -16, -37,
					-- layer=2 filter=104 channel=89
					6, -10, 20, 8, 15, -1, 34, 9, 6,
					-- layer=2 filter=104 channel=90
					-4, -2, 5, -4, 6, 10, 9, 8, 7,
					-- layer=2 filter=104 channel=91
					12, -9, -2, 11, -5, -15, 5, 0, 16,
					-- layer=2 filter=104 channel=92
					13, 0, 12, 13, 11, -6, 13, -14, -11,
					-- layer=2 filter=104 channel=93
					-54, -58, -52, -38, 37, 10, 17, -5, 73,
					-- layer=2 filter=104 channel=94
					32, -65, 5, 5, 59, 2, -2, -19, 49,
					-- layer=2 filter=104 channel=95
					0, -3, -1, -2, -10, -6, -13, 0, 0,
					-- layer=2 filter=104 channel=96
					-11, -55, 13, -28, 24, 72, -1, 10, 41,
					-- layer=2 filter=104 channel=97
					-7, 23, 9, -22, -24, -17, -8, 17, 5,
					-- layer=2 filter=104 channel=98
					5, -49, -7, 1, -18, -39, 16, 17, -11,
					-- layer=2 filter=104 channel=99
					-65, -46, 21, -4, -26, -5, 4, -24, 1,
					-- layer=2 filter=104 channel=100
					13, 45, 42, -19, 12, 0, -6, -9, 11,
					-- layer=2 filter=104 channel=101
					-16, -17, -42, 64, 41, -39, 14, 45, 64,
					-- layer=2 filter=104 channel=102
					3, -54, -12, 5, 10, 13, -16, -11, 3,
					-- layer=2 filter=104 channel=103
					-42, -23, -51, -33, 0, -9, 10, -40, -11,
					-- layer=2 filter=104 channel=104
					7, -36, -51, -19, 7, 1, -28, -28, 0,
					-- layer=2 filter=104 channel=105
					-66, -14, 23, 40, 36, 9, -8, -26, 8,
					-- layer=2 filter=104 channel=106
					1, -1, -56, 14, -10, -22, -5, 38, 28,
					-- layer=2 filter=104 channel=107
					79, 8, 12, 17, 25, 14, -40, -18, -22,
					-- layer=2 filter=104 channel=108
					30, -4, -33, -8, -53, 20, -1, -23, -7,
					-- layer=2 filter=104 channel=109
					12, -5, 7, 8, 8, -5, 19, 9, -5,
					-- layer=2 filter=104 channel=110
					-6, 13, 10, -40, -36, -38, -26, -40, -61,
					-- layer=2 filter=104 channel=111
					3, -3, 6, 6, 8, 8, 7, -8, 6,
					-- layer=2 filter=104 channel=112
					-52, -87, -64, 4, -7, -21, -6, 24, -2,
					-- layer=2 filter=104 channel=113
					40, 17, 9, 26, 1, -21, 17, -29, -17,
					-- layer=2 filter=104 channel=114
					-20, -10, -12, -11, 1, 10, -12, -8, 13,
					-- layer=2 filter=104 channel=115
					3, 3, -1, 7, 0, 4, 6, -7, 0,
					-- layer=2 filter=104 channel=116
					8, -20, -51, 7, 51, 19, 1, -5, 12,
					-- layer=2 filter=104 channel=117
					29, -65, 9, 34, 10, 11, 27, 12, 5,
					-- layer=2 filter=104 channel=118
					-20, -21, -49, -3, 3, 7, 12, -15, 13,
					-- layer=2 filter=104 channel=119
					14, 56, 30, -39, 21, -17, 29, 29, -11,
					-- layer=2 filter=104 channel=120
					7, -3, 3, 8, -7, -1, -2, 1, -5,
					-- layer=2 filter=104 channel=121
					-7, 3, -6, 10, -3, 0, 9, 3, 6,
					-- layer=2 filter=104 channel=122
					4, -10, 0, -7, -6, -4, 9, 1, -4,
					-- layer=2 filter=104 channel=123
					17, -6, 57, 5, 8, -18, 3, -9, 10,
					-- layer=2 filter=104 channel=124
					-11, 12, 30, 4, 27, -18, 12, 42, 23,
					-- layer=2 filter=104 channel=125
					-1, -4, -5, 0, 1, 2, -8, -3, -2,
					-- layer=2 filter=104 channel=126
					26, -16, -24, 3, 32, -21, -35, 66, 14,
					-- layer=2 filter=104 channel=127
					38, 36, 29, 12, -19, -18, -39, -17, 29,
					-- layer=2 filter=105 channel=0
					-28, -22, 6, -16, -21, -25, -1, -30, -8,
					-- layer=2 filter=105 channel=1
					-11, -12, -31, -7, -9, -12, -17, 0, 15,
					-- layer=2 filter=105 channel=2
					-7, -8, -8, -2, 5, -1, -4, -8, 6,
					-- layer=2 filter=105 channel=3
					-19, 11, -5, -29, -10, -1, -4, -22, -21,
					-- layer=2 filter=105 channel=4
					14, -15, -11, 12, 17, -28, -16, -11, -18,
					-- layer=2 filter=105 channel=5
					-3, 0, -23, -3, -2, -15, -16, -8, -26,
					-- layer=2 filter=105 channel=6
					-11, -10, -4, -1, 14, -11, -1, -20, -7,
					-- layer=2 filter=105 channel=7
					-1, -23, 31, -21, -6, -17, -11, -3, 4,
					-- layer=2 filter=105 channel=8
					-5, 7, 9, 2, -3, -1, -6, 8, -8,
					-- layer=2 filter=105 channel=9
					-22, -2, -19, -24, -3, -5, -6, 9, -11,
					-- layer=2 filter=105 channel=10
					-3, -1, -3, -14, -1, -4, -2, -19, -21,
					-- layer=2 filter=105 channel=11
					-19, -21, -16, -15, -16, -17, -19, -11, -26,
					-- layer=2 filter=105 channel=12
					-21, -20, -37, 2, -1, -18, -1, 17, 23,
					-- layer=2 filter=105 channel=13
					9, -6, -2, 7, 5, -4, -3, 1, -5,
					-- layer=2 filter=105 channel=14
					-29, -29, -25, -17, -7, -12, -21, -1, 0,
					-- layer=2 filter=105 channel=15
					23, -21, -12, 17, -7, -7, -7, 1, -17,
					-- layer=2 filter=105 channel=16
					-27, -16, -20, -31, -14, -13, -13, -20, -5,
					-- layer=2 filter=105 channel=17
					4, -5, 4, -2, 3, -2, -10, 8, 0,
					-- layer=2 filter=105 channel=18
					13, -6, -1, 9, 13, -12, -23, 6, -13,
					-- layer=2 filter=105 channel=19
					-7, 2, 14, -1, -6, -11, 0, -9, 5,
					-- layer=2 filter=105 channel=20
					0, 5, -9, -1, 1, 4, 8, -2, 3,
					-- layer=2 filter=105 channel=21
					-7, 1, -5, -6, -6, 3, -8, 8, 3,
					-- layer=2 filter=105 channel=22
					-6, -7, 1, 1, 10, 0, -6, -2, 9,
					-- layer=2 filter=105 channel=23
					-7, -29, -15, -10, -26, -17, -5, -13, -14,
					-- layer=2 filter=105 channel=24
					-7, 0, 8, -25, -7, -5, -21, -3, -8,
					-- layer=2 filter=105 channel=25
					-13, -19, -13, -19, -12, -11, -18, -12, -2,
					-- layer=2 filter=105 channel=26
					3, -4, 6, 0, 0, -4, 1, 5, 8,
					-- layer=2 filter=105 channel=27
					-14, -10, -19, -26, -11, -20, -7, -16, -11,
					-- layer=2 filter=105 channel=28
					-32, -11, -17, -23, -13, 0, -16, -16, -19,
					-- layer=2 filter=105 channel=29
					-8, -2, -8, 7, -1, -10, 0, -8, -10,
					-- layer=2 filter=105 channel=30
					-10, 0, -7, 7, -8, 15, -18, -12, -8,
					-- layer=2 filter=105 channel=31
					-5, 23, 4, -3, 10, -9, 6, 6, 9,
					-- layer=2 filter=105 channel=32
					-9, 11, 12, 1, 8, 8, 5, 2, 10,
					-- layer=2 filter=105 channel=33
					-14, -10, -18, -22, -13, 7, -10, 1, -6,
					-- layer=2 filter=105 channel=34
					-14, 8, 4, 0, 14, 7, -22, -12, -15,
					-- layer=2 filter=105 channel=35
					0, -12, 3, -27, -26, 2, -25, -22, 0,
					-- layer=2 filter=105 channel=36
					0, 4, -2, -3, -2, -8, -9, 1, -6,
					-- layer=2 filter=105 channel=37
					-9, -15, -18, -22, -20, -12, -14, -3, -30,
					-- layer=2 filter=105 channel=38
					-21, -8, -25, -27, -15, -4, -11, -18, -9,
					-- layer=2 filter=105 channel=39
					-28, -31, -12, -19, -2, -6, -11, -13, -2,
					-- layer=2 filter=105 channel=40
					10, -2, 12, 4, 24, -9, -1, 0, -19,
					-- layer=2 filter=105 channel=41
					9, -5, 0, 10, -6, 4, 0, 3, 5,
					-- layer=2 filter=105 channel=42
					-35, -20, -1, -19, 15, -34, 0, -1, 3,
					-- layer=2 filter=105 channel=43
					-18, 11, 0, -3, 8, -12, -15, -11, -20,
					-- layer=2 filter=105 channel=44
					2, 3, -8, -5, 3, 1, 5, -3, 4,
					-- layer=2 filter=105 channel=45
					-13, -7, -17, -12, -8, -13, 12, -14, -15,
					-- layer=2 filter=105 channel=46
					1, 10, 0, -3, 0, 16, -20, -32, -30,
					-- layer=2 filter=105 channel=47
					-14, -6, -23, -8, -15, -5, -20, -2, -26,
					-- layer=2 filter=105 channel=48
					6, -5, 9, 4, -7, -8, -10, -9, 7,
					-- layer=2 filter=105 channel=49
					24, 0, 0, 30, 20, -19, 4, 22, -14,
					-- layer=2 filter=105 channel=50
					-9, 5, 1, 7, -5, 2, 9, -4, -7,
					-- layer=2 filter=105 channel=51
					-26, 2, -12, -15, -3, -22, -8, -7, -22,
					-- layer=2 filter=105 channel=52
					-18, -7, -18, 9, 3, -15, -2, 2, -1,
					-- layer=2 filter=105 channel=53
					4, 5, 6, 25, 15, -29, 10, -11, -32,
					-- layer=2 filter=105 channel=54
					-4, -25, -6, 6, -4, -22, 10, -10, -8,
					-- layer=2 filter=105 channel=55
					-4, 4, 2, 6, -7, -4, 0, 1, -3,
					-- layer=2 filter=105 channel=56
					-8, -18, -5, -27, -3, -24, -15, -11, -30,
					-- layer=2 filter=105 channel=57
					3, -1, 1, 2, -3, -5, -11, 4, 3,
					-- layer=2 filter=105 channel=58
					-18, -30, -16, -15, -2, -11, -30, 0, 34,
					-- layer=2 filter=105 channel=59
					0, 3, -4, 1, -13, -32, -16, -6, 20,
					-- layer=2 filter=105 channel=60
					-26, -14, -24, -4, -15, 2, -15, -19, 7,
					-- layer=2 filter=105 channel=61
					-11, -16, 4, -31, -27, -8, 19, -22, -21,
					-- layer=2 filter=105 channel=62
					13, 2, -2, 0, 0, 0, -5, 2, -11,
					-- layer=2 filter=105 channel=63
					-28, -17, -9, -21, -25, 6, -8, -19, -17,
					-- layer=2 filter=105 channel=64
					-16, -1, -1, -20, -3, -1, -12, -4, -23,
					-- layer=2 filter=105 channel=65
					-23, 18, -20, -13, -12, 23, -7, -33, -5,
					-- layer=2 filter=105 channel=66
					-10, -17, -11, 6, 17, 15, -18, -5, 1,
					-- layer=2 filter=105 channel=67
					-5, -11, -13, 0, -11, -2, -6, -15, -7,
					-- layer=2 filter=105 channel=68
					-10, -5, 2, 3, -4, -5, 1, 8, 7,
					-- layer=2 filter=105 channel=69
					-17, -27, -24, -33, -20, -14, -30, -25, -1,
					-- layer=2 filter=105 channel=70
					-9, -19, -11, -18, -27, 20, -17, -11, -10,
					-- layer=2 filter=105 channel=71
					-10, -9, -23, -25, -15, -9, -17, -21, -10,
					-- layer=2 filter=105 channel=72
					-10, -11, -3, -23, -21, -16, -7, -27, -16,
					-- layer=2 filter=105 channel=73
					7, -15, 15, 5, -2, 0, 15, -10, -5,
					-- layer=2 filter=105 channel=74
					-6, -3, -6, 5, 16, -8, -3, -5, -13,
					-- layer=2 filter=105 channel=75
					-10, 0, -16, -2, -37, -26, -5, 4, 0,
					-- layer=2 filter=105 channel=76
					1, -16, 9, 17, -20, -8, 2, 15, -32,
					-- layer=2 filter=105 channel=77
					-10, 7, 3, -10, -6, -8, 6, 2, -9,
					-- layer=2 filter=105 channel=78
					-12, -5, -9, -10, 4, -23, -11, -9, -19,
					-- layer=2 filter=105 channel=79
					-6, 1, -7, -2, -9, 7, 5, -2, 9,
					-- layer=2 filter=105 channel=80
					-19, 17, -11, -14, 30, -8, -5, -1, -20,
					-- layer=2 filter=105 channel=81
					7, 0, 3, -5, -7, -6, -10, -4, -3,
					-- layer=2 filter=105 channel=82
					10, 0, -6, 1, 7, -7, 7, -8, 8,
					-- layer=2 filter=105 channel=83
					-13, -32, -28, -4, -28, -16, 1, -17, -17,
					-- layer=2 filter=105 channel=84
					2, -7, 1, 7, -9, -10, 2, -7, 0,
					-- layer=2 filter=105 channel=85
					0, 6, -2, -9, 8, 0, -6, 3, 7,
					-- layer=2 filter=105 channel=86
					0, 6, 0, 1, 8, -3, -1, -7, -1,
					-- layer=2 filter=105 channel=87
					-5, -6, 3, -8, -11, 1, -14, 5, -14,
					-- layer=2 filter=105 channel=88
					-10, -9, -25, -12, 0, -13, -2, -8, -13,
					-- layer=2 filter=105 channel=89
					-3, -5, -21, -20, -16, -25, -21, -11, 22,
					-- layer=2 filter=105 channel=90
					2, 6, 10, -3, -7, 0, -2, -6, 7,
					-- layer=2 filter=105 channel=91
					-30, -34, -37, 0, -23, -24, -35, 6, 21,
					-- layer=2 filter=105 channel=92
					-26, -28, -31, -21, 2, -10, -30, 1, 27,
					-- layer=2 filter=105 channel=93
					7, 23, -5, 16, 2, 23, 2, -15, 9,
					-- layer=2 filter=105 channel=94
					8, -25, 30, 7, -9, -7, 32, -9, -25,
					-- layer=2 filter=105 channel=95
					-1, -3, 4, -9, 5, 6, -9, 1, 0,
					-- layer=2 filter=105 channel=96
					0, -20, -21, -6, -24, -24, -2, -6, -3,
					-- layer=2 filter=105 channel=97
					-25, -8, -2, -29, -12, -15, -20, -4, -16,
					-- layer=2 filter=105 channel=98
					-26, -1, 4, -7, -14, 0, -7, -5, -23,
					-- layer=2 filter=105 channel=99
					-10, 7, -4, -2, -36, -10, 4, -6, -4,
					-- layer=2 filter=105 channel=100
					-25, -10, -13, -23, -3, -48, -8, -18, -5,
					-- layer=2 filter=105 channel=101
					-14, -24, -13, -13, -23, -2, -10, -4, 7,
					-- layer=2 filter=105 channel=102
					14, -3, -27, -2, -16, -21, -16, -5, -4,
					-- layer=2 filter=105 channel=103
					14, -24, -4, -11, 9, -6, -5, 57, 14,
					-- layer=2 filter=105 channel=104
					14, 15, -2, 26, 26, -12, 8, 24, -21,
					-- layer=2 filter=105 channel=105
					0, -29, 34, 2, -16, -4, -21, -2, 4,
					-- layer=2 filter=105 channel=106
					-9, -22, -15, -1, -24, 0, -22, 2, 4,
					-- layer=2 filter=105 channel=107
					-38, -13, 1, 29, -11, -26, 10, 4, -5,
					-- layer=2 filter=105 channel=108
					-11, -20, -22, -7, -18, -12, 3, 12, -19,
					-- layer=2 filter=105 channel=109
					-1, 9, -2, 3, 1, 9, 6, 5, -2,
					-- layer=2 filter=105 channel=110
					-17, -17, -2, -25, -21, 3, -17, -18, -11,
					-- layer=2 filter=105 channel=111
					-1, 7, 5, -3, 6, 10, 9, 4, -5,
					-- layer=2 filter=105 channel=112
					-7, -12, 7, -26, -34, 5, -28, -20, -7,
					-- layer=2 filter=105 channel=113
					-24, 12, -12, -4, -18, 29, -8, -22, 12,
					-- layer=2 filter=105 channel=114
					-4, -8, 0, 3, 5, -10, -6, 3, -2,
					-- layer=2 filter=105 channel=115
					-8, 10, 0, 7, 7, 7, 6, 4, 2,
					-- layer=2 filter=105 channel=116
					20, -9, 0, 13, -6, -2, -14, 10, -13,
					-- layer=2 filter=105 channel=117
					-4, -21, 28, -21, -4, -18, 18, 9, 8,
					-- layer=2 filter=105 channel=118
					4, 0, 1, 0, 14, -14, -14, -7, -23,
					-- layer=2 filter=105 channel=119
					4, -7, -24, 5, -10, -1, -25, -13, -7,
					-- layer=2 filter=105 channel=120
					-6, 5, -9, 0, -2, -3, -8, -9, -7,
					-- layer=2 filter=105 channel=121
					0, -7, 5, 5, -4, -4, -11, -3, 2,
					-- layer=2 filter=105 channel=122
					-2, -6, 4, 0, 3, 3, 8, -1, -3,
					-- layer=2 filter=105 channel=123
					-5, -4, -7, -8, -11, 0, -22, -30, 23,
					-- layer=2 filter=105 channel=124
					8, -27, -5, -1, 13, -3, -4, 5, 18,
					-- layer=2 filter=105 channel=125
					-3, -3, -6, -5, -2, 7, 6, 7, -9,
					-- layer=2 filter=105 channel=126
					-26, -18, 8, -15, 7, -14, 0, -4, -7,
					-- layer=2 filter=105 channel=127
					-30, -9, -35, 0, -20, 18, -6, -13, 0,
					-- layer=2 filter=106 channel=0
					21, -1, 21, 27, 0, 10, -23, 6, 1,
					-- layer=2 filter=106 channel=1
					-3, -8, 26, 5, 30, 2, -28, 2, -15,
					-- layer=2 filter=106 channel=2
					2, -1, 1, -5, -6, 3, 7, -3, -2,
					-- layer=2 filter=106 channel=3
					-39, -22, -64, -21, 1, -39, 46, 65, 62,
					-- layer=2 filter=106 channel=4
					4, 13, 11, -8, -18, 17, -23, 0, -13,
					-- layer=2 filter=106 channel=5
					37, 18, 20, 22, -9, -15, 18, 4, -11,
					-- layer=2 filter=106 channel=6
					-7, 20, 43, 43, 19, 40, -12, -80, -27,
					-- layer=2 filter=106 channel=7
					-35, 6, -25, 0, 26, 49, 24, 46, 50,
					-- layer=2 filter=106 channel=8
					-9, -4, -9, 6, 6, 8, -1, 0, 10,
					-- layer=2 filter=106 channel=9
					7, 16, -1, 0, 20, -3, 0, -13, -43,
					-- layer=2 filter=106 channel=10
					-6, 26, -10, -19, -29, -54, 17, 28, 28,
					-- layer=2 filter=106 channel=11
					14, 0, -3, 1, 4, 2, 4, -27, -11,
					-- layer=2 filter=106 channel=12
					-24, 29, 48, 7, 34, 31, 14, 42, 18,
					-- layer=2 filter=106 channel=13
					-2, -7, -7, -3, 5, 0, 7, 0, -8,
					-- layer=2 filter=106 channel=14
					-3, 7, 35, 0, 27, 28, -37, -9, -12,
					-- layer=2 filter=106 channel=15
					0, -4, 14, -77, -16, 23, -11, -4, 40,
					-- layer=2 filter=106 channel=16
					27, 7, -17, -8, 6, 0, -22, -24, -6,
					-- layer=2 filter=106 channel=17
					-7, 0, 6, 3, 9, -2, 10, 8, 1,
					-- layer=2 filter=106 channel=18
					-39, -43, -27, -41, -82, 14, 5, -12, -26,
					-- layer=2 filter=106 channel=19
					23, 20, -23, -3, 4, -12, -7, 14, 4,
					-- layer=2 filter=106 channel=20
					-2, -3, 10, -7, -4, 10, -5, 9, 3,
					-- layer=2 filter=106 channel=21
					14, -3, -3, 6, 9, 8, 6, 0, -5,
					-- layer=2 filter=106 channel=22
					6, 6, 8, -8, -1, -2, 7, -7, -5,
					-- layer=2 filter=106 channel=23
					-8, 10, 40, -26, -1, 0, 8, 8, -13,
					-- layer=2 filter=106 channel=24
					-11, -13, -31, -37, -28, -76, -12, -12, -19,
					-- layer=2 filter=106 channel=25
					12, 33, 6, 16, -24, -16, -14, -13, 3,
					-- layer=2 filter=106 channel=26
					-6, -10, -8, 8, 3, -7, -7, 0, -8,
					-- layer=2 filter=106 channel=27
					26, 25, 22, -5, 4, -18, -24, -32, -34,
					-- layer=2 filter=106 channel=28
					-15, 11, 5, -33, -28, -36, 4, 25, 18,
					-- layer=2 filter=106 channel=29
					6, -2, 5, -4, -1, 11, 0, 0, 2,
					-- layer=2 filter=106 channel=30
					8, 15, 2, -15, -28, -12, -10, -10, 28,
					-- layer=2 filter=106 channel=31
					-18, -39, 8, -18, -32, -24, -83, -46, -67,
					-- layer=2 filter=106 channel=32
					-4, 1, -8, -5, 10, -7, 1, -7, -2,
					-- layer=2 filter=106 channel=33
					-43, -13, -24, -31, 8, 4, 1, 30, 57,
					-- layer=2 filter=106 channel=34
					0, -11, -15, -51, 1, -32, -13, -35, -69,
					-- layer=2 filter=106 channel=35
					10, 13, 12, -10, 0, 1, 13, 39, 25,
					-- layer=2 filter=106 channel=36
					-7, 6, -1, 6, -6, 2, -4, 12, -1,
					-- layer=2 filter=106 channel=37
					19, 11, 4, 6, -12, 0, 2, -23, -6,
					-- layer=2 filter=106 channel=38
					24, 22, 19, 7, -29, -24, -33, -19, -42,
					-- layer=2 filter=106 channel=39
					0, -10, 12, -50, -3, -15, 4, -24, -45,
					-- layer=2 filter=106 channel=40
					-36, 3, 3, -18, -34, 18, 19, -28, 3,
					-- layer=2 filter=106 channel=41
					10, 6, 3, -6, -6, -7, -2, -4, 6,
					-- layer=2 filter=106 channel=42
					-8, 21, 10, 3, 42, 14, 0, 20, 24,
					-- layer=2 filter=106 channel=43
					25, -14, -23, -18, -13, -11, 44, 37, 34,
					-- layer=2 filter=106 channel=44
					0, 3, -3, -3, -3, -8, -7, 6, -5,
					-- layer=2 filter=106 channel=45
					31, 29, 33, -35, 21, 19, -38, 25, 29,
					-- layer=2 filter=106 channel=46
					24, 2, -18, -24, 34, -21, 6, -15, -20,
					-- layer=2 filter=106 channel=47
					-58, -36, -19, -17, -24, -13, -24, -2, -12,
					-- layer=2 filter=106 channel=48
					5, -5, -4, 4, -3, 4, 2, -8, -8,
					-- layer=2 filter=106 channel=49
					0, 3, -37, -36, -29, 28, -3, -28, -17,
					-- layer=2 filter=106 channel=50
					-2, -10, -3, 8, 9, 20, 0, 10, 18,
					-- layer=2 filter=106 channel=51
					13, 11, 6, 22, -4, 7, 0, -11, -10,
					-- layer=2 filter=106 channel=52
					6, -44, -16, 34, 18, 9, 2, -19, 16,
					-- layer=2 filter=106 channel=53
					-51, 0, -7, 5, 7, -9, -26, -37, -15,
					-- layer=2 filter=106 channel=54
					-55, 0, -12, -5, -22, -6, -19, -15, 23,
					-- layer=2 filter=106 channel=55
					0, 4, 5, 4, -5, -7, 2, 6, -4,
					-- layer=2 filter=106 channel=56
					37, 6, 24, 20, -21, -3, 14, -25, -24,
					-- layer=2 filter=106 channel=57
					-4, -6, -9, 6, 7, 3, -6, -6, -2,
					-- layer=2 filter=106 channel=58
					-11, 15, 62, 5, 32, 11, 0, 15, 35,
					-- layer=2 filter=106 channel=59
					16, -19, -15, 8, -7, -22, 3, 3, -25,
					-- layer=2 filter=106 channel=60
					-2, -24, -16, 27, 7, -5, 5, -24, -35,
					-- layer=2 filter=106 channel=61
					-51, -55, -98, 29, -39, 10, 7, -54, -32,
					-- layer=2 filter=106 channel=62
					5, -1, -12, 25, 8, 37, -35, -51, -37,
					-- layer=2 filter=106 channel=63
					14, -17, -15, 15, 5, 4, 3, 5, -17,
					-- layer=2 filter=106 channel=64
					-11, 0, -12, -17, -13, -4, -46, -23, -38,
					-- layer=2 filter=106 channel=65
					-19, -20, -70, 36, -5, 9, -12, -61, -57,
					-- layer=2 filter=106 channel=66
					-32, 27, -39, 43, 8, 28, -7, 42, -33,
					-- layer=2 filter=106 channel=67
					33, -3, -34, 9, 12, -70, -10, -31, -36,
					-- layer=2 filter=106 channel=68
					-4, 5, -2, 4, 1, -2, 5, 7, 8,
					-- layer=2 filter=106 channel=69
					-1, 0, -10, -14, 32, 19, -22, -2, -11,
					-- layer=2 filter=106 channel=70
					-7, 25, 29, -26, -36, -5, 12, 30, 31,
					-- layer=2 filter=106 channel=71
					43, 38, 12, 1, 19, 5, -31, -34, -33,
					-- layer=2 filter=106 channel=72
					-10, -3, -22, -2, 6, 30, 4, 60, 42,
					-- layer=2 filter=106 channel=73
					-21, -11, -37, -6, 7, -20, -38, -23, -32,
					-- layer=2 filter=106 channel=74
					9, 0, -1, 3, -11, -24, 8, -23, -49,
					-- layer=2 filter=106 channel=75
					-38, -11, 2, -17, 27, -20, -46, 12, -1,
					-- layer=2 filter=106 channel=76
					-73, -59, -40, 29, -30, 5, -12, -40, -70,
					-- layer=2 filter=106 channel=77
					-2, 6, -6, -6, 0, -8, 2, 4, -1,
					-- layer=2 filter=106 channel=78
					10, -28, -41, 8, -16, -9, -23, -23, -4,
					-- layer=2 filter=106 channel=79
					7, -5, 0, 0, -9, 6, 0, 4, -8,
					-- layer=2 filter=106 channel=80
					12, -14, -22, -32, -2, -21, 3, 0, 9,
					-- layer=2 filter=106 channel=81
					13, 5, -5, -2, 3, 8, 5, 5, -2,
					-- layer=2 filter=106 channel=82
					-2, -7, -7, 5, 5, 9, -6, -7, -7,
					-- layer=2 filter=106 channel=83
					8, 36, 19, -42, 3, -5, 7, 15, 8,
					-- layer=2 filter=106 channel=84
					-3, 0, 7, 4, 7, -5, -10, -5, 4,
					-- layer=2 filter=106 channel=85
					2, 1, 11, 6, 5, 9, -5, 16, 8,
					-- layer=2 filter=106 channel=86
					-6, 6, -17, 13, -5, 21, -3, -10, 5,
					-- layer=2 filter=106 channel=87
					-13, -30, -17, 10, -22, 41, 10, -35, -12,
					-- layer=2 filter=106 channel=88
					10, 17, 5, 10, -2, 12, 1, 25, -15,
					-- layer=2 filter=106 channel=89
					-8, 11, 7, 6, 22, 26, -4, 27, 24,
					-- layer=2 filter=106 channel=90
					-7, 0, 0, 2, -3, 0, 7, -2, 1,
					-- layer=2 filter=106 channel=91
					-4, 8, 34, 0, 30, 23, -7, 54, 29,
					-- layer=2 filter=106 channel=92
					-2, 26, 38, 2, 30, 13, 13, 31, 12,
					-- layer=2 filter=106 channel=93
					1, -30, -54, 46, 71, 33, 8, 3, -2,
					-- layer=2 filter=106 channel=94
					-16, 3, -1, 48, 1, -5, 18, -11, -2,
					-- layer=2 filter=106 channel=95
					11, -1, 1, 6, 0, -8, -1, -8, 4,
					-- layer=2 filter=106 channel=96
					45, 30, 13, 40, 19, 48, -35, 3, -57,
					-- layer=2 filter=106 channel=97
					-12, -14, -2, -26, 13, -11, -37, 13, -17,
					-- layer=2 filter=106 channel=98
					-34, 0, -34, -18, -22, -14, -2, 23, 9,
					-- layer=2 filter=106 channel=99
					-9, -6, -28, -4, 27, -13, -17, -37, -56,
					-- layer=2 filter=106 channel=100
					13, 29, 23, -7, -22, -27, 4, -10, 20,
					-- layer=2 filter=106 channel=101
					33, 42, -2, 3, 3, 25, 6, -16, 19,
					-- layer=2 filter=106 channel=102
					-5, 30, 8, 12, -7, 12, -7, 22, -58,
					-- layer=2 filter=106 channel=103
					-33, 1, 29, 38, 34, 2, 0, 3, -40,
					-- layer=2 filter=106 channel=104
					-1, 14, -18, 7, -43, 3, 5, -10, 6,
					-- layer=2 filter=106 channel=105
					-28, -9, -43, 36, -49, 9, 23, -40, -31,
					-- layer=2 filter=106 channel=106
					-1, 4, 16, 9, 2, 2, -7, -10, 1,
					-- layer=2 filter=106 channel=107
					15, -5, -26, 65, 14, -22, 19, 23, 8,
					-- layer=2 filter=106 channel=108
					17, 16, 4, -3, 10, 12, -35, -49, -69,
					-- layer=2 filter=106 channel=109
					-1, 0, 8, 4, -4, 10, 4, -7, -4,
					-- layer=2 filter=106 channel=110
					36, 44, -18, -8, 30, 7, 15, -11, 4,
					-- layer=2 filter=106 channel=111
					11, -2, 0, 1, 8, 2, 1, -1, -7,
					-- layer=2 filter=106 channel=112
					-14, -7, -39, 10, 12, -13, -8, 5, -17,
					-- layer=2 filter=106 channel=113
					-5, 1, -10, -21, 0, -45, -17, 9, 16,
					-- layer=2 filter=106 channel=114
					-10, 0, 4, -8, -1, -3, -7, -8, -12,
					-- layer=2 filter=106 channel=115
					6, 0, 2, -2, -5, -8, 7, -2, -14,
					-- layer=2 filter=106 channel=116
					-8, 0, -17, 0, -28, 24, 24, -28, -34,
					-- layer=2 filter=106 channel=117
					-39, 13, -23, 16, 18, 22, 25, 31, 38,
					-- layer=2 filter=106 channel=118
					-11, -32, -43, -14, -13, -17, 18, 23, 45,
					-- layer=2 filter=106 channel=119
					-21, -3, 5, -29, -34, 1, 38, -8, -39,
					-- layer=2 filter=106 channel=120
					0, 5, -4, -4, 3, 2, 6, 2, -3,
					-- layer=2 filter=106 channel=121
					6, 3, -7, 11, -4, 2, -4, 10, 9,
					-- layer=2 filter=106 channel=122
					8, -11, -6, 3, -4, 10, 0, -1, -8,
					-- layer=2 filter=106 channel=123
					-49, -18, -42, -1, -1, 19, -7, 36, 19,
					-- layer=2 filter=106 channel=124
					-59, -47, -58, -37, -3, 9, -33, 35, 26,
					-- layer=2 filter=106 channel=125
					-4, 0, -3, 4, 11, 4, -6, -1, 7,
					-- layer=2 filter=106 channel=126
					-78, -61, -28, -28, 46, 24, 20, 67, -47,
					-- layer=2 filter=106 channel=127
					14, -3, 18, -5, 15, -18, -3, 9, -11,
					-- layer=2 filter=107 channel=0
					-4, -15, 0, -10, 0, -4, -7, -10, 0,
					-- layer=2 filter=107 channel=1
					0, -6, -4, 3, -4, -9, -5, -3, -9,
					-- layer=2 filter=107 channel=2
					-7, 0, -3, 3, -2, -6, -9, 2, 5,
					-- layer=2 filter=107 channel=3
					3, -2, 0, -7, -10, -7, -7, -11, 5,
					-- layer=2 filter=107 channel=4
					-1, -12, -5, -17, 0, -3, -1, -8, -3,
					-- layer=2 filter=107 channel=5
					-9, -12, -6, -12, 0, 1, -10, 4, 0,
					-- layer=2 filter=107 channel=6
					-3, -4, 0, 6, -11, -10, -9, -9, -3,
					-- layer=2 filter=107 channel=7
					-3, 1, -10, 4, 4, 5, -1, -4, 10,
					-- layer=2 filter=107 channel=8
					1, -1, 8, -8, -6, 3, 0, -5, -1,
					-- layer=2 filter=107 channel=9
					-5, 2, -10, 1, -3, 3, 1, -4, -10,
					-- layer=2 filter=107 channel=10
					6, -2, 0, -11, 1, 1, -8, 1, -14,
					-- layer=2 filter=107 channel=11
					-11, -7, -14, -1, -8, -13, -1, -2, -8,
					-- layer=2 filter=107 channel=12
					7, -2, 6, -2, -6, -12, -12, -6, 7,
					-- layer=2 filter=107 channel=13
					7, -1, 8, -5, 6, -5, -6, -5, -7,
					-- layer=2 filter=107 channel=14
					-9, -11, 1, -5, -11, -11, -11, 0, 0,
					-- layer=2 filter=107 channel=15
					-7, 1, -5, -11, 3, 5, -3, -4, 0,
					-- layer=2 filter=107 channel=16
					7, 4, 5, -6, 4, -4, -9, 0, -1,
					-- layer=2 filter=107 channel=17
					9, -2, -8, 9, -9, 4, 0, -1, 8,
					-- layer=2 filter=107 channel=18
					0, 3, -9, -8, 8, 7, -14, -10, 0,
					-- layer=2 filter=107 channel=19
					7, -6, -3, -10, 4, -11, -6, -2, 8,
					-- layer=2 filter=107 channel=20
					0, 0, 6, -9, 1, -8, -10, -2, -5,
					-- layer=2 filter=107 channel=21
					4, 0, -1, 0, 3, 1, -4, -1, 3,
					-- layer=2 filter=107 channel=22
					-6, 7, -4, 9, -8, 5, 4, 7, 1,
					-- layer=2 filter=107 channel=23
					8, -7, -4, -1, -3, 3, 2, -1, -3,
					-- layer=2 filter=107 channel=24
					0, -2, 3, -3, -11, -7, 1, -9, -4,
					-- layer=2 filter=107 channel=25
					2, 0, 4, -9, -9, 1, 8, 6, 2,
					-- layer=2 filter=107 channel=26
					-2, 7, 9, -3, -5, -3, -3, -5, 0,
					-- layer=2 filter=107 channel=27
					-9, -1, -2, -5, -2, -1, -2, -15, -14,
					-- layer=2 filter=107 channel=28
					-7, -12, -2, -4, -10, -7, 8, -8, 2,
					-- layer=2 filter=107 channel=29
					-4, 2, -2, -4, -10, -1, -11, 0, 3,
					-- layer=2 filter=107 channel=30
					1, -4, -2, -8, -9, -6, -11, 0, 2,
					-- layer=2 filter=107 channel=31
					-6, -10, 0, 4, 3, 6, -7, 2, -4,
					-- layer=2 filter=107 channel=32
					-6, 5, 2, 5, 5, -6, -3, -2, 0,
					-- layer=2 filter=107 channel=33
					6, 7, -12, 0, 0, -8, 0, -3, -1,
					-- layer=2 filter=107 channel=34
					-4, 4, -15, -5, 7, -9, 2, -7, -9,
					-- layer=2 filter=107 channel=35
					-9, -3, -7, -1, -1, 7, 6, -1, 6,
					-- layer=2 filter=107 channel=36
					-1, -7, 3, 3, 2, 4, -6, -2, 3,
					-- layer=2 filter=107 channel=37
					-7, -18, -4, 2, -11, -17, -21, -14, 0,
					-- layer=2 filter=107 channel=38
					-4, -6, -2, -7, 0, -15, -2, 5, -7,
					-- layer=2 filter=107 channel=39
					-2, -1, 8, -9, 0, -12, -1, 4, -12,
					-- layer=2 filter=107 channel=40
					12, -6, 0, 9, 0, -3, 2, 0, 1,
					-- layer=2 filter=107 channel=41
					7, -8, 0, 6, -11, -9, -8, -4, 1,
					-- layer=2 filter=107 channel=42
					-10, -3, -9, -8, -10, 3, -11, -5, 1,
					-- layer=2 filter=107 channel=43
					-12, -3, 9, 3, 6, -4, -7, -4, 6,
					-- layer=2 filter=107 channel=44
					-1, 0, -3, -2, 1, 4, 5, 0, -7,
					-- layer=2 filter=107 channel=45
					0, -5, 1, -9, -4, -5, -7, -6, 6,
					-- layer=2 filter=107 channel=46
					-4, 5, 0, -9, -11, -7, 6, -8, 0,
					-- layer=2 filter=107 channel=47
					-1, -11, 0, -10, 4, 4, -2, -11, 1,
					-- layer=2 filter=107 channel=48
					9, 5, 5, 5, 5, -1, -4, 3, -7,
					-- layer=2 filter=107 channel=49
					-7, 5, 6, -15, 1, -2, -10, 3, -14,
					-- layer=2 filter=107 channel=50
					-2, 7, 1, 9, -4, 2, -2, -7, 9,
					-- layer=2 filter=107 channel=51
					-10, -18, -13, 0, -7, 4, 0, -1, -6,
					-- layer=2 filter=107 channel=52
					1, 6, -17, -1, -4, -14, 1, -8, -8,
					-- layer=2 filter=107 channel=53
					-2, -1, -3, -12, 0, -5, 4, -10, -12,
					-- layer=2 filter=107 channel=54
					-11, -10, 2, -12, 1, 2, -15, 10, -2,
					-- layer=2 filter=107 channel=55
					-2, 0, 8, -2, 10, -2, 1, -9, 2,
					-- layer=2 filter=107 channel=56
					-7, -6, -17, -9, -16, -13, -13, 5, 4,
					-- layer=2 filter=107 channel=57
					-6, -9, 9, -7, 3, 0, 0, -11, 4,
					-- layer=2 filter=107 channel=58
					-5, -12, -6, 0, -12, -7, -1, -7, 0,
					-- layer=2 filter=107 channel=59
					-10, -6, -5, -2, -10, -4, -6, -3, 7,
					-- layer=2 filter=107 channel=60
					4, -6, 2, 1, 2, -5, -4, -3, 6,
					-- layer=2 filter=107 channel=61
					-2, -6, -10, -8, -1, -2, -3, -4, 0,
					-- layer=2 filter=107 channel=62
					0, -2, 3, -3, -1, 0, -5, -9, -7,
					-- layer=2 filter=107 channel=63
					8, -8, 5, -10, 3, 3, 0, 0, 2,
					-- layer=2 filter=107 channel=64
					0, -4, -2, 0, 5, 2, -13, 3, 3,
					-- layer=2 filter=107 channel=65
					-12, -2, 2, -10, -2, -2, -5, -12, -12,
					-- layer=2 filter=107 channel=66
					-4, -12, -10, 0, -4, 5, -9, -11, 1,
					-- layer=2 filter=107 channel=67
					-7, 0, -5, 0, -8, 1, -9, 0, 4,
					-- layer=2 filter=107 channel=68
					0, -1, 3, -7, 0, -10, -11, -7, -11,
					-- layer=2 filter=107 channel=69
					-2, -9, -9, -2, 0, 0, -16, 0, 0,
					-- layer=2 filter=107 channel=70
					1, -9, -7, -6, 0, -8, -8, 0, -9,
					-- layer=2 filter=107 channel=71
					6, 8, -11, 4, 2, 2, -10, -2, 3,
					-- layer=2 filter=107 channel=72
					-3, 3, -10, 4, 7, -1, -12, -15, 4,
					-- layer=2 filter=107 channel=73
					4, 7, -10, -2, 6, -4, -1, 5, -6,
					-- layer=2 filter=107 channel=74
					4, -8, -3, -8, 1, 2, 5, 4, -8,
					-- layer=2 filter=107 channel=75
					2, 10, 10, 5, -12, 1, 2, 0, -3,
					-- layer=2 filter=107 channel=76
					-3, -9, -9, 4, -16, 4, -11, 1, 0,
					-- layer=2 filter=107 channel=77
					-11, -11, -3, -2, -6, 7, 0, 1, -11,
					-- layer=2 filter=107 channel=78
					-13, -14, -11, -4, 4, -10, 2, -12, -10,
					-- layer=2 filter=107 channel=79
					6, 0, 7, 4, -9, -2, -9, 3, 4,
					-- layer=2 filter=107 channel=80
					3, -4, -4, -8, 4, -2, 3, 5, -11,
					-- layer=2 filter=107 channel=81
					-9, -9, -4, -3, -9, 2, -2, 0, 5,
					-- layer=2 filter=107 channel=82
					1, 0, 0, 7, -8, 5, 6, -1, 9,
					-- layer=2 filter=107 channel=83
					6, 0, -5, -2, -14, 0, -4, -9, -1,
					-- layer=2 filter=107 channel=84
					10, 2, 5, 5, 4, -8, -12, -5, 7,
					-- layer=2 filter=107 channel=85
					0, -3, 7, -1, 4, 6, 5, 7, -7,
					-- layer=2 filter=107 channel=86
					-1, -4, -7, -4, -9, 4, 1, -8, 10,
					-- layer=2 filter=107 channel=87
					-12, -8, -11, -11, -4, -3, 6, -2, -9,
					-- layer=2 filter=107 channel=88
					-13, -7, -9, 5, -9, -7, 0, -10, 1,
					-- layer=2 filter=107 channel=89
					-3, -3, -12, -11, 3, -11, -2, 4, 5,
					-- layer=2 filter=107 channel=90
					-1, -6, 8, -7, 9, 4, -3, 8, 9,
					-- layer=2 filter=107 channel=91
					-9, 2, -13, 2, 6, -1, -13, 3, 9,
					-- layer=2 filter=107 channel=92
					-3, -7, -4, 0, -12, -10, 1, 3, 2,
					-- layer=2 filter=107 channel=93
					-4, -19, 0, 4, -8, -2, -10, 6, 5,
					-- layer=2 filter=107 channel=94
					2, -5, 7, 1, -4, -10, -10, -4, -14,
					-- layer=2 filter=107 channel=95
					-8, -9, 0, 0, -9, 6, 1, 4, 7,
					-- layer=2 filter=107 channel=96
					-11, -4, -4, 5, -11, 1, 2, -12, -3,
					-- layer=2 filter=107 channel=97
					-12, -4, -11, -3, 0, 5, 0, 4, -6,
					-- layer=2 filter=107 channel=98
					-10, 5, -2, -4, -8, -2, 0, -5, -15,
					-- layer=2 filter=107 channel=99
					-5, 1, 3, 7, 6, 6, 3, -2, 4,
					-- layer=2 filter=107 channel=100
					-6, -8, 0, 3, -2, -15, -2, -13, -12,
					-- layer=2 filter=107 channel=101
					1, -7, -7, 5, -7, -6, 9, 4, 11,
					-- layer=2 filter=107 channel=102
					-13, 6, 5, 1, -8, 5, -18, -16, 6,
					-- layer=2 filter=107 channel=103
					-11, -3, -8, -5, -2, -7, -8, 1, 2,
					-- layer=2 filter=107 channel=104
					-10, -4, 5, -12, -4, 4, -9, -6, -10,
					-- layer=2 filter=107 channel=105
					8, -4, 6, 2, -7, -11, -6, 4, -6,
					-- layer=2 filter=107 channel=106
					0, 1, -5, 6, -5, -10, 1, -12, -5,
					-- layer=2 filter=107 channel=107
					11, 0, 8, 7, 7, -8, 7, -4, -4,
					-- layer=2 filter=107 channel=108
					-14, 5, -5, -9, 2, 4, 0, -9, -7,
					-- layer=2 filter=107 channel=109
					-9, -11, 0, 2, -10, -4, -10, -12, 3,
					-- layer=2 filter=107 channel=110
					6, -5, 8, 0, -3, 7, -3, -4, 1,
					-- layer=2 filter=107 channel=111
					0, 4, 1, -10, 7, 0, 11, 0, -4,
					-- layer=2 filter=107 channel=112
					7, 4, 0, -4, -8, -1, 7, -5, 0,
					-- layer=2 filter=107 channel=113
					6, 0, 5, 0, -2, -7, -3, 2, -11,
					-- layer=2 filter=107 channel=114
					8, 3, -1, -2, 0, -4, 6, -4, 4,
					-- layer=2 filter=107 channel=115
					-6, -10, -9, -6, 5, -2, 1, -6, -7,
					-- layer=2 filter=107 channel=116
					-10, -12, -9, -14, 4, 7, -2, -3, -1,
					-- layer=2 filter=107 channel=117
					-2, -2, 4, 5, 0, 4, 0, -7, 4,
					-- layer=2 filter=107 channel=118
					-4, -10, 1, 1, -1, -10, -7, 4, -12,
					-- layer=2 filter=107 channel=119
					-13, 4, 1, -6, 4, 4, -4, 0, -4,
					-- layer=2 filter=107 channel=120
					9, -1, -7, -8, 3, -4, 5, 3, 3,
					-- layer=2 filter=107 channel=121
					9, 0, 7, 0, 7, -11, 5, -5, 1,
					-- layer=2 filter=107 channel=122
					1, 3, -3, -10, 6, 0, 6, 8, 8,
					-- layer=2 filter=107 channel=123
					4, 0, -5, 10, -1, 0, 3, -2, -11,
					-- layer=2 filter=107 channel=124
					8, -4, -8, -5, -11, 1, 3, -10, -7,
					-- layer=2 filter=107 channel=125
					7, 6, 3, 0, 0, -2, -9, -9, 4,
					-- layer=2 filter=107 channel=126
					0, 2, 0, 0, 5, -4, -6, -5, -1,
					-- layer=2 filter=107 channel=127
					-6, -2, -2, -6, -18, -9, -14, -9, -7,
					-- layer=2 filter=108 channel=0
					-12, -36, -2, -11, -20, -14, 17, -1, 10,
					-- layer=2 filter=108 channel=1
					-3, -23, -44, 34, -3, -8, -3, -30, 18,
					-- layer=2 filter=108 channel=2
					2, -8, -4, 7, -5, -1, 6, 5, 9,
					-- layer=2 filter=108 channel=3
					-50, -69, -79, -16, -24, 35, 23, -7, -5,
					-- layer=2 filter=108 channel=4
					-28, -24, -32, 23, 11, -34, 28, 16, 2,
					-- layer=2 filter=108 channel=5
					-4, 17, -34, -17, -11, 0, 14, -1, 0,
					-- layer=2 filter=108 channel=6
					15, 12, 10, 32, -15, 37, 25, 15, -8,
					-- layer=2 filter=108 channel=7
					9, -34, -36, 38, -24, -18, 4, -6, 12,
					-- layer=2 filter=108 channel=8
					2, 0, 8, 1, -2, 1, 6, 6, 2,
					-- layer=2 filter=108 channel=9
					-85, -47, -92, -87, -42, -51, 28, 13, -50,
					-- layer=2 filter=108 channel=10
					-4, -50, -67, 0, -28, 17, 46, 0, 50,
					-- layer=2 filter=108 channel=11
					-21, -11, -10, 4, -7, 14, -1, 15, 9,
					-- layer=2 filter=108 channel=12
					11, -29, -36, 0, -31, -10, 15, 5, -9,
					-- layer=2 filter=108 channel=13
					6, -3, 10, 6, 7, 6, -7, -2, 1,
					-- layer=2 filter=108 channel=14
					-44, -61, -30, -18, -21, -26, -4, -7, 12,
					-- layer=2 filter=108 channel=15
					32, 41, 6, 1, 38, -8, 29, 12, 19,
					-- layer=2 filter=108 channel=16
					-6, 24, -53, 24, -22, -62, -74, -76, -36,
					-- layer=2 filter=108 channel=17
					11, -3, 6, -1, 6, -7, 9, 0, -5,
					-- layer=2 filter=108 channel=18
					3, 13, -8, 35, 24, -31, 17, 10, -6,
					-- layer=2 filter=108 channel=19
					42, 14, -46, 46, 40, 19, 0, -13, 20,
					-- layer=2 filter=108 channel=20
					-9, -1, 1, -5, 7, 6, -12, 8, 0,
					-- layer=2 filter=108 channel=21
					-10, -7, -18, -1, 0, -3, -6, -2, 0,
					-- layer=2 filter=108 channel=22
					-4, -5, 4, 4, -7, 3, -4, 2, -8,
					-- layer=2 filter=108 channel=23
					3, 21, -7, -13, -17, 7, 10, -28, 35,
					-- layer=2 filter=108 channel=24
					-29, -35, 1, -4, -48, 22, 30, -4, 33,
					-- layer=2 filter=108 channel=25
					-23, -33, 39, -39, -74, 12, 12, -13, 27,
					-- layer=2 filter=108 channel=26
					-5, 3, 8, 9, -2, -7, -13, 3, 4,
					-- layer=2 filter=108 channel=27
					-21, -12, -22, -10, -8, -17, -23, -5, 9,
					-- layer=2 filter=108 channel=28
					-1, -63, -22, 28, -7, -15, -11, 32, 40,
					-- layer=2 filter=108 channel=29
					2, -9, 4, 0, 7, 3, 8, -8, -11,
					-- layer=2 filter=108 channel=30
					-70, -24, -68, 4, -26, -9, 2, -3, -7,
					-- layer=2 filter=108 channel=31
					-31, 57, -15, 11, 22, -32, 29, -16, -13,
					-- layer=2 filter=108 channel=32
					7, 10, 5, -4, 4, -1, -9, -1, 0,
					-- layer=2 filter=108 channel=33
					-33, -70, -54, -21, -17, -5, 0, 13, 17,
					-- layer=2 filter=108 channel=34
					54, 14, 0, 26, 13, -7, -25, 22, 57,
					-- layer=2 filter=108 channel=35
					-29, -86, -41, -2, -13, -13, 11, 12, 16,
					-- layer=2 filter=108 channel=36
					14, -1, -19, 9, 3, 5, 6, 7, 8,
					-- layer=2 filter=108 channel=37
					-28, 8, 0, 18, 10, 13, -8, 26, 7,
					-- layer=2 filter=108 channel=38
					-67, -26, -19, -7, 3, 6, -32, -21, 10,
					-- layer=2 filter=108 channel=39
					-64, -4, -50, 14, -97, -154, -72, -125, -15,
					-- layer=2 filter=108 channel=40
					-30, 10, 39, -3, -7, -1, 18, 10, -4,
					-- layer=2 filter=108 channel=41
					1, -5, 6, 1, 2, -9, -10, -6, 8,
					-- layer=2 filter=108 channel=42
					-17, 25, -49, -18, -73, -2, 2, -26, -20,
					-- layer=2 filter=108 channel=43
					-53, -43, -54, -24, -24, -3, -8, 8, 31,
					-- layer=2 filter=108 channel=44
					1, 1, -9, -9, 5, -7, -1, -1, 10,
					-- layer=2 filter=108 channel=45
					-16, 22, -38, 18, 26, 3, -14, -12, 2,
					-- layer=2 filter=108 channel=46
					-70, 50, -64, 25, -16, -10, 1, -4, 12,
					-- layer=2 filter=108 channel=47
					49, -52, -18, -14, -36, 13, -16, -1, 33,
					-- layer=2 filter=108 channel=48
					4, 0, 4, -11, -10, 3, -1, 4, 1,
					-- layer=2 filter=108 channel=49
					-4, 0, 4, 65, 9, -9, 24, -22, 3,
					-- layer=2 filter=108 channel=50
					4, 24, 14, 8, 19, 14, 1, 6, -32,
					-- layer=2 filter=108 channel=51
					-6, 0, 20, -8, -2, -4, 0, -1, 6,
					-- layer=2 filter=108 channel=52
					13, 2, 56, 26, 24, 29, 25, 36, -1,
					-- layer=2 filter=108 channel=53
					1, -14, -12, 8, 29, -23, 7, -6, 0,
					-- layer=2 filter=108 channel=54
					42, 10, -5, 33, 0, 0, 23, 14, 16,
					-- layer=2 filter=108 channel=55
					-10, -10, 0, 3, -6, -3, 5, 1, -9,
					-- layer=2 filter=108 channel=56
					-25, -3, -6, -12, -26, -19, -2, -9, 7,
					-- layer=2 filter=108 channel=57
					-18, 0, 22, 9, 10, 18, -1, -11, 4,
					-- layer=2 filter=108 channel=58
					-21, -11, -30, -34, -51, -34, 42, 6, -18,
					-- layer=2 filter=108 channel=59
					-21, -23, 29, 15, 21, -8, -6, -8, 36,
					-- layer=2 filter=108 channel=60
					-11, -3, 21, 11, 19, 33, 8, -7, 35,
					-- layer=2 filter=108 channel=61
					7, -6, 46, 13, -19, 15, 3, -9, 37,
					-- layer=2 filter=108 channel=62
					16, -3, -32, 21, 20, 3, -22, -16, -14,
					-- layer=2 filter=108 channel=63
					-52, 18, -18, -14, 34, -6, -25, 9, 18,
					-- layer=2 filter=108 channel=64
					15, 10, 10, 2, 1, 0, 6, 3, -3,
					-- layer=2 filter=108 channel=65
					-19, -11, 28, -5, 9, 34, 5, -3, -17,
					-- layer=2 filter=108 channel=66
					25, 7, -17, 3, -39, -21, 53, 20, -22,
					-- layer=2 filter=108 channel=67
					-12, 11, -60, -22, -37, -26, -1, -17, -32,
					-- layer=2 filter=108 channel=68
					-2, 2, -4, 5, -3, -10, -8, -11, -3,
					-- layer=2 filter=108 channel=69
					5, 5, -23, 18, -18, -21, 11, -52, -30,
					-- layer=2 filter=108 channel=70
					1, -41, -35, 13, 15, 9, -1, 31, 8,
					-- layer=2 filter=108 channel=71
					-9, 2, -12, -1, -35, -26, -12, -27, 29,
					-- layer=2 filter=108 channel=72
					10, -21, -23, 21, -21, 7, -11, 3, 15,
					-- layer=2 filter=108 channel=73
					24, 50, 16, 21, 29, 0, 48, 3, 14,
					-- layer=2 filter=108 channel=74
					-104, -33, -86, -55, -16, -31, 15, 48, 35,
					-- layer=2 filter=108 channel=75
					-7, -43, -67, -33, -48, -38, -46, 70, -30,
					-- layer=2 filter=108 channel=76
					-21, 17, -3, 48, 10, 5, 28, -10, 20,
					-- layer=2 filter=108 channel=77
					2, -2, 0, -2, 5, -12, -2, -11, 7,
					-- layer=2 filter=108 channel=78
					0, 22, -10, 17, -1, 27, 20, 14, -4,
					-- layer=2 filter=108 channel=79
					2, -8, 4, 8, -11, -5, -7, 2, -8,
					-- layer=2 filter=108 channel=80
					-63, 0, -29, -11, -26, 36, 12, 21, 6,
					-- layer=2 filter=108 channel=81
					0, -8, -1, -4, -2, -12, -14, -8, -9,
					-- layer=2 filter=108 channel=82
					6, -5, 0, 3, 8, 8, -4, 7, 12,
					-- layer=2 filter=108 channel=83
					-14, -22, -28, -5, -16, 2, 44, 21, 10,
					-- layer=2 filter=108 channel=84
					-6, 8, -4, -3, 1, 11, -1, -9, -1,
					-- layer=2 filter=108 channel=85
					12, -3, -11, -8, 1, -4, -4, 0, 22,
					-- layer=2 filter=108 channel=86
					-8, 12, 8, 7, -4, 9, -3, -8, 7,
					-- layer=2 filter=108 channel=87
					44, -11, -19, 4, 43, 14, 22, 22, 13,
					-- layer=2 filter=108 channel=88
					-61, -34, -83, -56, -7, -34, -40, -8, 0,
					-- layer=2 filter=108 channel=89
					-5, -43, -32, -3, -31, -16, -17, -8, -6,
					-- layer=2 filter=108 channel=90
					-7, -3, -1, 9, -2, 1, 5, -1, 7,
					-- layer=2 filter=108 channel=91
					-2, -46, -43, -31, -56, -60, -25, -24, -16,
					-- layer=2 filter=108 channel=92
					-15, -28, -25, -6, -30, -38, -20, -26, -8,
					-- layer=2 filter=108 channel=93
					45, 15, -28, 42, 0, -15, 41, -16, -3,
					-- layer=2 filter=108 channel=94
					21, 35, 18, 34, 12, 39, 26, 1, 11,
					-- layer=2 filter=108 channel=95
					-5, 4, 2, 2, 6, -25, 0, -10, -6,
					-- layer=2 filter=108 channel=96
					12, 44, 33, -22, 37, -10, 22, 0, -42,
					-- layer=2 filter=108 channel=97
					-44, -57, -35, -49, -51, -32, 25, 38, -8,
					-- layer=2 filter=108 channel=98
					28, -34, -3, 3, -6, 32, -1, 29, 36,
					-- layer=2 filter=108 channel=99
					32, 22, 42, 10, 21, 42, 31, 14, 13,
					-- layer=2 filter=108 channel=100
					-60, -7, -67, -16, -31, 30, 50, 0, 25,
					-- layer=2 filter=108 channel=101
					-46, -45, 2, -33, -48, -20, -4, 14, 31,
					-- layer=2 filter=108 channel=102
					27, 9, -1, 23, 1, -4, 32, 18, -45,
					-- layer=2 filter=108 channel=103
					-28, 3, -28, -13, 0, 40, -18, 5, -38,
					-- layer=2 filter=108 channel=104
					23, 26, -29, 45, 28, 9, 34, 7, 22,
					-- layer=2 filter=108 channel=105
					-12, -77, -48, 17, -47, -3, -12, 30, -43,
					-- layer=2 filter=108 channel=106
					-34, -53, 37, -72, -80, -27, -11, -37, 12,
					-- layer=2 filter=108 channel=107
					1, -2, 9, -1, 0, -43, -13, -89, -9,
					-- layer=2 filter=108 channel=108
					-22, -12, 26, 26, -40, -5, -31, -25, -4,
					-- layer=2 filter=108 channel=109
					4, -7, -14, -9, -14, -2, 8, 14, 6,
					-- layer=2 filter=108 channel=110
					42, 2, 61, -31, -19, -36, -1, 5, 15,
					-- layer=2 filter=108 channel=111
					-1, 6, 5, 1, -4, 9, -10, -2, 5,
					-- layer=2 filter=108 channel=112
					-39, -51, 15, 3, -11, 16, -26, -53, -6,
					-- layer=2 filter=108 channel=113
					-67, -35, 7, -6, 7, -28, -5, 4, -3,
					-- layer=2 filter=108 channel=114
					18, 16, -2, 24, 11, 18, 0, -5, 20,
					-- layer=2 filter=108 channel=115
					-4, 0, 6, 7, -2, -1, 3, -1, -6,
					-- layer=2 filter=108 channel=116
					36, 25, 4, 6, 44, -5, 9, -12, -8,
					-- layer=2 filter=108 channel=117
					48, 0, -4, 34, -22, -6, 31, 22, 0,
					-- layer=2 filter=108 channel=118
					-1, -9, -43, -4, 37, 24, 38, 45, 15,
					-- layer=2 filter=108 channel=119
					24, -17, -65, 24, 26, -27, -1, -9, -9,
					-- layer=2 filter=108 channel=120
					-8, -7, 0, 4, -5, -9, -5, -2, 7,
					-- layer=2 filter=108 channel=121
					-8, 9, 1, 1, 5, 2, 3, 6, -4,
					-- layer=2 filter=108 channel=122
					-5, 12, 0, 3, 1, 9, 0, 6, 0,
					-- layer=2 filter=108 channel=123
					16, -13, 2, 19, 4, 32, 26, 35, 2,
					-- layer=2 filter=108 channel=124
					11, 9, -13, 23, 8, -6, 60, 16, -22,
					-- layer=2 filter=108 channel=125
					-6, -5, -6, 7, -7, 10, 0, -7, -2,
					-- layer=2 filter=108 channel=126
					0, 11, -16, -46, 3, -5, 18, -17, 4,
					-- layer=2 filter=108 channel=127
					2, -21, -80, -17, 18, 11, 8, -17, -10,
					-- layer=2 filter=109 channel=0
					11, 39, 27, -7, 7, -6, 2, -8, 5,
					-- layer=2 filter=109 channel=1
					-19, -28, -40, -23, -22, 12, -26, 13, 16,
					-- layer=2 filter=109 channel=2
					-3, -7, 5, -2, -7, -2, 9, 8, -4,
					-- layer=2 filter=109 channel=3
					11, 20, -1, -6, -15, -28, -8, -38, -66,
					-- layer=2 filter=109 channel=4
					24, 5, 1, 21, 10, -4, -8, -5, 16,
					-- layer=2 filter=109 channel=5
					-4, -10, 13, -1, 14, -11, -17, -7, 4,
					-- layer=2 filter=109 channel=6
					11, -39, -4, -11, -22, -53, -7, -21, -37,
					-- layer=2 filter=109 channel=7
					-17, 33, 18, 23, -19, -9, -49, 0, 25,
					-- layer=2 filter=109 channel=8
					0, 0, -9, 7, 5, 8, -9, -4, -10,
					-- layer=2 filter=109 channel=9
					-21, -15, -10, 8, 0, -22, 14, -31, 20,
					-- layer=2 filter=109 channel=10
					-17, 37, 28, 16, -14, 3, 31, -5, 14,
					-- layer=2 filter=109 channel=11
					-5, -8, -2, 14, 17, 10, 4, 13, -16,
					-- layer=2 filter=109 channel=12
					18, -19, -17, -19, -10, 6, 13, 9, 21,
					-- layer=2 filter=109 channel=13
					7, 3, -7, -1, 0, 2, -3, 4, 6,
					-- layer=2 filter=109 channel=14
					19, -21, 3, -1, 23, 25, 10, 8, -5,
					-- layer=2 filter=109 channel=15
					-46, -25, -52, 48, -7, -54, 26, -61, -20,
					-- layer=2 filter=109 channel=16
					-38, -21, -36, 15, 10, -35, -12, 26, -11,
					-- layer=2 filter=109 channel=17
					-11, -3, 10, 4, 0, 8, 5, 0, 3,
					-- layer=2 filter=109 channel=18
					31, 24, 4, 60, 43, 23, 26, -6, 19,
					-- layer=2 filter=109 channel=19
					-3, -57, -36, 12, -19, -16, -24, 27, 34,
					-- layer=2 filter=109 channel=20
					6, 2, -6, 8, 4, -1, 8, -5, -4,
					-- layer=2 filter=109 channel=21
					-1, 20, 8, -5, 7, 11, 2, 12, 3,
					-- layer=2 filter=109 channel=22
					3, 0, 1, 8, 9, 5, 7, -6, -2,
					-- layer=2 filter=109 channel=23
					0, 33, 5, 3, -7, -5, 1, 21, 5,
					-- layer=2 filter=109 channel=24
					3, 4, -41, 42, 13, 11, 19, -45, -13,
					-- layer=2 filter=109 channel=25
					21, -16, -13, 37, 10, -14, 0, -41, -41,
					-- layer=2 filter=109 channel=26
					5, -1, 6, 5, 0, -10, -6, -4, -12,
					-- layer=2 filter=109 channel=27
					16, -19, 1, -28, -14, -12, -4, 13, -2,
					-- layer=2 filter=109 channel=28
					-15, 7, 34, 12, -6, -16, 2, -18, -10,
					-- layer=2 filter=109 channel=29
					-3, -7, -9, 5, -7, 5, -3, 0, 8,
					-- layer=2 filter=109 channel=30
					3, 12, -26, 0, 14, 32, 39, -13, -29,
					-- layer=2 filter=109 channel=31
					6, 0, -15, -31, 33, -42, -2, 11, -44,
					-- layer=2 filter=109 channel=32
					-2, -4, 7, 12, 9, 7, -8, 8, 4,
					-- layer=2 filter=109 channel=33
					26, 17, -16, 9, 21, -16, -20, -49, -41,
					-- layer=2 filter=109 channel=34
					-71, 19, -30, -10, 28, -28, -21, 14, -4,
					-- layer=2 filter=109 channel=35
					8, 4, 43, 32, -27, 0, 11, -14, -24,
					-- layer=2 filter=109 channel=36
					11, 4, 6, 3, -10, 0, -13, 7, -10,
					-- layer=2 filter=109 channel=37
					-2, -20, -7, 4, 10, -12, -15, 17, 5,
					-- layer=2 filter=109 channel=38
					6, -8, -15, -1, 25, 1, 14, 9, 5,
					-- layer=2 filter=109 channel=39
					-4, 5, -10, 2, 0, -13, 8, -3, -31,
					-- layer=2 filter=109 channel=40
					-29, 4, -28, 29, -59, -14, 14, -19, -2,
					-- layer=2 filter=109 channel=41
					4, 7, -3, -8, -9, 7, 4, 2, -3,
					-- layer=2 filter=109 channel=42
					1, 0, -7, -6, -2, 0, -7, 2, -4,
					-- layer=2 filter=109 channel=43
					-6, 0, -22, 33, -30, -48, 13, -17, -6,
					-- layer=2 filter=109 channel=44
					-11, -6, 1, -6, 3, 0, -9, -8, -3,
					-- layer=2 filter=109 channel=45
					37, -9, -20, 14, 3, -27, 58, 7, 33,
					-- layer=2 filter=109 channel=46
					19, 20, -7, 20, 16, -2, 28, -35, -19,
					-- layer=2 filter=109 channel=47
					-8, 5, 6, 5, -3, -4, 20, -5, 13,
					-- layer=2 filter=109 channel=48
					-6, 3, -8, -4, 3, 8, -6, -1, 9,
					-- layer=2 filter=109 channel=49
					-1, -12, -55, 28, 43, 11, 0, -31, 4,
					-- layer=2 filter=109 channel=50
					5, -6, 3, -15, -2, 1, 3, 8, -6,
					-- layer=2 filter=109 channel=51
					2, 7, 11, 17, 10, 12, -10, 3, 2,
					-- layer=2 filter=109 channel=52
					-20, -22, -10, -30, -52, 4, 0, -2, 0,
					-- layer=2 filter=109 channel=53
					12, -38, -9, 26, 14, 4, -4, -17, -45,
					-- layer=2 filter=109 channel=54
					8, 6, 9, 19, -13, -42, -17, -35, -27,
					-- layer=2 filter=109 channel=55
					-5, 4, 1, 0, -3, -5, -5, 0, 11,
					-- layer=2 filter=109 channel=56
					-4, -20, 2, 40, 28, 3, 29, 21, 1,
					-- layer=2 filter=109 channel=57
					1, -6, -1, 0, -7, -3, -3, 6, 6,
					-- layer=2 filter=109 channel=58
					27, 2, 30, -30, -18, -3, 41, 32, 1,
					-- layer=2 filter=109 channel=59
					13, 5, -25, -26, 0, 2, 30, 51, 1,
					-- layer=2 filter=109 channel=60
					-4, -35, 2, -30, 0, 13, -10, 29, 41,
					-- layer=2 filter=109 channel=61
					-24, -1, 59, 12, -11, 40, 16, 17, -8,
					-- layer=2 filter=109 channel=62
					-4, -19, -60, 7, 0, -59, -2, -32, -20,
					-- layer=2 filter=109 channel=63
					-15, 12, 5, 2, 6, 10, -3, -6, 2,
					-- layer=2 filter=109 channel=64
					21, 10, -21, -3, 23, 20, -10, 4, 1,
					-- layer=2 filter=109 channel=65
					6, -35, 6, 2, -15, 25, 26, 18, 6,
					-- layer=2 filter=109 channel=66
					-16, 8, -3, -10, -10, 11, 42, 9, 33,
					-- layer=2 filter=109 channel=67
					1, -21, -21, 0, 11, 9, 23, -10, 17,
					-- layer=2 filter=109 channel=68
					5, 4, -2, -7, 0, -1, 3, -8, 3,
					-- layer=2 filter=109 channel=69
					23, 15, -20, -8, 33, 14, -26, 0, -2,
					-- layer=2 filter=109 channel=70
					-11, 18, 48, -3, -8, -13, -5, -8, -15,
					-- layer=2 filter=109 channel=71
					2, -22, -1, 18, 6, 9, 36, 18, -27,
					-- layer=2 filter=109 channel=72
					-12, -13, -13, 6, 6, 29, -50, 19, 21,
					-- layer=2 filter=109 channel=73
					-31, 18, -6, 21, -4, -52, -17, 23, -40,
					-- layer=2 filter=109 channel=74
					31, -3, 12, -11, -19, 23, 13, 0, -1,
					-- layer=2 filter=109 channel=75
					0, -2, 21, -46, -2, 9, 62, 48, -36,
					-- layer=2 filter=109 channel=76
					-31, -22, -22, -36, 13, 13, 12, 52, 58,
					-- layer=2 filter=109 channel=77
					-3, 8, -5, 4, -5, -1, -4, -8, -6,
					-- layer=2 filter=109 channel=78
					6, -13, -25, 14, -9, -25, -5, -12, -42,
					-- layer=2 filter=109 channel=79
					-7, 4, 8, -8, 0, -5, 0, -7, -1,
					-- layer=2 filter=109 channel=80
					-6, -4, 9, -11, 6, 11, 17, 5, -43,
					-- layer=2 filter=109 channel=81
					-7, 4, -8, -14, -8, -8, -4, -1, -14,
					-- layer=2 filter=109 channel=82
					0, 5, -9, 1, 6, -6, -1, -7, -11,
					-- layer=2 filter=109 channel=83
					15, -17, 22, -31, -22, 4, 7, 10, -15,
					-- layer=2 filter=109 channel=84
					-4, -2, -2, -1, 7, 8, 1, 10, 10,
					-- layer=2 filter=109 channel=85
					-15, 10, 0, -11, -8, 3, 11, -7, 16,
					-- layer=2 filter=109 channel=86
					-6, -7, 9, -15, 0, -3, 6, -9, 4,
					-- layer=2 filter=109 channel=87
					9, -18, -5, 24, 4, -1, 38, 18, -10,
					-- layer=2 filter=109 channel=88
					13, -12, -6, 2, -6, 15, 24, -9, -9,
					-- layer=2 filter=109 channel=89
					-42, -39, -45, -18, -22, 5, 23, 13, 15,
					-- layer=2 filter=109 channel=90
					-10, 0, -13, 7, -2, -7, 5, -7, -1,
					-- layer=2 filter=109 channel=91
					-8, -46, -55, -33, -50, -5, -2, 28, 1,
					-- layer=2 filter=109 channel=92
					-4, -27, -3, -15, 12, 24, -3, 0, 34,
					-- layer=2 filter=109 channel=93
					-42, -19, -43, -8, 5, -51, 25, -14, -18,
					-- layer=2 filter=109 channel=94
					-21, -30, -10, -10, -9, -15, -10, -18, -28,
					-- layer=2 filter=109 channel=95
					3, 7, 0, -4, 9, -4, 14, 17, 15,
					-- layer=2 filter=109 channel=96
					-9, -89, -30, -76, -42, -1, -81, 29, 2,
					-- layer=2 filter=109 channel=97
					24, -6, -23, 27, 41, 5, 38, -7, -13,
					-- layer=2 filter=109 channel=98
					-14, 14, 35, 2, -44, 0, 8, -3, 2,
					-- layer=2 filter=109 channel=99
					-41, -65, 11, -49, -20, 57, 2, 26, 36,
					-- layer=2 filter=109 channel=100
					1, -10, 0, -16, -34, -27, 12, 37, 29,
					-- layer=2 filter=109 channel=101
					15, 21, -12, 43, 8, 23, 51, 10, -16,
					-- layer=2 filter=109 channel=102
					48, -17, -48, -21, -21, -12, -40, 24, 21,
					-- layer=2 filter=109 channel=103
					-29, 14, -17, -32, -11, 6, -61, 2, 42,
					-- layer=2 filter=109 channel=104
					16, -67, -5, 38, -2, 0, -6, -25, -35,
					-- layer=2 filter=109 channel=105
					-23, -33, 18, 8, -19, -23, 21, 12, 92,
					-- layer=2 filter=109 channel=106
					13, -4, -8, 26, 28, 0, 36, 5, -19,
					-- layer=2 filter=109 channel=107
					16, -18, -8, 35, 33, 2, -23, -18, 38,
					-- layer=2 filter=109 channel=108
					-15, -25, -21, -28, -33, -15, 1, 5, -12,
					-- layer=2 filter=109 channel=109
					1, 0, -4, 5, 0, 8, -2, 4, -1,
					-- layer=2 filter=109 channel=110
					-26, -40, -15, -2, -41, 14, 0, 15, 13,
					-- layer=2 filter=109 channel=111
					10, 6, 0, 9, -9, 5, -4, 0, 3,
					-- layer=2 filter=109 channel=112
					-13, 20, 21, 5, 17, 22, -3, -35, -11,
					-- layer=2 filter=109 channel=113
					-22, 30, 18, -12, -17, 49, 18, 14, -33,
					-- layer=2 filter=109 channel=114
					5, -7, -11, -15, 1, -3, -10, 1, 1,
					-- layer=2 filter=109 channel=115
					-5, 2, -3, -10, 4, -3, -4, 5, 0,
					-- layer=2 filter=109 channel=116
					-19, -14, 19, -18, -15, 0, -28, 15, -27,
					-- layer=2 filter=109 channel=117
					-53, -3, 2, 2, -41, -24, -38, 39, 29,
					-- layer=2 filter=109 channel=118
					14, 13, -1, 29, -19, -25, -18, -20, -24,
					-- layer=2 filter=109 channel=119
					-3, 8, -6, 32, 60, -25, 1, -4, -1,
					-- layer=2 filter=109 channel=120
					-1, -9, 6, 3, 10, 1, 0, 5, -4,
					-- layer=2 filter=109 channel=121
					-6, 6, 0, -1, -10, -7, -6, 10, 5,
					-- layer=2 filter=109 channel=122
					2, 1, -7, -4, -7, -7, 7, 3, 7,
					-- layer=2 filter=109 channel=123
					1, -18, -12, 9, -36, -19, -33, 1, 34,
					-- layer=2 filter=109 channel=124
					-22, 4, -29, 28, 40, -49, 21, -33, 33,
					-- layer=2 filter=109 channel=125
					11, 7, 7, 6, 9, -7, 5, 9, 8,
					-- layer=2 filter=109 channel=126
					16, 18, -27, 36, -51, 14, 16, -15, 14,
					-- layer=2 filter=109 channel=127
					13, -2, 15, -10, 19, 0, -5, -1, 3,
					-- layer=2 filter=110 channel=0
					-25, -11, -24, -18, -14, -24, 32, -3, 16,
					-- layer=2 filter=110 channel=1
					-12, 10, 31, 21, -22, 6, 32, 23, 18,
					-- layer=2 filter=110 channel=2
					-11, 4, -7, 5, 2, 1, 7, 2, -7,
					-- layer=2 filter=110 channel=3
					-14, -45, 7, -13, 14, -8, 13, 48, 57,
					-- layer=2 filter=110 channel=4
					17, -6, -23, 22, 11, -12, -9, 10, -7,
					-- layer=2 filter=110 channel=5
					-31, -51, -58, -42, -65, -61, -18, -3, -33,
					-- layer=2 filter=110 channel=6
					-45, -24, 10, 3, -45, 8, 9, -4, -25,
					-- layer=2 filter=110 channel=7
					12, 13, -17, -14, 16, -48, 6, 12, -3,
					-- layer=2 filter=110 channel=8
					-3, -2, 10, -1, 0, 2, 9, -8, -6,
					-- layer=2 filter=110 channel=9
					-30, -7, -18, -17, -10, -6, -23, -21, 12,
					-- layer=2 filter=110 channel=10
					4, -16, -16, -6, 23, -1, 33, 35, 17,
					-- layer=2 filter=110 channel=11
					-50, -47, -46, -59, -53, -52, 8, -1, 2,
					-- layer=2 filter=110 channel=12
					-3, -16, 16, 14, -31, -9, 9, 21, -21,
					-- layer=2 filter=110 channel=13
					4, 2, 1, 1, 8, -3, 7, -9, 8,
					-- layer=2 filter=110 channel=14
					-1, -7, 20, 0, -18, 3, 26, 30, 0,
					-- layer=2 filter=110 channel=15
					-19, -52, -38, 9, 33, 4, 48, 38, 56,
					-- layer=2 filter=110 channel=16
					2, -5, -15, -4, 5, 28, -62, -8, 0,
					-- layer=2 filter=110 channel=17
					-7, -6, -5, 0, -6, 8, -8, -8, 8,
					-- layer=2 filter=110 channel=18
					-2, -36, -21, 4, -16, -4, 21, 24, 10,
					-- layer=2 filter=110 channel=19
					-35, -43, -22, 19, -44, -12, 44, 21, -15,
					-- layer=2 filter=110 channel=20
					-4, -1, -6, 6, -5, 9, -9, -8, 2,
					-- layer=2 filter=110 channel=21
					-2, 6, -2, 24, 9, -5, 6, -4, 8,
					-- layer=2 filter=110 channel=22
					-10, 9, 8, 0, 10, -4, 0, -11, 0,
					-- layer=2 filter=110 channel=23
					-5, -4, 16, -8, 30, 31, -38, -9, 14,
					-- layer=2 filter=110 channel=24
					-26, 9, -27, -6, 8, -8, 46, 38, 27,
					-- layer=2 filter=110 channel=25
					6, 17, 7, -18, -17, 0, 39, 30, 5,
					-- layer=2 filter=110 channel=26
					7, 0, -5, -10, -3, 4, -3, -6, -3,
					-- layer=2 filter=110 channel=27
					18, -7, -10, 33, -29, -29, -2, -20, -9,
					-- layer=2 filter=110 channel=28
					27, 12, 17, -8, -20, 51, -10, 0, 19,
					-- layer=2 filter=110 channel=29
					9, -6, -7, 2, -7, 11, -7, -1, -4,
					-- layer=2 filter=110 channel=30
					2, -10, -23, 6, 9, -17, 0, 4, -11,
					-- layer=2 filter=110 channel=31
					-14, -27, 0, -60, -9, 40, 24, 12, 16,
					-- layer=2 filter=110 channel=32
					9, -3, -1, -4, 8, 6, 2, -8, 5,
					-- layer=2 filter=110 channel=33
					-40, -14, -16, 4, 46, -35, -2, -1, 0,
					-- layer=2 filter=110 channel=34
					31, -73, -44, 19, -4, 6, -24, 0, 29,
					-- layer=2 filter=110 channel=35
					12, 12, 24, 2, 24, 50, -19, -23, -10,
					-- layer=2 filter=110 channel=36
					-4, -11, 8, 4, 11, -2, -3, -6, 6,
					-- layer=2 filter=110 channel=37
					-41, -60, -60, -23, -59, -50, 12, 5, 0,
					-- layer=2 filter=110 channel=38
					20, 5, -34, 76, 5, -12, -10, -10, -23,
					-- layer=2 filter=110 channel=39
					-15, 9, 11, -17, 21, 16, -6, 5, 4,
					-- layer=2 filter=110 channel=40
					-65, -19, -16, 0, 23, 30, 11, 35, 40,
					-- layer=2 filter=110 channel=41
					0, -4, -5, -5, 3, 3, 3, -3, 4,
					-- layer=2 filter=110 channel=42
					5, 37, 30, -5, 40, 35, -32, 14, 30,
					-- layer=2 filter=110 channel=43
					-33, -12, -45, -17, -6, -10, -24, 42, 21,
					-- layer=2 filter=110 channel=44
					0, -5, 6, -9, -3, -8, -7, 4, -5,
					-- layer=2 filter=110 channel=45
					3, -5, -42, 31, -10, 24, -21, 28, 24,
					-- layer=2 filter=110 channel=46
					4, -37, -33, 6, 2, -10, 17, -1, 26,
					-- layer=2 filter=110 channel=47
					11, 3, -9, -5, 0, 10, -14, 10, 32,
					-- layer=2 filter=110 channel=48
					9, 1, -4, 7, -10, 7, 0, 14, 7,
					-- layer=2 filter=110 channel=49
					-28, -27, 14, 2, 23, 58, 30, 43, 44,
					-- layer=2 filter=110 channel=50
					14, -1, 7, 25, 20, 28, 7, 20, 22,
					-- layer=2 filter=110 channel=51
					-42, -26, -30, -41, -48, -51, 19, -13, -5,
					-- layer=2 filter=110 channel=52
					-73, -73, -13, -21, -34, -7, 47, -15, 13,
					-- layer=2 filter=110 channel=53
					47, 7, 7, 4, -16, -17, 59, 11, -2,
					-- layer=2 filter=110 channel=54
					-10, -13, 16, -9, -16, -10, 3, 14, -5,
					-- layer=2 filter=110 channel=55
					-1, -2, 0, -5, 0, 9, -1, 5, 9,
					-- layer=2 filter=110 channel=56
					-34, -5, -50, -31, -49, -62, 1, 0, -3,
					-- layer=2 filter=110 channel=57
					3, -15, 0, 9, -6, 0, 14, 0, 0,
					-- layer=2 filter=110 channel=58
					-6, -23, 24, 0, -23, -13, -6, 8, -19,
					-- layer=2 filter=110 channel=59
					26, 8, -38, 60, -9, -56, 33, 15, -26,
					-- layer=2 filter=110 channel=60
					41, 28, -22, 41, -54, -65, 26, -22, -46,
					-- layer=2 filter=110 channel=61
					-25, -16, -17, -7, -2, -60, 45, 0, -70,
					-- layer=2 filter=110 channel=62
					-23, -49, 12, 33, -17, 11, 42, -14, 26,
					-- layer=2 filter=110 channel=63
					-13, 16, -14, -10, 17, 4, -4, -3, 8,
					-- layer=2 filter=110 channel=64
					6, 19, 11, 2, 33, 16, -17, 8, 40,
					-- layer=2 filter=110 channel=65
					-14, 3, -49, -27, -49, -14, 10, -67, -30,
					-- layer=2 filter=110 channel=66
					-27, -41, 14, 10, -16, 27, -21, 16, 3,
					-- layer=2 filter=110 channel=67
					-14, -22, -28, -39, -11, -21, -19, 16, 21,
					-- layer=2 filter=110 channel=68
					-5, 6, 4, 6, -5, 6, 9, 4, -2,
					-- layer=2 filter=110 channel=69
					-9, 14, 12, -1, 19, 16, -21, 1, 24,
					-- layer=2 filter=110 channel=70
					-14, -21, -24, -11, 8, 38, -19, -5, 0,
					-- layer=2 filter=110 channel=71
					15, -3, -33, 9, -14, -33, -12, 28, 5,
					-- layer=2 filter=110 channel=72
					-1, 11, 1, 2, 0, -26, 0, -17, 5,
					-- layer=2 filter=110 channel=73
					19, -20, 6, -4, 7, -1, -6, 36, -25,
					-- layer=2 filter=110 channel=74
					6, 28, 1, 9, 6, -7, -12, 16, 20,
					-- layer=2 filter=110 channel=75
					-52, -54, -41, -78, -88, 16, 17, 41, 4,
					-- layer=2 filter=110 channel=76
					-30, -111, 14, -19, -51, -3, 3, 27, 10,
					-- layer=2 filter=110 channel=77
					7, 11, 9, -2, -5, 2, -6, 3, 0,
					-- layer=2 filter=110 channel=78
					-75, -68, -25, -50, -48, -29, 22, 14, 9,
					-- layer=2 filter=110 channel=79
					-9, -10, 9, -1, 2, -4, -4, 4, 2,
					-- layer=2 filter=110 channel=80
					-19, -7, 5, 5, 31, 35, -12, 5, 16,
					-- layer=2 filter=110 channel=81
					4, -8, 0, 1, -18, 2, -7, -5, -2,
					-- layer=2 filter=110 channel=82
					-11, 4, 8, 10, -9, -8, 10, -8, -6,
					-- layer=2 filter=110 channel=83
					-8, -18, -22, 0, 11, 20, -42, -18, -26,
					-- layer=2 filter=110 channel=84
					9, 9, 2, 0, -7, -8, 4, -6, 9,
					-- layer=2 filter=110 channel=85
					0, -8, 7, 1, 5, -2, 1, -17, 2,
					-- layer=2 filter=110 channel=86
					13, 5, 6, 0, 9, -6, 4, -5, -2,
					-- layer=2 filter=110 channel=87
					-31, -17, 18, 5, 22, 9, 14, 0, 68,
					-- layer=2 filter=110 channel=88
					14, 12, 13, 18, 9, -6, -21, 2, 3,
					-- layer=2 filter=110 channel=89
					8, 6, 19, 2, -2, 1, 33, 4, 12,
					-- layer=2 filter=110 channel=90
					0, 4, 4, 0, 8, 11, -5, -5, 5,
					-- layer=2 filter=110 channel=91
					5, 0, -3, 9, -18, 0, 31, 28, 20,
					-- layer=2 filter=110 channel=92
					-9, 16, 27, 42, -2, 17, 14, 12, 16,
					-- layer=2 filter=110 channel=93
					-17, -37, -29, -28, -24, -25, 15, 14, 33,
					-- layer=2 filter=110 channel=94
					-52, -36, 4, 21, -27, -28, 60, -1, -13,
					-- layer=2 filter=110 channel=95
					-8, 7, 6, -5, 7, 8, 0, -13, 2,
					-- layer=2 filter=110 channel=96
					18, -33, -22, -13, -38, -30, 41, -28, 21,
					-- layer=2 filter=110 channel=97
					-34, -9, -7, -64, 1, 7, -25, 31, 41,
					-- layer=2 filter=110 channel=98
					5, -5, 0, -22, -36, 41, 10, -11, 35,
					-- layer=2 filter=110 channel=99
					-28, -67, -38, -18, -46, 0, 40, -38, 13,
					-- layer=2 filter=110 channel=100
					9, -4, -5, 28, 4, -2, -39, 8, 0,
					-- layer=2 filter=110 channel=101
					7, -13, -4, -58, -29, -46, 3, -10, -1,
					-- layer=2 filter=110 channel=102
					19, -19, -38, -22, -36, -19, 6, -6, 44,
					-- layer=2 filter=110 channel=103
					13, 6, 37, -40, 23, -6, -3, 13, -41,
					-- layer=2 filter=110 channel=104
					-26, -9, 11, 23, -9, 8, 20, 22, 27,
					-- layer=2 filter=110 channel=105
					35, -6, -17, -45, -38, -4, -17, -2, 0,
					-- layer=2 filter=110 channel=106
					10, 2, -19, 14, -43, -16, 51, 28, 0,
					-- layer=2 filter=110 channel=107
					7, -5, -5, -18, 39, 2, -5, -45, -20,
					-- layer=2 filter=110 channel=108
					39, 11, -26, 10, -29, -30, 38, 14, -13,
					-- layer=2 filter=110 channel=109
					8, 10, 10, 16, -6, -22, 5, 16, -14,
					-- layer=2 filter=110 channel=110
					0, 15, 10, -14, -7, 27, -19, -12, 5,
					-- layer=2 filter=110 channel=111
					7, 1, -4, -6, 5, 5, 4, -3, 5,
					-- layer=2 filter=110 channel=112
					-9, -14, -7, -44, -39, -73, 39, -12, -13,
					-- layer=2 filter=110 channel=113
					-11, -7, -8, 5, 34, 15, -13, -36, -10,
					-- layer=2 filter=110 channel=114
					8, -1, 0, 9, 18, 10, 3, -11, -12,
					-- layer=2 filter=110 channel=115
					1, -5, 6, -5, 9, -8, 5, 2, -5,
					-- layer=2 filter=110 channel=116
					-38, -31, 24, -13, -10, 9, 10, 4, 63,
					-- layer=2 filter=110 channel=117
					-91, -43, -7, -10, -10, -35, 17, 19, -21,
					-- layer=2 filter=110 channel=118
					-41, -59, -32, -23, 10, 45, 10, 32, 33,
					-- layer=2 filter=110 channel=119
					24, -12, -11, 18, 16, -2, -25, 4, 8,
					-- layer=2 filter=110 channel=120
					0, 0, 9, 0, -10, 3, 6, -1, 4,
					-- layer=2 filter=110 channel=121
					-2, 1, 0, -7, -8, 12, 6, 6, -2,
					-- layer=2 filter=110 channel=122
					-5, 0, -11, 0, 0, 4, 7, -10, 6,
					-- layer=2 filter=110 channel=123
					-24, 5, 0, -35, -8, -30, 15, -5, 13,
					-- layer=2 filter=110 channel=124
					-64, -29, 23, 12, 33, 14, 33, 42, 33,
					-- layer=2 filter=110 channel=125
					1, 10, -3, -2, 6, -4, 8, 7, 1,
					-- layer=2 filter=110 channel=126
					53, 46, -19, 23, 10, -24, 33, -2, 24,
					-- layer=2 filter=110 channel=127
					10, 34, 18, 8, 8, 20, -14, -27, 1,
					-- layer=2 filter=111 channel=0
					-8, -10, 10, -6, -9, 11, 23, 1, 7,
					-- layer=2 filter=111 channel=1
					-5, -28, 23, 21, 0, -36, -38, -34, -11,
					-- layer=2 filter=111 channel=2
					10, 1, 6, -3, -1, 5, -6, -7, -5,
					-- layer=2 filter=111 channel=3
					-7, -28, -38, -16, -23, 13, 43, 53, 26,
					-- layer=2 filter=111 channel=4
					-12, -24, -27, -16, -57, -18, -5, 0, 13,
					-- layer=2 filter=111 channel=5
					-10, -26, -6, -13, -11, 14, 1, -9, 4,
					-- layer=2 filter=111 channel=6
					15, 13, -8, 12, 35, 33, -13, -35, -11,
					-- layer=2 filter=111 channel=7
					-7, 12, -9, 52, -6, -21, 49, 0, 11,
					-- layer=2 filter=111 channel=8
					5, 1, -5, -9, 14, -9, 3, -8, -2,
					-- layer=2 filter=111 channel=9
					8, -9, -24, -27, -16, -6, 12, 12, 6,
					-- layer=2 filter=111 channel=10
					0, 21, 9, -14, -2, -13, 18, 21, 21,
					-- layer=2 filter=111 channel=11
					2, -6, -5, 17, 13, -2, 9, -4, -1,
					-- layer=2 filter=111 channel=12
					-25, -6, 7, -4, -43, -38, 6, -36, -20,
					-- layer=2 filter=111 channel=13
					-3, 4, -10, -9, -7, 4, 0, 2, 0,
					-- layer=2 filter=111 channel=14
					24, 0, 11, 52, -4, -15, -2, -38, -39,
					-- layer=2 filter=111 channel=15
					21, 18, 35, -2, -9, 33, -19, -24, 2,
					-- layer=2 filter=111 channel=16
					-52, -31, 26, -45, -27, 9, 13, 38, 29,
					-- layer=2 filter=111 channel=17
					-11, 4, -2, -6, -5, -2, 0, -7, -5,
					-- layer=2 filter=111 channel=18
					40, 16, 12, 4, 39, 8, 15, -11, 5,
					-- layer=2 filter=111 channel=19
					9, 0, 18, -28, -26, -6, -43, 9, -17,
					-- layer=2 filter=111 channel=20
					-7, 3, -5, 4, -3, -7, -8, 1, -4,
					-- layer=2 filter=111 channel=21
					9, 17, 10, 3, 18, 2, -1, 4, -2,
					-- layer=2 filter=111 channel=22
					5, 4, -5, -4, 7, 0, -8, -6, -3,
					-- layer=2 filter=111 channel=23
					-27, -43, -18, 11, -21, 27, 2, 12, 18,
					-- layer=2 filter=111 channel=24
					9, -7, -13, -8, -45, -9, 14, 0, -16,
					-- layer=2 filter=111 channel=25
					-32, -27, -9, -26, -32, -41, -3, -31, -38,
					-- layer=2 filter=111 channel=26
					3, 9, -5, 0, -7, 6, -6, 1, 9,
					-- layer=2 filter=111 channel=27
					2, -9, -14, 12, -27, -6, 45, 30, 37,
					-- layer=2 filter=111 channel=28
					4, 13, 40, 19, 13, 4, 43, 4, -9,
					-- layer=2 filter=111 channel=29
					-10, -8, -9, 1, -5, -3, 10, -5, -9,
					-- layer=2 filter=111 channel=30
					-3, 4, -7, -36, -10, -4, -29, -25, 0,
					-- layer=2 filter=111 channel=31
					8, 0, -51, 10, -10, 25, -19, 45, -16,
					-- layer=2 filter=111 channel=32
					0, 2, 0, -3, -9, -10, -3, -5, 1,
					-- layer=2 filter=111 channel=33
					0, 17, 19, 25, -19, 8, 40, 4, 25,
					-- layer=2 filter=111 channel=34
					12, 20, -10, -26, 34, 6, -31, 1, -2,
					-- layer=2 filter=111 channel=35
					26, 6, -16, -11, 3, -13, 41, -1, -8,
					-- layer=2 filter=111 channel=36
					-14, 1, 0, -3, 1, 1, 14, 1, 6,
					-- layer=2 filter=111 channel=37
					17, -9, 3, 11, -10, -1, 2, -8, -10,
					-- layer=2 filter=111 channel=38
					9, -2, -10, 9, -4, 8, 9, 11, 2,
					-- layer=2 filter=111 channel=39
					-11, -12, -5, 25, -17, 27, 18, 14, 15,
					-- layer=2 filter=111 channel=40
					10, -20, -12, -3, 31, 35, -37, -19, 34,
					-- layer=2 filter=111 channel=41
					8, -5, 0, 0, 0, 4, 5, -10, -3,
					-- layer=2 filter=111 channel=42
					-7, 0, 26, 16, 7, 51, 11, 11, -18,
					-- layer=2 filter=111 channel=43
					7, -2, -15, -22, -8, 0, 4, 6, 21,
					-- layer=2 filter=111 channel=44
					2, 8, 7, -5, -4, 0, 5, 10, 7,
					-- layer=2 filter=111 channel=45
					-64, -39, -29, -39, -79, -35, 24, 19, 6,
					-- layer=2 filter=111 channel=46
					-13, 35, -26, -58, 0, -9, -22, 26, 1,
					-- layer=2 filter=111 channel=47
					-14, -24, 13, 10, -28, -16, 10, -29, -18,
					-- layer=2 filter=111 channel=48
					2, 9, -10, 3, 7, 2, -3, -9, -7,
					-- layer=2 filter=111 channel=49
					9, 35, 32, -6, 22, 0, -44, -38, -24,
					-- layer=2 filter=111 channel=50
					11, 8, -8, -1, -7, -24, 0, -6, -22,
					-- layer=2 filter=111 channel=51
					-7, -11, -5, 16, -4, 4, 0, 10, -7,
					-- layer=2 filter=111 channel=52
					0, 0, -6, -5, -9, 11, 13, 3, 8,
					-- layer=2 filter=111 channel=53
					17, 27, 43, -29, 32, 23, -11, 21, -41,
					-- layer=2 filter=111 channel=54
					9, -6, 24, 14, 5, 0, 24, -21, -6,
					-- layer=2 filter=111 channel=55
					0, -11, 11, 6, -4, -3, 5, 5, -4,
					-- layer=2 filter=111 channel=56
					-7, -18, -3, 11, 6, 0, 0, -5, -3,
					-- layer=2 filter=111 channel=57
					-8, 4, -4, -5, -12, -3, 3, -1, -3,
					-- layer=2 filter=111 channel=58
					4, -9, -5, 11, -50, -22, 14, -15, 3,
					-- layer=2 filter=111 channel=59
					-16, -1, -7, 7, -7, 10, -6, -10, -2,
					-- layer=2 filter=111 channel=60
					6, 9, 25, 16, 42, 20, -13, -37, -26,
					-- layer=2 filter=111 channel=61
					13, 18, 40, 33, 61, 23, 15, -17, 11,
					-- layer=2 filter=111 channel=62
					-6, -11, -16, -28, 13, 22, -66, -40, -2,
					-- layer=2 filter=111 channel=63
					-30, -11, 6, -6, -38, 1, 15, -17, 10,
					-- layer=2 filter=111 channel=64
					9, -11, -6, 23, 15, 22, 0, 18, 20,
					-- layer=2 filter=111 channel=65
					23, 36, 22, 27, 57, 22, -22, 2, 17,
					-- layer=2 filter=111 channel=66
					-22, 17, -8, 18, -14, -30, 3, -15, 0,
					-- layer=2 filter=111 channel=67
					-10, 24, -18, -24, -14, 10, -44, 21, 15,
					-- layer=2 filter=111 channel=68
					-2, 9, 7, 7, -4, -6, 1, -11, 0,
					-- layer=2 filter=111 channel=69
					-4, -13, 23, 17, -4, 23, -9, 0, 20,
					-- layer=2 filter=111 channel=70
					15, 4, 17, 15, 15, -24, 21, -22, -16,
					-- layer=2 filter=111 channel=71
					-7, -15, 0, 15, 15, 49, 35, 16, 29,
					-- layer=2 filter=111 channel=72
					-5, 23, 23, 35, 33, -4, 50, 6, -26,
					-- layer=2 filter=111 channel=73
					-24, 45, -13, -36, 18, 10, 15, -19, -12,
					-- layer=2 filter=111 channel=74
					-7, 38, -2, -19, -21, -19, -13, 37, 10,
					-- layer=2 filter=111 channel=75
					-17, 25, 14, 1, -3, -25, -11, -61, -65,
					-- layer=2 filter=111 channel=76
					-24, -47, -3, -42, 57, -34, 11, 0, 27,
					-- layer=2 filter=111 channel=77
					-4, 7, 4, 2, -2, 1, -1, -5, -4,
					-- layer=2 filter=111 channel=78
					14, -26, -13, -2, -12, -10, -21, -23, -13,
					-- layer=2 filter=111 channel=79
					9, 4, -4, 0, 1, -1, -1, 0, 1,
					-- layer=2 filter=111 channel=80
					7, 19, -4, -1, -12, 39, -16, 18, 46,
					-- layer=2 filter=111 channel=81
					-15, -7, -2, 6, -10, -3, 4, 0, 10,
					-- layer=2 filter=111 channel=82
					-7, -3, 7, -1, 8, 8, 7, 10, 5,
					-- layer=2 filter=111 channel=83
					-12, -42, -12, -31, -54, -23, -21, -27, 7,
					-- layer=2 filter=111 channel=84
					3, -6, 11, -7, 9, 9, -2, 2, -1,
					-- layer=2 filter=111 channel=85
					6, -5, -2, -6, -9, 7, -9, -4, -22,
					-- layer=2 filter=111 channel=86
					4, 7, 18, -8, 10, 8, -1, -6, -17,
					-- layer=2 filter=111 channel=87
					13, 7, -22, 0, 26, 33, 8, 16, 11,
					-- layer=2 filter=111 channel=88
					19, 14, -9, -8, -21, 13, -11, -4, 11,
					-- layer=2 filter=111 channel=89
					-38, -25, 14, 16, -7, -16, -31, -52, -37,
					-- layer=2 filter=111 channel=90
					3, -7, -6, 5, -3, -5, 9, -9, 10,
					-- layer=2 filter=111 channel=91
					-23, 19, 5, 9, -29, -4, 18, -43, -65,
					-- layer=2 filter=111 channel=92
					-20, -13, 11, 3, -9, -39, -28, -48, -57,
					-- layer=2 filter=111 channel=93
					26, 31, -56, 27, -13, -12, 6, -22, 39,
					-- layer=2 filter=111 channel=94
					-3, 4, 28, 0, 41, 16, -4, 0, 11,
					-- layer=2 filter=111 channel=95
					2, -8, -5, -4, -3, -1, -5, -9, -13,
					-- layer=2 filter=111 channel=96
					-35, -9, -24, -7, 17, 10, 3, -2, -14,
					-- layer=2 filter=111 channel=97
					11, -14, 13, 13, 0, 2, 12, 28, 2,
					-- layer=2 filter=111 channel=98
					8, -21, 14, 18, 16, -4, 17, -13, -7,
					-- layer=2 filter=111 channel=99
					33, -2, 1, 1, 40, 46, 35, 9, 18,
					-- layer=2 filter=111 channel=100
					-28, -40, -14, -25, -5, 5, 8, -12, 35,
					-- layer=2 filter=111 channel=101
					-13, 12, 10, 0, 7, 6, 21, -12, 11,
					-- layer=2 filter=111 channel=102
					11, 15, 2, 14, 52, 20, 10, -21, -1,
					-- layer=2 filter=111 channel=103
					-11, 18, -40, 10, 13, -11, -60, -19, -11,
					-- layer=2 filter=111 channel=104
					-13, 17, 38, 30, 33, 10, -6, 16, -27,
					-- layer=2 filter=111 channel=105
					-26, -24, 29, 4, -22, -15, -22, 1, 57,
					-- layer=2 filter=111 channel=106
					7, 34, -16, 30, -49, -37, 20, 0, -28,
					-- layer=2 filter=111 channel=107
					-36, 27, -3, -6, 17, 15, -14, -60, -40,
					-- layer=2 filter=111 channel=108
					26, -8, 1, 27, 9, 18, -6, -26, -6,
					-- layer=2 filter=111 channel=109
					-20, -17, -11, -9, -6, -12, -7, 6, 1,
					-- layer=2 filter=111 channel=110
					8, -22, 6, 26, 26, 15, 29, 8, 25,
					-- layer=2 filter=111 channel=111
					-7, 7, -5, 8, -5, 5, 3, -5, -1,
					-- layer=2 filter=111 channel=112
					8, 10, 8, 5, 7, 14, -31, -25, -3,
					-- layer=2 filter=111 channel=113
					-18, 12, 19, -22, -2, -20, 2, -27, 5,
					-- layer=2 filter=111 channel=114
					3, 0, -2, 0, -2, 0, 10, 6, 0,
					-- layer=2 filter=111 channel=115
					3, 8, 5, -3, -7, -2, 2, -10, 1,
					-- layer=2 filter=111 channel=116
					18, 20, 0, -22, 12, 22, -23, -16, 12,
					-- layer=2 filter=111 channel=117
					-8, 34, 14, 30, 14, -27, 20, -40, -49,
					-- layer=2 filter=111 channel=118
					11, -5, -8, -28, -28, 18, -13, 22, 11,
					-- layer=2 filter=111 channel=119
					8, 10, -23, -5, -4, 25, -9, -17, 36,
					-- layer=2 filter=111 channel=120
					5, 8, 6, 7, 4, -3, 2, 2, -10,
					-- layer=2 filter=111 channel=121
					4, 0, 3, 0, -9, 1, 3, -3, -10,
					-- layer=2 filter=111 channel=122
					-6, 0, 0, -12, 0, -10, 4, 18, -2,
					-- layer=2 filter=111 channel=123
					21, -3, 17, 53, 28, 1, 1, -14, 6,
					-- layer=2 filter=111 channel=124
					-34, -17, 8, 8, 30, 22, -28, -24, 6,
					-- layer=2 filter=111 channel=125
					-5, 3, 0, 7, -1, 13, -3, -10, 0,
					-- layer=2 filter=111 channel=126
					17, -54, -49, 20, -3, -5, 70, -38, -39,
					-- layer=2 filter=111 channel=127
					-22, -32, -11, -12, 4, 3, 2, -12, 3,
					-- layer=2 filter=112 channel=0
					-8, 7, 11, -17, 5, -18, -10, 20, -5,
					-- layer=2 filter=112 channel=1
					36, 35, 11, 11, -30, 16, 4, -23, -24,
					-- layer=2 filter=112 channel=2
					-12, -6, 10, -8, 0, 2, -3, 1, 0,
					-- layer=2 filter=112 channel=3
					18, 15, 11, 34, 15, -9, -50, -23, -33,
					-- layer=2 filter=112 channel=4
					-6, -25, -22, 3, -36, -1, -48, -74, -34,
					-- layer=2 filter=112 channel=5
					-12, -26, -9, 2, -14, 14, 8, 24, -22,
					-- layer=2 filter=112 channel=6
					-43, -24, -77, -25, -44, -12, 37, -35, 7,
					-- layer=2 filter=112 channel=7
					-20, -47, -41, -22, 7, -72, -4, -52, -9,
					-- layer=2 filter=112 channel=8
					-11, -6, 8, 0, 5, 1, -4, 5, 2,
					-- layer=2 filter=112 channel=9
					-17, 1, 10, -12, 5, 32, -32, 13, 45,
					-- layer=2 filter=112 channel=10
					4, 3, 6, -17, 3, 0, -45, -1, -21,
					-- layer=2 filter=112 channel=11
					-4, -19, -6, -5, 6, 7, 27, -4, -4,
					-- layer=2 filter=112 channel=12
					26, 12, -2, -13, -30, -31, -20, -24, -2,
					-- layer=2 filter=112 channel=13
					8, -8, 0, -7, 5, -1, -4, 2, -3,
					-- layer=2 filter=112 channel=14
					5, 42, 14, -11, -10, 11, 24, -1, 7,
					-- layer=2 filter=112 channel=15
					40, 34, 25, 60, 21, 28, 56, 46, -29,
					-- layer=2 filter=112 channel=16
					-37, -42, -23, 5, 10, 9, -17, -23, 8,
					-- layer=2 filter=112 channel=17
					-3, 5, 9, 3, -7, -7, -5, 4, 1,
					-- layer=2 filter=112 channel=18
					27, 31, 12, -19, 17, 15, 43, 0, 0,
					-- layer=2 filter=112 channel=19
					0, 5, -9, 29, 0, 21, 32, 23, -3,
					-- layer=2 filter=112 channel=20
					6, 7, 7, -9, 4, 7, -3, -6, -12,
					-- layer=2 filter=112 channel=21
					9, -2, 2, -13, -10, 5, -13, -1, -8,
					-- layer=2 filter=112 channel=22
					-3, -3, -6, 6, -3, -1, 4, -6, 1,
					-- layer=2 filter=112 channel=23
					40, -14, -2, 18, -34, 0, -11, -32, 23,
					-- layer=2 filter=112 channel=24
					12, 5, 1, 18, 19, 17, 1, -14, -5,
					-- layer=2 filter=112 channel=25
					-15, 8, -24, 37, 21, -4, 36, -5, -22,
					-- layer=2 filter=112 channel=26
					-7, 5, 9, 4, -1, -3, -5, -10, 0,
					-- layer=2 filter=112 channel=27
					-17, -6, 5, 0, 9, 0, 1, 17, -8,
					-- layer=2 filter=112 channel=28
					-56, -69, 4, 11, -28, -85, 1, -12, -18,
					-- layer=2 filter=112 channel=29
					-8, -5, -1, -5, 9, 3, 10, -4, 5,
					-- layer=2 filter=112 channel=30
					6, 9, 13, 31, -5, -5, 13, 23, 0,
					-- layer=2 filter=112 channel=31
					46, 11, -79, 9, 17, -32, 12, 31, -19,
					-- layer=2 filter=112 channel=32
					4, 7, -6, 0, -1, -2, 6, 6, 3,
					-- layer=2 filter=112 channel=33
					-4, 15, 15, 28, 2, -66, -8, -32, -72,
					-- layer=2 filter=112 channel=34
					31, -52, 17, 31, -34, -51, -3, 23, -15,
					-- layer=2 filter=112 channel=35
					-40, -74, -11, -14, -34, -83, -15, 3, -31,
					-- layer=2 filter=112 channel=36
					7, 6, 5, -4, 12, -5, -7, 7, 7,
					-- layer=2 filter=112 channel=37
					-7, 0, 0, -2, 1, 7, 34, 14, -20,
					-- layer=2 filter=112 channel=38
					-16, 12, -11, 0, -3, 3, 24, 22, -34,
					-- layer=2 filter=112 channel=39
					29, 20, 6, 22, 23, 19, -30, -9, 10,
					-- layer=2 filter=112 channel=40
					3, 7, 10, 31, -7, -84, 4, 39, -15,
					-- layer=2 filter=112 channel=41
					-1, -5, -9, -4, -9, -11, 9, -2, 6,
					-- layer=2 filter=112 channel=42
					23, 4, 45, 7, -5, 2, -44, 5, 38,
					-- layer=2 filter=112 channel=43
					44, -4, 14, 30, -14, 4, -5, 18, -22,
					-- layer=2 filter=112 channel=44
					5, 8, 11, 8, -6, 9, -11, 6, 4,
					-- layer=2 filter=112 channel=45
					-27, 14, -1, 18, -19, -42, 3, 3, -14,
					-- layer=2 filter=112 channel=46
					10, 7, 24, 3, 40, 6, -22, 46, -14,
					-- layer=2 filter=112 channel=47
					1, -8, 40, 20, 6, -96, 24, -28, 11,
					-- layer=2 filter=112 channel=48
					7, -6, -1, 9, -6, 3, -8, 6, -2,
					-- layer=2 filter=112 channel=49
					13, 49, 8, -43, 44, 73, 56, 46, 55,
					-- layer=2 filter=112 channel=50
					3, 4, -1, 30, 26, 17, 20, 0, 0,
					-- layer=2 filter=112 channel=51
					-26, -8, -3, 1, -6, -6, 18, 9, -6,
					-- layer=2 filter=112 channel=52
					-1, -19, 12, 0, -8, -23, 39, 5, 11,
					-- layer=2 filter=112 channel=53
					-11, 0, -40, -24, -5, 26, -28, 75, 50,
					-- layer=2 filter=112 channel=54
					-18, -58, -22, -45, -37, -40, 11, 0, 16,
					-- layer=2 filter=112 channel=55
					-6, 5, -1, 0, -5, 6, 0, 12, 2,
					-- layer=2 filter=112 channel=56
					3, -11, -13, 0, 10, 9, 9, 5, -9,
					-- layer=2 filter=112 channel=57
					2, 5, 2, 2, -3, 7, 1, -8, 2,
					-- layer=2 filter=112 channel=58
					19, 15, -16, -18, -43, -55, -12, -17, -11,
					-- layer=2 filter=112 channel=59
					22, 34, -53, -2, 21, -26, 35, 0, -14,
					-- layer=2 filter=112 channel=60
					7, 4, -51, -33, -29, -26, 2, -27, 2,
					-- layer=2 filter=112 channel=61
					-13, -36, -57, -20, 15, -24, 46, -4, 32,
					-- layer=2 filter=112 channel=62
					-16, -15, -8, -22, -56, 40, 14, -22, 14,
					-- layer=2 filter=112 channel=63
					41, 19, 9, 7, -7, 0, -7, 8, 16,
					-- layer=2 filter=112 channel=64
					14, 12, 34, 6, -4, 19, -6, -14, 44,
					-- layer=2 filter=112 channel=65
					-32, -18, -67, -5, -3, -33, 25, -50, 28,
					-- layer=2 filter=112 channel=66
					-19, -1, 4, 16, 7, 7, 9, 3, 9,
					-- layer=2 filter=112 channel=67
					-11, -1, 3, 1, 19, 12, -15, 2, -14,
					-- layer=2 filter=112 channel=68
					0, -9, 9, 3, 3, -3, 7, -3, -5,
					-- layer=2 filter=112 channel=69
					11, 15, 35, 25, -5, 5, -5, -29, 41,
					-- layer=2 filter=112 channel=70
					-35, -80, -7, 15, -70, -86, 13, 15, -40,
					-- layer=2 filter=112 channel=71
					-6, 12, -4, 4, 29, 17, -2, 42, -5,
					-- layer=2 filter=112 channel=72
					-15, 39, 15, 14, 3, -23, 11, -19, -62,
					-- layer=2 filter=112 channel=73
					39, 7, -83, 36, 35, 34, 61, 90, 28,
					-- layer=2 filter=112 channel=74
					-3, 0, 7, 10, 31, 2, -19, 15, -8,
					-- layer=2 filter=112 channel=75
					2, -28, -35, -11, -31, -58, 50, 25, 57,
					-- layer=2 filter=112 channel=76
					-13, 15, -101, 10, -34, -34, 39, 27, 12,
					-- layer=2 filter=112 channel=77
					3, -6, 2, 1, -2, 4, -1, -2, -8,
					-- layer=2 filter=112 channel=78
					-16, -12, -7, 4, 18, 21, 30, 6, 4,
					-- layer=2 filter=112 channel=79
					1, -8, 2, 4, 1, -3, -3, 11, 3,
					-- layer=2 filter=112 channel=80
					8, -4, 4, -16, -3, 14, -58, -36, -36,
					-- layer=2 filter=112 channel=81
					-1, -4, 3, -5, 12, 8, -5, 5, -1,
					-- layer=2 filter=112 channel=82
					-6, -8, 8, -9, 6, -4, 11, -5, -4,
					-- layer=2 filter=112 channel=83
					-6, -21, -14, -1, -40, -15, -29, -21, -27,
					-- layer=2 filter=112 channel=84
					0, 2, 7, -9, 6, 8, -1, 2, 0,
					-- layer=2 filter=112 channel=85
					-1, 3, 2, 10, 5, -5, 2, -10, -3,
					-- layer=2 filter=112 channel=86
					21, 16, 8, -2, 6, -20, 3, 25, 4,
					-- layer=2 filter=112 channel=87
					0, 15, 26, -42, -8, -4, -15, 0, -9,
					-- layer=2 filter=112 channel=88
					5, 21, 4, 12, 9, 2, 14, -7, -8,
					-- layer=2 filter=112 channel=89
					-17, 21, -5, -7, -33, 2, 20, 5, -1,
					-- layer=2 filter=112 channel=90
					0, -3, 7, 5, 9, -7, -9, 10, 0,
					-- layer=2 filter=112 channel=91
					7, 28, 10, -5, -27, -26, 28, 17, -6,
					-- layer=2 filter=112 channel=92
					23, 25, 8, 10, -28, -9, -27, -16, -43,
					-- layer=2 filter=112 channel=93
					34, -7, -18, 22, -22, 48, -1, -38, 0,
					-- layer=2 filter=112 channel=94
					-5, -22, -23, 8, 0, 7, 18, 3, 17,
					-- layer=2 filter=112 channel=95
					4, 2, 2, 17, -10, -6, 8, -6, -2,
					-- layer=2 filter=112 channel=96
					-52, -56, -12, -52, -32, 12, 35, 15, 31,
					-- layer=2 filter=112 channel=97
					11, 30, 13, 31, 16, 17, -25, 2, 0,
					-- layer=2 filter=112 channel=98
					10, -16, 26, 15, -17, -92, 13, 8, 2,
					-- layer=2 filter=112 channel=99
					-4, 5, -45, 9, -5, -36, 32, 1, 38,
					-- layer=2 filter=112 channel=100
					10, 19, -15, -35, -37, -15, -46, -24, -31,
					-- layer=2 filter=112 channel=101
					17, -13, -27, 8, 7, 5, 19, 11, 4,
					-- layer=2 filter=112 channel=102
					-23, 2, -14, -4, 10, 31, 34, 10, 74,
					-- layer=2 filter=112 channel=103
					-41, -37, -10, -2, -37, -5, -43, 40, -58,
					-- layer=2 filter=112 channel=104
					4, 29, 21, -19, 27, 43, 21, 41, 51,
					-- layer=2 filter=112 channel=105
					-20, 15, 7, -3, 2, 7, 31, 0, -8,
					-- layer=2 filter=112 channel=106
					-21, -23, -30, 9, -17, -20, 29, 0, -4,
					-- layer=2 filter=112 channel=107
					-14, -29, 20, -16, 13, 39, -45, 51, 7,
					-- layer=2 filter=112 channel=108
					-5, 20, 28, -3, 0, 22, 29, 31, 15,
					-- layer=2 filter=112 channel=109
					1, 4, -1, -4, 8, -17, 7, -12, 3,
					-- layer=2 filter=112 channel=110
					-25, 0, 19, 35, -23, 2, 20, -6, 63,
					-- layer=2 filter=112 channel=111
					-10, 0, -7, 4, 2, -2, -11, -1, -5,
					-- layer=2 filter=112 channel=112
					-14, -8, -31, -7, 24, -29, 14, 4, 11,
					-- layer=2 filter=112 channel=113
					14, 13, 17, 6, 9, -31, -37, 25, 47,
					-- layer=2 filter=112 channel=114
					11, 15, 6, 11, 17, 13, 0, 13, -2,
					-- layer=2 filter=112 channel=115
					7, 0, -12, -6, -4, -1, 1, 11, 9,
					-- layer=2 filter=112 channel=116
					8, -17, 25, 16, 0, 11, 10, -23, -7,
					-- layer=2 filter=112 channel=117
					-51, -69, -56, -18, 10, -39, -16, 9, -5,
					-- layer=2 filter=112 channel=118
					-2, -23, 8, -14, 6, 37, -35, 7, 12,
					-- layer=2 filter=112 channel=119
					-6, -46, -16, 3, -13, -13, 1, -13, -18,
					-- layer=2 filter=112 channel=120
					-1, 5, 5, 0, -8, 4, 0, 9, 6,
					-- layer=2 filter=112 channel=121
					-9, 4, 4, -10, 0, 5, -10, 2, 3,
					-- layer=2 filter=112 channel=122
					-5, -1, -5, 9, 0, 4, 16, 1, 7,
					-- layer=2 filter=112 channel=123
					-14, 11, 4, 8, -14, -66, 7, -15, -6,
					-- layer=2 filter=112 channel=124
					-38, 26, -27, 45, 19, -16, -26, -34, -22,
					-- layer=2 filter=112 channel=125
					0, 6, -4, 0, 2, 3, 12, -11, 11,
					-- layer=2 filter=112 channel=126
					-49, -112, 36, 15, 5, -30, 24, 72, -57,
					-- layer=2 filter=112 channel=127
					39, 34, 20, 23, -25, -25, -17, -33, 5,
					-- layer=2 filter=113 channel=0
					-11, -1, 4, 6, 7, 5, -9, -12, 9,
					-- layer=2 filter=113 channel=1
					1, 3, -12, -3, -9, -10, -6, 2, -10,
					-- layer=2 filter=113 channel=2
					-7, 1, 0, 8, 7, 8, -6, 0, -5,
					-- layer=2 filter=113 channel=3
					-3, 2, -3, -3, -4, -1, 7, 8, -5,
					-- layer=2 filter=113 channel=4
					9, -9, 2, 4, -7, -5, -2, -2, -2,
					-- layer=2 filter=113 channel=5
					2, 3, 2, 6, -9, -7, 5, 7, 8,
					-- layer=2 filter=113 channel=6
					-7, 4, -9, -10, 6, -6, 2, -10, -5,
					-- layer=2 filter=113 channel=7
					-8, 8, 5, -8, -5, -4, -1, 0, 3,
					-- layer=2 filter=113 channel=8
					3, -2, -4, 9, 4, -1, -5, -8, 7,
					-- layer=2 filter=113 channel=9
					-10, -11, 2, -1, 8, 5, 4, -10, 1,
					-- layer=2 filter=113 channel=10
					-5, 2, -7, -11, 3, -2, 8, -8, -5,
					-- layer=2 filter=113 channel=11
					1, -10, 3, 3, -1, 4, -6, -5, -15,
					-- layer=2 filter=113 channel=12
					-11, 3, 1, 5, -1, 4, 2, 6, 5,
					-- layer=2 filter=113 channel=13
					4, -1, 10, -3, 7, -2, 6, 3, -5,
					-- layer=2 filter=113 channel=14
					-10, 5, -8, 1, 1, -11, -9, 0, 0,
					-- layer=2 filter=113 channel=15
					-1, 0, -2, -9, 4, -2, 0, 3, -8,
					-- layer=2 filter=113 channel=16
					5, -6, -12, 5, -8, 4, -8, -6, -9,
					-- layer=2 filter=113 channel=17
					3, 8, 2, 0, -6, -7, -9, 5, 1,
					-- layer=2 filter=113 channel=18
					-4, -7, -7, 5, -12, 4, -6, -6, 3,
					-- layer=2 filter=113 channel=19
					-6, -1, -9, 1, 4, 1, 0, -12, 2,
					-- layer=2 filter=113 channel=20
					-5, 8, 1, 0, 9, -1, 8, 1, -11,
					-- layer=2 filter=113 channel=21
					-8, -11, 0, 3, -4, -4, 0, 5, -11,
					-- layer=2 filter=113 channel=22
					2, 4, -8, 5, -5, 1, 0, 0, 7,
					-- layer=2 filter=113 channel=23
					2, 5, -8, -10, -1, -6, -3, 0, -8,
					-- layer=2 filter=113 channel=24
					1, -6, -6, -8, 3, 6, 3, -10, -9,
					-- layer=2 filter=113 channel=25
					-9, -9, -14, 0, 2, -10, 7, 10, 6,
					-- layer=2 filter=113 channel=26
					5, 4, -5, 4, 1, -3, -9, -10, -10,
					-- layer=2 filter=113 channel=27
					2, -1, -8, -2, -5, -5, 6, -3, -5,
					-- layer=2 filter=113 channel=28
					-6, -2, -8, -8, -10, 1, -5, -11, -1,
					-- layer=2 filter=113 channel=29
					4, 5, 3, 8, 5, -7, -10, -11, 0,
					-- layer=2 filter=113 channel=30
					-12, 4, -7, 8, -8, -12, -11, 4, -7,
					-- layer=2 filter=113 channel=31
					8, -5, -4, -7, 2, 1, 5, 0, -11,
					-- layer=2 filter=113 channel=32
					7, -5, 0, 0, -1, -9, -3, -6, -3,
					-- layer=2 filter=113 channel=33
					-10, -9, -6, 1, 5, 3, 2, -11, -3,
					-- layer=2 filter=113 channel=34
					-9, 8, 0, 1, 9, -6, -3, 5, -11,
					-- layer=2 filter=113 channel=35
					-11, -8, -11, -12, 1, -3, 1, -5, 3,
					-- layer=2 filter=113 channel=36
					-2, -10, 3, 7, -8, -8, -9, 1, -11,
					-- layer=2 filter=113 channel=37
					-10, -9, 7, -1, -5, -12, -10, 5, -3,
					-- layer=2 filter=113 channel=38
					-9, -9, 5, 7, 1, 7, -7, 7, 4,
					-- layer=2 filter=113 channel=39
					3, -6, 5, -9, -10, -1, -9, -8, -9,
					-- layer=2 filter=113 channel=40
					-6, 3, 5, 2, 0, -6, -7, -6, -10,
					-- layer=2 filter=113 channel=41
					-4, -4, -5, -1, -1, 0, -2, 5, 0,
					-- layer=2 filter=113 channel=42
					-4, -1, -6, 8, 11, -8, -4, -7, -1,
					-- layer=2 filter=113 channel=43
					-8, -9, -9, -9, 0, 0, -3, -10, -9,
					-- layer=2 filter=113 channel=44
					-6, 8, 8, -6, 4, 6, 4, 8, -3,
					-- layer=2 filter=113 channel=45
					9, 8, 7, -4, -4, 5, 4, 4, 2,
					-- layer=2 filter=113 channel=46
					-7, 7, -2, -3, 2, -4, 6, 6, 3,
					-- layer=2 filter=113 channel=47
					-4, -9, 6, 1, -1, -7, 3, 4, -7,
					-- layer=2 filter=113 channel=48
					-1, -11, 0, -1, 1, -3, 5, 5, 7,
					-- layer=2 filter=113 channel=49
					6, 6, -10, -7, 1, -4, -10, -5, -4,
					-- layer=2 filter=113 channel=50
					-3, 8, -7, -2, 9, 9, -2, 11, -11,
					-- layer=2 filter=113 channel=51
					-6, 7, 3, -1, -3, 0, -8, 7, 0,
					-- layer=2 filter=113 channel=52
					-7, -9, -9, -5, -10, -2, -13, -2, -4,
					-- layer=2 filter=113 channel=53
					-5, -5, -2, 0, 0, 3, -2, 1, -10,
					-- layer=2 filter=113 channel=54
					5, -6, 7, -9, -12, 7, -2, -4, -6,
					-- layer=2 filter=113 channel=55
					-10, 0, 3, -8, -6, -8, -7, 6, 6,
					-- layer=2 filter=113 channel=56
					1, -10, 1, -4, -11, -2, -7, -10, -10,
					-- layer=2 filter=113 channel=57
					0, 4, 8, 9, -2, 3, -4, -2, -7,
					-- layer=2 filter=113 channel=58
					-9, -8, 9, 7, 4, 8, 3, -1, 0,
					-- layer=2 filter=113 channel=59
					-6, 10, 8, -4, -10, -7, 2, 3, -13,
					-- layer=2 filter=113 channel=60
					5, -10, -4, 5, -1, -1, 5, -8, 4,
					-- layer=2 filter=113 channel=61
					-5, -7, 5, -7, 6, -8, -2, 0, -3,
					-- layer=2 filter=113 channel=62
					-3, 8, -8, -1, 10, -2, -12, -4, 6,
					-- layer=2 filter=113 channel=63
					-4, -7, -5, -6, 0, -5, -4, 0, -9,
					-- layer=2 filter=113 channel=64
					-3, -8, -3, -11, -6, 8, -8, -6, -6,
					-- layer=2 filter=113 channel=65
					2, -10, 4, -11, -6, -6, 2, -2, 6,
					-- layer=2 filter=113 channel=66
					-11, 4, -5, -8, -6, 8, -3, -9, 5,
					-- layer=2 filter=113 channel=67
					-2, 0, -6, 5, -3, -7, -4, -4, 5,
					-- layer=2 filter=113 channel=68
					3, 0, 8, -8, -3, 5, 0, -8, -7,
					-- layer=2 filter=113 channel=69
					-8, -11, 7, 2, 3, -2, -11, -8, 0,
					-- layer=2 filter=113 channel=70
					-1, 9, 8, 2, -13, -8, -13, -1, -4,
					-- layer=2 filter=113 channel=71
					-6, -3, 5, 3, -2, 4, -5, -7, 0,
					-- layer=2 filter=113 channel=72
					0, 8, -2, -1, 2, -9, 3, -1, 1,
					-- layer=2 filter=113 channel=73
					-5, -4, -3, 1, 0, 3, -15, 6, 5,
					-- layer=2 filter=113 channel=74
					2, -2, -9, 1, 7, -7, 0, -5, 1,
					-- layer=2 filter=113 channel=75
					0, 0, -4, 9, 5, -5, -5, 6, 7,
					-- layer=2 filter=113 channel=76
					-2, -8, -11, 5, 5, -8, -12, -1, -5,
					-- layer=2 filter=113 channel=77
					0, -9, -10, -1, 5, -10, -1, -1, -2,
					-- layer=2 filter=113 channel=78
					-10, -7, 3, 0, 3, -1, -4, -9, 7,
					-- layer=2 filter=113 channel=79
					-6, -1, 6, 6, 5, -1, 5, 1, 2,
					-- layer=2 filter=113 channel=80
					-2, -10, -10, -8, -2, 6, -7, -7, -4,
					-- layer=2 filter=113 channel=81
					1, 8, 7, 8, -8, 5, 7, 2, 5,
					-- layer=2 filter=113 channel=82
					5, 1, 4, -5, 2, 3, 4, -8, 0,
					-- layer=2 filter=113 channel=83
					5, -3, -7, -7, -3, 2, -7, 7, 6,
					-- layer=2 filter=113 channel=84
					-10, -4, -9, -10, -6, 6, 4, 2, 6,
					-- layer=2 filter=113 channel=85
					-7, -4, 4, -9, -7, -6, -9, 6, 4,
					-- layer=2 filter=113 channel=86
					10, 8, -12, -3, -4, -4, -2, -4, 6,
					-- layer=2 filter=113 channel=87
					-4, -12, 1, 7, 5, -1, 4, 4, 0,
					-- layer=2 filter=113 channel=88
					0, 3, -1, -2, 5, -9, 8, 6, 6,
					-- layer=2 filter=113 channel=89
					3, 0, -11, -8, -9, -10, 0, -11, 6,
					-- layer=2 filter=113 channel=90
					-8, 2, -2, 7, -7, 9, 0, -4, 6,
					-- layer=2 filter=113 channel=91
					-10, -5, 5, 2, 8, 5, -10, -9, 9,
					-- layer=2 filter=113 channel=92
					-7, -7, 1, 6, 3, 0, 5, -8, -9,
					-- layer=2 filter=113 channel=93
					-10, -9, 8, -6, -2, 5, 5, -10, 8,
					-- layer=2 filter=113 channel=94
					4, 1, 5, -8, 2, -11, 4, -4, 5,
					-- layer=2 filter=113 channel=95
					-4, -10, 8, -7, -4, 5, -1, 7, 4,
					-- layer=2 filter=113 channel=96
					5, -11, -6, -10, -7, -2, -9, -1, 0,
					-- layer=2 filter=113 channel=97
					8, 7, -8, 2, 7, -5, 6, -11, 0,
					-- layer=2 filter=113 channel=98
					7, 1, -2, 0, 2, -7, -11, -8, 3,
					-- layer=2 filter=113 channel=99
					6, 0, 2, -12, 0, -1, -5, 6, 2,
					-- layer=2 filter=113 channel=100
					0, -2, 8, -9, -12, -5, 0, -7, 1,
					-- layer=2 filter=113 channel=101
					-1, -8, -6, 7, 1, -9, -4, -8, 5,
					-- layer=2 filter=113 channel=102
					0, -1, -12, 3, -8, 8, 6, 4, 3,
					-- layer=2 filter=113 channel=103
					-10, 0, 0, -10, -10, 2, 6, 3, 1,
					-- layer=2 filter=113 channel=104
					0, -2, -8, 1, -5, 3, -11, -8, -1,
					-- layer=2 filter=113 channel=105
					3, 2, 0, -6, -3, 10, -8, -6, -5,
					-- layer=2 filter=113 channel=106
					-2, -7, 4, 6, 2, -1, -5, 7, 7,
					-- layer=2 filter=113 channel=107
					7, -2, 6, 2, 7, 3, -1, -9, 6,
					-- layer=2 filter=113 channel=108
					-9, -9, -3, -4, -11, -7, -3, 8, -7,
					-- layer=2 filter=113 channel=109
					5, -11, 7, 2, 1, 4, -10, -9, 4,
					-- layer=2 filter=113 channel=110
					3, -11, -9, -3, 5, -5, 4, -1, -2,
					-- layer=2 filter=113 channel=111
					6, -10, -6, 2, -7, 5, -6, -7, -9,
					-- layer=2 filter=113 channel=112
					-5, -7, -2, -4, -9, 6, 5, -4, -9,
					-- layer=2 filter=113 channel=113
					-5, 3, 4, -7, -11, -5, 4, -5, 2,
					-- layer=2 filter=113 channel=114
					1, 3, 0, 0, -5, -2, 7, -6, -11,
					-- layer=2 filter=113 channel=115
					5, 0, 7, -8, 5, 6, -3, -3, -7,
					-- layer=2 filter=113 channel=116
					-1, -4, 5, -2, -10, -8, 6, 2, 0,
					-- layer=2 filter=113 channel=117
					-14, -3, -8, -10, -14, -12, 2, -9, 1,
					-- layer=2 filter=113 channel=118
					-10, 4, -7, 0, 3, 1, 7, -1, 6,
					-- layer=2 filter=113 channel=119
					-7, -9, -8, -5, -5, 4, 2, 2, 8,
					-- layer=2 filter=113 channel=120
					8, -10, 6, -6, 5, 3, -2, 0, 0,
					-- layer=2 filter=113 channel=121
					-9, 3, 4, -2, 2, 0, -11, 2, -3,
					-- layer=2 filter=113 channel=122
					-7, -9, 9, 8, 9, 6, 0, 5, 4,
					-- layer=2 filter=113 channel=123
					2, 1, -9, -3, 0, -3, 4, -5, 4,
					-- layer=2 filter=113 channel=124
					-5, 2, 1, 0, 6, 8, -11, -9, 6,
					-- layer=2 filter=113 channel=125
					-10, -3, -3, -7, 5, -3, -7, -1, -3,
					-- layer=2 filter=113 channel=126
					1, -11, -4, -5, -4, 0, 3, 8, 1,
					-- layer=2 filter=113 channel=127
					-9, 7, 9, -9, -10, 7, 6, 8, -5,
					-- layer=2 filter=114 channel=0
					-22, -9, 13, -35, -5, 0, 0, -20, 2,
					-- layer=2 filter=114 channel=1
					-9, -24, -24, -8, -2, 31, 0, -13, -66,
					-- layer=2 filter=114 channel=2
					-7, -7, 0, -6, 5, 7, 5, 6, -5,
					-- layer=2 filter=114 channel=3
					-5, -39, -30, -31, -25, -1, 11, 6, 35,
					-- layer=2 filter=114 channel=4
					1, 4, -35, -16, -10, 9, -18, -12, 30,
					-- layer=2 filter=114 channel=5
					26, 14, 34, -29, 6, 14, -18, -8, 3,
					-- layer=2 filter=114 channel=6
					-16, 8, -7, 3, 25, 31, 26, 9, -13,
					-- layer=2 filter=114 channel=7
					-2, 44, 36, -21, 30, 26, 14, -7, 16,
					-- layer=2 filter=114 channel=8
					3, -5, -5, -7, -3, 5, 3, 10, -7,
					-- layer=2 filter=114 channel=9
					-31, -9, -38, -14, -14, 6, -40, -23, -72,
					-- layer=2 filter=114 channel=10
					-15, -12, -3, -59, -30, -9, -7, -35, 24,
					-- layer=2 filter=114 channel=11
					-1, 23, 10, -12, 6, 3, -29, 25, 27,
					-- layer=2 filter=114 channel=12
					19, -6, 22, 3, 29, 6, 7, 26, -47,
					-- layer=2 filter=114 channel=13
					-2, -5, 1, 4, 5, -1, 10, 0, 4,
					-- layer=2 filter=114 channel=14
					16, 9, 23, -2, 0, 9, -24, -11, -55,
					-- layer=2 filter=114 channel=15
					-46, 10, 4, -48, -20, -34, -102, 0, -76,
					-- layer=2 filter=114 channel=16
					-14, 14, -31, -21, 4, -31, 27, 26, -17,
					-- layer=2 filter=114 channel=17
					4, -3, -10, -4, 5, -5, 6, 2, -10,
					-- layer=2 filter=114 channel=18
					0, 8, 9, -19, 6, -25, 3, -19, -31,
					-- layer=2 filter=114 channel=19
					-21, -18, -43, 3, 4, -1, -6, -16, -5,
					-- layer=2 filter=114 channel=20
					4, 6, -5, -12, -1, -10, -2, -7, 1,
					-- layer=2 filter=114 channel=21
					-5, -10, 0, 10, 2, 0, 19, 9, 12,
					-- layer=2 filter=114 channel=22
					5, -7, -2, -3, 0, -7, -5, 0, -9,
					-- layer=2 filter=114 channel=23
					-14, -7, -8, -4, -34, -21, 52, 49, 35,
					-- layer=2 filter=114 channel=24
					34, -14, -35, 22, -6, -38, 45, 44, 19,
					-- layer=2 filter=114 channel=25
					15, -31, -9, 32, -10, -36, 67, 67, 30,
					-- layer=2 filter=114 channel=26
					-4, -3, -9, 8, -6, -5, -7, -4, -3,
					-- layer=2 filter=114 channel=27
					-8, 1, -7, 36, 54, 43, -11, 21, 4,
					-- layer=2 filter=114 channel=28
					3, 34, 14, 37, 33, -14, 46, 3, 15,
					-- layer=2 filter=114 channel=29
					0, 10, 8, -9, -4, -5, -3, -6, 4,
					-- layer=2 filter=114 channel=30
					9, 4, -2, 45, -2, 3, -28, -12, -20,
					-- layer=2 filter=114 channel=31
					-24, -43, 11, 27, 19, -27, 18, 34, 18,
					-- layer=2 filter=114 channel=32
					-9, 6, -4, -5, -6, -3, -5, 2, -6,
					-- layer=2 filter=114 channel=33
					27, -10, -5, -25, -38, -10, 6, -19, 10,
					-- layer=2 filter=114 channel=34
					32, -9, 9, 36, 8, -37, 14, -13, -50,
					-- layer=2 filter=114 channel=35
					1, 42, -27, 12, 20, -94, 53, 10, 2,
					-- layer=2 filter=114 channel=36
					1, 0, -4, 1, -17, 8, -1, 0, -7,
					-- layer=2 filter=114 channel=37
					9, 20, 49, -6, -3, 26, -22, -2, 21,
					-- layer=2 filter=114 channel=38
					47, 24, 2, 6, 26, 5, -12, -4, -26,
					-- layer=2 filter=114 channel=39
					8, -1, 10, -23, -13, -3, -22, 21, -35,
					-- layer=2 filter=114 channel=40
					-11, 33, 11, -25, -59, 16, 16, -28, -17,
					-- layer=2 filter=114 channel=41
					3, -8, 0, -5, 9, 0, -5, 4, 5,
					-- layer=2 filter=114 channel=42
					-25, 18, 14, 32, -8, -6, 33, 38, 12,
					-- layer=2 filter=114 channel=43
					12, -42, -26, -62, 6, -17, 14, 6, 21,
					-- layer=2 filter=114 channel=44
					8, 8, -5, -2, 6, -6, -8, -5, -11,
					-- layer=2 filter=114 channel=45
					9, -27, -70, -9, 3, -24, 33, 71, 35,
					-- layer=2 filter=114 channel=46
					12, -29, 17, -15, -21, 0, -31, -22, 17,
					-- layer=2 filter=114 channel=47
					42, 63, 20, 4, 21, -3, 2, 0, -28,
					-- layer=2 filter=114 channel=48
					0, 0, 5, 3, 3, 3, -2, -10, 0,
					-- layer=2 filter=114 channel=49
					9, -9, -7, 1, 1, 18, -16, 19, -17,
					-- layer=2 filter=114 channel=50
					-2, -18, -1, 0, 14, 1, -5, -17, 4,
					-- layer=2 filter=114 channel=51
					-2, 4, 45, -10, -5, 4, -9, -5, 9,
					-- layer=2 filter=114 channel=52
					11, -8, 37, -44, 5, 25, -45, 4, 31,
					-- layer=2 filter=114 channel=53
					31, 2, 37, 0, 26, 35, -13, 11, -54,
					-- layer=2 filter=114 channel=54
					-22, -20, 22, -21, -29, -35, 35, 15, 9,
					-- layer=2 filter=114 channel=55
					-3, 0, 12, -1, 0, 6, -8, 12, -15,
					-- layer=2 filter=114 channel=56
					-3, 16, 18, -18, 15, 4, -23, 19, 7,
					-- layer=2 filter=114 channel=57
					3, -1, 3, 8, -2, 3, 19, -3, -4,
					-- layer=2 filter=114 channel=58
					32, 14, -2, 19, 16, 21, -28, 32, 9,
					-- layer=2 filter=114 channel=59
					46, -26, -46, 21, 5, -7, -12, -25, -63,
					-- layer=2 filter=114 channel=60
					-15, -43, -3, -22, -8, -42, -3, -77, -11,
					-- layer=2 filter=114 channel=61
					-23, 2, 30, 13, 27, -28, 24, -16, -4,
					-- layer=2 filter=114 channel=62
					-26, 2, -44, 8, -11, 20, -3, 19, -9,
					-- layer=2 filter=114 channel=63
					-12, -3, 36, -23, 26, -6, -9, 10, -36,
					-- layer=2 filter=114 channel=64
					-14, -11, -25, 17, -21, 0, 25, 23, 8,
					-- layer=2 filter=114 channel=65
					-15, -7, 34, 19, 15, 2, -3, -10, 0,
					-- layer=2 filter=114 channel=66
					19, 14, 25, -16, 14, -4, 17, -1, -21,
					-- layer=2 filter=114 channel=67
					-29, -11, -47, -8, -2, 12, -35, -25, -44,
					-- layer=2 filter=114 channel=68
					-3, -9, 5, -2, -2, 10, -4, -4, -5,
					-- layer=2 filter=114 channel=69
					-22, -1, -17, 0, 17, 0, 29, 28, -19,
					-- layer=2 filter=114 channel=70
					0, 27, 17, 0, -37, -33, 19, -20, 3,
					-- layer=2 filter=114 channel=71
					-13, 3, -45, 27, 52, 14, 3, -15, -1,
					-- layer=2 filter=114 channel=72
					-24, 34, 38, -30, 1, -11, 1, -23, -17,
					-- layer=2 filter=114 channel=73
					26, 13, -65, 80, 53, 22, 89, 68, 54,
					-- layer=2 filter=114 channel=74
					9, 0, -23, 20, 4, 9, -28, -29, -5,
					-- layer=2 filter=114 channel=75
					-43, 4, 13, -17, -27, -1, 10, 8, -12,
					-- layer=2 filter=114 channel=76
					-1, -29, 33, -27, -16, -23, 16, 28, 18,
					-- layer=2 filter=114 channel=77
					-8, -5, -4, 9, 0, -1, -1, 1, 3,
					-- layer=2 filter=114 channel=78
					20, -5, 7, 0, -18, 1, 10, 17, 45,
					-- layer=2 filter=114 channel=79
					11, -7, 7, 1, 6, -6, -9, 5, 0,
					-- layer=2 filter=114 channel=80
					-9, -13, -20, 7, -24, 11, -19, -18, 5,
					-- layer=2 filter=114 channel=81
					-5, 3, -2, -7, -8, -12, -1, -5, 6,
					-- layer=2 filter=114 channel=82
					-8, -9, -4, 9, -2, 6, 10, -6, 3,
					-- layer=2 filter=114 channel=83
					-19, -3, -6, 3, 8, -13, 16, 14, 9,
					-- layer=2 filter=114 channel=84
					-2, -5, 2, -4, 6, -4, 8, -8, 9,
					-- layer=2 filter=114 channel=85
					-5, 9, 6, 3, 7, -1, 4, -1, 0,
					-- layer=2 filter=114 channel=86
					-12, 2, 5, -7, 8, 8, -5, 1, 2,
					-- layer=2 filter=114 channel=87
					27, 14, -17, -4, -36, -52, 2, 16, 24,
					-- layer=2 filter=114 channel=88
					1, -22, -21, 17, 7, 20, -13, -35, -5,
					-- layer=2 filter=114 channel=89
					8, -18, -25, 4, -8, 2, -9, -5, -74,
					-- layer=2 filter=114 channel=90
					-4, 1, 0, -1, -4, -9, 1, -4, 9,
					-- layer=2 filter=114 channel=91
					-26, 10, -5, -12, -25, -21, 8, 8, -23,
					-- layer=2 filter=114 channel=92
					11, 12, 7, -4, 15, 21, 19, -6, -62,
					-- layer=2 filter=114 channel=93
					-38, -25, -20, 57, 8, 43, 27, -35, 20,
					-- layer=2 filter=114 channel=94
					-13, -12, 15, -15, 38, 7, 15, 5, -47,
					-- layer=2 filter=114 channel=95
					7, 9, 18, 7, 8, 17, 19, 14, 16,
					-- layer=2 filter=114 channel=96
					-22, -33, 15, 8, -7, 53, 17, 47, 23,
					-- layer=2 filter=114 channel=97
					4, 5, -3, -2, 0, 29, -34, -15, -13,
					-- layer=2 filter=114 channel=98
					-16, 48, 22, 1, 10, -38, 27, 1, 12,
					-- layer=2 filter=114 channel=99
					-11, -10, 15, 2, 23, -12, -51, -18, 41,
					-- layer=2 filter=114 channel=100
					44, -3, -2, 8, 18, 8, -20, 12, 0,
					-- layer=2 filter=114 channel=101
					7, -18, -9, 26, 44, -1, 38, 2, -9,
					-- layer=2 filter=114 channel=102
					0, -19, 33, -16, 36, 35, -25, 40, 6,
					-- layer=2 filter=114 channel=103
					-35, -7, 34, -36, -39, -26, -70, -17, -33,
					-- layer=2 filter=114 channel=104
					15, 5, -15, -20, 14, 22, -30, 17, -26,
					-- layer=2 filter=114 channel=105
					-2, 21, 6, -9, 2, -2, 16, 10, 34,
					-- layer=2 filter=114 channel=106
					6, -11, -74, 7, -8, -33, 32, 10, -28,
					-- layer=2 filter=114 channel=107
					-21, 22, 16, 58, 14, 2, -22, 9, -59,
					-- layer=2 filter=114 channel=108
					-22, 25, 19, 12, 26, 43, -38, 5, -43,
					-- layer=2 filter=114 channel=109
					19, -5, -6, -4, -7, 0, 11, -5, 3,
					-- layer=2 filter=114 channel=110
					17, -16, -10, 52, 1, -21, 75, 71, 11,
					-- layer=2 filter=114 channel=111
					-12, 7, -7, 9, 11, 3, -2, -5, -4,
					-- layer=2 filter=114 channel=112
					-47, -9, -16, 5, 1, -12, -9, -14, 1,
					-- layer=2 filter=114 channel=113
					-16, 9, 49, 16, 22, 7, -30, 2, 8,
					-- layer=2 filter=114 channel=114
					-6, 14, 22, 6, -9, 1, 2, 1, 11,
					-- layer=2 filter=114 channel=115
					-8, 5, 1, 9, -12, 9, 2, -9, 10,
					-- layer=2 filter=114 channel=116
					-5, -6, -33, -76, -32, -9, -8, 15, -19,
					-- layer=2 filter=114 channel=117
					-54, 63, 5, 17, 51, 9, 16, -8, 20,
					-- layer=2 filter=114 channel=118
					0, -18, -30, -1, -53, -10, 10, 14, 57,
					-- layer=2 filter=114 channel=119
					-7, 29, -50, -1, 34, -46, 35, 23, 3,
					-- layer=2 filter=114 channel=120
					3, 0, 9, -5, 1, 0, 2, 7, -9,
					-- layer=2 filter=114 channel=121
					-4, 5, 1, -4, -9, 4, 9, -1, -1,
					-- layer=2 filter=114 channel=122
					-11, -7, -10, 0, 1, 3, 2, -2, -8,
					-- layer=2 filter=114 channel=123
					-8, 5, 15, -50, 26, -22, 2, -12, -10,
					-- layer=2 filter=114 channel=124
					-36, -32, -50, -4, -24, -37, -7, -22, 13,
					-- layer=2 filter=114 channel=125
					10, -1, 6, -10, 0, -6, -6, 2, -3,
					-- layer=2 filter=114 channel=126
					46, 17, 9, 3, 61, -28, 17, -21, 3,
					-- layer=2 filter=114 channel=127
					-13, 10, 18, 17, 14, -22, 22, -5, -8,
					-- layer=2 filter=115 channel=0
					2, 12, 2, -29, 2, -4, -41, -13, 5,
					-- layer=2 filter=115 channel=1
					-2, 23, 20, 5, 5, -4, 26, 36, 26,
					-- layer=2 filter=115 channel=2
					-6, 0, 9, 0, -11, -3, -10, 7, -11,
					-- layer=2 filter=115 channel=3
					-31, -39, -28, 5, -25, 9, -15, -46, -13,
					-- layer=2 filter=115 channel=4
					21, -2, 7, -7, -5, -16, -25, -10, 13,
					-- layer=2 filter=115 channel=5
					9, 14, -19, -5, 3, 4, 30, -13, 19,
					-- layer=2 filter=115 channel=6
					-9, 5, 31, -12, 29, 2, 1, 7, 11,
					-- layer=2 filter=115 channel=7
					-10, -9, 8, 31, 9, 0, 5, 9, -49,
					-- layer=2 filter=115 channel=8
					2, 7, -6, -5, -6, -3, -9, -7, 7,
					-- layer=2 filter=115 channel=9
					3, -8, -42, 10, -6, -57, -38, -31, -23,
					-- layer=2 filter=115 channel=10
					-2, -4, -26, -11, -7, 12, -40, -23, 8,
					-- layer=2 filter=115 channel=11
					-18, -9, -9, -21, -18, -17, -20, -4, 2,
					-- layer=2 filter=115 channel=12
					-19, 40, 32, -31, -6, -12, 26, 52, 0,
					-- layer=2 filter=115 channel=13
					-3, 2, -3, -6, 7, 0, 2, 7, 10,
					-- layer=2 filter=115 channel=14
					-13, 2, -7, -10, -14, -27, 18, 44, 18,
					-- layer=2 filter=115 channel=15
					-26, -3, -32, -53, 13, 62, -10, -5, 41,
					-- layer=2 filter=115 channel=16
					58, 15, 18, 21, 16, -3, 1, -5, -40,
					-- layer=2 filter=115 channel=17
					-11, -9, -6, -6, 0, -1, 6, 10, 10,
					-- layer=2 filter=115 channel=18
					15, -7, 1, -16, 15, -9, -11, 23, 20,
					-- layer=2 filter=115 channel=19
					23, 18, 28, 1, 22, 23, 21, 30, -3,
					-- layer=2 filter=115 channel=20
					0, -8, -8, 7, -9, -11, -3, 0, -5,
					-- layer=2 filter=115 channel=21
					-7, -12, 0, 5, -5, -9, 5, 12, 6,
					-- layer=2 filter=115 channel=22
					7, 4, -2, -8, -14, 0, 1, -3, 0,
					-- layer=2 filter=115 channel=23
					-5, 20, -4, 14, -3, -2, -13, 6, 14,
					-- layer=2 filter=115 channel=24
					40, -12, -1, 37, -3, -14, -15, 10, -3,
					-- layer=2 filter=115 channel=25
					-16, -10, -6, -1, -22, -39, 0, -11, -8,
					-- layer=2 filter=115 channel=26
					-4, -7, -4, 1, 0, 1, 7, -3, -6,
					-- layer=2 filter=115 channel=27
					30, -3, 0, 22, 14, 2, -4, 1, -3,
					-- layer=2 filter=115 channel=28
					-26, 11, 58, -34, 7, -20, -1, -17, -11,
					-- layer=2 filter=115 channel=29
					1, -4, -1, 5, 0, -1, 2, -9, 7,
					-- layer=2 filter=115 channel=30
					19, -17, -9, 0, -14, -21, -37, -1, 14,
					-- layer=2 filter=115 channel=31
					-26, -44, -37, 30, -13, 47, -25, -5, 53,
					-- layer=2 filter=115 channel=32
					8, -1, -3, 7, 0, -1, -3, 8, -3,
					-- layer=2 filter=115 channel=33
					-33, -16, 22, 19, 12, 27, 37, -6, -14,
					-- layer=2 filter=115 channel=34
					4, -42, -38, -26, -2, -23, -41, -42, -51,
					-- layer=2 filter=115 channel=35
					-6, 26, 51, -7, 1, -10, 14, -13, -35,
					-- layer=2 filter=115 channel=36
					-16, -4, -2, -2, 1, 2, 10, 2, 2,
					-- layer=2 filter=115 channel=37
					-1, 19, -2, 0, 0, 20, -7, 14, 9,
					-- layer=2 filter=115 channel=38
					17, -8, -13, -17, -41, 14, -2, -6, -3,
					-- layer=2 filter=115 channel=39
					-17, -21, -13, 1, -1, -16, -9, -10, 5,
					-- layer=2 filter=115 channel=40
					-7, -12, -23, 2, -17, 48, -15, -19, 11,
					-- layer=2 filter=115 channel=41
					-8, -7, 2, 7, 11, 1, 1, -5, -1,
					-- layer=2 filter=115 channel=42
					-5, 10, 4, 2, -7, 9, -18, 21, -12,
					-- layer=2 filter=115 channel=43
					-16, 16, -10, -7, 1, 33, -15, 10, 2,
					-- layer=2 filter=115 channel=44
					2, -6, -7, -4, -5, 9, 9, -5, -10,
					-- layer=2 filter=115 channel=45
					8, 28, 49, 36, 2, 24, -24, -7, -5,
					-- layer=2 filter=115 channel=46
					-29, -25, -47, -17, 13, -16, -69, -5, 31,
					-- layer=2 filter=115 channel=47
					-18, -22, 18, -40, 11, -7, -18, -26, -43,
					-- layer=2 filter=115 channel=48
					-9, 2, 3, -1, 4, -1, -7, 1, -7,
					-- layer=2 filter=115 channel=49
					30, 7, -10, -35, 27, -22, -21, 17, 10,
					-- layer=2 filter=115 channel=50
					-3, 26, 4, -9, -16, -1, 13, 19, 30,
					-- layer=2 filter=115 channel=51
					0, -3, 9, -32, -23, -5, -11, -4, -4,
					-- layer=2 filter=115 channel=52
					-11, 35, 16, 11, 9, -3, -27, 29, 23,
					-- layer=2 filter=115 channel=53
					-16, -90, -11, -36, -36, -51, 25, 17, -30,
					-- layer=2 filter=115 channel=54
					-7, 13, 45, -2, 18, 9, 17, -5, 19,
					-- layer=2 filter=115 channel=55
					-9, 0, 0, 6, -5, -1, -6, -2, -5,
					-- layer=2 filter=115 channel=56
					-11, -11, 2, -1, -2, -8, -1, 17, 4,
					-- layer=2 filter=115 channel=57
					-10, -4, -2, -8, 12, 15, -5, -14, -4,
					-- layer=2 filter=115 channel=58
					-24, 32, 38, -28, -4, 10, 22, 26, 17,
					-- layer=2 filter=115 channel=59
					-25, 29, 49, -21, 24, 0, 14, 13, -28,
					-- layer=2 filter=115 channel=60
					0, -21, -3, -37, -6, -32, 28, -2, -43,
					-- layer=2 filter=115 channel=61
					10, 21, 23, -1, -17, -30, 5, -2, -76,
					-- layer=2 filter=115 channel=62
					-1, 13, -1, -10, 32, 10, -16, 4, 28,
					-- layer=2 filter=115 channel=63
					5, 3, 36, -7, -12, 3, -4, -13, -34,
					-- layer=2 filter=115 channel=64
					14, 5, -18, 47, 0, -20, 25, 22, -20,
					-- layer=2 filter=115 channel=65
					17, 13, 61, -12, -7, -12, -6, 24, -20,
					-- layer=2 filter=115 channel=66
					20, 9, -9, -5, 59, 39, -18, 14, 29,
					-- layer=2 filter=115 channel=67
					-20, -2, -52, -6, 0, -32, -43, -61, -1,
					-- layer=2 filter=115 channel=68
					-8, -5, -1, -10, 8, 4, -2, 3, -5,
					-- layer=2 filter=115 channel=69
					2, 0, 5, 24, -18, -6, 11, 37, -2,
					-- layer=2 filter=115 channel=70
					17, 29, 79, -1, 11, 33, -4, -13, -24,
					-- layer=2 filter=115 channel=71
					-19, -21, -29, 9, -18, -27, -26, -37, -3,
					-- layer=2 filter=115 channel=72
					8, -42, 0, -10, -2, 2, 26, 2, -10,
					-- layer=2 filter=115 channel=73
					-45, -17, -22, -24, -2, -28, -24, 24, 45,
					-- layer=2 filter=115 channel=74
					-7, -11, -30, 3, 17, 0, -13, -4, 28,
					-- layer=2 filter=115 channel=75
					15, -28, 11, -10, 3, -37, 13, 63, 17,
					-- layer=2 filter=115 channel=76
					-16, -18, 0, -75, -53, -43, -18, -20, -7,
					-- layer=2 filter=115 channel=77
					-5, 2, 4, 4, 0, -10, -3, 1, 8,
					-- layer=2 filter=115 channel=78
					-8, 0, -34, 16, -6, -16, -6, 3, 25,
					-- layer=2 filter=115 channel=79
					-10, -4, -3, 2, 8, -10, -8, 3, 6,
					-- layer=2 filter=115 channel=80
					7, -39, -30, -29, 12, -3, -27, -37, 14,
					-- layer=2 filter=115 channel=81
					-7, -7, -15, -6, 0, -1, -10, -3, 2,
					-- layer=2 filter=115 channel=82
					6, 6, 8, 0, -9, 4, 9, 4, -1,
					-- layer=2 filter=115 channel=83
					16, 23, 24, 12, 15, -2, -19, -24, -20,
					-- layer=2 filter=115 channel=84
					5, -1, 0, 4, 0, 3, 6, -2, -2,
					-- layer=2 filter=115 channel=85
					12, 0, -3, 16, 21, 14, 0, 3, -18,
					-- layer=2 filter=115 channel=86
					-2, 0, -1, -13, 27, -11, 7, -17, -11,
					-- layer=2 filter=115 channel=87
					-14, -49, -4, -38, -34, -6, -27, -46, -16,
					-- layer=2 filter=115 channel=88
					-8, 15, 11, -9, -15, -21, -5, -12, 27,
					-- layer=2 filter=115 channel=89
					-35, -10, 5, -22, 18, -4, 17, 25, 5,
					-- layer=2 filter=115 channel=90
					-5, -4, -7, -1, -5, -10, -7, 7, -2,
					-- layer=2 filter=115 channel=91
					-7, -13, 17, -23, 24, 1, 9, 12, -29,
					-- layer=2 filter=115 channel=92
					13, 28, 10, -3, 12, 18, 23, 0, 7,
					-- layer=2 filter=115 channel=93
					3, 26, 42, -13, 11, 50, 42, -8, -31,
					-- layer=2 filter=115 channel=94
					28, 11, 17, 19, 18, -25, 6, 28, -34,
					-- layer=2 filter=115 channel=95
					8, 10, 0, 14, 1, -9, -1, -4, 5,
					-- layer=2 filter=115 channel=96
					15, 62, 69, 31, 85, 22, 28, 6, -35,
					-- layer=2 filter=115 channel=97
					-2, -23, -4, 6, 16, 15, 7, -9, -2,
					-- layer=2 filter=115 channel=98
					1, -14, 30, -18, -12, 6, -15, -10, -22,
					-- layer=2 filter=115 channel=99
					-42, 46, 1, 22, 7, 1, -5, 36, -4,
					-- layer=2 filter=115 channel=100
					15, -8, -30, -15, -29, -11, -17, -2, -19,
					-- layer=2 filter=115 channel=101
					-50, -53, 16, 5, -24, 9, -7, -42, -49,
					-- layer=2 filter=115 channel=102
					22, 37, 15, -2, 39, -20, -11, 21, -12,
					-- layer=2 filter=115 channel=103
					36, 44, 52, 46, 10, -24, -11, 31, 31,
					-- layer=2 filter=115 channel=104
					0, -33, 1, -47, 19, -2, 5, 22, 12,
					-- layer=2 filter=115 channel=105
					11, 9, 13, 8, 43, 4, -7, 0, -46,
					-- layer=2 filter=115 channel=106
					-40, -32, 36, -21, -6, 8, 8, -2, -13,
					-- layer=2 filter=115 channel=107
					4, -22, -13, -13, -59, -13, 17, 36, -29,
					-- layer=2 filter=115 channel=108
					13, -3, -5, -7, -16, -6, -12, 12, 5,
					-- layer=2 filter=115 channel=109
					-7, -4, -8, 1, 7, -12, -7, 7, 6,
					-- layer=2 filter=115 channel=110
					27, 8, 10, 54, -10, -30, 23, 0, -27,
					-- layer=2 filter=115 channel=111
					11, -7, 4, 0, -4, 7, -3, 0, -8,
					-- layer=2 filter=115 channel=112
					6, 21, 11, -29, -42, -28, -40, -28, -13,
					-- layer=2 filter=115 channel=113
					13, 1, 36, -14, -21, -10, -41, -6, -18,
					-- layer=2 filter=115 channel=114
					12, 22, 24, -8, 9, 16, 11, 24, 24,
					-- layer=2 filter=115 channel=115
					10, -10, 2, 6, 0, 9, -11, 11, 7,
					-- layer=2 filter=115 channel=116
					-6, -10, 20, -24, -19, -13, -49, -22, 16,
					-- layer=2 filter=115 channel=117
					-28, -3, -15, -3, 32, -28, 38, 34, 0,
					-- layer=2 filter=115 channel=118
					4, -38, -10, 19, 28, 12, -45, -24, 19,
					-- layer=2 filter=115 channel=119
					19, 2, 21, 22, 13, -11, -20, -17, 7,
					-- layer=2 filter=115 channel=120
					6, -4, 2, 3, 7, -5, -2, -9, -1,
					-- layer=2 filter=115 channel=121
					0, 9, 2, 7, -5, 0, 10, 1, -3,
					-- layer=2 filter=115 channel=122
					8, 2, 0, -6, 10, -12, 3, 10, -5,
					-- layer=2 filter=115 channel=123
					0, -29, 6, 14, 11, 4, 13, 1, 3,
					-- layer=2 filter=115 channel=124
					5, 1, -19, 7, -12, 53, 5, -18, 64,
					-- layer=2 filter=115 channel=125
					-2, 1, 0, -10, 8, 12, 4, 4, 1,
					-- layer=2 filter=115 channel=126
					-26, -37, -22, -6, 11, -14, 29, -15, -7,
					-- layer=2 filter=115 channel=127
					11, -5, 17, -4, -2, -21, 0, 8, 17,
					-- layer=2 filter=116 channel=0
					19, -10, -13, -16, -13, -3, -9, 0, 18,
					-- layer=2 filter=116 channel=1
					44, 27, -33, -12, -6, -74, 4, 33, 15,
					-- layer=2 filter=116 channel=2
					4, -1, 5, 10, -6, 7, 0, -4, 1,
					-- layer=2 filter=116 channel=3
					26, 13, 12, -2, 29, 47, 3, 13, 23,
					-- layer=2 filter=116 channel=4
					6, 19, 40, -4, 16, 38, 2, -19, 9,
					-- layer=2 filter=116 channel=5
					0, -22, -20, 3, -20, -38, 9, 13, -5,
					-- layer=2 filter=116 channel=6
					-8, -22, -10, 34, 7, -11, 17, 29, 39,
					-- layer=2 filter=116 channel=7
					37, 18, -24, -9, 66, 77, 21, 31, 57,
					-- layer=2 filter=116 channel=8
					-8, -5, -6, 4, -9, 0, -11, 0, 7,
					-- layer=2 filter=116 channel=9
					2, 10, 5, 9, -18, -30, 3, -23, 12,
					-- layer=2 filter=116 channel=10
					12, 6, -17, -9, -3, -2, -13, -20, 13,
					-- layer=2 filter=116 channel=11
					2, -17, -16, -3, -10, -38, 32, -7, -6,
					-- layer=2 filter=116 channel=12
					58, 6, -3, -21, -1, -26, -7, 10, 16,
					-- layer=2 filter=116 channel=13
					12, 9, 7, 6, -6, -7, 9, -3, -2,
					-- layer=2 filter=116 channel=14
					43, 4, -25, -24, -32, -60, -23, 18, 31,
					-- layer=2 filter=116 channel=15
					-21, 24, -60, 0, -46, -15, -12, -34, -41,
					-- layer=2 filter=116 channel=16
					-53, -21, -23, -24, -10, 14, -29, -31, 2,
					-- layer=2 filter=116 channel=17
					0, -1, 8, 2, -7, -8, -4, -8, 3,
					-- layer=2 filter=116 channel=18
					-20, -7, 11, 0, -15, 0, 20, -61, -2,
					-- layer=2 filter=116 channel=19
					-12, -18, -59, 29, 9, -49, 14, 40, 35,
					-- layer=2 filter=116 channel=20
					-6, -8, -1, 2, -3, 5, 12, 9, 7,
					-- layer=2 filter=116 channel=21
					16, 14, 15, -2, 14, 4, -6, -13, -1,
					-- layer=2 filter=116 channel=22
					-6, 13, 0, 5, -1, -1, -1, 12, 6,
					-- layer=2 filter=116 channel=23
					35, 34, 9, 5, 19, 54, -28, 4, -10,
					-- layer=2 filter=116 channel=24
					-21, 5, 26, -39, -6, 39, 8, -13, 20,
					-- layer=2 filter=116 channel=25
					-13, -5, 6, -34, 15, 19, -10, 8, 19,
					-- layer=2 filter=116 channel=26
					-9, -8, -8, 2, -4, -2, -3, 0, 2,
					-- layer=2 filter=116 channel=27
					-18, -72, -66, 37, -21, -62, 43, 20, -26,
					-- layer=2 filter=116 channel=28
					37, -35, -22, -9, 56, 80, 1, 14, 15,
					-- layer=2 filter=116 channel=29
					-5, 3, -7, -4, -7, 7, 2, 7, -8,
					-- layer=2 filter=116 channel=30
					6, 20, -6, 28, -11, -36, 11, -28, -26,
					-- layer=2 filter=116 channel=31
					14, 14, -1, 47, -71, -30, 9, -9, 13,
					-- layer=2 filter=116 channel=32
					10, 5, 10, -8, 3, 0, 5, 0, -2,
					-- layer=2 filter=116 channel=33
					11, 2, -27, -26, 27, 20, -39, 71, 51,
					-- layer=2 filter=116 channel=34
					54, 25, -44, 2, -22, -29, 81, -27, -25,
					-- layer=2 filter=116 channel=35
					-15, -19, -9, -23, 36, 36, 5, -36, -12,
					-- layer=2 filter=116 channel=36
					-9, -6, -3, -1, -11, 3, -5, 8, 4,
					-- layer=2 filter=116 channel=37
					-8, -19, -31, 11, -24, -53, 9, 4, -25,
					-- layer=2 filter=116 channel=38
					20, -19, -96, 48, -19, -61, 48, 18, 6,
					-- layer=2 filter=116 channel=39
					47, 37, 2, 19, 23, 62, -72, -23, -22,
					-- layer=2 filter=116 channel=40
					31, -26, -64, 70, 33, -24, 26, -110, -56,
					-- layer=2 filter=116 channel=41
					5, -4, 0, 6, -4, 4, -8, 10, 6,
					-- layer=2 filter=116 channel=42
					10, 11, 24, -9, 16, 3, -31, 3, -7,
					-- layer=2 filter=116 channel=43
					-22, -50, -37, 4, -21, -45, -15, -32, -17,
					-- layer=2 filter=116 channel=44
					-8, 6, 4, 6, -2, -2, -12, -1, 10,
					-- layer=2 filter=116 channel=45
					-42, -49, -23, -22, 23, 7, -38, 23, 7,
					-- layer=2 filter=116 channel=46
					31, 14, -11, 5, 4, -22, -15, -25, -21,
					-- layer=2 filter=116 channel=47
					38, 13, -37, -5, 32, 76, -3, 49, 67,
					-- layer=2 filter=116 channel=48
					-7, -5, -8, -5, 1, 0, -10, 0, -1,
					-- layer=2 filter=116 channel=49
					16, -1, 39, 1, -8, -14, 13, 9, 39,
					-- layer=2 filter=116 channel=50
					5, -6, -3, 6, -7, -4, -30, -11, 9,
					-- layer=2 filter=116 channel=51
					7, -4, -28, 4, -14, -49, 30, 3, 15,
					-- layer=2 filter=116 channel=52
					8, 7, -29, 30, 37, -68, 53, 26, -4,
					-- layer=2 filter=116 channel=53
					13, 52, 20, 44, 5, -15, 41, -22, -4,
					-- layer=2 filter=116 channel=54
					10, 7, -17, -22, 42, 19, -12, 11, 22,
					-- layer=2 filter=116 channel=55
					-3, -3, -9, 2, -4, 0, 7, 12, -7,
					-- layer=2 filter=116 channel=56
					-5, -20, -5, 14, -11, -48, 6, 13, -19,
					-- layer=2 filter=116 channel=57
					-4, 9, -7, -1, -5, 3, -6, 14, 13,
					-- layer=2 filter=116 channel=58
					40, 11, -11, -6, 5, 22, -1, -16, 14,
					-- layer=2 filter=116 channel=59
					15, -9, -48, 16, -10, -52, 42, -20, -12,
					-- layer=2 filter=116 channel=60
					32, 41, -38, -38, -24, -25, 0, -1, -11,
					-- layer=2 filter=116 channel=61
					10, 33, -16, -48, 15, 0, -32, -55, 13,
					-- layer=2 filter=116 channel=62
					6, -3, -4, 19, 7, -37, 34, -3, -24,
					-- layer=2 filter=116 channel=63
					36, 19, -12, -7, 25, 15, -14, 6, 25,
					-- layer=2 filter=116 channel=64
					-14, 5, 3, -37, -8, 22, -70, -71, -47,
					-- layer=2 filter=116 channel=65
					11, 8, -43, -4, 2, -8, -13, -2, 3,
					-- layer=2 filter=116 channel=66
					29, 6, 5, -11, 7, 10, 34, 20, -30,
					-- layer=2 filter=116 channel=67
					7, 25, 19, 13, 8, -26, 11, -27, -20,
					-- layer=2 filter=116 channel=68
					9, -3, 0, -1, 8, 3, -7, 3, -9,
					-- layer=2 filter=116 channel=69
					-13, 12, 10, -18, 3, 13, -64, -31, 0,
					-- layer=2 filter=116 channel=70
					4, -6, -54, 26, 39, 32, -5, -8, 2,
					-- layer=2 filter=116 channel=71
					-14, -11, 14, 42, 0, -61, 44, 15, -28,
					-- layer=2 filter=116 channel=72
					31, -5, -39, -9, -6, 4, -44, 0, -7,
					-- layer=2 filter=116 channel=73
					-10, -18, 17, 3, -44, 36, 45, -25, 59,
					-- layer=2 filter=116 channel=74
					14, 22, -7, 10, 7, -9, -22, -30, -29,
					-- layer=2 filter=116 channel=75
					-18, 38, -2, -12, 13, 16, 9, 3, 22,
					-- layer=2 filter=116 channel=76
					-34, 15, 40, 24, -87, -1, 0, -49, 9,
					-- layer=2 filter=116 channel=77
					-11, -5, 5, 6, -5, 7, 8, -3, 11,
					-- layer=2 filter=116 channel=78
					-12, 2, 20, -23, 13, -5, -9, -10, -10,
					-- layer=2 filter=116 channel=79
					4, -7, 0, 0, 11, -12, 10, 1, -6,
					-- layer=2 filter=116 channel=80
					2, 35, 18, -1, 10, 20, -11, -22, -15,
					-- layer=2 filter=116 channel=81
					3, 3, 16, 3, 1, 2, 1, -10, -13,
					-- layer=2 filter=116 channel=82
					-7, 3, -6, 5, 12, -3, 2, -3, -3,
					-- layer=2 filter=116 channel=83
					-6, 12, 26, -18, 24, 44, -23, -5, -37,
					-- layer=2 filter=116 channel=84
					6, -3, 8, -6, 0, 8, 0, -5, -5,
					-- layer=2 filter=116 channel=85
					4, -10, -6, -2, -9, -8, -8, -10, 4,
					-- layer=2 filter=116 channel=86
					-17, 4, 1, 8, 10, 1, -10, 9, 8,
					-- layer=2 filter=116 channel=87
					-4, 21, 12, 5, -35, -20, 9, -21, -53,
					-- layer=2 filter=116 channel=88
					31, 13, 3, 2, -46, -14, -39, -3, -15,
					-- layer=2 filter=116 channel=89
					7, -1, -28, -27, -35, -45, -6, -8, -1,
					-- layer=2 filter=116 channel=90
					-5, -6, 5, -2, 5, -4, -7, -1, -1,
					-- layer=2 filter=116 channel=91
					39, 18, 2, -8, -6, -5, 13, 2, -4,
					-- layer=2 filter=116 channel=92
					35, 0, -43, -25, -23, -52, 0, 45, -2,
					-- layer=2 filter=116 channel=93
					-7, 11, -11, -3, 34, -41, -56, 34, -21,
					-- layer=2 filter=116 channel=94
					12, 21, 21, 7, 42, -23, -1, 3, 8,
					-- layer=2 filter=116 channel=95
					2, -6, 13, -4, 9, 4, 10, -2, 15,
					-- layer=2 filter=116 channel=96
					19, 30, 25, -14, 8, -8, 8, 36, -5,
					-- layer=2 filter=116 channel=97
					-36, -1, 26, 0, -12, 56, -31, -34, 27,
					-- layer=2 filter=116 channel=98
					32, -17, -38, -21, 40, 70, -23, 3, 43,
					-- layer=2 filter=116 channel=99
					5, 27, -19, 10, 0, -51, 61, -21, -6,
					-- layer=2 filter=116 channel=100
					25, -5, 2, 25, 0, 8, -4, -15, -52,
					-- layer=2 filter=116 channel=101
					22, -15, 11, 22, -12, -36, 34, -1, -2,
					-- layer=2 filter=116 channel=102
					-6, -4, 21, 32, 20, -5, 11, 13, 1,
					-- layer=2 filter=116 channel=103
					28, -4, -39, -1, -17, -49, 41, 34, 70,
					-- layer=2 filter=116 channel=104
					36, 30, 83, 3, -23, -27, -3, 24, 15,
					-- layer=2 filter=116 channel=105
					-14, -22, -33, 43, -36, -28, 46, -23, -1,
					-- layer=2 filter=116 channel=106
					7, 3, 21, -9, 12, -4, -4, -7, 8,
					-- layer=2 filter=116 channel=107
					-4, -26, -16, 14, 5, -33, 71, 39, 64,
					-- layer=2 filter=116 channel=108
					-9, 23, -26, 26, -5, -70, 46, 45, 16,
					-- layer=2 filter=116 channel=109
					15, -14, -5, 6, -14, 6, 1, 7, 2,
					-- layer=2 filter=116 channel=110
					-62, 20, 10, -71, -28, -10, -75, -22, 5,
					-- layer=2 filter=116 channel=111
					5, 10, -2, 2, -2, 6, -1, 2, 0,
					-- layer=2 filter=116 channel=112
					30, 10, -8, -15, -11, -22, 15, -21, 13,
					-- layer=2 filter=116 channel=113
					9, 29, -12, -8, 22, -11, -9, -37, -27,
					-- layer=2 filter=116 channel=114
					4, -6, -13, 12, 1, 8, 0, 9, 6,
					-- layer=2 filter=116 channel=115
					3, 8, -7, 8, -2, 10, -5, 2, 8,
					-- layer=2 filter=116 channel=116
					19, 26, -17, 16, 1, -23, 24, -59, -50,
					-- layer=2 filter=116 channel=117
					42, -7, -42, 0, 44, 4, 13, 22, 12,
					-- layer=2 filter=116 channel=118
					-5, -15, 13, -6, -12, 6, 3, -17, -10,
					-- layer=2 filter=116 channel=119
					-20, -14, 0, -7, 45, 47, 19, 0, 37,
					-- layer=2 filter=116 channel=120
					2, 0, 8, 5, -1, -3, -6, 8, 7,
					-- layer=2 filter=116 channel=121
					-1, 5, -7, -4, 2, -1, 6, -1, -6,
					-- layer=2 filter=116 channel=122
					-8, -2, -11, -14, 13, -10, 4, 4, -9,
					-- layer=2 filter=116 channel=123
					21, -10, -35, 11, 34, 54, -36, 2, 20,
					-- layer=2 filter=116 channel=124
					-30, -3, -65, -2, -28, 6, -36, 7, -61,
					-- layer=2 filter=116 channel=125
					4, 2, 11, 0, -4, -1, 8, -2, 8,
					-- layer=2 filter=116 channel=126
					-35, 37, 32, -54, 7, -19, 26, -43, -13,
					-- layer=2 filter=116 channel=127
					18, 19, -18, -4, 7, -22, -13, 56, 1,
					-- layer=2 filter=117 channel=0
					13, 35, 15, 14, 18, 29, -30, -4, -45,
					-- layer=2 filter=117 channel=1
					26, 5, -30, -11, -18, -15, 35, 15, 36,
					-- layer=2 filter=117 channel=2
					9, 0, 3, 11, 3, 9, 0, 9, -1,
					-- layer=2 filter=117 channel=3
					5, 15, 12, -31, -34, 3, 14, 11, 18,
					-- layer=2 filter=117 channel=4
					0, 15, -7, -39, -24, -13, -46, -26, -32,
					-- layer=2 filter=117 channel=5
					14, 26, 17, 9, 17, 30, -8, 37, -35,
					-- layer=2 filter=117 channel=6
					27, 57, 33, 9, 37, 21, -30, 41, 48,
					-- layer=2 filter=117 channel=7
					0, -61, -8, 33, -4, -40, 0, -3, -2,
					-- layer=2 filter=117 channel=8
					5, -5, -9, -2, 6, -8, -7, -3, 9,
					-- layer=2 filter=117 channel=9
					27, 15, 23, -12, -11, 26, -6, 0, 7,
					-- layer=2 filter=117 channel=10
					24, 32, 30, -22, 32, 6, -4, -15, -33,
					-- layer=2 filter=117 channel=11
					-11, -17, -23, -7, -11, -12, -9, -18, 8,
					-- layer=2 filter=117 channel=12
					20, -4, -13, -26, -11, 20, 48, 50, 53,
					-- layer=2 filter=117 channel=13
					2, 7, 2, -2, -9, 2, 8, -5, -9,
					-- layer=2 filter=117 channel=14
					16, -7, -13, 6, -13, -1, 25, 25, 42,
					-- layer=2 filter=117 channel=15
					-40, -42, -9, -30, 36, -13, -27, 35, 64,
					-- layer=2 filter=117 channel=16
					22, -6, -26, -32, -44, -60, -11, 14, -9,
					-- layer=2 filter=117 channel=17
					-9, -7, -4, 5, -6, 6, 9, 3, -9,
					-- layer=2 filter=117 channel=18
					13, 30, 31, 39, -45, -15, 28, -11, -27,
					-- layer=2 filter=117 channel=19
					-48, -52, -48, -14, -29, -34, 7, -19, 1,
					-- layer=2 filter=117 channel=20
					-7, -7, 8, 2, -8, -7, 2, 3, -5,
					-- layer=2 filter=117 channel=21
					15, 6, 15, -3, 0, 4, 13, 7, -2,
					-- layer=2 filter=117 channel=22
					-7, 0, 9, -1, 0, 4, 11, 0, 2,
					-- layer=2 filter=117 channel=23
					0, 7, -17, -22, -25, -41, -15, -19, -7,
					-- layer=2 filter=117 channel=24
					0, 0, 15, 0, 5, -32, 13, 25, -2,
					-- layer=2 filter=117 channel=25
					-53, -68, 0, -22, -10, -21, 15, 19, 6,
					-- layer=2 filter=117 channel=26
					5, 1, -5, -9, 9, -7, 9, 2, 5,
					-- layer=2 filter=117 channel=27
					23, 17, -10, 14, 18, 5, 4, -19, -28,
					-- layer=2 filter=117 channel=28
					14, -19, -5, -18, 0, -7, 29, -62, -47,
					-- layer=2 filter=117 channel=29
					10, 2, -10, -6, 0, -6, -2, -9, -2,
					-- layer=2 filter=117 channel=30
					33, -9, 12, 7, 11, -12, -30, 12, -4,
					-- layer=2 filter=117 channel=31
					-7, -66, 47, -6, -26, 36, 16, -7, -72,
					-- layer=2 filter=117 channel=32
					7, 3, -2, 0, -8, -3, -8, 3, 6,
					-- layer=2 filter=117 channel=33
					-10, 46, -4, -43, -1, 21, 6, -5, 16,
					-- layer=2 filter=117 channel=34
					-5, -1, 7, 46, -24, 5, 15, 2, -27,
					-- layer=2 filter=117 channel=35
					-15, -13, -39, -20, -19, -10, 0, -58, 9,
					-- layer=2 filter=117 channel=36
					1, 12, 11, -2, 3, -1, 12, 12, 9,
					-- layer=2 filter=117 channel=37
					-6, 7, -23, -10, 9, 8, 5, -12, -2,
					-- layer=2 filter=117 channel=38
					29, 17, 0, 3, 0, -7, -6, 13, -29,
					-- layer=2 filter=117 channel=39
					-3, -16, -22, -6, 6, -58, -33, 36, -14,
					-- layer=2 filter=117 channel=40
					-37, -39, -60, -32, 7, 0, -57, 48, -14,
					-- layer=2 filter=117 channel=41
					-7, -4, -5, 5, -9, -3, 2, -7, -2,
					-- layer=2 filter=117 channel=42
					5, -4, -8, -12, 4, -4, 25, 23, 39,
					-- layer=2 filter=117 channel=43
					5, 34, 0, -9, 30, 19, -5, -46, 2,
					-- layer=2 filter=117 channel=44
					10, 2, 4, 7, 2, 6, -3, -4, 3,
					-- layer=2 filter=117 channel=45
					46, 23, 20, 15, 14, 37, -49, -53, -85,
					-- layer=2 filter=117 channel=46
					26, 10, 7, -29, 15, 11, -49, 1, -51,
					-- layer=2 filter=117 channel=47
					-5, -14, 4, -42, -11, -6, -21, -17, -14,
					-- layer=2 filter=117 channel=48
					5, 7, 5, -7, -7, 6, 0, -2, -7,
					-- layer=2 filter=117 channel=49
					38, 53, 34, 11, 6, -5, 21, 6, 27,
					-- layer=2 filter=117 channel=50
					-11, -4, -17, 12, -16, -23, -11, -20, -18,
					-- layer=2 filter=117 channel=51
					0, 7, -5, -18, -15, 2, -23, -14, -19,
					-- layer=2 filter=117 channel=52
					20, -17, -17, 7, -19, -21, 0, -38, 2,
					-- layer=2 filter=117 channel=53
					39, -13, 7, 32, -43, -52, -25, -22, -6,
					-- layer=2 filter=117 channel=54
					12, 1, -26, 5, -24, -2, 13, -8, -9,
					-- layer=2 filter=117 channel=55
					0, 1, -8, -12, 0, -6, -9, -2, -5,
					-- layer=2 filter=117 channel=56
					-12, -3, 2, -11, -5, -28, -8, -2, 6,
					-- layer=2 filter=117 channel=57
					-3, 8, -5, -4, 3, 9, -4, -10, -6,
					-- layer=2 filter=117 channel=58
					12, 10, 1, 4, 0, 26, 35, 38, 44,
					-- layer=2 filter=117 channel=59
					20, -22, -7, 5, -29, -44, 37, -2, 10,
					-- layer=2 filter=117 channel=60
					-22, 10, -22, 15, 13, -2, 14, 46, -11,
					-- layer=2 filter=117 channel=61
					-5, 1, -14, 4, -15, -70, 8, 2, -61,
					-- layer=2 filter=117 channel=62
					7, 21, 33, 19, -18, 2, -36, -29, 44,
					-- layer=2 filter=117 channel=63
					10, 3, -12, -1, -5, -43, -8, -5, -13,
					-- layer=2 filter=117 channel=64
					9, -10, -4, 10, -4, -16, 0, 7, 2,
					-- layer=2 filter=117 channel=65
					-3, -4, -11, -12, -10, -30, -37, -1, -37,
					-- layer=2 filter=117 channel=66
					1, 48, 10, 5, 15, 19, 44, 37, 13,
					-- layer=2 filter=117 channel=67
					18, 29, 5, -12, 31, -19, -56, 4, -7,
					-- layer=2 filter=117 channel=68
					2, 9, -5, 3, 6, -5, -8, -1, 5,
					-- layer=2 filter=117 channel=69
					0, -24, -36, -1, 14, -20, -13, 6, 10,
					-- layer=2 filter=117 channel=70
					-18, 0, -8, -20, -23, 20, -44, -71, -30,
					-- layer=2 filter=117 channel=71
					0, 21, -6, 22, 19, 12, -25, -53, -29,
					-- layer=2 filter=117 channel=72
					-17, -22, -14, 9, -35, -12, 54, 22, 33,
					-- layer=2 filter=117 channel=73
					21, -41, -22, -29, -22, -51, -31, -29, -50,
					-- layer=2 filter=117 channel=74
					6, -1, -25, -24, -2, -2, -30, 1, 3,
					-- layer=2 filter=117 channel=75
					-5, -9, 21, -6, 1, 14, 0, 62, 59,
					-- layer=2 filter=117 channel=76
					-42, -49, 7, 22, 4, -55, -80, -47, 20,
					-- layer=2 filter=117 channel=77
					-6, -3, -6, 0, 5, 9, -12, 1, -9,
					-- layer=2 filter=117 channel=78
					-32, -18, -40, 6, -9, -5, -20, -34, 18,
					-- layer=2 filter=117 channel=79
					-8, 5, 4, -4, -4, 7, 5, -3, -5,
					-- layer=2 filter=117 channel=80
					-1, -10, -6, -33, 9, -4, -25, 31, -5,
					-- layer=2 filter=117 channel=81
					-12, -6, -5, -9, -7, -14, -13, 0, -4,
					-- layer=2 filter=117 channel=82
					-12, 6, 0, 0, -6, -1, -6, 10, 0,
					-- layer=2 filter=117 channel=83
					-1, 0, -21, -25, -19, 0, -30, -43, -12,
					-- layer=2 filter=117 channel=84
					1, 3, -8, 3, 10, -3, 5, 6, 8,
					-- layer=2 filter=117 channel=85
					7, 11, 0, -5, 8, -1, 12, -8, -4,
					-- layer=2 filter=117 channel=86
					12, -14, 0, 14, 9, 9, 0, -1, 8,
					-- layer=2 filter=117 channel=87
					-3, 30, 57, -39, -8, -47, 11, -4, 4,
					-- layer=2 filter=117 channel=88
					25, -4, -9, -6, 4, -11, -23, 20, 18,
					-- layer=2 filter=117 channel=89
					-15, -49, -22, -5, -8, 4, 36, 21, 58,
					-- layer=2 filter=117 channel=90
					9, 10, 0, 8, -2, -8, 2, -2, 7,
					-- layer=2 filter=117 channel=91
					-18, -9, -28, -17, 5, 20, 58, 46, 48,
					-- layer=2 filter=117 channel=92
					26, -16, -22, -14, -10, 5, 57, 35, 42,
					-- layer=2 filter=117 channel=93
					10, -14, 30, 61, 63, 99, -25, 48, 30,
					-- layer=2 filter=117 channel=94
					3, -16, -7, -9, -50, -63, -22, -33, -41,
					-- layer=2 filter=117 channel=95
					19, 6, 5, 8, 22, 8, 11, 8, 15,
					-- layer=2 filter=117 channel=96
					-5, 91, 35, 41, 49, 34, 0, 16, 2,
					-- layer=2 filter=117 channel=97
					-7, 0, 3, -6, 0, 12, -11, -10, -6,
					-- layer=2 filter=117 channel=98
					-23, -36, -28, -42, -12, -26, -22, -43, -17,
					-- layer=2 filter=117 channel=99
					-58, -40, -38, -35, -31, -54, -14, -27, 0,
					-- layer=2 filter=117 channel=100
					15, 7, -4, 1, 2, 10, 0, -4, -16,
					-- layer=2 filter=117 channel=101
					-28, -17, -4, -38, -1, 12, -23, -1, -8,
					-- layer=2 filter=117 channel=102
					-4, 29, 37, 26, -3, 32, -2, -26, 8,
					-- layer=2 filter=117 channel=103
					30, 22, 15, -2, 66, 60, 27, -28, -13,
					-- layer=2 filter=117 channel=104
					19, 21, -11, 11, -48, -21, -26, -24, 22,
					-- layer=2 filter=117 channel=105
					-68, -35, -12, -64, -44, -34, 15, -18, 26,
					-- layer=2 filter=117 channel=106
					-43, 1, 13, -22, 16, 28, 12, 17, 19,
					-- layer=2 filter=117 channel=107
					-23, -63, 2, 44, 18, 16, 1, -17, 68,
					-- layer=2 filter=117 channel=108
					28, 36, 31, 40, 17, 3, -27, -9, 4,
					-- layer=2 filter=117 channel=109
					-10, -2, 10, -8, -13, 0, -10, -4, 14,
					-- layer=2 filter=117 channel=110
					11, -1, -10, 14, 24, 20, 23, 33, 50,
					-- layer=2 filter=117 channel=111
					6, 3, 6, -4, 4, 0, -4, 7, 5,
					-- layer=2 filter=117 channel=112
					-6, -6, 5, -21, 57, -6, -22, 15, -53,
					-- layer=2 filter=117 channel=113
					16, 14, -9, -9, -22, -18, -1, -2, -15,
					-- layer=2 filter=117 channel=114
					21, -6, -8, -8, -4, 0, 3, 4, -5,
					-- layer=2 filter=117 channel=115
					-2, -6, -4, -8, 0, 4, 0, 10, 1,
					-- layer=2 filter=117 channel=116
					-11, 15, 12, -21, 32, -30, -5, 3, -1,
					-- layer=2 filter=117 channel=117
					-19, -7, -36, 19, 13, 18, 12, 4, 18,
					-- layer=2 filter=117 channel=118
					39, 70, 33, -9, 23, 29, 8, -31, -3,
					-- layer=2 filter=117 channel=119
					13, 11, 37, 20, -27, -16, 18, -53, -55,
					-- layer=2 filter=117 channel=120
					7, -9, -10, -4, -4, 6, -4, 8, 7,
					-- layer=2 filter=117 channel=121
					-3, -4, -2, 0, 1, -8, -6, -5, -4,
					-- layer=2 filter=117 channel=122
					5, -7, 9, 13, 1, 7, -12, 3, 5,
					-- layer=2 filter=117 channel=123
					-13, -60, -28, -14, -36, -49, -11, 7, 7,
					-- layer=2 filter=117 channel=124
					-1, 0, 18, 21, 13, -15, 0, 21, 99,
					-- layer=2 filter=117 channel=125
					-3, 1, -8, -6, -4, 6, -2, -5, 10,
					-- layer=2 filter=117 channel=126
					-4, 48, 0, 21, 66, -72, 4, 11, 11,
					-- layer=2 filter=117 channel=127
					-7, 8, -12, 6, -18, -19, 16, -23, 7,
					-- layer=2 filter=118 channel=0
					1, 14, 10, 2, -19, -24, -21, -33, 0,
					-- layer=2 filter=118 channel=1
					-14, 8, 1, -11, 24, 20, 23, 4, 14,
					-- layer=2 filter=118 channel=2
					8, -2, 3, -5, -2, 9, -7, 0, 7,
					-- layer=2 filter=118 channel=3
					-10, 1, -18, -41, -3, -39, -41, -33, -9,
					-- layer=2 filter=118 channel=4
					2, 10, 28, 4, 12, 22, -21, -33, 10,
					-- layer=2 filter=118 channel=5
					7, 8, 17, -1, -5, -12, 11, 1, -16,
					-- layer=2 filter=118 channel=6
					-2, -13, 0, 31, 45, -49, 49, 56, 67,
					-- layer=2 filter=118 channel=7
					24, 11, 16, -58, -39, -13, 0, -27, 3,
					-- layer=2 filter=118 channel=8
					-2, 4, -3, 9, -3, -7, -9, -7, 0,
					-- layer=2 filter=118 channel=9
					-8, 13, 0, -38, 27, -2, -73, -16, -26,
					-- layer=2 filter=118 channel=10
					2, -4, 12, -46, -14, -24, -27, -57, -42,
					-- layer=2 filter=118 channel=11
					-1, -5, -5, -3, -8, 5, 4, 1, 9,
					-- layer=2 filter=118 channel=12
					-8, 18, 31, -24, -2, -5, 23, 1, 8,
					-- layer=2 filter=118 channel=13
					-2, 8, -5, -2, 7, -2, 0, -2, -8,
					-- layer=2 filter=118 channel=14
					-8, 0, 1, 12, 11, 18, 17, 20, 15,
					-- layer=2 filter=118 channel=15
					16, 46, -27, 19, 26, 20, -22, 3, 22,
					-- layer=2 filter=118 channel=16
					44, 44, 29, 34, 35, 14, 11, -15, -21,
					-- layer=2 filter=118 channel=17
					-5, 2, -9, 7, 2, -7, 10, 0, -2,
					-- layer=2 filter=118 channel=18
					-3, 15, 14, 3, 19, 38, -8, 0, -8,
					-- layer=2 filter=118 channel=19
					-26, -39, -24, 6, 42, -2, 24, 15, -1,
					-- layer=2 filter=118 channel=20
					6, -4, 1, -1, -8, -6, 7, 5, 3,
					-- layer=2 filter=118 channel=21
					-4, -14, 2, -16, -14, 0, -13, -5, 7,
					-- layer=2 filter=118 channel=22
					-2, 11, 2, 10, -9, 8, 2, -5, -5,
					-- layer=2 filter=118 channel=23
					5, 19, 10, 5, 5, 26, 22, 13, 14,
					-- layer=2 filter=118 channel=24
					21, 5, -10, -1, 0, -3, -3, -30, -8,
					-- layer=2 filter=118 channel=25
					43, 12, 13, 43, 4, -20, 9, -1, -5,
					-- layer=2 filter=118 channel=26
					-8, 2, 0, 0, 0, -9, -13, -6, 5,
					-- layer=2 filter=118 channel=27
					-3, -8, -9, 27, 24, 5, 17, 17, -30,
					-- layer=2 filter=118 channel=28
					-17, 18, 20, -31, -8, -47, 3, -5, 11,
					-- layer=2 filter=118 channel=29
					0, -5, 0, -6, -8, 0, 0, -7, 6,
					-- layer=2 filter=118 channel=30
					-12, 0, 13, 4, -2, -5, 8, -27, -11,
					-- layer=2 filter=118 channel=31
					-15, 27, 31, -127, 17, -27, -69, -19, -105,
					-- layer=2 filter=118 channel=32
					3, 1, -3, -3, -1, -7, -1, -11, -3,
					-- layer=2 filter=118 channel=33
					-1, 16, -31, 0, -7, -7, 1, -7, 25,
					-- layer=2 filter=118 channel=34
					26, -26, -20, -3, -11, 6, -4, 33, -29,
					-- layer=2 filter=118 channel=35
					-8, 10, 1, -28, -53, -35, 14, 21, -2,
					-- layer=2 filter=118 channel=36
					-8, -2, 13, -3, 0, -2, 0, 0, -15,
					-- layer=2 filter=118 channel=37
					3, 12, -2, 14, 2, 8, 10, 1, 2,
					-- layer=2 filter=118 channel=38
					-24, -24, -6, 21, 1, 6, 2, 8, -20,
					-- layer=2 filter=118 channel=39
					18, 9, -9, -4, 16, -16, -9, -41, -23,
					-- layer=2 filter=118 channel=40
					-22, -27, 6, -17, -17, 1, -51, 17, -21,
					-- layer=2 filter=118 channel=41
					7, 0, 11, -8, -13, 0, 3, -2, 0,
					-- layer=2 filter=118 channel=42
					-4, 30, 9, 16, -1, 8, 26, 30, -11,
					-- layer=2 filter=118 channel=43
					-15, 2, -39, -49, -16, -53, -44, -39, -39,
					-- layer=2 filter=118 channel=44
					7, -6, 8, 3, 10, 0, -7, -8, 6,
					-- layer=2 filter=118 channel=45
					46, 33, -12, 32, 18, -32, 0, -3, -18,
					-- layer=2 filter=118 channel=46
					-12, 0, -3, -29, -9, 0, -14, -42, -43,
					-- layer=2 filter=118 channel=47
					50, 67, 41, -2, 18, -65, 0, 3, 30,
					-- layer=2 filter=118 channel=48
					9, 0, 6, 8, -7, 3, -6, 0, 7,
					-- layer=2 filter=118 channel=49
					28, 13, 14, 4, 29, 27, -3, -23, -20,
					-- layer=2 filter=118 channel=50
					23, 1, -2, -9, -13, 11, 15, 9, 13,
					-- layer=2 filter=118 channel=51
					-1, -11, 8, 6, -20, -4, -21, 0, 10,
					-- layer=2 filter=118 channel=52
					-38, -38, -34, 2, 37, -14, 7, 19, 24,
					-- layer=2 filter=118 channel=53
					16, -62, -88, -7, -2, -31, 7, 30, 4,
					-- layer=2 filter=118 channel=54
					-3, -8, 8, 9, -1, -15, 42, 4, 39,
					-- layer=2 filter=118 channel=55
					4, -1, -4, 8, -10, -7, 6, -11, -4,
					-- layer=2 filter=118 channel=56
					1, 11, 14, 0, 0, 1, 0, 17, 0,
					-- layer=2 filter=118 channel=57
					-13, 10, -5, 0, 4, 5, 0, -2, 3,
					-- layer=2 filter=118 channel=58
					6, 24, 36, -4, -6, -19, 15, 7, 3,
					-- layer=2 filter=118 channel=59
					-8, -32, -41, 31, -10, 9, 17, 22, -5,
					-- layer=2 filter=118 channel=60
					-11, -53, -27, -4, 1, -16, 22, 36, 10,
					-- layer=2 filter=118 channel=61
					-48, -90, -15, 3, -14, -8, 6, -15, 37,
					-- layer=2 filter=118 channel=62
					13, -25, -15, 7, 27, -7, -9, -5, -17,
					-- layer=2 filter=118 channel=63
					9, -4, 0, -24, 31, -1, -2, 10, 18,
					-- layer=2 filter=118 channel=64
					8, 9, 1, 14, 13, 1, 8, -15, -17,
					-- layer=2 filter=118 channel=65
					-25, -78, -11, 6, -24, -17, 34, 12, 36,
					-- layer=2 filter=118 channel=66
					-7, 5, 26, 32, -4, 15, 35, 24, -41,
					-- layer=2 filter=118 channel=67
					-10, 5, -5, -47, 37, 7, -17, -39, -18,
					-- layer=2 filter=118 channel=68
					5, -4, 3, -10, 7, 8, -3, -11, 11,
					-- layer=2 filter=118 channel=69
					8, 8, 25, 11, 17, -3, 0, 16, -3,
					-- layer=2 filter=118 channel=70
					19, 37, 39, -8, -23, -45, -2, -9, -26,
					-- layer=2 filter=118 channel=71
					-13, -33, -19, 26, 26, 27, 31, 22, 17,
					-- layer=2 filter=118 channel=72
					-26, -21, -16, -15, -8, 17, 16, 1, -1,
					-- layer=2 filter=118 channel=73
					21, -19, -56, -46, 5, 4, -36, -20, -62,
					-- layer=2 filter=118 channel=74
					-26, -24, -4, -6, 13, -3, -50, -14, -24,
					-- layer=2 filter=118 channel=75
					-16, -41, -8, -12, 25, -53, 69, 49, -10,
					-- layer=2 filter=118 channel=76
					44, -31, -39, -89, -55, -34, -34, -1, 43,
					-- layer=2 filter=118 channel=77
					8, -4, 6, 4, 0, 6, 0, 1, -7,
					-- layer=2 filter=118 channel=78
					-7, 0, -12, -1, 18, -22, 14, -8, 0,
					-- layer=2 filter=118 channel=79
					8, 0, 2, 5, 0, -1, -5, -6, -11,
					-- layer=2 filter=118 channel=80
					-6, 6, 10, -35, -9, -19, -25, -8, -36,
					-- layer=2 filter=118 channel=81
					-8, -9, 3, -16, -5, -8, -10, -5, -11,
					-- layer=2 filter=118 channel=82
					-3, -5, 6, 7, 4, -8, -6, 0, -2,
					-- layer=2 filter=118 channel=83
					-1, 9, 38, 27, -8, 6, 36, -9, -24,
					-- layer=2 filter=118 channel=84
					-7, 9, 2, 8, 1, -12, 3, 5, 0,
					-- layer=2 filter=118 channel=85
					0, -14, 0, 2, 9, -5, 0, 9, -20,
					-- layer=2 filter=118 channel=86
					-13, 18, 0, -7, 12, 7, -6, 6, 12,
					-- layer=2 filter=118 channel=87
					29, -30, -22, 7, -36, -22, 27, 0, 22,
					-- layer=2 filter=118 channel=88
					3, 0, -2, 7, 8, 13, -23, -14, -7,
					-- layer=2 filter=118 channel=89
					-22, -22, -16, -19, -4, 4, 34, 17, 4,
					-- layer=2 filter=118 channel=90
					1, -1, 7, -2, 0, 8, -5, 0, 9,
					-- layer=2 filter=118 channel=91
					-31, -6, -6, 8, -13, -18, 35, 20, -37,
					-- layer=2 filter=118 channel=92
					5, 9, 22, -20, 7, 24, 16, -7, 5,
					-- layer=2 filter=118 channel=93
					10, -24, -27, 9, 3, -20, 2, 40, 10,
					-- layer=2 filter=118 channel=94
					-25, -68, -15, 8, 34, -18, 38, 46, 45,
					-- layer=2 filter=118 channel=95
					9, -4, 2, 6, -14, -9, -2, 1, -3,
					-- layer=2 filter=118 channel=96
					-7, -51, -14, 41, 5, 35, 56, 46, 23,
					-- layer=2 filter=118 channel=97
					-7, 32, -15, -22, -2, -15, -43, -15, -28,
					-- layer=2 filter=118 channel=98
					6, 30, 19, -48, -20, -49, -16, -11, 1,
					-- layer=2 filter=118 channel=99
					-63, -79, -38, 0, 41, 9, 26, 49, 75,
					-- layer=2 filter=118 channel=100
					-16, -13, 0, 6, -31, -14, 1, 35, -97,
					-- layer=2 filter=118 channel=101
					-10, -18, -32, 24, 1, 37, 22, 10, 36,
					-- layer=2 filter=118 channel=102
					-13, -25, 9, 31, -3, 28, 65, 53, -4,
					-- layer=2 filter=118 channel=103
					-4, -27, -19, -49, -53, -13, -39, -47, -13,
					-- layer=2 filter=118 channel=104
					30, -40, -13, 9, 35, 43, 7, -5, 20,
					-- layer=2 filter=118 channel=105
					-2, -33, -3, -49, -8, 25, 1, -11, 13,
					-- layer=2 filter=118 channel=106
					21, 24, 22, 41, 13, 14, 20, 11, -2,
					-- layer=2 filter=118 channel=107
					-26, 41, 13, -38, 12, 21, -18, -50, -30,
					-- layer=2 filter=118 channel=108
					-11, -16, -25, 7, 19, 17, 31, 9, -24,
					-- layer=2 filter=118 channel=109
					3, 5, -2, -5, -13, -6, -7, 7, 1,
					-- layer=2 filter=118 channel=110
					25, 16, 1, 31, 52, 8, 49, 15, 8,
					-- layer=2 filter=118 channel=111
					9, -10, -8, -10, 1, 4, 0, 1, -6,
					-- layer=2 filter=118 channel=112
					-24, -11, 9, -34, -5, 1, -15, -28, 2,
					-- layer=2 filter=118 channel=113
					0, -10, 23, 1, 29, 15, -5, -5, -5,
					-- layer=2 filter=118 channel=114
					-9, 12, 0, -3, -2, -12, -2, -12, -10,
					-- layer=2 filter=118 channel=115
					12, -9, 4, -5, 2, 6, -4, -12, -7,
					-- layer=2 filter=118 channel=116
					8, 0, 17, 38, -2, 6, 19, 37, -11,
					-- layer=2 filter=118 channel=117
					-57, -45, -34, -70, -43, 9, 26, 30, 43,
					-- layer=2 filter=118 channel=118
					20, 21, -4, -33, 18, -53, -57, -30, -8,
					-- layer=2 filter=118 channel=119
					16, 16, 16, 29, 22, 6, -5, 12, -4,
					-- layer=2 filter=118 channel=120
					3, -6, 3, -9, 0, 0, 9, 1, -2,
					-- layer=2 filter=118 channel=121
					-8, 6, 3, 7, -1, 8, -7, 8, 3,
					-- layer=2 filter=118 channel=122
					0, -8, 1, 9, -13, -12, 12, 4, 9,
					-- layer=2 filter=118 channel=123
					-2, -5, -26, -58, 10, -43, 11, 21, 14,
					-- layer=2 filter=118 channel=124
					2, -2, -26, -51, 0, -18, -3, -9, 27,
					-- layer=2 filter=118 channel=125
					-7, 0, -11, 1, -3, 2, 7, -1, -14,
					-- layer=2 filter=118 channel=126
					47, -35, -68, -36, 0, 4, 27, 75, 20,
					-- layer=2 filter=118 channel=127
					-21, -24, 0, -2, 4, 0, 12, 37, -21,
					-- layer=2 filter=119 channel=0
					30, 16, 34, 19, -17, -2, 1, -4, -20,
					-- layer=2 filter=119 channel=1
					28, 37, 10, 15, 26, 18, -16, 14, 25,
					-- layer=2 filter=119 channel=2
					0, 3, 8, -8, -5, -9, 3, -11, 5,
					-- layer=2 filter=119 channel=3
					-37, -22, -3, -4, 1, 12, 40, 17, 31,
					-- layer=2 filter=119 channel=4
					-6, 27, 4, -14, -30, -12, -11, -78, -3,
					-- layer=2 filter=119 channel=5
					44, 20, 35, 0, -2, -4, 19, -43, -13,
					-- layer=2 filter=119 channel=6
					-30, 6, 8, -39, -69, -59, -59, -70, -28,
					-- layer=2 filter=119 channel=7
					17, 6, -2, 52, 28, 38, 49, 64, 34,
					-- layer=2 filter=119 channel=8
					7, 10, -11, 7, 2, -1, 0, 10, 10,
					-- layer=2 filter=119 channel=9
					7, 27, -2, -8, 32, 5, 27, 27, 20,
					-- layer=2 filter=119 channel=10
					-1, -6, 20, -13, -26, -7, 42, 11, 10,
					-- layer=2 filter=119 channel=11
					25, 40, 16, -24, 1, -9, -28, -15, -10,
					-- layer=2 filter=119 channel=12
					20, 28, 0, 47, 52, 15, 4, 19, 52,
					-- layer=2 filter=119 channel=13
					3, -10, 1, -12, -2, 4, 8, -10, -11,
					-- layer=2 filter=119 channel=14
					18, 22, -9, 40, 27, 35, -12, 25, 25,
					-- layer=2 filter=119 channel=15
					71, -9, 9, -44, -5, -5, -22, 15, -1,
					-- layer=2 filter=119 channel=16
					-9, 15, 3, -11, -2, -29, -6, -40, -9,
					-- layer=2 filter=119 channel=17
					-8, -9, 2, -7, -3, -10, 4, -2, 10,
					-- layer=2 filter=119 channel=18
					-4, 1, -27, 19, -5, -30, -15, -31, -15,
					-- layer=2 filter=119 channel=19
					31, 54, 39, -16, -1, -21, -12, -12, 25,
					-- layer=2 filter=119 channel=20
					-1, -11, -11, 2, -6, -4, -7, 9, 9,
					-- layer=2 filter=119 channel=21
					11, 0, -15, 10, 4, 4, 18, 3, 2,
					-- layer=2 filter=119 channel=22
					9, -6, 2, -4, -7, -9, 7, -9, 3,
					-- layer=2 filter=119 channel=23
					1, 17, -8, 0, -15, 7, 24, -12, 25,
					-- layer=2 filter=119 channel=24
					-48, -6, 4, -36, 19, 20, 0, 22, 37,
					-- layer=2 filter=119 channel=25
					-52, -11, -8, -14, 17, 5, -37, -4, -12,
					-- layer=2 filter=119 channel=26
					7, 0, 4, 0, 8, 2, 0, 3, 0,
					-- layer=2 filter=119 channel=27
					15, 43, 40, -22, -16, -14, -23, -46, -22,
					-- layer=2 filter=119 channel=28
					-29, -2, -4, 39, 29, 33, 15, -2, -20,
					-- layer=2 filter=119 channel=29
					0, 5, 8, -9, 2, -6, 5, -5, -5,
					-- layer=2 filter=119 channel=30
					-1, 1, 5, -7, -13, -32, -37, -17, -19,
					-- layer=2 filter=119 channel=31
					32, -11, -4, 14, -18, 7, 0, -39, -7,
					-- layer=2 filter=119 channel=32
					2, 1, 5, 0, -3, -5, 4, 0, 9,
					-- layer=2 filter=119 channel=33
					4, 33, 6, -16, -57, 12, -21, -3, -2,
					-- layer=2 filter=119 channel=34
					28, -3, 46, -47, -30, -95, -108, -78, -90,
					-- layer=2 filter=119 channel=35
					26, 30, 34, 4, -3, 0, -42, 1, -9,
					-- layer=2 filter=119 channel=36
					-3, -5, 0, 1, -9, 10, 15, 1, -1,
					-- layer=2 filter=119 channel=37
					32, 42, 11, -29, 6, -18, -3, 0, -2,
					-- layer=2 filter=119 channel=38
					19, -8, 19, -36, -18, -18, -70, -83, -48,
					-- layer=2 filter=119 channel=39
					-23, -2, 0, -14, 1, 17, -4, 9, 10,
					-- layer=2 filter=119 channel=40
					67, 7, -10, 9, 1, -13, -67, -22, -19,
					-- layer=2 filter=119 channel=41
					-3, 7, 6, -9, 4, 0, 2, 2, -6,
					-- layer=2 filter=119 channel=42
					-18, -6, -31, 24, 15, 11, 18, -4, 35,
					-- layer=2 filter=119 channel=43
					6, 27, -34, -13, -41, -9, 0, 14, 18,
					-- layer=2 filter=119 channel=44
					-8, 4, 7, -11, -10, 0, 6, 5, 2,
					-- layer=2 filter=119 channel=45
					-11, -21, -12, -26, 0, 9, -16, -29, 3,
					-- layer=2 filter=119 channel=46
					-25, -25, 6, -57, -27, -33, -42, -57, -24,
					-- layer=2 filter=119 channel=47
					-10, 15, 11, 3, 26, 27, -9, -26, -40,
					-- layer=2 filter=119 channel=48
					8, -8, 4, 8, 4, 2, 9, 8, 7,
					-- layer=2 filter=119 channel=49
					16, 33, -27, 37, -4, -4, 14, 35, 47,
					-- layer=2 filter=119 channel=50
					-19, 0, 3, 0, 5, -3, -9, -10, 3,
					-- layer=2 filter=119 channel=51
					18, 36, 18, -3, -5, -6, -10, 0, -19,
					-- layer=2 filter=119 channel=52
					9, 18, 0, -25, 8, -6, -35, -8, 3,
					-- layer=2 filter=119 channel=53
					-28, -70, 17, -28, -34, -69, -22, -75, -25,
					-- layer=2 filter=119 channel=54
					19, 12, -12, 16, 21, -13, -1, 4, 7,
					-- layer=2 filter=119 channel=55
					-8, 3, -3, -4, -9, 11, -5, -4, 1,
					-- layer=2 filter=119 channel=56
					25, 33, 6, -35, 0, -2, -24, -17, -17,
					-- layer=2 filter=119 channel=57
					6, -1, -7, 8, -5, -8, 6, 1, -11,
					-- layer=2 filter=119 channel=58
					15, 29, 15, 21, 51, 12, 8, 4, 33,
					-- layer=2 filter=119 channel=59
					22, 3, 0, -6, -65, 3, -19, -62, 5,
					-- layer=2 filter=119 channel=60
					40, -3, -4, 16, 26, -22, 17, 2, 5,
					-- layer=2 filter=119 channel=61
					15, 11, -39, 14, 12, -44, 26, 1, 12,
					-- layer=2 filter=119 channel=62
					22, 7, 3, -30, -34, 3, -67, -54, 11,
					-- layer=2 filter=119 channel=63
					19, 1, -8, 8, 17, 6, 32, 5, 14,
					-- layer=2 filter=119 channel=64
					-11, 4, -28, -5, 5, 4, 15, 3, 8,
					-- layer=2 filter=119 channel=65
					8, 6, -33, -27, -3, -65, -26, -27, -36,
					-- layer=2 filter=119 channel=66
					-41, 3, -2, 22, 23, 10, 43, 10, 2,
					-- layer=2 filter=119 channel=67
					21, 8, 5, -41, -7, -47, 17, -35, 9,
					-- layer=2 filter=119 channel=68
					-6, 3, -6, 4, -8, 0, 8, -13, 4,
					-- layer=2 filter=119 channel=69
					1, 9, -8, 14, -2, 24, 12, 2, 31,
					-- layer=2 filter=119 channel=70
					1, -5, 33, 23, 2, -6, -19, -18, -24,
					-- layer=2 filter=119 channel=71
					34, 31, 3, -16, 25, -6, -29, 3, 1,
					-- layer=2 filter=119 channel=72
					3, -8, -11, 40, 24, 43, 53, 62, 57,
					-- layer=2 filter=119 channel=73
					13, -48, -7, 16, 22, -20, 23, -20, 12,
					-- layer=2 filter=119 channel=74
					11, -7, 7, -18, -2, -23, -30, -29, -20,
					-- layer=2 filter=119 channel=75
					-12, 7, -6, 20, 12, -15, -23, -33, 5,
					-- layer=2 filter=119 channel=76
					-29, 15, 11, -6, -25, -40, -26, -69, 10,
					-- layer=2 filter=119 channel=77
					-4, -6, 7, -4, -12, 5, -12, 0, -5,
					-- layer=2 filter=119 channel=78
					-7, 17, -3, -22, -14, -7, -62, 16, 5,
					-- layer=2 filter=119 channel=79
					-6, 6, 0, -3, -5, -5, -7, -7, -5,
					-- layer=2 filter=119 channel=80
					-11, 2, 14, -26, -30, -20, 22, -16, 1,
					-- layer=2 filter=119 channel=81
					-1, -3, 15, -1, 0, -1, 12, 0, 6,
					-- layer=2 filter=119 channel=82
					0, 4, -8, 2, 5, -9, 1, 7, 6,
					-- layer=2 filter=119 channel=83
					14, 10, 1, -25, 7, -22, 24, -23, 12,
					-- layer=2 filter=119 channel=84
					1, -8, -2, 8, 7, 8, -4, 0, -11,
					-- layer=2 filter=119 channel=85
					-2, 3, -9, -8, -5, -4, 13, -8, -6,
					-- layer=2 filter=119 channel=86
					3, -13, -7, 19, 0, -1, 9, -10, 4,
					-- layer=2 filter=119 channel=87
					4, -33, 52, -34, -44, -8, -70, -50, -15,
					-- layer=2 filter=119 channel=88
					24, 38, 14, 0, 24, -3, -7, -12, -5,
					-- layer=2 filter=119 channel=89
					13, 13, 1, 25, -12, 28, -9, -5, 16,
					-- layer=2 filter=119 channel=90
					-7, 8, 7, -4, 11, -8, 5, 4, 4,
					-- layer=2 filter=119 channel=91
					11, 17, 23, 18, 11, 31, 5, 21, 32,
					-- layer=2 filter=119 channel=92
					12, 14, 4, 23, 41, 34, 16, 12, 43,
					-- layer=2 filter=119 channel=93
					-15, 12, -61, -65, 16, 8, -69, 30, 44,
					-- layer=2 filter=119 channel=94
					34, 5, 5, 26, -14, -49, 20, -43, 32,
					-- layer=2 filter=119 channel=95
					-10, -2, -2, -6, -8, 0, -12, -14, 1,
					-- layer=2 filter=119 channel=96
					32, 6, -17, 33, 2, -2, -17, -31, -40,
					-- layer=2 filter=119 channel=97
					-25, 0, 15, -21, -29, 2, -2, -4, 18,
					-- layer=2 filter=119 channel=98
					-7, 20, 13, 20, 35, 31, 0, 18, -13,
					-- layer=2 filter=119 channel=99
					-2, 43, 21, -3, -29, -27, 20, 18, -18,
					-- layer=2 filter=119 channel=100
					38, 21, 3, 4, -2, -23, 1, -49, -19,
					-- layer=2 filter=119 channel=101
					5, 33, 8, -15, 24, 11, -31, -1, 0,
					-- layer=2 filter=119 channel=102
					-18, 15, -14, -26, -51, -3, -39, -2, 10,
					-- layer=2 filter=119 channel=103
					-20, 20, 10, -15, -3, -26, 20, 0, -16,
					-- layer=2 filter=119 channel=104
					6, -20, -6, -39, -13, -35, -19, -69, 27,
					-- layer=2 filter=119 channel=105
					39, 23, -42, 27, -73, -27, -8, -42, -14,
					-- layer=2 filter=119 channel=106
					-52, -5, 9, -35, -1, 8, -18, -37, -34,
					-- layer=2 filter=119 channel=107
					9, -10, -16, 44, -3, -2, 16, -6, 19,
					-- layer=2 filter=119 channel=108
					21, 25, 9, 0, -10, -2, -28, -16, -26,
					-- layer=2 filter=119 channel=109
					0, 4, -10, -3, 0, -7, -10, 1, 11,
					-- layer=2 filter=119 channel=110
					-11, 0, -22, 36, 32, -13, 3, 22, -25,
					-- layer=2 filter=119 channel=111
					1, -1, 3, -9, -7, 0, 1, -8, -2,
					-- layer=2 filter=119 channel=112
					9, -2, 5, -23, -21, -36, 46, 30, 10,
					-- layer=2 filter=119 channel=113
					6, 0, 12, 0, 33, -3, 11, 32, -9,
					-- layer=2 filter=119 channel=114
					-6, 1, -15, -7, -8, -18, -10, -13, -13,
					-- layer=2 filter=119 channel=115
					0, 0, -6, 2, 3, 11, 3, 1, 7,
					-- layer=2 filter=119 channel=116
					18, -16, 16, -30, -14, -48, -46, -24, -52,
					-- layer=2 filter=119 channel=117
					41, 7, 1, 25, 36, 16, 63, 73, 68,
					-- layer=2 filter=119 channel=118
					23, 17, 41, -6, -50, -19, 5, 5, 11,
					-- layer=2 filter=119 channel=119
					-10, 19, 4, -10, -12, 0, -34, -59, -11,
					-- layer=2 filter=119 channel=120
					-3, -4, 7, 1, -6, 5, 10, -6, 3,
					-- layer=2 filter=119 channel=121
					10, 6, 7, 4, 7, -5, 11, -1, 10,
					-- layer=2 filter=119 channel=122
					-2, -11, -1, -3, 0, 0, -14, -4, -18,
					-- layer=2 filter=119 channel=123
					-9, 5, 0, 16, 0, 12, 6, 13, 36,
					-- layer=2 filter=119 channel=124
					33, -15, -4, -35, -47, 8, -18, -28, 19,
					-- layer=2 filter=119 channel=125
					10, 8, 4, -15, -3, -7, -5, -3, 3,
					-- layer=2 filter=119 channel=126
					7, -2, -24, 12, -40, 50, -43, -44, -92,
					-- layer=2 filter=119 channel=127
					6, 11, 2, 18, 1, -2, 0, -2, -2,
					-- layer=2 filter=120 channel=0
					-61, -50, -46, -52, 2, -29, -23, -10, 23,
					-- layer=2 filter=120 channel=1
					19, 16, 3, -27, 21, 13, -3, 1, 33,
					-- layer=2 filter=120 channel=2
					-6, -9, 5, -8, 5, -8, 2, -8, -8,
					-- layer=2 filter=120 channel=3
					-45, -7, -10, -4, 11, -15, -26, 23, 6,
					-- layer=2 filter=120 channel=4
					7, 0, 1, -94, -16, -32, -64, -10, -11,
					-- layer=2 filter=120 channel=5
					-17, -37, -45, -57, -12, -60, -24, -66, 5,
					-- layer=2 filter=120 channel=6
					-5, 27, -13, 56, 37, 8, 6, 31, 19,
					-- layer=2 filter=120 channel=7
					30, 31, -3, -52, -7, -23, 47, -11, 2,
					-- layer=2 filter=120 channel=8
					-7, 0, -4, -1, 5, 2, -2, -1, 1,
					-- layer=2 filter=120 channel=9
					-68, -11, -17, 8, -48, -37, -53, -37, 3,
					-- layer=2 filter=120 channel=10
					-38, -23, -28, 2, 23, -8, -15, 0, 18,
					-- layer=2 filter=120 channel=11
					-43, -20, -27, -64, -45, -48, -30, -48, -1,
					-- layer=2 filter=120 channel=12
					43, 22, 0, 4, 17, 9, 6, 3, 18,
					-- layer=2 filter=120 channel=13
					-1, -11, -3, -8, -3, 1, -3, -5, 0,
					-- layer=2 filter=120 channel=14
					17, 20, 9, -19, 17, 12, -18, 0, 6,
					-- layer=2 filter=120 channel=15
					14, -52, -47, 14, -9, 17, -1, 0, 29,
					-- layer=2 filter=120 channel=16
					-15, 7, 34, -16, 9, 1, -12, -16, 15,
					-- layer=2 filter=120 channel=17
					-7, -7, -8, -1, 0, 1, 1, -7, 10,
					-- layer=2 filter=120 channel=18
					11, -23, -25, -57, -4, -21, -11, -3, 0,
					-- layer=2 filter=120 channel=19
					0, -10, 16, 6, 39, 13, 28, 32, 18,
					-- layer=2 filter=120 channel=20
					-1, 3, -11, -2, -7, 11, -9, 0, 7,
					-- layer=2 filter=120 channel=21
					-13, -5, -15, -9, -22, -17, -6, 4, -9,
					-- layer=2 filter=120 channel=22
					-4, 7, 10, 5, -3, -3, -7, -3, 0,
					-- layer=2 filter=120 channel=23
					34, 43, 32, 8, -2, 21, -23, 1, -1,
					-- layer=2 filter=120 channel=24
					-35, 7, -9, -36, -34, -12, -22, -13, -17,
					-- layer=2 filter=120 channel=25
					-65, -57, -38, -70, -38, 11, -51, -23, -20,
					-- layer=2 filter=120 channel=26
					1, 2, -6, -4, -7, -7, -5, 0, -3,
					-- layer=2 filter=120 channel=27
					-22, 3, -6, -14, 4, 5, -22, -8, -1,
					-- layer=2 filter=120 channel=28
					-12, 4, 32, -20, -51, -61, 40, 19, 29,
					-- layer=2 filter=120 channel=29
					-9, 4, 0, 3, -1, -1, -7, 0, 6,
					-- layer=2 filter=120 channel=30
					-33, -13, -16, 5, -17, -4, -30, -62, -9,
					-- layer=2 filter=120 channel=31
					40, -27, -59, 37, -25, -29, 71, -1, -4,
					-- layer=2 filter=120 channel=32
					6, -10, 8, -3, -9, 6, 6, 4, 0,
					-- layer=2 filter=120 channel=33
					-13, -5, 5, 3, 12, -25, -2, 14, 31,
					-- layer=2 filter=120 channel=34
					-56, 6, 2, 7, -25, 23, 14, 4, -2,
					-- layer=2 filter=120 channel=35
					-35, -22, -56, -60, -39, -39, 21, -6, 13,
					-- layer=2 filter=120 channel=36
					6, -7, -5, -9, 9, 1, -2, -3, -2,
					-- layer=2 filter=120 channel=37
					-8, -40, -28, -48, -43, -36, -4, -29, -6,
					-- layer=2 filter=120 channel=38
					-40, 0, -14, -27, -7, -14, -50, -20, 0,
					-- layer=2 filter=120 channel=39
					-11, 32, 25, -20, -14, 42, -11, -41, 19,
					-- layer=2 filter=120 channel=40
					-15, 1, -21, -45, 5, -55, -9, 18, -28,
					-- layer=2 filter=120 channel=41
					-9, 4, 2, -1, -3, 0, 0, -5, 9,
					-- layer=2 filter=120 channel=42
					18, 36, 34, 34, 29, 11, -2, 27, 28,
					-- layer=2 filter=120 channel=43
					-35, -72, -9, 23, 23, -45, -14, 2, 0,
					-- layer=2 filter=120 channel=44
					-6, 4, 7, 5, -6, 5, 4, -1, 4,
					-- layer=2 filter=120 channel=45
					23, 10, 8, -2, 11, 21, 23, 30, 36,
					-- layer=2 filter=120 channel=46
					-40, 9, -18, 18, 24, 0, -16, 10, -26,
					-- layer=2 filter=120 channel=47
					-11, 20, 20, -54, -88, -71, 28, -9, 15,
					-- layer=2 filter=120 channel=48
					-11, -5, 7, 0, 6, 9, -8, -8, -8,
					-- layer=2 filter=120 channel=49
					29, -22, 26, -17, 19, -13, -30, 9, 27,
					-- layer=2 filter=120 channel=50
					13, 9, 1, 12, 0, -21, -13, -1, 13,
					-- layer=2 filter=120 channel=51
					-44, -36, -48, -38, -50, -57, -19, -41, -31,
					-- layer=2 filter=120 channel=52
					-48, 15, -8, -40, -54, -21, -19, -33, 9,
					-- layer=2 filter=120 channel=53
					24, 0, -8, 11, -14, -3, -39, -26, -21,
					-- layer=2 filter=120 channel=54
					32, 40, -38, -17, 4, 19, 12, 7, 1,
					-- layer=2 filter=120 channel=55
					1, 0, -3, 7, -4, 0, 9, 3, 2,
					-- layer=2 filter=120 channel=56
					0, 9, -17, -62, -37, -44, -32, -54, -19,
					-- layer=2 filter=120 channel=57
					-1, 2, 8, 5, 9, -8, -6, 3, 0,
					-- layer=2 filter=120 channel=58
					29, 16, 15, 23, -20, 10, -10, 5, 7,
					-- layer=2 filter=120 channel=59
					35, 19, -3, -41, -19, 62, 4, 6, -5,
					-- layer=2 filter=120 channel=60
					8, -15, -15, -10, 22, -20, 16, 4, -53,
					-- layer=2 filter=120 channel=61
					6, -37, -53, 11, 10, -57, 13, -21, -62,
					-- layer=2 filter=120 channel=62
					-26, 11, 6, 34, 21, 17, -48, 6, 29,
					-- layer=2 filter=120 channel=63
					18, -10, 1, -4, -18, 0, -4, -30, -42,
					-- layer=2 filter=120 channel=64
					-19, 10, 20, -9, 4, 14, -12, -6, 16,
					-- layer=2 filter=120 channel=65
					-11, -14, -52, 55, 3, -2, -13, -14, 2,
					-- layer=2 filter=120 channel=66
					44, -7, 18, 8, 12, 25, -11, 13, -12,
					-- layer=2 filter=120 channel=67
					-65, -14, -32, -3, -29, -22, 7, -39, -90,
					-- layer=2 filter=120 channel=68
					10, -5, -5, 0, -1, -1, 2, 4, 2,
					-- layer=2 filter=120 channel=69
					-6, 25, 20, -5, 24, 36, -1, -6, 40,
					-- layer=2 filter=120 channel=70
					1, -1, -18, -48, -36, -29, 16, 16, 11,
					-- layer=2 filter=120 channel=71
					0, -15, -10, 27, 63, 40, -12, 12, -8,
					-- layer=2 filter=120 channel=72
					41, 29, 42, -32, -17, -1, 18, 0, 12,
					-- layer=2 filter=120 channel=73
					15, 58, -57, -25, 0, -12, 13, 41, 15,
					-- layer=2 filter=120 channel=74
					-43, -36, -28, -12, -57, 11, 11, 14, -62,
					-- layer=2 filter=120 channel=75
					19, 6, 22, -14, -17, -10, 24, 2, -9,
					-- layer=2 filter=120 channel=76
					-6, -7, -45, -78, -42, -24, -41, -21, -21,
					-- layer=2 filter=120 channel=77
					9, 1, -7, 6, 0, 3, -13, -1, 9,
					-- layer=2 filter=120 channel=78
					-74, -36, -17, -56, -57, -6, -59, -35, 24,
					-- layer=2 filter=120 channel=79
					7, 3, 1, -9, -10, -7, 4, -6, 0,
					-- layer=2 filter=120 channel=80
					-16, 7, -3, -16, 39, 15, -48, -37, -18,
					-- layer=2 filter=120 channel=81
					-1, 0, 6, 5, 4, 7, -8, 1, 0,
					-- layer=2 filter=120 channel=82
					-8, 0, 0, -6, -3, 0, 0, 1, 2,
					-- layer=2 filter=120 channel=83
					23, -3, 27, 4, 23, 24, -36, -1, -2,
					-- layer=2 filter=120 channel=84
					-4, 3, 0, -8, 2, -6, -4, -4, -5,
					-- layer=2 filter=120 channel=85
					4, -8, 13, 6, 4, -4, 0, 12, 2,
					-- layer=2 filter=120 channel=86
					3, 13, 7, -2, 8, -2, -13, 9, -1,
					-- layer=2 filter=120 channel=87
					7, -6, 8, -39, 5, 6, -36, 7, 52,
					-- layer=2 filter=120 channel=88
					-23, -12, -5, -16, -41, -24, -19, -15, -32,
					-- layer=2 filter=120 channel=89
					25, 19, 39, -24, -2, 16, -15, 4, 24,
					-- layer=2 filter=120 channel=90
					7, -9, 9, -11, 1, 9, 5, 6, 0,
					-- layer=2 filter=120 channel=91
					22, 24, 24, -12, 18, 35, 24, 56, 28,
					-- layer=2 filter=120 channel=92
					41, 2, 10, -15, 25, 27, -25, 17, 21,
					-- layer=2 filter=120 channel=93
					-116, -32, -42, 49, 87, 38, 6, 73, 15,
					-- layer=2 filter=120 channel=94
					48, 24, -36, 30, 16, -3, -16, 13, -27,
					-- layer=2 filter=120 channel=95
					1, 6, 5, -15, 7, -8, -10, -4, 3,
					-- layer=2 filter=120 channel=96
					47, -1, -29, 29, 63, 77, 39, 37, 22,
					-- layer=2 filter=120 channel=97
					-59, -18, -5, 1, -4, 0, -12, -25, -8,
					-- layer=2 filter=120 channel=98
					-19, 0, -3, -56, -93, -46, 38, 12, 10,
					-- layer=2 filter=120 channel=99
					19, -5, -5, 15, -46, -9, -3, -41, -47,
					-- layer=2 filter=120 channel=100
					-14, -3, -23, -7, -8, 3, -16, -10, -5,
					-- layer=2 filter=120 channel=101
					-15, -12, -10, 15, 28, 7, 16, 21, -51,
					-- layer=2 filter=120 channel=102
					27, 4, -23, 28, 60, 58, 31, 32, 27,
					-- layer=2 filter=120 channel=103
					-1, 19, 14, -36, -38, -26, -10, -9, 15,
					-- layer=2 filter=120 channel=104
					22, 1, -34, -8, 4, -19, -69, 3, 10,
					-- layer=2 filter=120 channel=105
					52, 11, 35, -65, -49, 13, -39, 2, 42,
					-- layer=2 filter=120 channel=106
					-38, -32, -47, -34, -27, 20, 24, 24, 25,
					-- layer=2 filter=120 channel=107
					-34, 24, 1, 22, 4, 8, -13, 13, 73,
					-- layer=2 filter=120 channel=108
					-7, -8, 0, 8, 60, 22, 3, -19, 3,
					-- layer=2 filter=120 channel=109
					10, 0, -6, 16, 14, 10, 8, 10, -16,
					-- layer=2 filter=120 channel=110
					19, -4, 17, -13, -16, 0, -4, 12, -26,
					-- layer=2 filter=120 channel=111
					6, 11, 2, 11, 0, 5, 3, 10, -7,
					-- layer=2 filter=120 channel=112
					-38, -13, -27, -56, -33, -80, -60, -51, -26,
					-- layer=2 filter=120 channel=113
					13, 10, 24, 11, -23, -28, -28, -30, -45,
					-- layer=2 filter=120 channel=114
					8, 8, -1, 10, 2, -8, 15, 12, 14,
					-- layer=2 filter=120 channel=115
					-6, 0, 3, 6, -4, 8, 7, 9, 3,
					-- layer=2 filter=120 channel=116
					19, -54, -46, -30, 6, 35, -26, 7, 34,
					-- layer=2 filter=120 channel=117
					5, -5, -19, -18, -15, -44, 22, -12, -3,
					-- layer=2 filter=120 channel=118
					-22, 0, 14, -30, -10, -23, -43, 0, 9,
					-- layer=2 filter=120 channel=119
					5, 31, -9, -69, 30, -20, -21, 5, 11,
					-- layer=2 filter=120 channel=120
					0, -9, 8, 4, 1, 4, 6, 2, -3,
					-- layer=2 filter=120 channel=121
					-6, 3, -5, -6, 1, 7, -5, 8, -7,
					-- layer=2 filter=120 channel=122
					-5, -18, -2, 3, 0, 3, 0, 20, 9,
					-- layer=2 filter=120 channel=123
					36, 39, 24, -31, -41, -10, 34, 11, 9,
					-- layer=2 filter=120 channel=124
					7, -6, -9, 4, 39, 50, -35, 12, 62,
					-- layer=2 filter=120 channel=125
					9, -5, -1, -9, -5, -1, -4, 10, 1,
					-- layer=2 filter=120 channel=126
					24, -20, -1, 15, 4, 49, 32, 28, -28,
					-- layer=2 filter=120 channel=127
					30, 18, 38, -5, -16, 21, -71, -16, -3,
					-- layer=2 filter=121 channel=0
					6, -32, -12, 13, 22, 32, 0, 21, 9,
					-- layer=2 filter=121 channel=1
					-15, -16, -58, -3, -57, -12, -36, -39, -64,
					-- layer=2 filter=121 channel=2
					2, -2, -2, -8, 3, 8, -4, -4, 8,
					-- layer=2 filter=121 channel=3
					-12, -4, 13, 24, 4, 21, 28, 14, 26,
					-- layer=2 filter=121 channel=4
					-48, -47, -64, -11, 14, -49, 4, 9, -11,
					-- layer=2 filter=121 channel=5
					4, -14, -1, 23, 19, 13, 6, 17, 3,
					-- layer=2 filter=121 channel=6
					-11, 47, 21, 5, 18, 12, -20, -19, 0,
					-- layer=2 filter=121 channel=7
					-23, -30, -9, -3, -38, -26, -29, 19, -28,
					-- layer=2 filter=121 channel=8
					-8, 4, -6, 0, -4, -1, 0, 5, 7,
					-- layer=2 filter=121 channel=9
					-32, -47, -9, 2, -1, -16, -6, -12, -7,
					-- layer=2 filter=121 channel=10
					18, -19, -16, 13, 4, 24, 11, 31, 40,
					-- layer=2 filter=121 channel=11
					-5, 12, 5, 3, 16, 26, 34, 31, 18,
					-- layer=2 filter=121 channel=12
					8, -12, -35, -47, 5, -4, -8, -50, -30,
					-- layer=2 filter=121 channel=13
					1, 0, 1, -7, 0, 7, -3, 2, 3,
					-- layer=2 filter=121 channel=14
					3, -10, -10, -14, -11, 2, -8, -12, -19,
					-- layer=2 filter=121 channel=15
					25, -15, 11, 19, -14, 17, 1, -22, -25,
					-- layer=2 filter=121 channel=16
					-17, -46, -24, 25, -12, -38, -74, -36, 15,
					-- layer=2 filter=121 channel=17
					-10, -3, -5, 8, 3, -7, 4, -8, 1,
					-- layer=2 filter=121 channel=18
					-78, -67, -26, -26, 12, -25, -2, -9, -38,
					-- layer=2 filter=121 channel=19
					-25, -29, -63, -35, -54, -26, -46, -18, -15,
					-- layer=2 filter=121 channel=20
					-10, 7, 8, 0, 12, -8, -7, -6, 8,
					-- layer=2 filter=121 channel=21
					9, 6, 20, 8, 3, 10, 0, 11, 9,
					-- layer=2 filter=121 channel=22
					-8, 8, 10, 2, -8, 5, 2, -6, 2,
					-- layer=2 filter=121 channel=23
					21, -13, -17, -39, 3, -65, 14, -35, -40,
					-- layer=2 filter=121 channel=24
					17, 15, 28, 24, -4, 7, -13, 14, 24,
					-- layer=2 filter=121 channel=25
					15, 25, 35, 6, -11, 0, -7, 11, 12,
					-- layer=2 filter=121 channel=26
					-4, 6, -5, 4, 6, -4, 10, 4, -5,
					-- layer=2 filter=121 channel=27
					5, -25, -24, 11, -22, -27, 5, 0, -1,
					-- layer=2 filter=121 channel=28
					28, -21, 4, -21, -41, -8, -26, 22, 36,
					-- layer=2 filter=121 channel=29
					-7, -6, -7, 0, 2, -6, -8, -7, 6,
					-- layer=2 filter=121 channel=30
					-14, -13, -11, 7, -27, -34, -8, -5, -3,
					-- layer=2 filter=121 channel=31
					11, 16, 35, 33, 31, 57, 13, 7, 47,
					-- layer=2 filter=121 channel=32
					0, 6, -9, 0, -8, -6, -10, 6, -6,
					-- layer=2 filter=121 channel=33
					37, 19, 5, 12, -9, 0, 22, 3, -16,
					-- layer=2 filter=121 channel=34
					-15, -7, 24, 18, 18, 18, -28, -12, 2,
					-- layer=2 filter=121 channel=35
					10, -39, 3, -9, -20, -22, -5, 34, 4,
					-- layer=2 filter=121 channel=36
					4, -2, -5, 4, 7, -8, -14, -9, -3,
					-- layer=2 filter=121 channel=37
					9, 13, 7, 20, -1, 10, 13, 0, 13,
					-- layer=2 filter=121 channel=38
					-4, -17, -42, -19, -12, -9, 25, 12, -6,
					-- layer=2 filter=121 channel=39
					16, -15, -3, -66, -97, -70, -95, -84, -67,
					-- layer=2 filter=121 channel=40
					-15, -12, 18, 4, 30, 7, 51, -9, 10,
					-- layer=2 filter=121 channel=41
					-9, 5, 8, -7, 7, -7, 11, 0, -9,
					-- layer=2 filter=121 channel=42
					10, -16, -18, -27, -50, -28, -28, -25, -2,
					-- layer=2 filter=121 channel=43
					-2, -8, 23, -10, 24, 48, 38, 44, 59,
					-- layer=2 filter=121 channel=44
					3, 2, 0, 6, -6, -9, 0, 7, -9,
					-- layer=2 filter=121 channel=45
					-44, -30, -36, -31, -74, -42, -103, -68, -50,
					-- layer=2 filter=121 channel=46
					-30, -22, -55, 14, 16, 0, 41, 24, 21,
					-- layer=2 filter=121 channel=47
					12, 17, 35, 7, -19, 4, -12, -26, 11,
					-- layer=2 filter=121 channel=48
					-7, -5, -1, -3, -10, 9, -8, -7, 7,
					-- layer=2 filter=121 channel=49
					-73, -51, -42, -47, -12, 1, 4, -18, -31,
					-- layer=2 filter=121 channel=50
					11, 4, 14, -8, 27, -6, 9, 0, 1,
					-- layer=2 filter=121 channel=51
					2, 6, 20, 6, 21, 34, 14, 14, 27,
					-- layer=2 filter=121 channel=52
					-3, 1, 29, 12, 7, -5, 17, 2, -8,
					-- layer=2 filter=121 channel=53
					-77, -33, 7, -34, -10, 46, -42, -12, -23,
					-- layer=2 filter=121 channel=54
					0, 32, 14, 2, 21, -1, -5, 22, 7,
					-- layer=2 filter=121 channel=55
					0, 2, 0, 9, 3, -5, -9, 8, 8,
					-- layer=2 filter=121 channel=56
					3, -4, -7, 1, 9, 19, 45, 14, 16,
					-- layer=2 filter=121 channel=57
					-7, -2, -6, -4, 3, 7, -16, 5, 4,
					-- layer=2 filter=121 channel=58
					34, -3, -21, -48, 11, -3, -16, -20, -16,
					-- layer=2 filter=121 channel=59
					-10, -26, -67, -61, -8, 17, -87, -29, -62,
					-- layer=2 filter=121 channel=60
					11, -1, -34, -62, -15, -21, -50, -68, -7,
					-- layer=2 filter=121 channel=61
					-41, -48, -49, -37, 0, -21, -18, -44, 0,
					-- layer=2 filter=121 channel=62
					-16, 3, 42, -19, 11, 11, 0, 11, -23,
					-- layer=2 filter=121 channel=63
					-3, -42, -44, -36, -23, -33, -45, -3, -16,
					-- layer=2 filter=121 channel=64
					18, 21, 28, 28, -8, -30, 15, -22, -33,
					-- layer=2 filter=121 channel=65
					-41, 8, -38, -21, -18, -18, 19, 20, -5,
					-- layer=2 filter=121 channel=66
					-22, -17, 23, 8, -29, -2, -28, -9, 40,
					-- layer=2 filter=121 channel=67
					-9, -9, -40, 5, 12, -19, 0, -25, 15,
					-- layer=2 filter=121 channel=68
					-5, 0, -5, -7, 7, 0, 0, -8, 3,
					-- layer=2 filter=121 channel=69
					26, 39, 21, 5, 5, -20, 12, -26, -30,
					-- layer=2 filter=121 channel=70
					26, -11, 16, -2, -12, 6, 10, 25, 21,
					-- layer=2 filter=121 channel=71
					-27, 3, 13, -20, 4, 2, 1, -20, 3,
					-- layer=2 filter=121 channel=72
					30, 7, 21, -7, -7, -20, -1, 39, 54,
					-- layer=2 filter=121 channel=73
					27, 37, 25, 33, 17, 20, 6, 55, 64,
					-- layer=2 filter=121 channel=74
					-37, -46, -43, -26, 24, -10, 1, 25, 19,
					-- layer=2 filter=121 channel=75
					-19, 17, 41, -43, 13, 19, 2, 27, 21,
					-- layer=2 filter=121 channel=76
					-30, 18, -18, 66, 24, -2, 6, -22, -48,
					-- layer=2 filter=121 channel=77
					1, -2, 6, -2, 3, -7, -3, 3, 10,
					-- layer=2 filter=121 channel=78
					-22, 7, 13, 11, 7, 22, 11, 19, 6,
					-- layer=2 filter=121 channel=79
					5, -10, -6, 2, 8, 0, -3, 0, 0,
					-- layer=2 filter=121 channel=80
					-28, 1, -27, -20, 9, -8, -22, -19, 8,
					-- layer=2 filter=121 channel=81
					-4, -3, -2, 1, -2, 5, -10, -6, -3,
					-- layer=2 filter=121 channel=82
					-2, 9, 0, 9, -2, 0, -3, 9, -8,
					-- layer=2 filter=121 channel=83
					-12, -69, -12, 10, -20, -45, -10, -6, -25,
					-- layer=2 filter=121 channel=84
					-11, -10, 1, 7, 4, -4, -6, 4, 7,
					-- layer=2 filter=121 channel=85
					1, -2, 2, -3, 0, -4, -3, -1, 0,
					-- layer=2 filter=121 channel=86
					4, -12, -10, 9, 9, -8, -1, 4, -9,
					-- layer=2 filter=121 channel=87
					33, 13, 33, -13, 7, -24, 21, 13, -57,
					-- layer=2 filter=121 channel=88
					40, -12, -16, -15, -25, -60, -12, -28, 0,
					-- layer=2 filter=121 channel=89
					30, 12, -10, -23, 5, -4, -36, -11, -61,
					-- layer=2 filter=121 channel=90
					-3, 9, 7, -10, -3, -3, -1, 8, -10,
					-- layer=2 filter=121 channel=91
					26, -2, -5, -43, -23, -20, -25, -36, -17,
					-- layer=2 filter=121 channel=92
					10, 12, -32, -45, -16, -4, -21, -46, -61,
					-- layer=2 filter=121 channel=93
					19, -17, 7, 21, 31, 28, 34, -1, 15,
					-- layer=2 filter=121 channel=94
					8, -45, -3, -21, 15, -36, -1, -6, -13,
					-- layer=2 filter=121 channel=95
					-8, -9, -15, -13, 7, -17, -14, 1, -5,
					-- layer=2 filter=121 channel=96
					23, 40, 83, 87, 11, 22, 34, -6, -17,
					-- layer=2 filter=121 channel=97
					-14, -26, 3, -1, -7, -11, 16, -13, -5,
					-- layer=2 filter=121 channel=98
					30, 11, 29, 0, -7, 5, 7, 28, 21,
					-- layer=2 filter=121 channel=99
					-27, -1, 44, 30, -14, 22, -2, 13, 0,
					-- layer=2 filter=121 channel=100
					0, -58, -31, -19, 12, 1, -9, 23, 25,
					-- layer=2 filter=121 channel=101
					6, 23, 36, -11, 9, 20, 0, -1, 5,
					-- layer=2 filter=121 channel=102
					-80, 15, 25, 35, 37, -21, 58, -17, -50,
					-- layer=2 filter=121 channel=103
					-14, 33, 11, -16, -4, 21, -4, 0, 17,
					-- layer=2 filter=121 channel=104
					-42, -12, -23, -39, 0, -41, -9, 1, -64,
					-- layer=2 filter=121 channel=105
					-22, -2, -32, -11, 0, -6, -39, 8, 6,
					-- layer=2 filter=121 channel=106
					7, -12, -23, -23, -8, -14, -24, 3, -24,
					-- layer=2 filter=121 channel=107
					6, 1, 17, -26, 10, 37, 21, 31, -33,
					-- layer=2 filter=121 channel=108
					-79, -61, 3, -15, -42, -24, -9, -29, -65,
					-- layer=2 filter=121 channel=109
					-1, -19, -17, 8, 0, 1, 7, 3, 11,
					-- layer=2 filter=121 channel=110
					28, -1, -1, 29, 0, -39, -24, 4, -29,
					-- layer=2 filter=121 channel=111
					-5, -9, 1, -6, 1, 1, 0, 2, 4,
					-- layer=2 filter=121 channel=112
					-3, 8, -20, -25, -6, 7, 19, 0, 10,
					-- layer=2 filter=121 channel=113
					-10, -43, -46, -52, -72, -6, 13, 0, -55,
					-- layer=2 filter=121 channel=114
					-3, -8, -4, -6, -17, -10, -4, 0, 0,
					-- layer=2 filter=121 channel=115
					-7, 5, 0, -1, -3, -1, 3, -3, 6,
					-- layer=2 filter=121 channel=116
					34, -5, 27, 27, 6, -34, 29, -8, -10,
					-- layer=2 filter=121 channel=117
					-24, 36, 26, 12, -19, -2, 21, 54, 13,
					-- layer=2 filter=121 channel=118
					-4, 15, 20, 33, 13, 19, 44, 22, 42,
					-- layer=2 filter=121 channel=119
					-42, -64, -20, -22, -45, -67, 11, 8, -61,
					-- layer=2 filter=121 channel=120
					10, -8, -5, 8, 2, 1, -10, 9, -7,
					-- layer=2 filter=121 channel=121
					2, -2, 6, 5, 5, -2, -10, 1, -11,
					-- layer=2 filter=121 channel=122
					13, -4, 14, -1, -2, -12, -8, -3, 10,
					-- layer=2 filter=121 channel=123
					-15, 6, 13, -4, -33, -17, -37, 37, -10,
					-- layer=2 filter=121 channel=124
					13, 22, -30, 49, 34, -8, 58, 23, -17,
					-- layer=2 filter=121 channel=125
					0, 0, -1, -4, 6, -7, 14, 6, -10,
					-- layer=2 filter=121 channel=126
					14, -108, -7, -17, 57, -47, -115, 29, -60,
					-- layer=2 filter=121 channel=127
					8, -4, -23, -10, -60, -14, 19, -23, -61,
					-- layer=2 filter=122 channel=0
					-18, 0, -4, 1, -40, -39, 17, -11, -30,
					-- layer=2 filter=122 channel=1
					28, -44, -14, 7, -13, 13, -31, -35, -63,
					-- layer=2 filter=122 channel=2
					-3, 4, 9, -3, -2, -1, -3, 2, 5,
					-- layer=2 filter=122 channel=3
					-26, 4, 7, -10, 8, -10, 14, -10, -23,
					-- layer=2 filter=122 channel=4
					19, -48, -46, -51, -59, 6, 8, -6, -2,
					-- layer=2 filter=122 channel=5
					7, -7, 0, 23, 2, 10, 0, -24, -10,
					-- layer=2 filter=122 channel=6
					-22, -40, 41, 22, -20, 36, 18, 50, 2,
					-- layer=2 filter=122 channel=7
					-13, -64, -64, 44, 30, 57, 31, 8, 0,
					-- layer=2 filter=122 channel=8
					0, -2, 1, -6, -2, 0, 0, 10, 0,
					-- layer=2 filter=122 channel=9
					-8, -4, -11, 25, 39, 15, 7, -2, 11,
					-- layer=2 filter=122 channel=10
					-32, 24, -3, -13, -16, -31, 22, -17, -4,
					-- layer=2 filter=122 channel=11
					1, 8, -4, 0, 2, 18, -6, 9, -4,
					-- layer=2 filter=122 channel=12
					-22, -13, -11, 14, 35, 20, -26, -8, -10,
					-- layer=2 filter=122 channel=13
					5, -3, -9, -6, -5, 6, 7, -4, -6,
					-- layer=2 filter=122 channel=14
					24, -10, -5, -13, -16, 5, -29, -47, -26,
					-- layer=2 filter=122 channel=15
					-66, -83, 2, -29, 10, 34, -13, -27, -22,
					-- layer=2 filter=122 channel=16
					-21, -20, -57, 31, 2, 25, 5, -4, 29,
					-- layer=2 filter=122 channel=17
					1, 6, 0, 0, -1, -9, 7, 5, 7,
					-- layer=2 filter=122 channel=18
					26, -62, -33, -25, 19, -3, -1, -1, -2,
					-- layer=2 filter=122 channel=19
					0, -15, -3, 52, -10, 39, -15, 47, -16,
					-- layer=2 filter=122 channel=20
					9, -8, -6, -3, -7, 8, 5, -10, 6,
					-- layer=2 filter=122 channel=21
					-16, -5, -5, -1, -3, -15, -9, -1, -1,
					-- layer=2 filter=122 channel=22
					7, 7, -3, 6, 0, -6, 7, 7, -1,
					-- layer=2 filter=122 channel=23
					-7, -33, -27, -18, -35, -9, 37, 6, 3,
					-- layer=2 filter=122 channel=24
					3, 18, 4, -20, 27, -23, 0, 5, 2,
					-- layer=2 filter=122 channel=25
					13, 23, 12, -2, 30, 0, -11, 5, 9,
					-- layer=2 filter=122 channel=26
					-3, -4, 4, 8, -4, -3, -5, 10, 4,
					-- layer=2 filter=122 channel=27
					13, -8, -4, 37, -13, -21, -25, -53, -38,
					-- layer=2 filter=122 channel=28
					0, 22, 53, -35, -24, 1, 3, 41, 45,
					-- layer=2 filter=122 channel=29
					4, 0, 3, 9, -5, -6, 2, 0, -9,
					-- layer=2 filter=122 channel=30
					8, -56, -19, -6, -63, -17, 31, -90, -5,
					-- layer=2 filter=122 channel=31
					-49, -36, 6, -9, -35, -5, 52, 15, 0,
					-- layer=2 filter=122 channel=32
					-5, -4, -8, -2, -1, 9, -7, -2, 3,
					-- layer=2 filter=122 channel=33
					41, 26, -22, 1, -15, 46, -7, -49, -17,
					-- layer=2 filter=122 channel=34
					28, -53, -21, 25, -25, -33, 38, 26, 32,
					-- layer=2 filter=122 channel=35
					15, -20, 22, -26, -48, -15, 28, 30, 16,
					-- layer=2 filter=122 channel=36
					-11, -7, -4, 0, -19, 1, 3, 8, -2,
					-- layer=2 filter=122 channel=37
					20, -15, 18, -3, -22, -14, -9, -20, -9,
					-- layer=2 filter=122 channel=38
					0, -18, 9, 9, -12, 0, -30, -35, -82,
					-- layer=2 filter=122 channel=39
					-39, -46, -31, 25, 33, 24, -10, 10, 7,
					-- layer=2 filter=122 channel=40
					12, -15, -7, -93, -16, 58, -4, 9, -8,
					-- layer=2 filter=122 channel=41
					11, 8, -6, 8, -1, 0, -4, 5, 4,
					-- layer=2 filter=122 channel=42
					2, -3, -14, -7, 7, 15, -43, -4, -11,
					-- layer=2 filter=122 channel=43
					7, 20, 47, -7, -28, -8, -25, -27, 0,
					-- layer=2 filter=122 channel=44
					-5, -7, -1, -8, 8, 0, 5, 5, -6,
					-- layer=2 filter=122 channel=45
					-30, -25, 28, -35, -33, 4, -2, -24, -44,
					-- layer=2 filter=122 channel=46
					-47, -42, -51, 17, 9, -21, -8, -46, 0,
					-- layer=2 filter=122 channel=47
					-5, 26, -11, -19, -53, -5, 17, 28, 18,
					-- layer=2 filter=122 channel=48
					0, -7, -10, -5, -7, 4, -8, -1, -9,
					-- layer=2 filter=122 channel=49
					-9, -56, -42, -19, -2, 1, -68, 13, -2,
					-- layer=2 filter=122 channel=50
					-18, -2, 22, 11, -1, 8, -2, -9, -7,
					-- layer=2 filter=122 channel=51
					26, 17, 8, -14, -13, 1, -6, -9, -20,
					-- layer=2 filter=122 channel=52
					34, -50, 35, 30, 2, 36, 41, -51, -29,
					-- layer=2 filter=122 channel=53
					-40, -74, 1, -26, 2, 1, -27, -11, 64,
					-- layer=2 filter=122 channel=54
					11, -23, -49, -9, 2, 24, 31, 47, 46,
					-- layer=2 filter=122 channel=55
					0, 0, 8, 0, 8, -3, -4, 8, -9,
					-- layer=2 filter=122 channel=56
					6, -3, -4, 15, -10, -11, -29, -29, -16,
					-- layer=2 filter=122 channel=57
					-8, -1, -4, -5, -4, 0, 3, -12, 3,
					-- layer=2 filter=122 channel=58
					-39, -4, -15, 21, 48, 38, 10, -24, -1,
					-- layer=2 filter=122 channel=59
					-3, -47, 19, 10, 19, 32, -23, 10, -40,
					-- layer=2 filter=122 channel=60
					4, -41, 10, 16, 1, -15, 10, 35, -48,
					-- layer=2 filter=122 channel=61
					-35, -31, 28, 22, -40, -55, 24, 22, -48,
					-- layer=2 filter=122 channel=62
					8, -32, -25, 26, -18, 29, -7, 30, 17,
					-- layer=2 filter=122 channel=63
					-49, -28, 6, -34, -33, -24, 14, -12, -2,
					-- layer=2 filter=122 channel=64
					-2, -38, -41, -26, -25, -55, 28, -28, -31,
					-- layer=2 filter=122 channel=65
					-21, -48, 59, -3, -22, 9, 17, 0, -50,
					-- layer=2 filter=122 channel=66
					-4, -21, 5, 3, 22, 13, 2, -6, 16,
					-- layer=2 filter=122 channel=67
					-30, 16, -18, 24, 60, -60, 38, -8, -26,
					-- layer=2 filter=122 channel=68
					3, -11, 4, 0, -5, -8, -3, 5, 5,
					-- layer=2 filter=122 channel=69
					5, -25, -37, -13, -23, -46, 34, -16, -31,
					-- layer=2 filter=122 channel=70
					-6, -31, -8, -33, -48, 0, 35, 30, 22,
					-- layer=2 filter=122 channel=71
					12, 20, 27, 28, 5, -13, -5, -41, -36,
					-- layer=2 filter=122 channel=72
					49, 4, 5, -2, -20, 12, -28, 11, 20,
					-- layer=2 filter=122 channel=73
					-36, -15, 13, 10, -4, 4, 13, 37, -16,
					-- layer=2 filter=122 channel=74
					-70, 17, -30, -41, 1, 7, 12, -43, -23,
					-- layer=2 filter=122 channel=75
					-58, -2, 18, -36, -21, 46, -36, -56, 7,
					-- layer=2 filter=122 channel=76
					41, -23, 20, 14, -29, 2, 59, 26, -23,
					-- layer=2 filter=122 channel=77
					-6, -8, 4, 0, -3, 0, -10, -10, -4,
					-- layer=2 filter=122 channel=78
					18, -5, -4, 23, -11, -6, 19, 3, 3,
					-- layer=2 filter=122 channel=79
					0, 4, -10, 0, 3, -3, -3, 7, 0,
					-- layer=2 filter=122 channel=80
					-61, -56, -38, -55, -69, 3, -34, -34, -50,
					-- layer=2 filter=122 channel=81
					11, 6, 2, 0, -5, 11, 2, 12, 2,
					-- layer=2 filter=122 channel=82
					-7, 5, -3, 5, -8, 8, -8, 4, 6,
					-- layer=2 filter=122 channel=83
					-51, -15, 20, 14, -35, 10, -10, -44, -5,
					-- layer=2 filter=122 channel=84
					9, 5, 3, -1, 3, -11, -5, -4, -5,
					-- layer=2 filter=122 channel=85
					10, 1, 0, -1, -4, 9, 4, -10, 1,
					-- layer=2 filter=122 channel=86
					-1, 4, -4, 1, 1, 5, -10, -10, 6,
					-- layer=2 filter=122 channel=87
					-17, -51, -36, -57, -49, 33, -22, -15, -42,
					-- layer=2 filter=122 channel=88
					-15, -9, -4, -60, -64, -18, 20, -36, -34,
					-- layer=2 filter=122 channel=89
					1, -12, 0, 1, 13, 44, -26, -31, -20,
					-- layer=2 filter=122 channel=90
					-9, -6, 6, 7, -1, -2, 7, 0, -8,
					-- layer=2 filter=122 channel=91
					5, 35, 22, 19, 43, 18, -44, -5, -12,
					-- layer=2 filter=122 channel=92
					19, -3, -15, 15, 4, 24, -69, 0, -17,
					-- layer=2 filter=122 channel=93
					1, -42, 23, 40, 34, 6, 14, 25, -35,
					-- layer=2 filter=122 channel=94
					-55, -43, 0, 65, -46, 18, 10, 39, -4,
					-- layer=2 filter=122 channel=95
					18, -17, 16, 0, -3, -16, -6, 18, 2,
					-- layer=2 filter=122 channel=96
					43, 43, 43, -20, 1, 9, -6, 12, -35,
					-- layer=2 filter=122 channel=97
					-8, -21, -35, -10, 40, 23, -25, -40, 3,
					-- layer=2 filter=122 channel=98
					-48, 3, 19, -42, -73, -20, 29, 27, 7,
					-- layer=2 filter=122 channel=99
					16, -13, 59, 9, 5, -4, 5, 6, -16,
					-- layer=2 filter=122 channel=100
					-16, 6, -23, 52, -49, -8, 47, -42, 0,
					-- layer=2 filter=122 channel=101
					15, 29, 27, 3, 24, 8, -17, 0, -14,
					-- layer=2 filter=122 channel=102
					68, 33, 12, 13, 5, -20, 2, -41, -56,
					-- layer=2 filter=122 channel=103
					25, 30, -5, 55, 1, -45, -40, -24, -67,
					-- layer=2 filter=122 channel=104
					-52, -62, -46, -25, -41, 4, -50, 24, -6,
					-- layer=2 filter=122 channel=105
					65, -1, -12, -16, -5, 1, 18, 74, -5,
					-- layer=2 filter=122 channel=106
					3, 33, 15, 3, 29, 23, -8, 17, 20,
					-- layer=2 filter=122 channel=107
					29, -19, -2, -22, -38, -4, -59, -32, 29,
					-- layer=2 filter=122 channel=108
					43, -24, 19, -2, -12, 2, -18, -38, -47,
					-- layer=2 filter=122 channel=109
					-3, -18, 17, -12, 0, -22, 5, 12, 12,
					-- layer=2 filter=122 channel=110
					36, 26, 11, 24, 24, -16, 18, -12, 1,
					-- layer=2 filter=122 channel=111
					2, -3, -6, 0, 6, -4, 8, 0, 9,
					-- layer=2 filter=122 channel=112
					-1, -23, 28, 4, -8, -55, 22, -25, -71,
					-- layer=2 filter=122 channel=113
					-23, -69, 22, -35, -111, -41, 26, -50, -16,
					-- layer=2 filter=122 channel=114
					0, -6, 2, 12, 4, -9, -1, -2, 6,
					-- layer=2 filter=122 channel=115
					-6, -6, -1, -8, -10, 0, -3, 6, -1,
					-- layer=2 filter=122 channel=116
					22, -52, -35, -44, -17, 2, 0, -26, -19,
					-- layer=2 filter=122 channel=117
					-32, 0, -26, 33, 0, 20, 29, 31, 20,
					-- layer=2 filter=122 channel=118
					-9, 16, 30, -8, -14, 1, -17, -42, -22,
					-- layer=2 filter=122 channel=119
					62, -32, -39, -1, -32, -34, -15, -5, 9,
					-- layer=2 filter=122 channel=120
					-5, 8, 6, 0, 2, -3, 3, -2, 7,
					-- layer=2 filter=122 channel=121
					8, 5, -8, 2, -2, 3, 5, -5, -1,
					-- layer=2 filter=122 channel=122
					-5, -10, 10, -2, 9, 4, 8, -10, 0,
					-- layer=2 filter=122 channel=123
					28, -24, -30, 13, -2, 40, 20, 21, 13,
					-- layer=2 filter=122 channel=124
					-21, -74, -15, 17, 7, 60, 19, -1, 11,
					-- layer=2 filter=122 channel=125
					3, 0, -9, 3, 8, -10, -2, -7, 3,
					-- layer=2 filter=122 channel=126
					-19, -39, 63, 33, 6, -24, -23, 0, -45,
					-- layer=2 filter=122 channel=127
					30, -55, 29, -92, -84, -38, 29, -68, -11,
					-- layer=2 filter=123 channel=0
					-9, -1, 7, -8, 6, -9, 4, -5, 6,
					-- layer=2 filter=123 channel=1
					-5, 4, -14, -11, -5, -2, -9, -7, -8,
					-- layer=2 filter=123 channel=2
					1, 4, 1, -6, -3, -1, 3, 7, -10,
					-- layer=2 filter=123 channel=3
					2, 8, -4, 6, 5, -4, 0, 9, 5,
					-- layer=2 filter=123 channel=4
					-1, 3, 2, 0, 0, 1, -10, 7, 9,
					-- layer=2 filter=123 channel=5
					4, 0, 5, -1, 3, -3, 8, -10, 0,
					-- layer=2 filter=123 channel=6
					1, -9, -2, -12, 4, 9, -13, 0, 0,
					-- layer=2 filter=123 channel=7
					2, -7, -6, 6, -1, -9, 4, 0, 1,
					-- layer=2 filter=123 channel=8
					2, 0, -3, -1, -2, 6, 11, 8, -9,
					-- layer=2 filter=123 channel=9
					0, -2, -11, 6, 8, 6, -5, 0, -1,
					-- layer=2 filter=123 channel=10
					-13, -1, -3, -12, -4, -6, -6, -10, -4,
					-- layer=2 filter=123 channel=11
					1, 7, -12, -8, -2, -2, 3, 2, 6,
					-- layer=2 filter=123 channel=12
					5, 3, 6, -3, -11, 4, 0, -3, -10,
					-- layer=2 filter=123 channel=13
					3, -7, 0, -4, -11, -2, -9, -3, 7,
					-- layer=2 filter=123 channel=14
					0, 0, -8, -2, 1, -15, -7, -11, -6,
					-- layer=2 filter=123 channel=15
					-2, -5, -5, -6, -10, -3, 0, 5, -12,
					-- layer=2 filter=123 channel=16
					0, 6, -1, -5, 0, 1, 4, -1, -6,
					-- layer=2 filter=123 channel=17
					10, -4, 2, 6, -7, 2, -8, 8, -2,
					-- layer=2 filter=123 channel=18
					-6, -11, -9, 2, -6, -10, -8, -7, -7,
					-- layer=2 filter=123 channel=19
					5, -3, 7, -10, -1, -16, -15, -2, -14,
					-- layer=2 filter=123 channel=20
					3, -9, 6, -10, 7, 8, -8, -3, 0,
					-- layer=2 filter=123 channel=21
					2, 2, 6, -8, 8, -8, 5, -10, -5,
					-- layer=2 filter=123 channel=22
					-3, 3, 2, -4, -1, -9, -8, 8, 1,
					-- layer=2 filter=123 channel=23
					8, 6, -13, -7, -1, 0, -7, -11, -2,
					-- layer=2 filter=123 channel=24
					0, 0, -5, -2, 4, -9, -5, -11, 4,
					-- layer=2 filter=123 channel=25
					-14, -19, -11, 1, -1, 0, 5, 3, 0,
					-- layer=2 filter=123 channel=26
					1, 1, -5, -6, -7, 10, 2, 0, 2,
					-- layer=2 filter=123 channel=27
					3, 4, -3, 4, -2, -3, 1, -1, 15,
					-- layer=2 filter=123 channel=28
					-7, 6, -2, -6, 0, 9, -2, 10, -2,
					-- layer=2 filter=123 channel=29
					0, -8, -3, 2, 3, -10, 0, 2, -10,
					-- layer=2 filter=123 channel=30
					7, -8, -12, 6, -4, 4, 0, 4, -11,
					-- layer=2 filter=123 channel=31
					-1, 5, 3, -8, -2, -11, 0, -9, -2,
					-- layer=2 filter=123 channel=32
					-9, -2, 5, 6, -4, 6, -9, -9, -9,
					-- layer=2 filter=123 channel=33
					-6, -10, -10, -1, -5, 4, -11, 4, -1,
					-- layer=2 filter=123 channel=34
					-10, -9, 0, -9, -9, -11, -10, -10, -7,
					-- layer=2 filter=123 channel=35
					2, -8, -5, -9, -7, -10, 4, -3, 1,
					-- layer=2 filter=123 channel=36
					-7, 3, 0, -8, 0, -9, 3, -7, 6,
					-- layer=2 filter=123 channel=37
					-14, -1, -9, -4, -15, -18, -2, -8, -2,
					-- layer=2 filter=123 channel=38
					-11, -2, -6, -13, 4, -3, -3, -9, 5,
					-- layer=2 filter=123 channel=39
					9, 8, -5, 7, 3, 7, -8, -7, -2,
					-- layer=2 filter=123 channel=40
					2, -17, -4, -3, -8, -7, 1, 5, -12,
					-- layer=2 filter=123 channel=41
					0, -2, 6, -3, -3, -3, 3, 0, -7,
					-- layer=2 filter=123 channel=42
					10, -3, 6, -8, -12, 0, -11, -11, 1,
					-- layer=2 filter=123 channel=43
					8, 5, -8, 8, 2, -8, 8, 0, -11,
					-- layer=2 filter=123 channel=44
					7, -1, 1, -2, 0, -9, 2, 2, 10,
					-- layer=2 filter=123 channel=45
					-8, -10, -5, 3, -6, 1, -3, -13, 0,
					-- layer=2 filter=123 channel=46
					7, 1, -13, 3, -10, -8, 1, 0, 0,
					-- layer=2 filter=123 channel=47
					-3, -7, -13, 10, -3, 6, -11, 7, 0,
					-- layer=2 filter=123 channel=48
					-9, -9, 9, 6, 6, 7, -9, -7, -1,
					-- layer=2 filter=123 channel=49
					-3, 3, 3, -10, 0, 0, 8, -5, -13,
					-- layer=2 filter=123 channel=50
					3, 7, -11, 0, 1, 9, 3, -5, 8,
					-- layer=2 filter=123 channel=51
					-13, -10, -10, 2, -3, -9, -8, -12, 1,
					-- layer=2 filter=123 channel=52
					-1, 6, -11, -1, -8, -3, -5, 4, -7,
					-- layer=2 filter=123 channel=53
					-7, 8, -8, 2, -10, -3, 7, 4, -7,
					-- layer=2 filter=123 channel=54
					-14, 0, -18, -7, -15, -2, 0, -2, -11,
					-- layer=2 filter=123 channel=55
					2, 4, -3, -9, -6, 2, 9, -5, 0,
					-- layer=2 filter=123 channel=56
					-14, 0, -13, -12, 3, -5, -2, -2, -3,
					-- layer=2 filter=123 channel=57
					2, -5, 8, 8, 7, 5, 9, -3, 6,
					-- layer=2 filter=123 channel=58
					-4, -7, -6, -3, 4, -10, -7, 0, 7,
					-- layer=2 filter=123 channel=59
					3, -11, -11, -5, -2, 2, -2, -9, -7,
					-- layer=2 filter=123 channel=60
					-11, -7, -1, -5, -15, 3, 4, 1, 0,
					-- layer=2 filter=123 channel=61
					-1, -12, 5, -4, -2, -12, 7, 1, 7,
					-- layer=2 filter=123 channel=62
					-1, -6, -2, -2, -4, 1, 0, 7, 3,
					-- layer=2 filter=123 channel=63
					-7, -11, -4, -9, -2, 2, 4, 5, -4,
					-- layer=2 filter=123 channel=64
					-1, 1, 7, -6, -3, 0, 8, -7, -8,
					-- layer=2 filter=123 channel=65
					1, -6, -6, 4, 1, -3, 0, 1, -10,
					-- layer=2 filter=123 channel=66
					8, -11, 6, 7, -10, -7, 0, -4, -3,
					-- layer=2 filter=123 channel=67
					1, -11, 4, -8, 6, -11, -6, -7, -1,
					-- layer=2 filter=123 channel=68
					9, 1, 1, -5, 0, -9, 0, -3, 2,
					-- layer=2 filter=123 channel=69
					1, -11, -10, 9, -11, 2, -11, -8, 4,
					-- layer=2 filter=123 channel=70
					-13, -7, -3, -5, 0, 3, -6, -9, -1,
					-- layer=2 filter=123 channel=71
					-12, 2, 4, -1, 4, -1, 10, -5, -6,
					-- layer=2 filter=123 channel=72
					-11, -13, 1, 9, 4, -5, 0, 6, 0,
					-- layer=2 filter=123 channel=73
					-7, -1, 6, 0, 4, 2, 10, 1, -7,
					-- layer=2 filter=123 channel=74
					-7, -4, -10, 7, -8, 3, 3, -7, -9,
					-- layer=2 filter=123 channel=75
					4, 2, -2, -4, 4, 1, 7, -9, 5,
					-- layer=2 filter=123 channel=76
					5, -10, 4, 5, 0, -10, 9, -4, -3,
					-- layer=2 filter=123 channel=77
					2, -1, 4, -9, 2, 8, -10, -11, -6,
					-- layer=2 filter=123 channel=78
					3, 6, 0, -8, -11, 6, -12, -2, -11,
					-- layer=2 filter=123 channel=79
					-4, 2, -2, -9, 3, 6, -6, -8, 5,
					-- layer=2 filter=123 channel=80
					-9, 6, -2, 3, -2, 0, -4, 2, 0,
					-- layer=2 filter=123 channel=81
					-1, -4, -3, 7, 0, 0, 7, 1, -1,
					-- layer=2 filter=123 channel=82
					7, 11, -7, 0, 7, 7, -11, -4, -3,
					-- layer=2 filter=123 channel=83
					7, 5, -4, 3, -2, 7, -10, -7, -9,
					-- layer=2 filter=123 channel=84
					7, 4, -9, 10, -5, 6, 7, 7, 6,
					-- layer=2 filter=123 channel=85
					-8, 3, 5, -6, 0, 8, 1, 4, 10,
					-- layer=2 filter=123 channel=86
					-7, -7, 3, 0, 7, -7, 6, -6, 4,
					-- layer=2 filter=123 channel=87
					7, -1, 2, 0, 4, 2, -10, 5, -8,
					-- layer=2 filter=123 channel=88
					2, 0, 5, 5, 0, -11, 2, 6, -7,
					-- layer=2 filter=123 channel=89
					-3, -2, -9, -6, 1, -6, -10, -8, -16,
					-- layer=2 filter=123 channel=90
					-3, -3, -2, 3, 5, -10, 6, -4, -1,
					-- layer=2 filter=123 channel=91
					-7, -12, -13, 1, 2, 0, -14, -16, -10,
					-- layer=2 filter=123 channel=92
					-2, 3, -3, -5, 5, 5, -14, 4, -6,
					-- layer=2 filter=123 channel=93
					-7, -14, 1, -8, -1, -11, -5, -1, -7,
					-- layer=2 filter=123 channel=94
					-9, 6, -3, -4, -9, -9, -9, -6, 6,
					-- layer=2 filter=123 channel=95
					-1, -11, -10, 6, -10, 4, 1, -4, 3,
					-- layer=2 filter=123 channel=96
					-4, -7, -9, -7, 2, -13, 14, 4, 0,
					-- layer=2 filter=123 channel=97
					-6, -8, -10, 1, 0, 4, -3, -3, 7,
					-- layer=2 filter=123 channel=98
					-7, 1, -2, 3, 0, -4, -14, 4, -6,
					-- layer=2 filter=123 channel=99
					-15, -1, 3, -14, 2, 0, 4, -7, -9,
					-- layer=2 filter=123 channel=100
					-10, 5, -5, -13, -9, 2, 0, -8, 3,
					-- layer=2 filter=123 channel=101
					-7, -16, -10, -4, -1, -18, -11, -2, 0,
					-- layer=2 filter=123 channel=102
					-3, -4, -2, -3, -7, -13, 10, 0, 0,
					-- layer=2 filter=123 channel=103
					-3, -3, -5, -9, 1, 6, -8, -5, 5,
					-- layer=2 filter=123 channel=104
					5, -11, 4, -11, 0, -15, 0, 1, 4,
					-- layer=2 filter=123 channel=105
					-2, 10, 8, -1, 13, 9, 8, -6, -6,
					-- layer=2 filter=123 channel=106
					-9, -22, -1, -19, -14, -11, -9, -19, 3,
					-- layer=2 filter=123 channel=107
					3, 0, -2, -4, 2, -9, -4, 0, -9,
					-- layer=2 filter=123 channel=108
					2, -12, -2, -7, 2, 0, 7, 1, -3,
					-- layer=2 filter=123 channel=109
					2, -8, 8, 1, -4, -1, -9, 2, 7,
					-- layer=2 filter=123 channel=110
					-5, 4, 1, -8, 5, 3, -13, -3, -5,
					-- layer=2 filter=123 channel=111
					8, -5, 8, -8, -4, 1, -4, -3, -2,
					-- layer=2 filter=123 channel=112
					-4, -5, 6, -6, -7, -2, -9, -1, -7,
					-- layer=2 filter=123 channel=113
					1, 5, -14, 2, -3, 4, -6, -5, -9,
					-- layer=2 filter=123 channel=114
					7, 8, 9, 0, 3, -6, 5, -2, -6,
					-- layer=2 filter=123 channel=115
					-4, -7, 5, 6, 6, 1, -11, 8, -7,
					-- layer=2 filter=123 channel=116
					8, -11, -11, 0, -9, -12, 1, -3, -7,
					-- layer=2 filter=123 channel=117
					-3, -11, -7, -7, -21, -6, -3, -4, -2,
					-- layer=2 filter=123 channel=118
					4, 3, 1, -8, -3, -4, 8, 7, -3,
					-- layer=2 filter=123 channel=119
					-9, -9, 0, -5, 6, -9, 2, -9, 6,
					-- layer=2 filter=123 channel=120
					2, 6, -1, 7, -2, -5, -9, 5, 5,
					-- layer=2 filter=123 channel=121
					-8, 12, 2, 4, -2, 7, -2, 7, 10,
					-- layer=2 filter=123 channel=122
					-7, -9, -6, -8, -2, 0, 5, 4, 10,
					-- layer=2 filter=123 channel=123
					-8, 0, 1, 6, 0, -2, -3, -3, 0,
					-- layer=2 filter=123 channel=124
					-6, -6, 1, -11, -5, -6, 0, 2, 0,
					-- layer=2 filter=123 channel=125
					6, 9, -9, 9, -10, 9, 11, 9, 0,
					-- layer=2 filter=123 channel=126
					-4, -10, -7, -3, 7, -8, 12, -7, -3,
					-- layer=2 filter=123 channel=127
					0, 0, -11, 2, -9, -6, -2, -6, 4,
					-- layer=2 filter=124 channel=0
					-5, 5, -6, -10, -11, -12, 6, -2, 5,
					-- layer=2 filter=124 channel=1
					-11, 0, -10, 0, -8, -1, 1, -18, -4,
					-- layer=2 filter=124 channel=2
					7, 0, -1, 2, 10, 11, -7, 7, 6,
					-- layer=2 filter=124 channel=3
					-9, -3, -9, -4, 4, -2, -6, -6, 5,
					-- layer=2 filter=124 channel=4
					-8, 3, -11, -8, -7, -7, -3, -10, -10,
					-- layer=2 filter=124 channel=5
					-7, 3, 3, -10, -5, -6, -3, 3, -6,
					-- layer=2 filter=124 channel=6
					10, 4, 1, -3, 0, 7, 7, 5, 22,
					-- layer=2 filter=124 channel=7
					-3, -21, 8, 3, 14, -14, 0, -5, -16,
					-- layer=2 filter=124 channel=8
					4, -2, 8, -1, -6, 4, 0, 4, -1,
					-- layer=2 filter=124 channel=9
					-8, 0, 0, -6, 7, 5, 1, -11, 8,
					-- layer=2 filter=124 channel=10
					-7, -12, -10, -9, -5, -9, -1, -10, -9,
					-- layer=2 filter=124 channel=11
					4, 7, 6, -16, -1, -5, 1, -5, -4,
					-- layer=2 filter=124 channel=12
					-6, -10, -17, -11, -5, -18, 0, -10, 6,
					-- layer=2 filter=124 channel=13
					-7, 0, 7, -12, 0, 10, -8, -5, -5,
					-- layer=2 filter=124 channel=14
					-16, -14, -16, 0, -2, -12, 3, -2, 0,
					-- layer=2 filter=124 channel=15
					-2, 0, 7, 4, 3, -10, -6, -4, -10,
					-- layer=2 filter=124 channel=16
					6, 8, 6, 3, 4, -8, 0, -10, -9,
					-- layer=2 filter=124 channel=17
					3, -8, -1, 2, 1, -8, 7, -8, 2,
					-- layer=2 filter=124 channel=18
					-16, 5, -14, -23, -5, -2, -6, 0, -6,
					-- layer=2 filter=124 channel=19
					-9, 0, -4, -10, -13, -15, -13, -4, -6,
					-- layer=2 filter=124 channel=20
					11, 0, -2, -6, 10, 9, -4, 9, 12,
					-- layer=2 filter=124 channel=21
					9, 1, -10, 1, -3, 0, 0, -4, 9,
					-- layer=2 filter=124 channel=22
					4, -3, 2, -6, 3, -8, -10, 4, 3,
					-- layer=2 filter=124 channel=23
					-5, -11, -7, -6, 1, -6, -16, -9, 0,
					-- layer=2 filter=124 channel=24
					-18, -1, -3, -10, -13, -4, 2, -8, -11,
					-- layer=2 filter=124 channel=25
					-9, 3, 0, -5, -15, -6, 8, -12, 0,
					-- layer=2 filter=124 channel=26
					-7, -4, -3, 9, -5, -7, 9, 7, 1,
					-- layer=2 filter=124 channel=27
					-10, -1, -15, -11, -15, -10, -14, -9, -8,
					-- layer=2 filter=124 channel=28
					-18, -14, 1, 8, -4, -14, -10, -12, -23,
					-- layer=2 filter=124 channel=29
					0, 2, 4, 1, -1, 9, 10, 0, 9,
					-- layer=2 filter=124 channel=30
					-9, 2, 2, -5, -3, -3, 6, 3, -6,
					-- layer=2 filter=124 channel=31
					-10, 2, -12, 3, -8, -1, -12, -6, -4,
					-- layer=2 filter=124 channel=32
					2, -1, 1, -9, 9, -4, 5, -9, -1,
					-- layer=2 filter=124 channel=33
					-8, -11, -9, 4, -5, 0, -15, -12, -4,
					-- layer=2 filter=124 channel=34
					-5, -13, 1, -1, -9, -5, -4, 4, -12,
					-- layer=2 filter=124 channel=35
					-21, -9, -13, 0, 0, -11, -9, 1, -15,
					-- layer=2 filter=124 channel=36
					-10, 4, -1, 7, -11, 5, 1, -6, 6,
					-- layer=2 filter=124 channel=37
					0, 6, -1, -13, -3, 0, -9, 6, -10,
					-- layer=2 filter=124 channel=38
					3, -26, -5, -20, -11, -18, -5, -17, 2,
					-- layer=2 filter=124 channel=39
					-9, 7, -6, -11, -4, -5, 4, -10, 0,
					-- layer=2 filter=124 channel=40
					-9, -2, -5, 8, 2, -14, -21, -9, -10,
					-- layer=2 filter=124 channel=41
					5, 3, 2, -2, 1, -5, 3, 11, 7,
					-- layer=2 filter=124 channel=42
					-13, 0, -3, -12, -6, -1, -14, 0, 1,
					-- layer=2 filter=124 channel=43
					-16, -14, 9, -1, 1, -12, -1, 0, -9,
					-- layer=2 filter=124 channel=44
					4, -4, 4, -4, -9, -1, 0, -4, -8,
					-- layer=2 filter=124 channel=45
					-7, 0, -6, 4, 0, -3, -13, 1, -1,
					-- layer=2 filter=124 channel=46
					-3, 0, -2, -6, 2, -9, -12, -11, -12,
					-- layer=2 filter=124 channel=47
					3, -10, 10, -4, -8, -19, -3, -9, -33,
					-- layer=2 filter=124 channel=48
					-1, 8, 6, 1, 3, -7, 9, 0, 11,
					-- layer=2 filter=124 channel=49
					-10, 4, -15, -6, -1, -2, -6, -13, 3,
					-- layer=2 filter=124 channel=50
					-10, -6, 2, -3, 5, 3, -9, -10, -7,
					-- layer=2 filter=124 channel=51
					-10, -6, -4, -16, -2, 4, -7, 0, 5,
					-- layer=2 filter=124 channel=52
					-3, -1, 3, -6, -8, 3, 0, -6, -9,
					-- layer=2 filter=124 channel=53
					4, 1, -13, -7, -1, -9, -16, -13, 7,
					-- layer=2 filter=124 channel=54
					-7, -20, -22, -31, -7, -6, -4, -24, -6,
					-- layer=2 filter=124 channel=55
					7, -2, 5, 3, -8, 13, 4, 1, 4,
					-- layer=2 filter=124 channel=56
					-2, -8, 7, -4, 5, 7, -3, 3, 0,
					-- layer=2 filter=124 channel=57
					-7, -5, 12, -1, -7, 2, 4, -4, -8,
					-- layer=2 filter=124 channel=58
					2, -17, -9, -2, -10, -15, -4, -16, -12,
					-- layer=2 filter=124 channel=59
					-13, -12, -11, -20, -11, 5, 0, -23, 0,
					-- layer=2 filter=124 channel=60
					0, -12, 0, -16, -29, 15, -4, -26, -2,
					-- layer=2 filter=124 channel=61
					5, -6, 6, -2, 1, 5, -3, -15, 5,
					-- layer=2 filter=124 channel=62
					-17, -7, 0, -9, -5, -12, 0, 2, 8,
					-- layer=2 filter=124 channel=63
					7, 0, -1, -15, -3, -6, -5, -8, 0,
					-- layer=2 filter=124 channel=64
					0, 2, -5, 0, -9, -1, -12, -6, -9,
					-- layer=2 filter=124 channel=65
					5, -13, -13, -10, -3, 8, -9, -11, -2,
					-- layer=2 filter=124 channel=66
					4, 5, -8, 8, -7, -9, 9, 3, -2,
					-- layer=2 filter=124 channel=67
					-11, -8, -1, -9, 0, 2, -4, -6, -5,
					-- layer=2 filter=124 channel=68
					-1, -10, -8, -7, -2, -2, 4, 0, -7,
					-- layer=2 filter=124 channel=69
					4, 1, 4, -6, 0, 0, 2, -2, -6,
					-- layer=2 filter=124 channel=70
					-18, -2, -12, -7, -6, -9, -9, 0, -13,
					-- layer=2 filter=124 channel=71
					-1, -10, 1, -10, -5, -2, -3, 1, 0,
					-- layer=2 filter=124 channel=72
					-13, 7, -8, -14, 0, -11, -13, -17, -22,
					-- layer=2 filter=124 channel=73
					-6, -22, -18, -15, -15, -22, 4, -31, -10,
					-- layer=2 filter=124 channel=74
					-5, -4, -11, -6, -8, -1, 6, 2, 1,
					-- layer=2 filter=124 channel=75
					-10, -11, 2, -1, -10, -6, -12, 6, -2,
					-- layer=2 filter=124 channel=76
					5, 0, 1, -5, -6, 2, -5, -7, -1,
					-- layer=2 filter=124 channel=77
					-2, 5, -9, 3, -5, -6, 1, -3, -1,
					-- layer=2 filter=124 channel=78
					0, -3, -2, -2, 7, 2, -7, -5, -4,
					-- layer=2 filter=124 channel=79
					-5, -3, 6, 5, 2, 0, 5, 7, 0,
					-- layer=2 filter=124 channel=80
					-12, -1, -6, 2, -6, -8, 2, -6, -7,
					-- layer=2 filter=124 channel=81
					-1, -3, -2, -4, 0, 6, -1, -3, 4,
					-- layer=2 filter=124 channel=82
					-1, -3, 2, -6, 2, -5, -6, 8, 0,
					-- layer=2 filter=124 channel=83
					-13, -2, 7, -13, 4, -7, 3, -1, 0,
					-- layer=2 filter=124 channel=84
					-5, -6, 7, 1, 11, 2, -3, -2, 4,
					-- layer=2 filter=124 channel=85
					5, -5, 6, -1, 10, 1, -7, -10, 9,
					-- layer=2 filter=124 channel=86
					-6, 8, -5, 9, 6, -7, 8, 5, 1,
					-- layer=2 filter=124 channel=87
					-11, -1, -3, 0, 19, 0, -15, -15, 10,
					-- layer=2 filter=124 channel=88
					6, -10, -16, 2, -6, 2, -6, -12, 2,
					-- layer=2 filter=124 channel=89
					-2, -9, 0, -6, -14, -13, 4, -8, -7,
					-- layer=2 filter=124 channel=90
					4, -7, 0, 8, 3, -7, 2, 7, -10,
					-- layer=2 filter=124 channel=91
					-19, -3, -22, -9, -23, -18, 2, -3, -11,
					-- layer=2 filter=124 channel=92
					-6, -10, -14, -2, -14, -6, -13, -21, -5,
					-- layer=2 filter=124 channel=93
					10, -11, 9, -9, -4, 6, 11, 0, 16,
					-- layer=2 filter=124 channel=94
					-5, 5, -3, -23, 4, -10, 1, -3, 12,
					-- layer=2 filter=124 channel=95
					-10, -11, -1, 1, 6, -8, -4, 6, 4,
					-- layer=2 filter=124 channel=96
					3, 7, -5, -15, -5, -5, -2, -8, 9,
					-- layer=2 filter=124 channel=97
					1, -2, 4, -9, 3, -9, -13, 0, -6,
					-- layer=2 filter=124 channel=98
					-11, -11, -9, 12, 0, -24, -21, -10, -27,
					-- layer=2 filter=124 channel=99
					-6, -2, 0, -1, 0, 8, -6, -6, -7,
					-- layer=2 filter=124 channel=100
					3, -14, -25, -7, -1, -12, 1, 2, -2,
					-- layer=2 filter=124 channel=101
					-9, -13, -6, -14, 0, -9, -3, -12, -14,
					-- layer=2 filter=124 channel=102
					-4, 0, -9, -7, -2, -4, -4, 0, -10,
					-- layer=2 filter=124 channel=103
					7, 1, 6, -3, 8, 1, 0, -5, 0,
					-- layer=2 filter=124 channel=104
					-1, 14, -8, -12, 0, -15, 7, -3, 6,
					-- layer=2 filter=124 channel=105
					1, -9, -9, 6, -2, 0, -11, 3, -5,
					-- layer=2 filter=124 channel=106
					-16, -8, -4, -5, -5, -14, -2, -8, -9,
					-- layer=2 filter=124 channel=107
					7, 2, -6, 1, -6, 5, 12, -5, 8,
					-- layer=2 filter=124 channel=108
					-13, -1, -9, -2, -10, -12, -6, 1, 0,
					-- layer=2 filter=124 channel=109
					7, 9, -5, 1, 10, 8, 10, 7, -1,
					-- layer=2 filter=124 channel=110
					-14, 1, -2, -7, -10, -12, -14, -16, 0,
					-- layer=2 filter=124 channel=111
					-8, 5, -7, 8, 8, 4, 4, 7, 0,
					-- layer=2 filter=124 channel=112
					8, 5, 6, -14, -12, -10, -7, -6, 6,
					-- layer=2 filter=124 channel=113
					6, -14, 0, -2, -12, 2, -10, -8, -8,
					-- layer=2 filter=124 channel=114
					3, -7, 10, 5, -8, -7, 3, -2, 7,
					-- layer=2 filter=124 channel=115
					8, 4, -9, -10, 9, -2, -1, 5, 3,
					-- layer=2 filter=124 channel=116
					-22, -14, -13, -17, 11, -8, -11, -7, -3,
					-- layer=2 filter=124 channel=117
					-13, -22, 1, -26, -17, -15, 0, -11, 3,
					-- layer=2 filter=124 channel=118
					0, 2, -4, -13, -6, 6, 5, -10, -14,
					-- layer=2 filter=124 channel=119
					-11, -3, -7, 0, -2, 2, -4, 6, -6,
					-- layer=2 filter=124 channel=120
					4, 10, -1, 0, 9, -7, -3, -1, 2,
					-- layer=2 filter=124 channel=121
					9, -8, 12, 6, 3, 2, 8, -5, 6,
					-- layer=2 filter=124 channel=122
					-6, -1, -10, 9, 1, 11, -5, -1, -10,
					-- layer=2 filter=124 channel=123
					-18, -12, -2, -6, -2, -1, -3, -9, -20,
					-- layer=2 filter=124 channel=124
					-7, -6, 10, 0, 3, -8, -9, -3, 14,
					-- layer=2 filter=124 channel=125
					8, 5, -6, -6, 0, -7, 0, 8, -9,
					-- layer=2 filter=124 channel=126
					9, -3, -5, -1, 6, -7, 5, -1, -8,
					-- layer=2 filter=124 channel=127
					5, -11, -11, 3, -15, 3, -14, -15, -10,
					-- layer=2 filter=125 channel=0
					-28, -20, -26, -18, -22, 8, 7, -6, -17,
					-- layer=2 filter=125 channel=1
					-16, -16, -38, -16, -26, -10, 5, -29, 16,
					-- layer=2 filter=125 channel=2
					11, -4, -5, -2, 2, 4, -3, 7, 9,
					-- layer=2 filter=125 channel=3
					-9, -6, 5, -14, -44, -5, -20, -12, -19,
					-- layer=2 filter=125 channel=4
					-14, -11, -3, 15, 12, 7, 3, 10, 11,
					-- layer=2 filter=125 channel=5
					-30, -6, -22, 6, 16, 1, 3, -7, 1,
					-- layer=2 filter=125 channel=6
					-14, 15, 5, -19, -3, -26, -58, 2, 21,
					-- layer=2 filter=125 channel=7
					20, -3, 9, 12, -16, -13, -24, -18, -14,
					-- layer=2 filter=125 channel=8
					-6, -1, 5, 1, 8, 0, 0, -4, 0,
					-- layer=2 filter=125 channel=9
					-43, -38, -22, -7, -26, -14, 3, 16, 3,
					-- layer=2 filter=125 channel=10
					-9, -16, -14, -5, -11, 22, 6, -16, -6,
					-- layer=2 filter=125 channel=11
					-2, -1, -20, -6, -11, -21, -3, -27, -28,
					-- layer=2 filter=125 channel=12
					0, -14, -56, -16, -21, 0, 0, 0, -1,
					-- layer=2 filter=125 channel=13
					8, 7, -9, 5, -1, -7, 7, 11, 11,
					-- layer=2 filter=125 channel=14
					-17, -14, -77, -19, -42, -30, -12, -22, -27,
					-- layer=2 filter=125 channel=15
					44, 14, -41, 6, -14, 10, -17, -14, -28,
					-- layer=2 filter=125 channel=16
					-41, -35, -42, 6, -11, -34, -29, -31, -16,
					-- layer=2 filter=125 channel=17
					-6, 0, 3, 6, 0, 7, -8, 9, -3,
					-- layer=2 filter=125 channel=18
					-7, 5, 7, 14, -10, -31, -8, -9, 2,
					-- layer=2 filter=125 channel=19
					-5, -9, -19, -9, -32, -3, -27, -27, -9,
					-- layer=2 filter=125 channel=20
					-7, 0, 12, 6, 3, 5, 0, 1, 8,
					-- layer=2 filter=125 channel=21
					2, -6, 0, 0, 9, 2, 8, -3, -3,
					-- layer=2 filter=125 channel=22
					8, 5, 6, -8, 5, 2, 2, -8, 4,
					-- layer=2 filter=125 channel=23
					-4, -7, -18, -17, -28, -20, -6, -25, -40,
					-- layer=2 filter=125 channel=24
					-22, -37, -49, -14, -26, -39, 0, -32, -37,
					-- layer=2 filter=125 channel=25
					-18, 0, -34, -5, -29, -33, -12, -17, -32,
					-- layer=2 filter=125 channel=26
					5, 3, 4, 3, 0, -5, -3, 0, 2,
					-- layer=2 filter=125 channel=27
					-3, 2, -6, -5, 3, 32, 8, 5, 16,
					-- layer=2 filter=125 channel=28
					-22, 25, 48, 30, 30, -27, -23, -28, -14,
					-- layer=2 filter=125 channel=29
					4, 0, 3, 10, 2, 9, -2, 0, -4,
					-- layer=2 filter=125 channel=30
					-30, 16, -35, 0, 5, 4, 0, 4, -13,
					-- layer=2 filter=125 channel=31
					27, -19, -15, 3, -2, -17, -12, -20, -16,
					-- layer=2 filter=125 channel=32
					6, -1, 7, -9, 12, 1, -12, 4, -3,
					-- layer=2 filter=125 channel=33
					12, 17, 2, -2, -23, -2, 6, 10, 4,
					-- layer=2 filter=125 channel=34
					-46, 19, 17, 22, -5, 7, -10, -31, 8,
					-- layer=2 filter=125 channel=35
					-19, 13, 27, 22, 0, -25, -7, -35, -2,
					-- layer=2 filter=125 channel=36
					-5, -5, 5, -9, -10, 4, -6, 0, 0,
					-- layer=2 filter=125 channel=37
					-11, -2, 2, -3, 1, 0, -5, 7, -7,
					-- layer=2 filter=125 channel=38
					-2, -29, -47, -18, -6, 11, 9, 23, 19,
					-- layer=2 filter=125 channel=39
					0, -28, -44, 15, -3, -4, -5, -5, 1,
					-- layer=2 filter=125 channel=40
					30, 45, -2, 9, -12, -13, 19, -8, -5,
					-- layer=2 filter=125 channel=41
					-6, 3, -3, -3, 4, 8, -8, 1, 11,
					-- layer=2 filter=125 channel=42
					-25, -28, -28, -23, -50, -48, 2, -40, -42,
					-- layer=2 filter=125 channel=43
					0, 8, 48, 44, 28, 26, -2, 0, 9,
					-- layer=2 filter=125 channel=44
					9, 7, 6, -11, -2, 0, 9, -4, -8,
					-- layer=2 filter=125 channel=45
					6, -13, -6, 12, 11, 15, -7, -5, 1,
					-- layer=2 filter=125 channel=46
					-35, -46, -42, -16, 7, 48, 41, 31, 24,
					-- layer=2 filter=125 channel=47
					-7, 25, 15, 26, -2, -4, -1, -7, -6,
					-- layer=2 filter=125 channel=48
					-2, 11, 1, 3, 2, -10, -8, 8, 2,
					-- layer=2 filter=125 channel=49
					3, -32, -28, -11, -36, -36, -17, -3, 4,
					-- layer=2 filter=125 channel=50
					-3, 2, 2, -3, -4, -5, 3, 2, 0,
					-- layer=2 filter=125 channel=51
					-4, 2, -25, -13, -1, -36, -8, -11, -33,
					-- layer=2 filter=125 channel=52
					8, 12, -37, -9, 0, -39, -10, -7, -2,
					-- layer=2 filter=125 channel=53
					11, -31, -6, 7, 25, -25, -9, 5, -35,
					-- layer=2 filter=125 channel=54
					-16, 15, -9, 11, -16, -25, -10, -21, -19,
					-- layer=2 filter=125 channel=55
					4, -11, -6, -4, 6, -2, 0, -9, -8,
					-- layer=2 filter=125 channel=56
					-22, 8, 25, 9, 18, -9, 0, 1, -10,
					-- layer=2 filter=125 channel=57
					-5, 1, -8, 4, 4, 7, -4, 9, -8,
					-- layer=2 filter=125 channel=58
					-9, 0, -59, -37, -22, 6, 12, 2, -6,
					-- layer=2 filter=125 channel=59
					27, -30, -42, -43, -23, 0, -20, 15, 10,
					-- layer=2 filter=125 channel=60
					-6, -39, -31, -21, -32, 0, -29, 18, -13,
					-- layer=2 filter=125 channel=61
					-1, -26, -18, -32, -30, -22, -25, 16, -4,
					-- layer=2 filter=125 channel=62
					-3, 5, 8, -15, -8, -24, -29, -22, 7,
					-- layer=2 filter=125 channel=63
					2, -21, -12, -32, 5, 13, -32, 9, -16,
					-- layer=2 filter=125 channel=64
					-56, -40, -50, -19, -42, -37, -13, -35, -26,
					-- layer=2 filter=125 channel=65
					-6, 7, -5, -14, -31, -3, -52, 14, 25,
					-- layer=2 filter=125 channel=66
					-8, -11, -8, 0, -14, 9, 8, -4, -18,
					-- layer=2 filter=125 channel=67
					-7, -50, -36, -23, 4, 4, 8, 23, -7,
					-- layer=2 filter=125 channel=68
					2, 0, -7, 9, -5, -1, -8, -3, 4,
					-- layer=2 filter=125 channel=69
					-51, -43, -29, -25, -49, -52, -26, -34, -10,
					-- layer=2 filter=125 channel=70
					-27, 23, 38, 34, 18, 0, 7, -12, 13,
					-- layer=2 filter=125 channel=71
					-27, -8, -33, -23, -5, -1, -28, -15, -17,
					-- layer=2 filter=125 channel=72
					-14, 6, 9, -12, -33, -54, -32, -10, -32,
					-- layer=2 filter=125 channel=73
					5, -16, -50, -8, -18, -50, -13, -25, -8,
					-- layer=2 filter=125 channel=74
					-19, -36, -30, -16, -1, 21, 12, 22, 24,
					-- layer=2 filter=125 channel=75
					6, -13, 8, -28, 2, 0, -32, -7, -16,
					-- layer=2 filter=125 channel=76
					47, -21, -16, 20, 2, -11, -23, -12, 14,
					-- layer=2 filter=125 channel=77
					0, -7, 6, -2, -9, -4, 4, 8, -10,
					-- layer=2 filter=125 channel=78
					7, -10, -13, 3, -26, -48, -19, -36, -34,
					-- layer=2 filter=125 channel=79
					6, -2, 8, 2, 0, 8, -7, 11, -1,
					-- layer=2 filter=125 channel=80
					-15, -36, -29, -7, 13, 6, 1, 7, 8,
					-- layer=2 filter=125 channel=81
					6, -7, 0, 4, 5, 0, 2, -2, -6,
					-- layer=2 filter=125 channel=82
					-7, 5, 1, 2, 1, 9, 7, 11, -1,
					-- layer=2 filter=125 channel=83
					-29, -11, -8, 22, -4, -35, 1, 4, -12,
					-- layer=2 filter=125 channel=84
					4, 1, 7, 2, 8, -6, -9, 11, -3,
					-- layer=2 filter=125 channel=85
					3, -1, 1, 4, -2, -11, -11, 6, 0,
					-- layer=2 filter=125 channel=86
					-5, 6, 1, 10, -8, -8, -9, -11, 6,
					-- layer=2 filter=125 channel=87
					4, 1, 19, 4, 0, -25, -23, 9, -23,
					-- layer=2 filter=125 channel=88
					-35, -53, -20, -5, -24, -15, -13, -18, 2,
					-- layer=2 filter=125 channel=89
					-16, -4, -73, -15, -50, -38, -34, -21, -29,
					-- layer=2 filter=125 channel=90
					1, -9, 4, -10, -3, 2, 5, 0, 3,
					-- layer=2 filter=125 channel=91
					-14, -25, -30, 1, -42, -21, -19, -26, -18,
					-- layer=2 filter=125 channel=92
					-13, -4, -63, -8, -38, -24, -6, -22, -9,
					-- layer=2 filter=125 channel=93
					-23, 4, 26, -14, -22, 22, -34, 7, 5,
					-- layer=2 filter=125 channel=94
					-6, 1, -6, -44, 12, -27, -27, 0, -10,
					-- layer=2 filter=125 channel=95
					3, -2, 2, -8, 6, -3, -4, 6, -11,
					-- layer=2 filter=125 channel=96
					-2, 49, -6, -3, 14, -38, -27, 4, -16,
					-- layer=2 filter=125 channel=97
					-27, -45, 4, -32, -13, -10, -13, -22, -17,
					-- layer=2 filter=125 channel=98
					-7, 20, 28, 16, 3, 3, -3, 0, -6,
					-- layer=2 filter=125 channel=99
					4, -12, -35, -24, -59, -8, -49, -9, 5,
					-- layer=2 filter=125 channel=100
					2, 2, -35, 24, 7, 31, 25, 41, 50,
					-- layer=2 filter=125 channel=101
					-10, 25, -5, 25, -17, -10, 2, -29, -23,
					-- layer=2 filter=125 channel=102
					-21, 14, -8, -16, -34, -46, -15, -8, -4,
					-- layer=2 filter=125 channel=103
					-2, 8, 4, -5, -28, 10, 7, 9, -4,
					-- layer=2 filter=125 channel=104
					-7, -22, -15, 0, -13, -18, -4, -10, 9,
					-- layer=2 filter=125 channel=105
					16, 1, 25, 12, -35, -19, 6, -5, -4,
					-- layer=2 filter=125 channel=106
					12, -37, -14, -20, -22, -27, -14, -20, -37,
					-- layer=2 filter=125 channel=107
					0, -16, -24, -7, 8, 12, 2, -27, 12,
					-- layer=2 filter=125 channel=108
					-26, -31, -36, -18, -19, -14, -29, 2, -4,
					-- layer=2 filter=125 channel=109
					-1, 3, -1, 1, -6, -9, -5, -4, -10,
					-- layer=2 filter=125 channel=110
					-37, -47, -37, -22, -24, -63, -24, -39, -55,
					-- layer=2 filter=125 channel=111
					-1, -8, 0, -4, -6, -8, 0, 1, 3,
					-- layer=2 filter=125 channel=112
					-24, -37, -19, -8, 0, 10, -7, -4, 11,
					-- layer=2 filter=125 channel=113
					-5, -5, -14, -7, -7, -37, -1, -12, 1,
					-- layer=2 filter=125 channel=114
					5, -3, 3, 5, 11, -6, 1, -8, 8,
					-- layer=2 filter=125 channel=115
					4, 0, 9, 3, 0, -9, -4, -1, 0,
					-- layer=2 filter=125 channel=116
					-6, 7, -6, 0, 2, -36, -12, 22, -6,
					-- layer=2 filter=125 channel=117
					3, -12, -3, 18, -22, -4, -44, -24, -42,
					-- layer=2 filter=125 channel=118
					9, 4, 28, 3, -11, 5, -5, -10, -11,
					-- layer=2 filter=125 channel=119
					5, 12, 14, 24, -3, 11, -24, -28, 30,
					-- layer=2 filter=125 channel=120
					0, 0, 0, 0, -3, -10, 1, 6, -10,
					-- layer=2 filter=125 channel=121
					3, -6, -8, 2, 10, 8, 6, 7, 0,
					-- layer=2 filter=125 channel=122
					8, 5, -9, 8, 5, -3, 4, 5, 8,
					-- layer=2 filter=125 channel=123
					11, 0, 15, -17, -30, -24, -32, -1, -22,
					-- layer=2 filter=125 channel=124
					31, -6, -24, -26, -35, 3, -11, -11, -30,
					-- layer=2 filter=125 channel=125
					7, -3, -2, -4, 1, 8, -6, 0, 4,
					-- layer=2 filter=125 channel=126
					-6, 15, -19, -22, 4, -27, -15, 3, -10,
					-- layer=2 filter=125 channel=127
					-23, -7, -47, -12, -7, -44, -21, -30, -3,
					-- layer=2 filter=126 channel=0
					-59, 0, -21, -16, -34, -56, 0, -11, -54,
					-- layer=2 filter=126 channel=1
					-10, -8, 36, -12, 13, 9, -8, -23, -22,
					-- layer=2 filter=126 channel=2
					-8, -4, -5, -3, 6, -11, -6, -4, -7,
					-- layer=2 filter=126 channel=3
					27, 28, -30, 48, 40, 3, -13, -6, 1,
					-- layer=2 filter=126 channel=4
					-13, 15, 37, -6, 1, -48, -36, -35, -87,
					-- layer=2 filter=126 channel=5
					-16, -14, -36, -9, 1, -14, 2, -43, -44,
					-- layer=2 filter=126 channel=6
					7, 19, -14, 15, -21, -2, -1, 22, -19,
					-- layer=2 filter=126 channel=7
					-1, -23, -54, -3, -11, -21, 11, -43, -27,
					-- layer=2 filter=126 channel=8
					6, -2, 6, 4, 10, 5, -5, 8, -9,
					-- layer=2 filter=126 channel=9
					-25, -23, -41, 23, -4, -12, -2, -6, 7,
					-- layer=2 filter=126 channel=10
					37, -7, 7, -5, -8, -42, -33, -19, -4,
					-- layer=2 filter=126 channel=11
					-2, -16, -30, 13, -26, -10, 0, -24, -11,
					-- layer=2 filter=126 channel=12
					-17, -27, 30, -19, 25, 24, -31, -26, -10,
					-- layer=2 filter=126 channel=13
					7, -5, 0, 3, -7, -7, -4, 4, 8,
					-- layer=2 filter=126 channel=14
					-23, -52, 20, -35, -6, -14, -28, -17, -34,
					-- layer=2 filter=126 channel=15
					81, 22, 23, 23, 41, -10, 4, 0, -21,
					-- layer=2 filter=126 channel=16
					-52, -2, 40, -29, -38, 46, -15, -26, 42,
					-- layer=2 filter=126 channel=17
					-6, 1, 8, -9, -5, -10, 3, -3, 4,
					-- layer=2 filter=126 channel=18
					17, 6, 4, 3, 9, -33, -26, -26, -100,
					-- layer=2 filter=126 channel=19
					27, -16, 30, 0, 25, 19, 20, 36, 31,
					-- layer=2 filter=126 channel=20
					0, 0, 2, 0, 1, 5, -6, -10, -4,
					-- layer=2 filter=126 channel=21
					-8, 8, 6, -6, -5, 9, -2, 12, -7,
					-- layer=2 filter=126 channel=22
					0, 2, 10, -1, -4, -3, 3, -7, -8,
					-- layer=2 filter=126 channel=23
					-13, -8, 0, -27, 16, -4, -20, -39, -56,
					-- layer=2 filter=126 channel=24
					2, 2, 4, -12, 1, 36, 2, 14, 50,
					-- layer=2 filter=126 channel=25
					0, 0, 32, -3, -15, 17, 9, 11, 39,
					-- layer=2 filter=126 channel=26
					3, -6, 9, 0, 3, -7, -5, -10, 10,
					-- layer=2 filter=126 channel=27
					-21, -16, -8, -50, -30, 5, -55, -43, -22,
					-- layer=2 filter=126 channel=28
					15, -29, -49, -47, -8, -61, -50, -62, -49,
					-- layer=2 filter=126 channel=29
					0, -3, -3, 1, 1, 8, 0, -8, -10,
					-- layer=2 filter=126 channel=30
					-2, -17, -11, 13, -30, 21, -11, -57, -29,
					-- layer=2 filter=126 channel=31
					3, 26, -43, -1, 87, -18, 22, 54, 23,
					-- layer=2 filter=126 channel=32
					5, 3, 0, -10, -7, 0, -3, -6, -7,
					-- layer=2 filter=126 channel=33
					24, -36, 2, -34, -27, -28, -59, -57, -26,
					-- layer=2 filter=126 channel=34
					-1, 16, -2, 53, 5, 21, 22, 17, 18,
					-- layer=2 filter=126 channel=35
					-19, -25, 8, -26, -37, -36, -57, -63, -64,
					-- layer=2 filter=126 channel=36
					4, -2, 3, 7, 7, 3, 7, 2, -6,
					-- layer=2 filter=126 channel=37
					-12, -22, -29, 31, -7, -36, 3, -17, -9,
					-- layer=2 filter=126 channel=38
					-15, -66, -26, -57, -38, 24, -44, -63, -9,
					-- layer=2 filter=126 channel=39
					-22, -51, -1, -14, -3, 8, -42, -49, -2,
					-- layer=2 filter=126 channel=40
					11, 6, 82, 4, -3, 22, -47, -16, 15,
					-- layer=2 filter=126 channel=41
					-2, -2, 9, 0, 2, -5, 3, 3, -3,
					-- layer=2 filter=126 channel=42
					-21, -3, 42, 2, 37, 35, -18, 21, 6,
					-- layer=2 filter=126 channel=43
					18, -17, -3, 41, -10, -89, -27, -24, -76,
					-- layer=2 filter=126 channel=44
					5, 3, -4, -7, -4, 0, 9, 7, -3,
					-- layer=2 filter=126 channel=45
					15, 14, 18, 0, 1, -29, -28, -11, -21,
					-- layer=2 filter=126 channel=46
					13, -70, 0, -9, -43, -27, -32, -63, -62,
					-- layer=2 filter=126 channel=47
					5, -35, -33, -29, 3, -90, -66, -71, -34,
					-- layer=2 filter=126 channel=48
					-10, 0, -9, 0, 0, 0, 4, 3, -1,
					-- layer=2 filter=126 channel=49
					13, 23, 38, 25, 23, -50, 27, 3, -44,
					-- layer=2 filter=126 channel=50
					18, 27, 15, 1, 8, -7, -8, 8, 24,
					-- layer=2 filter=126 channel=51
					-24, -28, -29, 7, -5, -11, 13, 3, -6,
					-- layer=2 filter=126 channel=52
					-5, -23, 7, 16, -21, -4, 30, 5, 0,
					-- layer=2 filter=126 channel=53
					4, 19, 31, -15, 16, -6, 7, 54, -15,
					-- layer=2 filter=126 channel=54
					-11, 3, 34, -5, 32, 0, 4, -19, -44,
					-- layer=2 filter=126 channel=55
					-8, 0, -8, 8, 2, 3, 7, 5, 2,
					-- layer=2 filter=126 channel=56
					-23, -62, -47, 18, -26, -11, -11, -51, -44,
					-- layer=2 filter=126 channel=57
					-8, 13, 0, 5, -12, 0, 4, 3, -3,
					-- layer=2 filter=126 channel=58
					-22, -28, 29, -26, 2, 15, -32, -4, -21,
					-- layer=2 filter=126 channel=59
					-18, -74, -1, -6, -15, -7, -39, 8, 15,
					-- layer=2 filter=126 channel=60
					4, 6, 9, -32, 13, 33, 20, 14, 62,
					-- layer=2 filter=126 channel=61
					-2, -8, -29, -19, -10, 22, 14, -9, 17,
					-- layer=2 filter=126 channel=62
					21, 25, -9, -3, 25, 14, 15, 28, -30,
					-- layer=2 filter=126 channel=63
					-33, -18, 5, -19, 14, -33, -11, -47, -34,
					-- layer=2 filter=126 channel=64
					-42, -10, 28, -24, -31, 37, -38, -2, 12,
					-- layer=2 filter=126 channel=65
					-6, -7, -15, 2, 1, 23, -6, 0, 21,
					-- layer=2 filter=126 channel=66
					-2, -19, 47, -5, -30, -24, -4, 7, -17,
					-- layer=2 filter=126 channel=67
					-2, -28, -31, -48, 4, -25, -43, -5, -31,
					-- layer=2 filter=126 channel=68
					5, -2, -1, -9, 0, 8, 6, -4, 8,
					-- layer=2 filter=126 channel=69
					-57, 7, 16, -21, -20, 26, -22, -9, -25,
					-- layer=2 filter=126 channel=70
					-13, -31, 7, -4, 6, -37, -26, -26, -56,
					-- layer=2 filter=126 channel=71
					7, -24, -38, -21, -22, 9, -40, -52, -41,
					-- layer=2 filter=126 channel=72
					39, -28, -16, -23, 26, 14, 32, -22, 7,
					-- layer=2 filter=126 channel=73
					59, 59, -27, 50, 19, 13, 61, 35, 8,
					-- layer=2 filter=126 channel=74
					11, -28, -16, 14, -23, -17, -55, -44, -15,
					-- layer=2 filter=126 channel=75
					59, 21, 27, 19, -16, 0, -47, 14, -8,
					-- layer=2 filter=126 channel=76
					-20, 62, 5, -12, 20, -58, -12, 44, -12,
					-- layer=2 filter=126 channel=77
					4, 4, 4, -10, -1, -6, -8, -7, -3,
					-- layer=2 filter=126 channel=78
					6, 0, -2, 17, -21, -22, 37, -2, -6,
					-- layer=2 filter=126 channel=79
					-2, 5, 4, 8, -11, -7, -6, 1, 1,
					-- layer=2 filter=126 channel=80
					12, 27, 15, 6, 29, 5, -7, 34, 23,
					-- layer=2 filter=126 channel=81
					-12, -2, 2, 5, -8, -5, 3, 4, -12,
					-- layer=2 filter=126 channel=82
					-3, -8, 6, -5, -3, -9, -6, -4, -2,
					-- layer=2 filter=126 channel=83
					-2, -10, 48, -35, 16, 37, -40, -42, -11,
					-- layer=2 filter=126 channel=84
					3, -6, 0, -9, 6, 7, 0, -7, -7,
					-- layer=2 filter=126 channel=85
					-1, 6, 12, -3, 8, 14, 0, 8, 3,
					-- layer=2 filter=126 channel=86
					10, 0, 7, -13, 0, 6, -2, 5, 12,
					-- layer=2 filter=126 channel=87
					33, 49, 10, 0, 35, -21, -19, 21, -53,
					-- layer=2 filter=126 channel=88
					-30, -6, 18, 1, -29, -1, -60, -50, -24,
					-- layer=2 filter=126 channel=89
					-2, -35, 9, -4, 8, -10, -27, -6, -12,
					-- layer=2 filter=126 channel=90
					-6, -2, 3, -1, 0, 8, -4, 3, -6,
					-- layer=2 filter=126 channel=91
					18, -27, 15, 21, 14, 29, -49, -29, 40,
					-- layer=2 filter=126 channel=92
					-15, -48, 10, -5, 30, 7, -46, 4, -2,
					-- layer=2 filter=126 channel=93
					25, 28, 47, 33, 8, -11, -10, 33, 32,
					-- layer=2 filter=126 channel=94
					3, 8, -33, -14, 15, -17, 31, 9, -38,
					-- layer=2 filter=126 channel=95
					-5, -9, -4, -6, 2, -12, -10, 4, -10,
					-- layer=2 filter=126 channel=96
					0, 45, 32, 36, -10, -34, 33, 3, -11,
					-- layer=2 filter=126 channel=97
					24, -2, -17, -23, -56, -42, -29, -22, -32,
					-- layer=2 filter=126 channel=98
					11, 5, -8, -22, 4, -24, -11, -49, -26,
					-- layer=2 filter=126 channel=99
					14, 1, -3, -8, -15, 11, 22, 22, 36,
					-- layer=2 filter=126 channel=100
					31, 6, 31, 2, -13, 27, -36, -23, 3,
					-- layer=2 filter=126 channel=101
					60, 7, -10, 24, -24, 14, -29, -17, 12,
					-- layer=2 filter=126 channel=102
					4, 32, 13, 58, -9, -35, 30, 4, -51,
					-- layer=2 filter=126 channel=103
					-31, 46, 11, -1, 96, 48, 37, -20, 56,
					-- layer=2 filter=126 channel=104
					1, 2, 17, -12, 56, -24, 25, 10, -77,
					-- layer=2 filter=126 channel=105
					20, -60, -1, -6, -48, -57, 29, -9, -36,
					-- layer=2 filter=126 channel=106
					48, 1, 5, -32, 5, 4, -43, -14, 56,
					-- layer=2 filter=126 channel=107
					59, 19, 22, -36, 70, -22, -47, 14, 61,
					-- layer=2 filter=126 channel=108
					-3, 2, -18, 30, -33, 16, -17, -39, -38,
					-- layer=2 filter=126 channel=109
					11, 13, -6, 14, -8, -11, 2, 8, -14,
					-- layer=2 filter=126 channel=110
					-42, -15, 42, -19, -10, 40, -48, 0, 27,
					-- layer=2 filter=126 channel=111
					-3, 0, -3, 7, -4, 4, 5, 10, -5,
					-- layer=2 filter=126 channel=112
					29, -23, -27, -37, 0, 4, -6, 2, 26,
					-- layer=2 filter=126 channel=113
					-24, -41, 4, -16, 18, 13, -19, -31, -13,
					-- layer=2 filter=126 channel=114
					13, -1, -3, 6, 4, -5, 1, -6, -3,
					-- layer=2 filter=126 channel=115
					-7, -9, -1, -2, 0, 9, -8, 0, 4,
					-- layer=2 filter=126 channel=116
					37, 49, 7, 11, 6, -16, 17, 2, -68,
					-- layer=2 filter=126 channel=117
					33, 20, 14, 6, 11, 4, 54, 8, -14,
					-- layer=2 filter=126 channel=118
					44, 31, -27, 64, 32, -45, 27, 28, -37,
					-- layer=2 filter=126 channel=119
					-16, 31, 8, -48, 5, -31, -56, -39, -48,
					-- layer=2 filter=126 channel=120
					-1, 2, -10, 8, -6, 2, 0, -10, -10,
					-- layer=2 filter=126 channel=121
					-1, -9, -7, 2, 5, -7, 7, -8, -10,
					-- layer=2 filter=126 channel=122
					0, -11, -4, 3, 11, 2, 3, 10, 4,
					-- layer=2 filter=126 channel=123
					24, -12, -24, -44, 0, -52, 33, -31, -28,
					-- layer=2 filter=126 channel=124
					37, 24, 40, 1, 45, 1, -8, 16, -58,
					-- layer=2 filter=126 channel=125
					-9, -1, -2, 1, -4, 9, -7, 0, -9,
					-- layer=2 filter=126 channel=126
					37, 0, 1, 36, 0, -4, 46, 23, 65,
					-- layer=2 filter=126 channel=127
					-43, -23, 17, 9, -5, 24, -84, -55, -31,
					-- layer=2 filter=127 channel=0
					1, 5, 15, -18, -38, -15, -6, -11, -18,
					-- layer=2 filter=127 channel=1
					27, 0, 16, 11, 28, 7, 13, 23, 11,
					-- layer=2 filter=127 channel=2
					-1, -9, -10, 8, -12, -3, -8, 3, 2,
					-- layer=2 filter=127 channel=3
					-21, 4, -3, -11, -43, -34, 25, 13, 17,
					-- layer=2 filter=127 channel=4
					0, 37, 4, -21, -11, -39, -25, -1, -23,
					-- layer=2 filter=127 channel=5
					13, -4, 7, -8, -31, 0, 0, -20, 1,
					-- layer=2 filter=127 channel=6
					-9, 7, 20, 33, 0, 40, -40, -5, 16,
					-- layer=2 filter=127 channel=7
					-29, -28, 15, 14, -8, -13, 5, 16, -4,
					-- layer=2 filter=127 channel=8
					-11, 7, -4, 0, -5, 2, 6, 0, 5,
					-- layer=2 filter=127 channel=9
					-5, -24, -68, -78, -75, -95, -55, -34, -37,
					-- layer=2 filter=127 channel=10
					-5, 30, 13, -35, -34, -13, 15, -25, -13,
					-- layer=2 filter=127 channel=11
					7, 4, -10, 17, 1, -5, 8, 0, 10,
					-- layer=2 filter=127 channel=12
					14, -2, 27, 14, 16, 26, 18, 31, 27,
					-- layer=2 filter=127 channel=13
					7, -2, 7, -5, 0, 1, -1, 8, 0,
					-- layer=2 filter=127 channel=14
					17, -3, -7, 10, 21, 15, 10, 36, 26,
					-- layer=2 filter=127 channel=15
					7, -33, 14, -54, -21, 11, -24, -74, 4,
					-- layer=2 filter=127 channel=16
					13, 33, 14, -2, 21, -28, 5, -36, -65,
					-- layer=2 filter=127 channel=17
					-3, 8, 3, -5, 0, 2, 8, 10, -3,
					-- layer=2 filter=127 channel=18
					-9, -49, -20, -8, -25, -38, -49, -46, -13,
					-- layer=2 filter=127 channel=19
					12, -10, 14, -3, 26, -2, 26, -1, 30,
					-- layer=2 filter=127 channel=20
					6, 0, 7, -10, 5, -1, -6, 6, 1,
					-- layer=2 filter=127 channel=21
					-3, 18, 8, 11, -1, -2, 21, 20, 6,
					-- layer=2 filter=127 channel=22
					2, -11, 4, -2, -9, 0, -1, -1, 4,
					-- layer=2 filter=127 channel=23
					-5, 29, 1, 17, 25, 2, 0, 5, 9,
					-- layer=2 filter=127 channel=24
					13, 0, -17, -5, -11, -16, 19, 12, 15,
					-- layer=2 filter=127 channel=25
					18, 0, -16, 6, 15, -9, 28, 26, 17,
					-- layer=2 filter=127 channel=26
					9, -2, 2, 8, -1, -6, -3, 8, 6,
					-- layer=2 filter=127 channel=27
					19, 30, 37, -16, -10, 27, -10, -22, -2,
					-- layer=2 filter=127 channel=28
					-21, -10, -17, -27, -31, -19, -18, -2, 22,
					-- layer=2 filter=127 channel=29
					-5, 2, -3, 7, -6, -9, 3, 7, -10,
					-- layer=2 filter=127 channel=30
					0, 0, -7, -40, -1, -13, -30, -44, -30,
					-- layer=2 filter=127 channel=31
					16, 9, -33, -14, -84, -11, 3, -20, -69,
					-- layer=2 filter=127 channel=32
					-6, -5, -4, -12, 1, 6, -5, 8, -4,
					-- layer=2 filter=127 channel=33
					-33, -27, 2, -42, -58, -32, -42, -33, -13,
					-- layer=2 filter=127 channel=34
					9, -20, -3, 6, 2, 21, -9, 3, 30,
					-- layer=2 filter=127 channel=35
					-27, -29, 5, -22, -24, -7, -18, -24, 20,
					-- layer=2 filter=127 channel=36
					-5, 3, 5, 6, 6, 2, 11, 17, -7,
					-- layer=2 filter=127 channel=37
					25, 0, 8, -8, 6, 17, 3, -8, -12,
					-- layer=2 filter=127 channel=38
					13, -18, 24, -3, -18, 3, -8, -42, -21,
					-- layer=2 filter=127 channel=39
					24, 38, 11, 4, -34, -24, 8, -27, -64,
					-- layer=2 filter=127 channel=40
					-52, -37, 17, -18, -6, -34, 36, -12, 20,
					-- layer=2 filter=127 channel=41
					-6, 3, 3, 6, 6, -8, 11, -2, 5,
					-- layer=2 filter=127 channel=42
					20, 15, -6, 7, 50, -16, 11, 18, -22,
					-- layer=2 filter=127 channel=43
					-25, -17, -19, -45, -46, -25, -56, -37, -6,
					-- layer=2 filter=127 channel=44
					-9, -7, 2, 3, -9, -1, 11, -2, -9,
					-- layer=2 filter=127 channel=45
					34, 46, 48, -22, -22, 46, -63, -18, -47,
					-- layer=2 filter=127 channel=46
					-10, 37, 16, -44, -29, -15, -71, -66, -48,
					-- layer=2 filter=127 channel=47
					-72, 16, 25, -56, -48, -46, -33, -19, 2,
					-- layer=2 filter=127 channel=48
					-4, -5, 7, 0, 3, 5, 10, -3, 0,
					-- layer=2 filter=127 channel=49
					21, -28, 0, 20, 0, -30, -2, -51, -42,
					-- layer=2 filter=127 channel=50
					-10, -4, 12, -15, -10, -11, -19, -3, -14,
					-- layer=2 filter=127 channel=51
					14, -7, -4, 6, -12, -17, 14, 6, -8,
					-- layer=2 filter=127 channel=52
					4, 2, 2, 9, 14, -2, 12, 5, 9,
					-- layer=2 filter=127 channel=53
					-21, -19, -9, -22, -59, -3, 1, -100, -32,
					-- layer=2 filter=127 channel=54
					-13, -7, 7, 35, 46, 15, 30, 33, 43,
					-- layer=2 filter=127 channel=55
					-14, 0, -7, -2, 3, -2, -2, 4, 5,
					-- layer=2 filter=127 channel=56
					10, -5, 4, -15, -11, 1, -8, -27, -19,
					-- layer=2 filter=127 channel=57
					0, 1, 12, -8, -7, 3, 4, -5, 2,
					-- layer=2 filter=127 channel=58
					3, 23, 16, 4, 10, 59, 32, 23, 34,
					-- layer=2 filter=127 channel=59
					14, 20, 14, -6, -8, 8, 27, -1, 17,
					-- layer=2 filter=127 channel=60
					9, -10, 11, 52, 6, 15, 46, 27, 20,
					-- layer=2 filter=127 channel=61
					-12, -16, -38, 45, -42, -32, 19, -11, -39,
					-- layer=2 filter=127 channel=62
					8, -7, -2, 32, 15, 14, -5, 1, 9,
					-- layer=2 filter=127 channel=63
					7, 36, 8, -18, 22, 21, -16, -15, -11,
					-- layer=2 filter=127 channel=64
					4, 29, 4, -36, 33, -2, -25, 19, 18,
					-- layer=2 filter=127 channel=65
					-2, -9, 1, 16, -30, -4, 0, -30, -9,
					-- layer=2 filter=127 channel=66
					13, 6, -33, -55, -16, -14, -28, 30, 5,
					-- layer=2 filter=127 channel=67
					-34, -22, -47, -90, -75, -81, -46, -47, -44,
					-- layer=2 filter=127 channel=68
					7, -6, -2, -6, -4, -7, 5, -3, 1,
					-- layer=2 filter=127 channel=69
					33, 26, -1, 4, 43, 6, -2, 33, -13,
					-- layer=2 filter=127 channel=70
					-3, -13, 8, -3, -14, 8, 7, -7, 28,
					-- layer=2 filter=127 channel=71
					12, 7, 5, -18, 1, 23, -25, 5, -7,
					-- layer=2 filter=127 channel=72
					4, -4, -7, 49, 16, -5, 21, 24, 36,
					-- layer=2 filter=127 channel=73
					25, 14, -33, -9, -43, -28, -33, -29, -34,
					-- layer=2 filter=127 channel=74
					-33, 10, -3, -40, -8, 5, -29, -11, -58,
					-- layer=2 filter=127 channel=75
					-12, -12, 3, -5, -13, 5, -44, -27, -12,
					-- layer=2 filter=127 channel=76
					-44, 1, -37, -47, -45, -62, -19, -45, -64,
					-- layer=2 filter=127 channel=77
					-5, 4, -6, 7, 0, -7, 7, -10, 8,
					-- layer=2 filter=127 channel=78
					-3, -22, -5, 3, 2, -16, 1, 6, -13,
					-- layer=2 filter=127 channel=79
					3, -7, 8, -9, 4, -10, 8, -9, -10,
					-- layer=2 filter=127 channel=80
					1, 48, 9, -36, 5, -12, -17, -32, -78,
					-- layer=2 filter=127 channel=81
					1, 1, 12, 6, -4, 9, -5, 0, -3,
					-- layer=2 filter=127 channel=82
					-6, -4, 5, 5, 4, -6, 11, -2, -10,
					-- layer=2 filter=127 channel=83
					21, 37, 26, -15, 9, 8, -19, -14, 6,
					-- layer=2 filter=127 channel=84
					-2, 7, 5, -1, -8, 8, 5, -1, -1,
					-- layer=2 filter=127 channel=85
					-6, 5, 11, 0, 3, -8, 8, 0, 1,
					-- layer=2 filter=127 channel=86
					-2, 6, -6, -14, -5, 15, 5, 1, 5,
					-- layer=2 filter=127 channel=87
					-20, 0, 33, 0, 10, -15, 15, -3, 8,
					-- layer=2 filter=127 channel=88
					8, 18, 42, -23, 14, 28, -36, 3, 11,
					-- layer=2 filter=127 channel=89
					1, -18, 9, -9, 5, 12, -2, 26, 33,
					-- layer=2 filter=127 channel=90
					3, 8, -9, -6, -10, -11, 2, 4, -1,
					-- layer=2 filter=127 channel=91
					-1, -4, -1, 20, 8, 24, 3, -2, 22,
					-- layer=2 filter=127 channel=92
					22, 20, 25, 3, 12, 11, 7, 16, 11,
					-- layer=2 filter=127 channel=93
					-50, -28, -38, -9, -11, -22, -41, 16, 2,
					-- layer=2 filter=127 channel=94
					-28, -24, -58, 43, -13, -25, 37, 14, 3,
					-- layer=2 filter=127 channel=95
					-4, 6, 1, 17, 12, 9, 14, 7, -2,
					-- layer=2 filter=127 channel=96
					-2, -17, 6, 27, 13, 17, 47, 43, 31,
					-- layer=2 filter=127 channel=97
					-6, 12, -11, -61, -29, -52, -49, -49, -54,
					-- layer=2 filter=127 channel=98
					-11, 23, 23, 25, 12, 3, 0, 29, 21,
					-- layer=2 filter=127 channel=99
					0, 32, 2, 9, 32, 23, 35, 25, 25,
					-- layer=2 filter=127 channel=100
					4, -9, 19, -30, -40, -15, 14, -15, -11,
					-- layer=2 filter=127 channel=101
					-10, -1, -15, 3, 7, 0, 1, 11, 4,
					-- layer=2 filter=127 channel=102
					20, -17, -28, -13, -7, -74, 16, 47, -17,
					-- layer=2 filter=127 channel=103
					5, -58, -17, -24, -1, -50, -13, 9, 21,
					-- layer=2 filter=127 channel=104
					7, -56, 15, 9, -18, -39, 12, -60, -28,
					-- layer=2 filter=127 channel=105
					-50, 51, 8, 5, 32, 30, 14, -18, -34,
					-- layer=2 filter=127 channel=106
					-11, -5, -34, 6, -11, 6, 20, 9, -10,
					-- layer=2 filter=127 channel=107
					-49, -14, -21, -1, 11, -54, 6, -9, -14,
					-- layer=2 filter=127 channel=108
					22, 2, -5, 0, 2, -6, 7, 14, -24,
					-- layer=2 filter=127 channel=109
					0, 2, -5, 10, -2, -9, -4, -11, -3,
					-- layer=2 filter=127 channel=110
					18, 0, -6, -2, 28, 8, 9, 22, 29,
					-- layer=2 filter=127 channel=111
					-1, 2, 0, 9, -11, 5, 0, 6, -5,
					-- layer=2 filter=127 channel=112
					-10, -10, -7, 8, -44, -56, 5, -9, -19,
					-- layer=2 filter=127 channel=113
					-2, 15, -6, 10, 15, 39, 0, -37, 0,
					-- layer=2 filter=127 channel=114
					1, -11, 8, 8, 18, -6, -1, -2, -3,
					-- layer=2 filter=127 channel=115
					-5, 4, -8, 0, -2, 13, 4, -3, 3,
					-- layer=2 filter=127 channel=116
					-23, -23, 1, -4, -24, -27, 9, -12, 6,
					-- layer=2 filter=127 channel=117
					0, -53, -1, 42, 26, -9, 30, 47, -6,
					-- layer=2 filter=127 channel=118
					31, 50, 39, -33, -26, -16, -50, -45, -32,
					-- layer=2 filter=127 channel=119
					-10, 0, -28, 8, -16, -41, -72, -23, 10,
					-- layer=2 filter=127 channel=120
					8, -8, -5, -3, -7, 0, 6, 8, 10,
					-- layer=2 filter=127 channel=121
					0, 6, 5, 1, 4, -5, -5, -3, 4,
					-- layer=2 filter=127 channel=122
					17, -9, 6, -5, 0, -11, 4, 1, -9,
					-- layer=2 filter=127 channel=123
					11, 28, 8, 34, 3, -15, 9, 12, 4,
					-- layer=2 filter=127 channel=124
					-56, -30, 16, -44, -37, -2, -30, 4, 21,
					-- layer=2 filter=127 channel=125
					8, 0, -1, 3, -8, -10, 3, 4, -12,
					-- layer=2 filter=127 channel=126
					3, -20, -98, -77, -75, -78, -44, -23, -13,
					-- layer=2 filter=127 channel=127
					13, 19, 12, 12, 8, 12, 13, 10, -2,
					-- layer=2 filter=128 channel=0
					-4, 7, -11, 8, 7, -11, 5, -3, 6,
					-- layer=2 filter=128 channel=1
					3, -11, 5, -6, -15, 2, -7, -14, -10,
					-- layer=2 filter=128 channel=2
					-2, 1, 5, 0, 4, -1, 8, 0, -1,
					-- layer=2 filter=128 channel=3
					10, 0, -1, -4, -10, -5, -10, -11, 0,
					-- layer=2 filter=128 channel=4
					-1, -7, -7, -2, 2, -7, -3, 0, -6,
					-- layer=2 filter=128 channel=5
					5, -2, -4, -5, 3, -9, -9, 0, 4,
					-- layer=2 filter=128 channel=6
					-10, -8, -7, -5, 0, 7, -3, 0, 4,
					-- layer=2 filter=128 channel=7
					-6, -8, -3, 0, 1, -8, 3, -4, -10,
					-- layer=2 filter=128 channel=8
					-8, 7, -5, -8, -8, 9, 5, 2, -2,
					-- layer=2 filter=128 channel=9
					-4, -8, 7, -11, 0, -4, -7, 7, -10,
					-- layer=2 filter=128 channel=10
					-7, -11, -4, -6, -2, 6, -1, -7, 6,
					-- layer=2 filter=128 channel=11
					-14, -12, -13, -3, 1, -5, 1, -16, -7,
					-- layer=2 filter=128 channel=12
					-10, 3, 0, -8, -3, -3, -11, 0, 3,
					-- layer=2 filter=128 channel=13
					7, 0, 0, 7, 2, -8, 0, 9, -4,
					-- layer=2 filter=128 channel=14
					3, 8, -10, -2, 7, 7, -3, -9, -2,
					-- layer=2 filter=128 channel=15
					-11, -4, 7, -4, -11, 2, -1, -6, -4,
					-- layer=2 filter=128 channel=16
					-5, -6, -1, 0, -6, -1, -1, 0, 0,
					-- layer=2 filter=128 channel=17
					4, 8, 6, -10, -6, 5, 6, 9, -7,
					-- layer=2 filter=128 channel=18
					6, -12, 3, 2, -10, -15, -4, -10, -11,
					-- layer=2 filter=128 channel=19
					-1, 1, 1, 2, -11, 5, 0, 0, -2,
					-- layer=2 filter=128 channel=20
					-3, 0, 8, 7, -6, -10, -4, -6, 3,
					-- layer=2 filter=128 channel=21
					-6, -7, 8, -1, -6, -3, -4, 1, -2,
					-- layer=2 filter=128 channel=22
					1, -1, -1, -8, -8, 8, 1, -9, 6,
					-- layer=2 filter=128 channel=23
					6, -12, 3, -2, -12, 1, 1, 4, -8,
					-- layer=2 filter=128 channel=24
					3, -11, 0, -12, 6, 5, -10, -12, 4,
					-- layer=2 filter=128 channel=25
					-4, -11, -10, 8, 1, -6, 0, -11, -10,
					-- layer=2 filter=128 channel=26
					9, 6, -2, -1, 7, -2, -5, -9, -2,
					-- layer=2 filter=128 channel=27
					5, -12, 2, 0, 0, -2, 0, 1, -6,
					-- layer=2 filter=128 channel=28
					-8, -2, -6, -1, 2, -14, 2, -5, 0,
					-- layer=2 filter=128 channel=29
					-1, 4, 7, -4, 0, 5, 6, -5, 8,
					-- layer=2 filter=128 channel=30
					2, 1, -6, -9, -4, -4, 8, -8, 0,
					-- layer=2 filter=128 channel=31
					0, 0, 8, -5, 9, 7, 0, -11, 8,
					-- layer=2 filter=128 channel=32
					-7, 3, -8, 8, 7, 6, -8, -6, 1,
					-- layer=2 filter=128 channel=33
					-12, -9, -8, 3, -5, 3, -3, -5, -4,
					-- layer=2 filter=128 channel=34
					-9, 5, 8, -12, 0, -6, 5, 2, 1,
					-- layer=2 filter=128 channel=35
					3, 5, -11, -1, 1, -4, 3, -3, -2,
					-- layer=2 filter=128 channel=36
					10, -1, -8, -12, -5, -10, -10, 0, 7,
					-- layer=2 filter=128 channel=37
					-4, -8, -1, -10, 6, 2, 0, 0, 2,
					-- layer=2 filter=128 channel=38
					1, -3, -10, 8, 2, 3, 0, 4, 2,
					-- layer=2 filter=128 channel=39
					4, -2, -10, 0, -2, -1, 8, -2, -12,
					-- layer=2 filter=128 channel=40
					5, -12, -2, 4, 4, 1, 6, 6, 12,
					-- layer=2 filter=128 channel=41
					1, -10, -4, -9, -9, 7, -1, 3, -11,
					-- layer=2 filter=128 channel=42
					-11, 7, 2, -3, -4, -10, -16, -1, -13,
					-- layer=2 filter=128 channel=43
					-1, -9, -8, -3, 7, -4, -9, -7, -12,
					-- layer=2 filter=128 channel=44
					3, 3, 6, -6, 4, -4, 1, 7, -6,
					-- layer=2 filter=128 channel=45
					-9, -3, -8, -11, 3, -3, -5, -10, -11,
					-- layer=2 filter=128 channel=46
					-2, -7, 7, -10, 0, -9, -10, 1, 4,
					-- layer=2 filter=128 channel=47
					-8, 7, -2, 1, -9, -4, 9, -13, 5,
					-- layer=2 filter=128 channel=48
					-8, -6, -5, 0, 5, 7, 6, 0, -8,
					-- layer=2 filter=128 channel=49
					1, 4, -5, -2, -12, 6, 1, 4, -10,
					-- layer=2 filter=128 channel=50
					4, -1, 4, -7, -5, -1, -5, -4, -7,
					-- layer=2 filter=128 channel=51
					1, -9, -6, 3, 0, 5, -12, -5, -2,
					-- layer=2 filter=128 channel=52
					-8, 0, 4, 0, 7, -5, 7, 1, -8,
					-- layer=2 filter=128 channel=53
					-9, 0, -2, 7, -2, -11, -12, 6, -13,
					-- layer=2 filter=128 channel=54
					-12, -18, -7, 0, -5, -4, -4, 0, -19,
					-- layer=2 filter=128 channel=55
					-8, -9, 8, 6, 1, 2, 1, -7, 10,
					-- layer=2 filter=128 channel=56
					0, -9, 7, -9, -4, 0, -8, -9, -3,
					-- layer=2 filter=128 channel=57
					-1, 6, 8, -8, -11, 3, 9, -10, 6,
					-- layer=2 filter=128 channel=58
					-13, -7, -3, -10, -6, -8, 5, 4, -13,
					-- layer=2 filter=128 channel=59
					0, -8, -1, 6, -10, -4, 0, -17, 1,
					-- layer=2 filter=128 channel=60
					3, -13, 3, 0, -12, -11, -3, 2, -9,
					-- layer=2 filter=128 channel=61
					0, -6, 0, -12, -2, -4, 7, -3, -9,
					-- layer=2 filter=128 channel=62
					7, 0, -13, -3, -1, -4, -5, -11, -2,
					-- layer=2 filter=128 channel=63
					-8, -7, -11, -7, -3, -5, 4, 6, 2,
					-- layer=2 filter=128 channel=64
					-5, -7, 2, 1, -2, 1, -11, -6, 4,
					-- layer=2 filter=128 channel=65
					7, 3, 0, -1, 3, -1, -13, 0, -3,
					-- layer=2 filter=128 channel=66
					5, 4, 2, -2, 7, -1, 0, -10, -9,
					-- layer=2 filter=128 channel=67
					0, -7, 0, -12, 1, 5, -12, -8, 3,
					-- layer=2 filter=128 channel=68
					7, -2, -8, -9, -1, -3, -8, 2, 7,
					-- layer=2 filter=128 channel=69
					4, -4, -14, 1, -12, -3, 3, -7, -1,
					-- layer=2 filter=128 channel=70
					10, 7, -4, -11, -5, -1, -1, 7, -5,
					-- layer=2 filter=128 channel=71
					-7, -7, 6, 5, 3, 2, -6, -4, 6,
					-- layer=2 filter=128 channel=72
					-10, 8, 2, -2, -9, -4, 8, 1, -2,
					-- layer=2 filter=128 channel=73
					-13, -8, -8, -9, 0, -3, -8, 3, 5,
					-- layer=2 filter=128 channel=74
					-2, -4, -8, 0, -9, -10, -8, -8, -5,
					-- layer=2 filter=128 channel=75
					0, 0, -2, -10, -4, 7, 6, -10, 3,
					-- layer=2 filter=128 channel=76
					9, 3, 6, -8, -3, -6, -2, -5, 1,
					-- layer=2 filter=128 channel=77
					6, 8, 0, -7, 3, 5, -10, -5, 1,
					-- layer=2 filter=128 channel=78
					-6, 1, 7, 1, 1, 6, -2, 0, 0,
					-- layer=2 filter=128 channel=79
					-7, -4, 1, -1, -3, -2, 5, -11, -2,
					-- layer=2 filter=128 channel=80
					-2, -9, 1, -7, 4, -5, -7, -2, 7,
					-- layer=2 filter=128 channel=81
					1, 2, -2, 0, -10, 0, -9, -7, -11,
					-- layer=2 filter=128 channel=82
					0, 4, 1, -10, -2, 0, -5, 6, 0,
					-- layer=2 filter=128 channel=83
					-2, -3, 7, 0, 5, 6, -11, -10, -4,
					-- layer=2 filter=128 channel=84
					2, -11, 6, -7, 0, 2, 0, 0, 8,
					-- layer=2 filter=128 channel=85
					0, 5, 0, 1, 5, 0, 3, 4, 6,
					-- layer=2 filter=128 channel=86
					2, -2, 2, -8, -5, -8, -4, -12, -10,
					-- layer=2 filter=128 channel=87
					-1, -3, 6, -10, 2, -9, -1, 2, 0,
					-- layer=2 filter=128 channel=88
					-7, -8, -10, -11, 0, 2, -4, 0, -7,
					-- layer=2 filter=128 channel=89
					0, -12, 0, 3, -9, -4, 7, -6, -13,
					-- layer=2 filter=128 channel=90
					-6, 1, -5, -9, 7, -2, 1, 1, -10,
					-- layer=2 filter=128 channel=91
					0, -1, -15, -7, -6, -10, -9, -2, 3,
					-- layer=2 filter=128 channel=92
					-5, -9, 0, 2, -4, -5, -11, 4, -8,
					-- layer=2 filter=128 channel=93
					-10, 3, -6, -3, 4, -5, -6, -16, -2,
					-- layer=2 filter=128 channel=94
					3, -2, -14, -3, -21, 6, -10, -20, 5,
					-- layer=2 filter=128 channel=95
					-5, -7, 1, 6, -6, -5, -1, -9, 4,
					-- layer=2 filter=128 channel=96
					-6, -12, 0, -9, 0, -7, -3, 0, -12,
					-- layer=2 filter=128 channel=97
					-8, -3, -10, 1, 8, 5, 0, 7, -5,
					-- layer=2 filter=128 channel=98
					4, 1, 7, -2, -12, 0, -7, 6, -5,
					-- layer=2 filter=128 channel=99
					-1, 1, -12, 3, -4, -9, -6, -16, -3,
					-- layer=2 filter=128 channel=100
					5, -7, -3, -11, -8, 8, 3, -10, -7,
					-- layer=2 filter=128 channel=101
					4, -5, 2, 8, -10, -8, -3, -8, 5,
					-- layer=2 filter=128 channel=102
					-13, 3, 0, -12, 4, -12, 0, -5, 5,
					-- layer=2 filter=128 channel=103
					-8, -2, -4, 6, 8, 0, -2, -8, -7,
					-- layer=2 filter=128 channel=104
					7, -12, -10, 9, -8, -4, 0, -3, -1,
					-- layer=2 filter=128 channel=105
					-5, -8, -3, 0, -4, 0, 1, 5, -11,
					-- layer=2 filter=128 channel=106
					5, -2, 6, 3, -8, 0, 2, -1, -7,
					-- layer=2 filter=128 channel=107
					-2, 2, -8, -1, -4, -9, -2, 2, 0,
					-- layer=2 filter=128 channel=108
					-8, -1, 5, -6, -1, 0, -11, -2, -4,
					-- layer=2 filter=128 channel=109
					7, -7, 0, -7, -2, -9, -4, 4, 4,
					-- layer=2 filter=128 channel=110
					-4, 5, 4, -7, -2, -16, -8, -9, 1,
					-- layer=2 filter=128 channel=111
					-4, 0, 1, 8, -7, 4, 11, -9, 0,
					-- layer=2 filter=128 channel=112
					-1, -11, -5, -6, 3, 1, -3, -12, -3,
					-- layer=2 filter=128 channel=113
					2, 2, -12, 5, -9, -16, -7, 4, -6,
					-- layer=2 filter=128 channel=114
					-2, -3, -8, 0, 5, 6, 0, -1, -3,
					-- layer=2 filter=128 channel=115
					5, -7, 0, -9, 1, -5, 2, -3, -8,
					-- layer=2 filter=128 channel=116
					1, 5, -14, 1, -7, -5, 4, -6, 0,
					-- layer=2 filter=128 channel=117
					10, -1, -1, -4, -5, -3, -1, -11, 3,
					-- layer=2 filter=128 channel=118
					-8, 2, -11, -10, -1, 0, 1, 4, -6,
					-- layer=2 filter=128 channel=119
					-5, 2, -4, 8, -8, 6, -1, 2, 0,
					-- layer=2 filter=128 channel=120
					-4, 8, 10, -8, 8, 3, -3, -6, 1,
					-- layer=2 filter=128 channel=121
					-9, 6, -2, -11, -8, 2, -5, 0, 6,
					-- layer=2 filter=128 channel=122
					7, 3, 3, -2, 1, 3, 0, -10, -3,
					-- layer=2 filter=128 channel=123
					-7, -1, 0, -3, -4, -4, -3, 4, 2,
					-- layer=2 filter=128 channel=124
					8, -10, -2, -5, 7, 0, -1, 5, -2,
					-- layer=2 filter=128 channel=125
					0, 1, 2, -10, -9, 10, -5, -8, -8,
					-- layer=2 filter=128 channel=126
					-9, -9, 9, 1, -4, -6, -9, 0, 7,
					-- layer=2 filter=128 channel=127
					-4, 7, 2, -13, 3, -11, -6, -7, -17,
					-- layer=2 filter=129 channel=0
					28, -11, -4, 31, 5, -33, 8, 12, -24,
					-- layer=2 filter=129 channel=1
					-5, 25, 21, -42, 5, 31, 18, -6, 10,
					-- layer=2 filter=129 channel=2
					-6, 0, 7, 9, 5, 3, 11, 5, -7,
					-- layer=2 filter=129 channel=3
					-4, 3, 1, 36, -2, -38, 7, 7, -53,
					-- layer=2 filter=129 channel=4
					-24, -39, 5, -21, -57, 14, -2, -42, -10,
					-- layer=2 filter=129 channel=5
					26, 1, -4, 27, -1, -21, 14, 2, 0,
					-- layer=2 filter=129 channel=6
					-26, 5, -43, -32, 25, -9, -14, -49, -48,
					-- layer=2 filter=129 channel=7
					-14, -7, -17, -25, 6, 37, -22, -8, 3,
					-- layer=2 filter=129 channel=8
					-1, 4, -3, 6, -3, -8, -4, -8, 0,
					-- layer=2 filter=129 channel=9
					-22, 11, 37, -11, -36, -32, -7, 7, -36,
					-- layer=2 filter=129 channel=10
					5, -1, 16, 15, 10, 3, 47, 21, 0,
					-- layer=2 filter=129 channel=11
					25, 9, -19, 14, 7, -7, 8, -17, -11,
					-- layer=2 filter=129 channel=12
					5, 40, -14, -60, 2, 42, -13, 17, 3,
					-- layer=2 filter=129 channel=13
					-11, -4, 4, -2, -6, 0, -6, -8, -10,
					-- layer=2 filter=129 channel=14
					-4, 16, -6, -9, -18, 31, -18, -4, 0,
					-- layer=2 filter=129 channel=15
					4, -5, 64, -84, 29, 12, -74, 16, -2,
					-- layer=2 filter=129 channel=16
					-41, -20, -5, -27, -66, 12, -69, -86, -15,
					-- layer=2 filter=129 channel=17
					6, 4, -3, 2, -3, 2, 6, -2, 3,
					-- layer=2 filter=129 channel=18
					35, -34, 11, -4, -41, 25, -8, -10, -6,
					-- layer=2 filter=129 channel=19
					25, 27, 35, -34, 3, 46, -21, -1, 10,
					-- layer=2 filter=129 channel=20
					2, -7, -9, 7, -10, -7, -6, 4, 1,
					-- layer=2 filter=129 channel=21
					17, 8, 19, 24, 28, 12, 0, 4, 6,
					-- layer=2 filter=129 channel=22
					4, 2, -10, 6, -3, 5, 1, 8, 0,
					-- layer=2 filter=129 channel=23
					-58, -26, 18, -20, 29, 11, -10, 15, 0,
					-- layer=2 filter=129 channel=24
					-26, 11, 18, 13, -19, -15, 28, -13, -17,
					-- layer=2 filter=129 channel=25
					14, 9, -2, -1, -17, 8, -4, -27, -28,
					-- layer=2 filter=129 channel=26
					5, 9, -3, 6, 9, -3, -4, 6, -6,
					-- layer=2 filter=129 channel=27
					8, 26, 26, 6, 6, 17, 31, 18, 10,
					-- layer=2 filter=129 channel=28
					5, 36, 6, -8, 7, -28, -37, 9, -4,
					-- layer=2 filter=129 channel=29
					4, -8, -1, 4, 3, -6, -12, -10, -6,
					-- layer=2 filter=129 channel=30
					-35, -18, 23, 10, -50, -2, 0, 1, 26,
					-- layer=2 filter=129 channel=31
					-26, -7, 39, -14, 6, -31, -23, 15, -35,
					-- layer=2 filter=129 channel=32
					-2, -8, 4, -4, 7, -10, -6, -8, 7,
					-- layer=2 filter=129 channel=33
					-25, -3, -48, -64, -19, -7, -68, -3, -1,
					-- layer=2 filter=129 channel=34
					65, -5, 1, -36, -12, 16, -45, 30, -4,
					-- layer=2 filter=129 channel=35
					38, 18, 8, -33, -10, -22, -42, 10, 11,
					-- layer=2 filter=129 channel=36
					7, -14, 0, 0, -2, -12, 8, 24, 4,
					-- layer=2 filter=129 channel=37
					2, 3, -3, 2, -9, -27, 5, 1, -17,
					-- layer=2 filter=129 channel=38
					-14, -1, 4, 6, -12, -2, 21, -11, 2,
					-- layer=2 filter=129 channel=39
					-66, 7, 16, -18, -58, -4, -37, 0, 35,
					-- layer=2 filter=129 channel=40
					18, 16, 63, -39, 49, -9, -17, 100, 13,
					-- layer=2 filter=129 channel=41
					-11, 0, 0, 7, -11, 4, -3, -7, -3,
					-- layer=2 filter=129 channel=42
					-42, 2, 17, -86, -22, 8, -21, 42, 39,
					-- layer=2 filter=129 channel=43
					22, 23, 6, 18, -37, -48, 5, -22, -33,
					-- layer=2 filter=129 channel=44
					-6, 4, 3, -8, 1, -6, -8, 5, 5,
					-- layer=2 filter=129 channel=45
					-33, 40, -11, -30, -47, -19, -35, -24, 10,
					-- layer=2 filter=129 channel=46
					15, -45, -31, -5, -19, 5, -13, 22, 7,
					-- layer=2 filter=129 channel=47
					-30, -16, -15, -52, 1, -23, -46, -17, -12,
					-- layer=2 filter=129 channel=48
					6, 0, -11, -3, -2, -6, -6, 2, -4,
					-- layer=2 filter=129 channel=49
					10, -29, 54, 0, -18, 35, -15, 18, -44,
					-- layer=2 filter=129 channel=50
					-27, -1, 12, 18, -23, -6, -16, 3, 14,
					-- layer=2 filter=129 channel=51
					39, 8, -24, 40, -6, -32, 20, 1, -27,
					-- layer=2 filter=129 channel=52
					54, 33, 7, 26, -4, -5, -34, -15, 0,
					-- layer=2 filter=129 channel=53
					-46, -44, -12, -20, -46, -20, -32, 30, 5,
					-- layer=2 filter=129 channel=54
					45, 34, 29, 0, 30, 19, -40, -28, 21,
					-- layer=2 filter=129 channel=55
					0, -8, 3, 2, -12, 3, 7, 6, -5,
					-- layer=2 filter=129 channel=56
					27, 5, -31, 19, 1, -32, 39, 12, -12,
					-- layer=2 filter=129 channel=57
					10, 2, 16, 8, 10, 9, 5, 3, -5,
					-- layer=2 filter=129 channel=58
					14, 65, 12, -73, 1, 20, 12, -8, 6,
					-- layer=2 filter=129 channel=59
					-29, -14, -24, -14, 55, 71, 8, -6, 41,
					-- layer=2 filter=129 channel=60
					54, -2, 27, 28, 47, 44, 7, 36, 50,
					-- layer=2 filter=129 channel=61
					31, -15, -8, 56, 36, -2, 13, 37, 30,
					-- layer=2 filter=129 channel=62
					0, -8, 16, -69, -9, -11, -28, 0, -28,
					-- layer=2 filter=129 channel=63
					-47, -29, 8, -31, -7, -8, -9, 4, 22,
					-- layer=2 filter=129 channel=64
					-37, 0, 29, -5, -42, 22, -6, 6, 24,
					-- layer=2 filter=129 channel=65
					20, -19, -28, 10, 17, 13, -22, 41, 29,
					-- layer=2 filter=129 channel=66
					55, -1, -11, -29, -20, -3, 43, 21, 10,
					-- layer=2 filter=129 channel=67
					5, 0, -13, -37, -45, -56, 12, 0, -22,
					-- layer=2 filter=129 channel=68
					-2, 6, -7, -6, -8, -2, 10, -3, -7,
					-- layer=2 filter=129 channel=69
					-32, 15, 31, -12, -19, 33, -24, 9, 28,
					-- layer=2 filter=129 channel=70
					41, 43, 4, 1, 7, -15, -36, 20, -6,
					-- layer=2 filter=129 channel=71
					6, 14, -9, 17, 3, 12, 17, 25, -1,
					-- layer=2 filter=129 channel=72
					-26, 29, -1, -23, 17, 20, -12, 13, 4,
					-- layer=2 filter=129 channel=73
					6, 30, -4, -7, -10, -42, 9, 11, -7,
					-- layer=2 filter=129 channel=74
					-23, 11, 25, -26, 12, -9, 19, -17, 15,
					-- layer=2 filter=129 channel=75
					-66, -32, -47, -60, -35, -25, -67, -34, -11,
					-- layer=2 filter=129 channel=76
					41, 6, 29, -33, 13, -76, -11, 11, 0,
					-- layer=2 filter=129 channel=77
					-1, -5, -4, -5, -5, -4, 8, -7, -6,
					-- layer=2 filter=129 channel=78
					40, 5, 24, -3, -1, -17, -8, -32, -28,
					-- layer=2 filter=129 channel=79
					1, -3, 4, 1, 1, 7, -10, 8, -5,
					-- layer=2 filter=129 channel=80
					-10, -6, 27, -39, -20, 17, 3, -5, 7,
					-- layer=2 filter=129 channel=81
					0, -3, 2, 0, -2, -7, 14, -7, -6,
					-- layer=2 filter=129 channel=82
					-13, 9, 0, -8, 9, 13, 0, 0, 1,
					-- layer=2 filter=129 channel=83
					-72, -14, 21, -39, -45, 33, -6, -20, -5,
					-- layer=2 filter=129 channel=84
					8, -2, 1, 7, 0, 10, -6, -8, 0,
					-- layer=2 filter=129 channel=85
					-15, -1, 14, 3, 12, -15, 1, 14, -6,
					-- layer=2 filter=129 channel=86
					13, 6, 3, 5, 6, 5, -10, 0, 5,
					-- layer=2 filter=129 channel=87
					18, -6, 40, 8, 27, 5, -44, 8, -2,
					-- layer=2 filter=129 channel=88
					-28, 18, 13, -36, 0, 4, -2, -12, -1,
					-- layer=2 filter=129 channel=89
					-13, 15, 0, -57, -16, 44, -36, 9, -14,
					-- layer=2 filter=129 channel=90
					8, -9, 5, 6, -10, -8, 7, -2, 11,
					-- layer=2 filter=129 channel=91
					-4, 28, 5, -72, 8, 17, -4, -4, 6,
					-- layer=2 filter=129 channel=92
					-13, 26, 13, -51, -15, 52, -23, 3, 4,
					-- layer=2 filter=129 channel=93
					-17, 40, 2, -56, 11, -37, -80, 33, -19,
					-- layer=2 filter=129 channel=94
					-16, -4, -10, 47, 22, 29, 6, -28, 19,
					-- layer=2 filter=129 channel=95
					-16, 15, 1, -9, -1, 7, -10, 6, -6,
					-- layer=2 filter=129 channel=96
					10, -18, -27, 19, 12, -35, -47, 0, -33,
					-- layer=2 filter=129 channel=97
					19, -5, 25, 2, -42, -39, -2, -29, -69,
					-- layer=2 filter=129 channel=98
					44, 28, 28, -8, 35, 11, -12, 30, 3,
					-- layer=2 filter=129 channel=99
					34, 21, 0, 12, 24, 17, 14, 3, 25,
					-- layer=2 filter=129 channel=100
					-55, -9, -16, -41, 2, 0, 28, 5, 15,
					-- layer=2 filter=129 channel=101
					52, 34, -29, 2, -2, -20, 12, 16, -24,
					-- layer=2 filter=129 channel=102
					48, -63, 9, 11, -45, 3, -35, -37, -56,
					-- layer=2 filter=129 channel=103
					10, 9, 16, -3, 1, -35, -12, 0, 1,
					-- layer=2 filter=129 channel=104
					-35, -16, 16, 17, -29, 21, 4, 0, -18,
					-- layer=2 filter=129 channel=105
					-15, -16, -10, -9, 26, 2, -5, -7, 21,
					-- layer=2 filter=129 channel=106
					-4, 36, 3, -34, -21, -23, 15, -20, -22,
					-- layer=2 filter=129 channel=107
					2, -22, 0, 32, -17, 29, 38, 16, 78,
					-- layer=2 filter=129 channel=108
					-3, -25, 36, -3, -28, 13, -6, -25, -38,
					-- layer=2 filter=129 channel=109
					2, 0, 13, -3, -14, -5, 14, -3, -16,
					-- layer=2 filter=129 channel=110
					-43, 14, 10, -9, -19, 16, -12, 12, 26,
					-- layer=2 filter=129 channel=111
					0, 1, 4, -6, -10, 4, 8, 5, 5,
					-- layer=2 filter=129 channel=112
					45, -22, -5, 16, 15, -17, 22, -1, -2,
					-- layer=2 filter=129 channel=113
					-11, -15, -9, 25, -45, 35, -11, 39, 16,
					-- layer=2 filter=129 channel=114
					7, -10, 9, 7, -9, 2, -7, 11, -19,
					-- layer=2 filter=129 channel=115
					8, 0, -2, 7, 8, -2, 10, 9, 8,
					-- layer=2 filter=129 channel=116
					44, -30, 53, -48, 9, -2, -64, 0, -11,
					-- layer=2 filter=129 channel=117
					61, 26, 13, -26, -23, 29, -68, -19, 36,
					-- layer=2 filter=129 channel=118
					7, 7, 7, -2, 0, -19, 0, -1, -43,
					-- layer=2 filter=129 channel=119
					-10, -11, 18, -12, -54, 6, -24, -28, -18,
					-- layer=2 filter=129 channel=120
					-8, 1, 4, -9, 6, 8, 0, 9, -2,
					-- layer=2 filter=129 channel=121
					-2, -2, 0, -1, -7, 0, 5, 5, 9,
					-- layer=2 filter=129 channel=122
					9, 1, -4, 20, 7, 6, 2, 2, 0,
					-- layer=2 filter=129 channel=123
					4, 23, -28, -30, 25, 7, -51, 2, 16,
					-- layer=2 filter=129 channel=124
					27, -3, 68, -45, 16, 29, -24, 40, 11,
					-- layer=2 filter=129 channel=125
					-2, -1, -3, 11, 3, 5, 7, 0, 3,
					-- layer=2 filter=129 channel=126
					1, -16, -19, 11, -36, 31, -63, -57, -43,
					-- layer=2 filter=129 channel=127
					-19, 15, -3, 1, -5, 14, -16, -24, -31,
					-- layer=2 filter=130 channel=0
					28, 6, 17, 15, -1, 23, -9, -19, -14,
					-- layer=2 filter=130 channel=1
					-43, 11, -14, 26, 2, -11, 17, 2, -6,
					-- layer=2 filter=130 channel=2
					-7, 1, -10, -7, -3, 3, -7, 0, 0,
					-- layer=2 filter=130 channel=3
					-1, -2, -14, 3, 11, 5, 4, -8, 10,
					-- layer=2 filter=130 channel=4
					9, 0, -19, -4, 18, 16, 1, -28, -28,
					-- layer=2 filter=130 channel=5
					21, 20, 31, -3, 7, -3, -10, -31, 22,
					-- layer=2 filter=130 channel=6
					-65, -35, -1, -75, -19, -64, 20, 52, 28,
					-- layer=2 filter=130 channel=7
					-16, -45, 0, 1, 62, 39, -11, -13, -51,
					-- layer=2 filter=130 channel=8
					-11, -8, 5, 3, 6, -7, -7, 2, 2,
					-- layer=2 filter=130 channel=9
					-10, -18, 0, -30, 10, -8, 8, -13, -24,
					-- layer=2 filter=130 channel=10
					22, 7, 0, 17, 15, 18, -13, -6, -18,
					-- layer=2 filter=130 channel=11
					9, 7, 0, -10, -17, -10, 5, 20, 15,
					-- layer=2 filter=130 channel=12
					-19, 16, -4, 32, 25, 1, -2, 6, -19,
					-- layer=2 filter=130 channel=13
					-1, 11, 0, -6, 0, -8, -7, 1, 1,
					-- layer=2 filter=130 channel=14
					-37, -11, -3, 7, 3, 1, 35, 5, 0,
					-- layer=2 filter=130 channel=15
					-11, -94, 5, -29, -23, -2, -27, -4, -52,
					-- layer=2 filter=130 channel=16
					7, 1, -24, -2, -1, -1, -13, -27, -35,
					-- layer=2 filter=130 channel=17
					-3, -10, -2, 8, 0, -3, -4, 2, 8,
					-- layer=2 filter=130 channel=18
					-67, 19, 6, -32, 1, -31, 7, 0, -7,
					-- layer=2 filter=130 channel=19
					-62, -39, -24, -21, -16, -7, 12, -28, -6,
					-- layer=2 filter=130 channel=20
					4, -5, 5, -9, -8, 6, 0, 4, 0,
					-- layer=2 filter=130 channel=21
					0, -5, 11, -1, 0, -10, -22, -9, -5,
					-- layer=2 filter=130 channel=22
					-8, -2, 5, -1, -2, -11, 0, -1, 2,
					-- layer=2 filter=130 channel=23
					26, 22, 21, 14, 2, 5, 6, -23, -23,
					-- layer=2 filter=130 channel=24
					8, -3, -31, 4, 15, -6, 31, 45, 39,
					-- layer=2 filter=130 channel=25
					-21, -28, -52, -5, -7, -6, 23, 42, 38,
					-- layer=2 filter=130 channel=26
					-7, 6, 2, -5, -6, 0, -6, 10, -8,
					-- layer=2 filter=130 channel=27
					27, 32, 49, 16, 18, 25, 3, -16, 11,
					-- layer=2 filter=130 channel=28
					6, 33, 38, 16, 27, 19, -1, -3, 19,
					-- layer=2 filter=130 channel=29
					5, 12, -8, 2, 5, 8, 0, 4, 0,
					-- layer=2 filter=130 channel=30
					-3, 9, 0, 2, -12, 2, -30, 6, -12,
					-- layer=2 filter=130 channel=31
					-20, 16, -21, -36, 12, -52, 28, 48, 0,
					-- layer=2 filter=130 channel=32
					4, 4, 9, -4, 1, 6, 0, -4, -2,
					-- layer=2 filter=130 channel=33
					-6, -20, 5, -12, 29, 36, 10, -1, -23,
					-- layer=2 filter=130 channel=34
					-67, 36, 15, 0, -17, -8, 6, 36, 17,
					-- layer=2 filter=130 channel=35
					8, 31, 22, -22, 1, -6, -12, 0, 20,
					-- layer=2 filter=130 channel=36
					3, 10, 1, 11, -3, -6, 5, -3, -10,
					-- layer=2 filter=130 channel=37
					2, 14, 12, 5, -9, 4, 6, 13, 6,
					-- layer=2 filter=130 channel=38
					12, 32, 36, 13, 17, 12, -2, -9, 3,
					-- layer=2 filter=130 channel=39
					16, 13, -5, 19, 21, 37, -28, -22, -29,
					-- layer=2 filter=130 channel=40
					-7, -2, 3, -28, -45, -48, -26, 71, 28,
					-- layer=2 filter=130 channel=41
					1, 6, 8, 7, -10, 6, -9, 2, -10,
					-- layer=2 filter=130 channel=42
					22, 20, 5, 22, -4, 12, 0, -2, -7,
					-- layer=2 filter=130 channel=43
					16, 25, 49, -8, -28, 0, -67, -32, -11,
					-- layer=2 filter=130 channel=44
					4, -4, 0, 6, -6, -3, 7, 4, -8,
					-- layer=2 filter=130 channel=45
					-14, -18, -37, -3, -6, -15, -12, -19, -7,
					-- layer=2 filter=130 channel=46
					19, 3, 21, 30, 4, 24, -28, -24, -30,
					-- layer=2 filter=130 channel=47
					15, 28, 6, 28, 44, 75, -7, 42, 9,
					-- layer=2 filter=130 channel=48
					3, 8, -8, 7, 0, -5, 4, -8, -5,
					-- layer=2 filter=130 channel=49
					-65, -31, -17, -53, -30, -23, 12, 11, 30,
					-- layer=2 filter=130 channel=50
					0, -20, -3, 0, 0, 2, 0, -27, -12,
					-- layer=2 filter=130 channel=51
					13, 6, 4, -14, -9, -2, 15, 2, 17,
					-- layer=2 filter=130 channel=52
					-44, -39, -3, -27, -60, -70, 6, 12, -2,
					-- layer=2 filter=130 channel=53
					-24, -64, -13, 6, 19, 32, -19, -5, -67,
					-- layer=2 filter=130 channel=54
					-48, -10, -17, -32, -18, -5, -1, 16, 34,
					-- layer=2 filter=130 channel=55
					1, -1, -6, 6, -12, 10, -6, 0, 8,
					-- layer=2 filter=130 channel=56
					5, 38, 24, 6, -2, -5, 20, 0, 12,
					-- layer=2 filter=130 channel=57
					7, 11, -7, 1, 11, -7, 13, 1, -3,
					-- layer=2 filter=130 channel=58
					-22, 38, 22, 22, 19, 8, -21, -13, -13,
					-- layer=2 filter=130 channel=59
					-13, -4, 38, 34, 20, 25, -30, 6, -14,
					-- layer=2 filter=130 channel=60
					-26, 39, 5, 13, -3, -11, -27, -10, 12,
					-- layer=2 filter=130 channel=61
					-5, -67, -9, -65, -66, -113, -5, 0, -1,
					-- layer=2 filter=130 channel=62
					-58, -32, -24, -43, -42, -44, 12, 33, 28,
					-- layer=2 filter=130 channel=63
					13, -9, -5, 7, 3, -10, -8, -15, -7,
					-- layer=2 filter=130 channel=64
					7, 19, -12, 23, 12, 16, 4, 20, 18,
					-- layer=2 filter=130 channel=65
					-60, -25, -2, -67, -98, -72, -9, -7, -38,
					-- layer=2 filter=130 channel=66
					45, 16, -2, -10, 37, 18, -20, -3, 14,
					-- layer=2 filter=130 channel=67
					33, 26, 31, 44, 12, 28, -25, -3, -42,
					-- layer=2 filter=130 channel=68
					0, -7, 6, 1, 6, 5, -2, 3, -8,
					-- layer=2 filter=130 channel=69
					10, 12, -16, 28, 6, 20, 6, 15, 23,
					-- layer=2 filter=130 channel=70
					-12, 38, 43, -9, 1, -4, 0, -3, 18,
					-- layer=2 filter=130 channel=71
					24, 36, 34, 4, 26, 3, 2, -7, 19,
					-- layer=2 filter=130 channel=72
					8, -35, 17, -18, 31, 8, 26, -18, -19,
					-- layer=2 filter=130 channel=73
					-10, 20, 9, 19, 19, -29, 12, 66, 41,
					-- layer=2 filter=130 channel=74
					13, 3, 5, 36, 1, 11, -21, 1, -2,
					-- layer=2 filter=130 channel=75
					0, -12, -22, 16, -27, -26, -17, -29, -38,
					-- layer=2 filter=130 channel=76
					-33, -34, -16, -36, -51, -76, -38, -22, -51,
					-- layer=2 filter=130 channel=77
					6, -9, 5, -1, 7, -3, 10, 8, -3,
					-- layer=2 filter=130 channel=78
					9, 22, -8, -20, -31, 2, 23, 40, 32,
					-- layer=2 filter=130 channel=79
					-9, 7, 5, 2, 11, 0, -7, 7, -2,
					-- layer=2 filter=130 channel=80
					25, -5, -18, 26, 22, 39, -28, -40, -25,
					-- layer=2 filter=130 channel=81
					-4, -11, -7, 5, 2, -6, -14, -12, 0,
					-- layer=2 filter=130 channel=82
					2, 2, 0, -4, 3, -4, 12, -9, -2,
					-- layer=2 filter=130 channel=83
					9, 11, 3, 20, 17, -14, -15, -20, -2,
					-- layer=2 filter=130 channel=84
					2, -11, -3, 4, 8, 7, -3, 7, 7,
					-- layer=2 filter=130 channel=85
					11, 0, 20, 3, 2, -9, 0, -8, 6,
					-- layer=2 filter=130 channel=86
					-14, -28, -4, -3, 8, -2, -8, 1, -15,
					-- layer=2 filter=130 channel=87
					10, -8, 10, -57, 1, -24, -21, 19, -54,
					-- layer=2 filter=130 channel=88
					0, -4, -16, 29, -18, -7, -10, 23, 2,
					-- layer=2 filter=130 channel=89
					-33, 10, 13, 18, 9, 10, 12, -4, -35,
					-- layer=2 filter=130 channel=90
					5, -9, 0, -8, -9, 4, 5, -9, -6,
					-- layer=2 filter=130 channel=91
					-22, 27, 10, 14, 8, -4, -1, -1, -34,
					-- layer=2 filter=130 channel=92
					-17, 11, -15, 0, 20, -4, 5, -3, 0,
					-- layer=2 filter=130 channel=93
					-135, -18, 20, -94, -37, -9, 6, 39, 15,
					-- layer=2 filter=130 channel=94
					-12, -93, -38, -59, -24, -84, 11, 0, -20,
					-- layer=2 filter=130 channel=95
					-17, -7, -1, -1, -12, -11, 4, -10, 8,
					-- layer=2 filter=130 channel=96
					-38, -20, -32, -4, -91, -30, 27, -29, -32,
					-- layer=2 filter=130 channel=97
					7, -15, -21, 0, 23, 16, 6, 46, 28,
					-- layer=2 filter=130 channel=98
					-5, -2, 15, -1, 19, 27, 14, 42, 25,
					-- layer=2 filter=130 channel=99
					-19, -6, 42, -32, -53, 11, -17, 43, 37,
					-- layer=2 filter=130 channel=100
					12, 35, 7, 13, 0, 15, -35, -18, -9,
					-- layer=2 filter=130 channel=101
					12, 10, -10, -12, -1, 1, 0, -33, -28,
					-- layer=2 filter=130 channel=102
					-39, -24, -44, -45, -74, -43, 16, -21, 4,
					-- layer=2 filter=130 channel=103
					1, 0, -10, -27, -11, 15, -23, -8, 0,
					-- layer=2 filter=130 channel=104
					-18, 31, -20, -41, -25, -101, 35, -46, -35,
					-- layer=2 filter=130 channel=105
					-7, 22, 22, -58, -7, -25, -67, -21, -18,
					-- layer=2 filter=130 channel=106
					-10, 0, -14, 5, 25, 5, 15, 4, -16,
					-- layer=2 filter=130 channel=107
					-3, -7, -53, 56, 38, 48, 48, 13, 30,
					-- layer=2 filter=130 channel=108
					-9, 44, 12, 0, 25, 25, 0, -28, 33,
					-- layer=2 filter=130 channel=109
					-1, 4, 0, -4, 6, -3, -3, 6, -3,
					-- layer=2 filter=130 channel=110
					4, -8, 13, -1, 7, 32, -4, -18, -24,
					-- layer=2 filter=130 channel=111
					0, -3, 4, -8, 2, -8, 7, 5, 9,
					-- layer=2 filter=130 channel=112
					-9, 5, 16, -20, -26, -26, 20, 1, -17,
					-- layer=2 filter=130 channel=113
					-23, 30, 12, 3, -28, -22, -29, -21, -13,
					-- layer=2 filter=130 channel=114
					-4, 0, 1, -4, 7, 8, -1, 5, 7,
					-- layer=2 filter=130 channel=115
					-2, -2, -3, 10, 7, -2, -7, 6, 1,
					-- layer=2 filter=130 channel=116
					-18, -1, -3, -85, -31, -31, -1, -12, -77,
					-- layer=2 filter=130 channel=117
					-40, -19, -26, -9, -14, -21, 5, 12, 8,
					-- layer=2 filter=130 channel=118
					10, 33, 33, 25, 16, 14, -2, -16, -12,
					-- layer=2 filter=130 channel=119
					-46, -20, -46, -20, 2, 3, -19, -36, -13,
					-- layer=2 filter=130 channel=120
					9, 10, -7, -4, 8, 2, -9, 5, -5,
					-- layer=2 filter=130 channel=121
					9, 2, 1, 4, -3, 1, -1, 7, -9,
					-- layer=2 filter=130 channel=122
					-12, -7, -6, -8, 8, 0, -4, 15, 12,
					-- layer=2 filter=130 channel=123
					-7, -40, 25, 3, 28, 30, -1, -9, -11,
					-- layer=2 filter=130 channel=124
					2, -60, -4, -15, 2, 22, -72, -61, -51,
					-- layer=2 filter=130 channel=125
					-11, 8, 2, -6, 1, 1, -4, 7, 3,
					-- layer=2 filter=130 channel=126
					-11, -5, 20, -7, -18, -52, -91, 29, 28,
					-- layer=2 filter=130 channel=127
					-19, 16, -17, 36, -19, -5, 14, -21, -15,
					-- layer=2 filter=131 channel=0
					-6, 13, 9, 0, 27, 17, 18, 5, 18,
					-- layer=2 filter=131 channel=1
					-21, 0, -44, -42, -38, -57, 5, -7, 46,
					-- layer=2 filter=131 channel=2
					1, -9, -4, 7, 6, -8, -6, 4, 2,
					-- layer=2 filter=131 channel=3
					-28, -3, 35, -2, 18, 23, -11, -5, 0,
					-- layer=2 filter=131 channel=4
					-1, -14, 20, 4, -12, 18, 21, 20, 23,
					-- layer=2 filter=131 channel=5
					-4, -8, -16, 0, 8, 26, 38, 19, 8,
					-- layer=2 filter=131 channel=6
					-18, -39, 0, -20, 39, 41, -1, 59, 72,
					-- layer=2 filter=131 channel=7
					-15, -8, 1, -74, -9, 73, -29, -52, -42,
					-- layer=2 filter=131 channel=8
					8, -1, 8, -1, 0, -3, -5, 0, 6,
					-- layer=2 filter=131 channel=9
					14, 11, -18, 0, 18, -9, 22, 26, -18,
					-- layer=2 filter=131 channel=10
					4, 2, 8, 21, 20, 26, 27, -17, 16,
					-- layer=2 filter=131 channel=11
					-37, -25, 13, -17, -20, 22, -17, 5, 8,
					-- layer=2 filter=131 channel=12
					-24, 12, -54, -69, -56, 1, -1, -20, 19,
					-- layer=2 filter=131 channel=13
					2, 0, 2, -7, 9, -6, 6, -10, 5,
					-- layer=2 filter=131 channel=14
					-40, -29, -45, -55, -63, -54, 17, -27, 23,
					-- layer=2 filter=131 channel=15
					2, -24, -3, -15, -9, 16, -29, -23, -6,
					-- layer=2 filter=131 channel=16
					-11, -9, -28, 5, 5, -32, 36, 27, -21,
					-- layer=2 filter=131 channel=17
					7, 8, 9, 5, 6, -6, 5, 5, -2,
					-- layer=2 filter=131 channel=18
					-32, -16, -38, -21, -57, 40, -71, -35, 8,
					-- layer=2 filter=131 channel=19
					-25, -25, -45, -21, 0, -5, -35, -34, 30,
					-- layer=2 filter=131 channel=20
					-4, 2, -6, -4, -7, -3, 1, -2, 7,
					-- layer=2 filter=131 channel=21
					-12, -2, -12, 14, -2, -6, -5, -6, -4,
					-- layer=2 filter=131 channel=22
					-9, 1, 9, 10, -7, -6, -5, -5, 6,
					-- layer=2 filter=131 channel=23
					38, 17, 21, 9, 28, 39, 7, 26, 13,
					-- layer=2 filter=131 channel=24
					-18, 7, 15, -20, 5, 14, 0, 15, 13,
					-- layer=2 filter=131 channel=25
					-47, -9, 14, -37, -10, 28, -8, 4, 34,
					-- layer=2 filter=131 channel=26
					-5, 6, 0, 0, 5, 5, 4, 7, 6,
					-- layer=2 filter=131 channel=27
					-31, -35, -37, 14, 10, -24, -13, -4, -11,
					-- layer=2 filter=131 channel=28
					-8, 14, -15, -53, -16, -26, -30, -1, 0,
					-- layer=2 filter=131 channel=29
					9, 6, 3, 8, 6, -9, 9, 3, -7,
					-- layer=2 filter=131 channel=30
					11, 3, 1, 19, 8, -32, 12, -20, 6,
					-- layer=2 filter=131 channel=31
					12, -5, 33, 27, 19, 21, -7, 40, 31,
					-- layer=2 filter=131 channel=32
					-6, -4, 11, -8, 3, -2, -4, -10, 3,
					-- layer=2 filter=131 channel=33
					-11, -11, 65, -17, -18, 22, -22, -31, -17,
					-- layer=2 filter=131 channel=34
					27, -15, 13, -52, -34, 65, -101, 45, 65,
					-- layer=2 filter=131 channel=35
					-23, 2, -36, -64, -49, -25, -17, -18, 41,
					-- layer=2 filter=131 channel=36
					9, 2, -5, 4, 4, -1, 6, -2, -4,
					-- layer=2 filter=131 channel=37
					-11, 1, 1, 6, -2, 13, 6, 20, 0,
					-- layer=2 filter=131 channel=38
					-16, -13, -5, 16, -6, 18, -21, -20, 39,
					-- layer=2 filter=131 channel=39
					-10, -3, 3, -6, 1, -10, -1, 7, -38,
					-- layer=2 filter=131 channel=40
					-16, 1, 5, -38, -11, 22, -31, 6, 24,
					-- layer=2 filter=131 channel=41
					7, -1, -3, 7, 4, -7, -9, -5, -1,
					-- layer=2 filter=131 channel=42
					9, 30, 18, 7, -10, -8, 27, 15, 3,
					-- layer=2 filter=131 channel=43
					-9, -23, -34, 19, 13, 15, 31, 41, 49,
					-- layer=2 filter=131 channel=44
					1, 8, 7, 0, -4, 0, 0, 6, 0,
					-- layer=2 filter=131 channel=45
					-32, -84, -71, -24, -5, -10, -4, 15, 8,
					-- layer=2 filter=131 channel=46
					8, 10, 7, 8, 11, -12, 5, -19, 0,
					-- layer=2 filter=131 channel=47
					27, 9, 27, -34, 15, 34, -11, 11, 29,
					-- layer=2 filter=131 channel=48
					-8, 1, -4, -4, 4, -3, 0, 8, -3,
					-- layer=2 filter=131 channel=49
					7, -41, -65, -8, -72, 2, -27, -13, -11,
					-- layer=2 filter=131 channel=50
					3, -9, 0, 0, 6, -6, -1, -12, -7,
					-- layer=2 filter=131 channel=51
					-14, 2, 35, 7, -3, 33, 19, 31, 21,
					-- layer=2 filter=131 channel=52
					-32, -49, 2, 1, -47, 1, -11, -18, -31,
					-- layer=2 filter=131 channel=53
					-26, 13, -32, 5, 37, 1, -18, 20, 29,
					-- layer=2 filter=131 channel=54
					-5, -7, -12, -77, -23, 39, -7, -9, 52,
					-- layer=2 filter=131 channel=55
					10, -6, 4, 4, -5, -4, 11, 2, -6,
					-- layer=2 filter=131 channel=56
					-22, 14, 13, -21, 5, -3, -5, -5, -13,
					-- layer=2 filter=131 channel=57
					-7, 1, 2, 0, 5, -7, 6, 3, 4,
					-- layer=2 filter=131 channel=58
					-43, -5, -40, -42, -21, 6, -8, -29, 41,
					-- layer=2 filter=131 channel=59
					-55, -42, -35, -75, -7, -69, -54, -39, 11,
					-- layer=2 filter=131 channel=60
					-4, -12, -22, -33, -59, -21, -70, -55, 4,
					-- layer=2 filter=131 channel=61
					5, -45, -21, -59, -41, -21, -38, -39, -55,
					-- layer=2 filter=131 channel=62
					32, -51, 13, -28, -19, 29, -44, 20, 51,
					-- layer=2 filter=131 channel=63
					1, -15, -28, 1, 14, 0, -4, 5, -37,
					-- layer=2 filter=131 channel=64
					21, 7, 28, 14, -3, 6, 3, -1, -11,
					-- layer=2 filter=131 channel=65
					39, -31, 22, -9, -29, 24, -13, -29, 13,
					-- layer=2 filter=131 channel=66
					15, 18, 1, -7, 21, -22, 9, 31, -29,
					-- layer=2 filter=131 channel=67
					30, 12, 12, 9, 9, -1, 29, 19, 7,
					-- layer=2 filter=131 channel=68
					2, -9, 2, 0, 0, -4, 11, 9, 4,
					-- layer=2 filter=131 channel=69
					2, 15, 25, 12, 15, -2, 10, 15, -2,
					-- layer=2 filter=131 channel=70
					-8, 0, -39, -55, -6, -14, -52, -5, 35,
					-- layer=2 filter=131 channel=71
					-72, -47, -41, -40, -36, -41, -21, 10, -10,
					-- layer=2 filter=131 channel=72
					-41, 1, 21, -66, -35, 0, -23, -32, -30,
					-- layer=2 filter=131 channel=73
					7, -28, -57, 72, 60, -33, 39, 54, -33,
					-- layer=2 filter=131 channel=74
					7, 7, -12, 10, 7, -3, 9, 10, -1,
					-- layer=2 filter=131 channel=75
					-17, -13, -31, -32, -14, -16, 46, 9, 6,
					-- layer=2 filter=131 channel=76
					-81, -23, 20, -31, 22, 5, -54, 51, -34,
					-- layer=2 filter=131 channel=77
					1, 2, -12, 7, 9, 5, 3, -5, -1,
					-- layer=2 filter=131 channel=78
					-55, -49, 1, -6, 5, 30, -19, 13, -5,
					-- layer=2 filter=131 channel=79
					8, -6, -6, -7, 10, -4, 0, 5, -7,
					-- layer=2 filter=131 channel=80
					6, -2, 0, 17, 3, -5, 18, 12, 5,
					-- layer=2 filter=131 channel=81
					3, 7, 9, 11, 7, 2, 3, -9, -3,
					-- layer=2 filter=131 channel=82
					9, 8, 3, 0, -5, -2, 3, 2, -3,
					-- layer=2 filter=131 channel=83
					4, -1, -13, 8, 0, -6, 25, -1, 13,
					-- layer=2 filter=131 channel=84
					-4, -6, -1, -6, 1, 8, 0, 3, 4,
					-- layer=2 filter=131 channel=85
					4, -1, -9, 11, 10, 4, 13, 7, 14,
					-- layer=2 filter=131 channel=86
					16, -9, 15, 6, 0, 10, -2, 19, -14,
					-- layer=2 filter=131 channel=87
					-9, 12, -13, -4, -26, 20, -57, 18, 2,
					-- layer=2 filter=131 channel=88
					5, 0, 0, 8, -6, -25, 2, 10, 1,
					-- layer=2 filter=131 channel=89
					-57, -2, -27, -54, -5, -37, 26, -2, 25,
					-- layer=2 filter=131 channel=90
					0, 11, 0, -4, -6, 0, -5, 1, 4,
					-- layer=2 filter=131 channel=91
					-27, -9, -13, -7, 0, 16, 46, 29, 64,
					-- layer=2 filter=131 channel=92
					-22, -4, -53, -67, -56, -57, -1, -25, 24,
					-- layer=2 filter=131 channel=93
					12, -59, -1, 52, -17, -12, -19, -36, 23,
					-- layer=2 filter=131 channel=94
					4, -35, -31, -86, 51, -12, -31, 25, 6,
					-- layer=2 filter=131 channel=95
					-1, 4, 6, 3, 1, 4, 2, -11, 10,
					-- layer=2 filter=131 channel=96
					-8, -66, 12, 21, -17, 3, 55, 0, 10,
					-- layer=2 filter=131 channel=97
					-1, 0, 14, 6, 1, 16, 29, 14, 20,
					-- layer=2 filter=131 channel=98
					0, -6, -14, -86, -6, 13, -26, 22, -2,
					-- layer=2 filter=131 channel=99
					-60, -78, -10, -4, -37, -84, -52, -32, -34,
					-- layer=2 filter=131 channel=100
					13, 12, -11, -9, 14, -19, 7, -27, 34,
					-- layer=2 filter=131 channel=101
					-51, -43, -11, -39, -25, 8, -5, 4, 38,
					-- layer=2 filter=131 channel=102
					-4, -50, -22, 12, -64, -12, -2, -46, -43,
					-- layer=2 filter=131 channel=103
					15, 2, -6, 7, 5, -25, 32, 15, 23,
					-- layer=2 filter=131 channel=104
					-10, -16, -45, -8, 4, 13, -6, 14, 0,
					-- layer=2 filter=131 channel=105
					-5, -39, 18, -42, 8, 5, -12, -11, 13,
					-- layer=2 filter=131 channel=106
					-27, 7, 37, -27, -5, 27, 4, 14, 79,
					-- layer=2 filter=131 channel=107
					36, -21, -51, -11, -3, -68, -16, -35, 7,
					-- layer=2 filter=131 channel=108
					-43, -48, -67, -20, -23, -59, 1, -16, -35,
					-- layer=2 filter=131 channel=109
					-2, 8, -8, -2, 0, -7, -1, -4, 3,
					-- layer=2 filter=131 channel=110
					9, 13, 24, -8, 5, -24, 4, -4, -2,
					-- layer=2 filter=131 channel=111
					-4, 0, -7, 0, -9, 7, 7, -5, 2,
					-- layer=2 filter=131 channel=112
					-11, 17, 35, -29, 4, 33, 8, -28, 20,
					-- layer=2 filter=131 channel=113
					32, -7, 11, 4, 8, -24, 15, -36, 10,
					-- layer=2 filter=131 channel=114
					-5, 7, 3, 4, 5, 5, 3, 5, -2,
					-- layer=2 filter=131 channel=115
					-3, 4, 7, 6, 10, -4, -7, 8, -7,
					-- layer=2 filter=131 channel=116
					-25, 42, -44, -20, -26, 19, -36, 6, -8,
					-- layer=2 filter=131 channel=117
					-4, -6, -17, -84, -4, 47, 16, 4, -29,
					-- layer=2 filter=131 channel=118
					8, -9, 8, 14, 12, 18, 29, 25, 11,
					-- layer=2 filter=131 channel=119
					-12, -22, -33, -15, -25, 21, 2, 7, 17,
					-- layer=2 filter=131 channel=120
					-4, 1, 7, 7, 9, 5, -9, 0, 8,
					-- layer=2 filter=131 channel=121
					4, -7, -4, -4, 0, 4, 8, -8, 5,
					-- layer=2 filter=131 channel=122
					8, 7, 3, -3, 6, 0, -5, -7, 6,
					-- layer=2 filter=131 channel=123
					-13, -17, 26, -72, 11, 44, -24, -27, -32,
					-- layer=2 filter=131 channel=124
					-3, 1, 46, -98, 5, 33, -22, -7, -13,
					-- layer=2 filter=131 channel=125
					0, -3, -1, -7, 0, -5, -6, 1, 9,
					-- layer=2 filter=131 channel=126
					21, 9, -18, 66, 14, -11, 2, 25, -8,
					-- layer=2 filter=131 channel=127
					-16, -20, 21, -9, -13, -15, -23, 11, 0,
					-- layer=2 filter=132 channel=0
					-11, -2, 2, 5, -5, 4, -9, 3, -2,
					-- layer=2 filter=132 channel=1
					-5, 2, -4, 2, 2, 0, 0, -4, 5,
					-- layer=2 filter=132 channel=2
					-6, 6, -9, 5, -4, -6, -5, -4, 6,
					-- layer=2 filter=132 channel=3
					-9, -10, -2, -3, -10, 0, -3, -8, 5,
					-- layer=2 filter=132 channel=4
					-2, 5, 8, -2, -7, -3, 6, 5, -4,
					-- layer=2 filter=132 channel=5
					-7, -15, -6, -8, 0, -12, 0, -5, 2,
					-- layer=2 filter=132 channel=6
					1, 5, -8, -11, 4, 1, -1, -6, 4,
					-- layer=2 filter=132 channel=7
					2, 0, -9, -6, -14, -8, -8, 0, -3,
					-- layer=2 filter=132 channel=8
					2, 10, 0, 4, 8, 8, -8, 3, 9,
					-- layer=2 filter=132 channel=9
					-5, -2, 4, -11, 4, -7, -1, 2, 4,
					-- layer=2 filter=132 channel=10
					0, 0, -5, -6, -4, -8, 3, -1, -13,
					-- layer=2 filter=132 channel=11
					0, 0, -11, -9, 0, 1, -9, 4, -14,
					-- layer=2 filter=132 channel=12
					-5, -15, -7, -1, -13, -9, 7, -8, -5,
					-- layer=2 filter=132 channel=13
					-3, -2, -3, -5, 8, -4, 0, -4, -4,
					-- layer=2 filter=132 channel=14
					5, 2, -8, -8, -12, 9, -8, 0, -9,
					-- layer=2 filter=132 channel=15
					4, -10, -3, 3, 0, -12, -11, 6, -8,
					-- layer=2 filter=132 channel=16
					-14, 4, 4, -11, 3, 1, -2, 0, -8,
					-- layer=2 filter=132 channel=17
					-3, -6, 6, 7, 5, 0, -7, 0, 3,
					-- layer=2 filter=132 channel=18
					-4, -6, -3, 0, 0, -10, -1, -3, 4,
					-- layer=2 filter=132 channel=19
					-12, 5, -3, 5, -9, -4, -1, -7, 5,
					-- layer=2 filter=132 channel=20
					-11, -8, -9, -1, 10, -3, 4, 2, 3,
					-- layer=2 filter=132 channel=21
					7, 4, -1, -11, 1, -1, -7, 2, 4,
					-- layer=2 filter=132 channel=22
					3, 6, -8, -6, 8, -5, -7, -10, -10,
					-- layer=2 filter=132 channel=23
					0, 7, 1, -7, -1, 2, -14, 5, -5,
					-- layer=2 filter=132 channel=24
					-3, 4, -3, 2, -4, -15, 5, 7, -10,
					-- layer=2 filter=132 channel=25
					-4, 2, -5, 3, -6, 5, 3, 4, -12,
					-- layer=2 filter=132 channel=26
					4, -4, 5, 0, 5, 2, -4, 3, -7,
					-- layer=2 filter=132 channel=27
					-1, -9, 6, 1, -10, 7, -5, -3, 0,
					-- layer=2 filter=132 channel=28
					-1, 0, 9, 0, -4, -10, -15, -1, 5,
					-- layer=2 filter=132 channel=29
					4, 2, -1, -1, 4, -1, 8, 4, -7,
					-- layer=2 filter=132 channel=30
					-9, -4, 5, -16, -11, -3, -2, 3, -11,
					-- layer=2 filter=132 channel=31
					0, -5, -9, 7, -11, 2, -5, -3, -7,
					-- layer=2 filter=132 channel=32
					-6, -5, 1, 1, -9, 9, 3, -5, -7,
					-- layer=2 filter=132 channel=33
					-13, -3, 3, -1, -14, 5, -6, -1, -10,
					-- layer=2 filter=132 channel=34
					-4, 2, -4, 6, 0, 0, 1, -1, 7,
					-- layer=2 filter=132 channel=35
					-12, -2, 4, -4, -6, -4, -3, 1, -14,
					-- layer=2 filter=132 channel=36
					-11, -2, -5, -9, -5, -5, -2, -2, -10,
					-- layer=2 filter=132 channel=37
					-2, 4, 2, 0, -2, -8, -5, 0, -9,
					-- layer=2 filter=132 channel=38
					0, -5, -12, -4, -9, -4, -14, -2, -9,
					-- layer=2 filter=132 channel=39
					-12, -10, 7, -3, -9, 3, -10, -11, -5,
					-- layer=2 filter=132 channel=40
					5, 7, 0, -6, 1, 3, 6, -3, -8,
					-- layer=2 filter=132 channel=41
					1, -7, 0, 7, -5, -3, 0, -1, -6,
					-- layer=2 filter=132 channel=42
					-10, 6, 4, 4, 4, 0, -12, 8, -6,
					-- layer=2 filter=132 channel=43
					-16, 0, -4, -9, -1, 1, -7, -6, -14,
					-- layer=2 filter=132 channel=44
					6, 8, 8, 7, 9, 3, -7, 2, -3,
					-- layer=2 filter=132 channel=45
					0, -8, 0, -9, 0, 5, -8, -7, 8,
					-- layer=2 filter=132 channel=46
					-11, -10, -8, -5, 2, -8, 6, -8, 7,
					-- layer=2 filter=132 channel=47
					1, -3, -2, -7, 0, -11, 0, 3, -7,
					-- layer=2 filter=132 channel=48
					8, 1, -10, 7, 3, -4, 5, -5, -10,
					-- layer=2 filter=132 channel=49
					-15, 0, 4, -6, 3, -7, -8, -7, -11,
					-- layer=2 filter=132 channel=50
					6, -9, -10, 7, -7, -5, -6, 9, 0,
					-- layer=2 filter=132 channel=51
					-4, -3, -5, -12, -9, 1, -11, -2, -9,
					-- layer=2 filter=132 channel=52
					-16, -4, -3, -7, -5, -14, -8, -9, 3,
					-- layer=2 filter=132 channel=53
					5, -7, 3, 4, -8, -6, -10, 6, -9,
					-- layer=2 filter=132 channel=54
					1, -17, 5, -1, -7, -4, 4, 5, -14,
					-- layer=2 filter=132 channel=55
					-10, 0, 8, -6, 8, 4, -8, 5, -3,
					-- layer=2 filter=132 channel=56
					-11, -12, 1, 4, 6, -7, 6, 0, -1,
					-- layer=2 filter=132 channel=57
					7, -5, 8, 8, -8, 4, 1, 0, -2,
					-- layer=2 filter=132 channel=58
					-5, 2, 0, 0, -15, 0, 6, 2, 0,
					-- layer=2 filter=132 channel=59
					0, 9, 0, -14, -6, 11, -3, 7, -3,
					-- layer=2 filter=132 channel=60
					-7, -12, -12, -7, -6, -6, 0, -9, -5,
					-- layer=2 filter=132 channel=61
					-9, -10, -8, 0, 0, -7, -5, -2, 0,
					-- layer=2 filter=132 channel=62
					-9, 1, -2, -3, -11, -11, 8, 7, 8,
					-- layer=2 filter=132 channel=63
					-3, -1, -12, 1, -11, 7, 0, -3, -6,
					-- layer=2 filter=132 channel=64
					-13, -11, -6, -1, 6, -11, -11, 2, -10,
					-- layer=2 filter=132 channel=65
					3, -8, -10, -13, -15, -10, -11, -3, -9,
					-- layer=2 filter=132 channel=66
					-7, 6, 0, 2, 5, 2, 6, 4, -5,
					-- layer=2 filter=132 channel=67
					7, 2, 6, -12, -6, 4, -7, -6, -13,
					-- layer=2 filter=132 channel=68
					-2, 9, -8, -7, 8, -4, 5, 5, -11,
					-- layer=2 filter=132 channel=69
					0, 3, 3, 0, -4, -11, -3, 3, -2,
					-- layer=2 filter=132 channel=70
					-2, -13, 0, 5, -6, -14, 4, -14, -1,
					-- layer=2 filter=132 channel=71
					10, 1, 0, 0, -1, 1, -7, 4, 6,
					-- layer=2 filter=132 channel=72
					2, 8, -13, -13, 4, -10, 3, -11, -5,
					-- layer=2 filter=132 channel=73
					-6, -3, 0, -6, 5, -4, 2, -2, 2,
					-- layer=2 filter=132 channel=74
					3, -7, 3, 2, -5, 5, 5, 6, -3,
					-- layer=2 filter=132 channel=75
					-11, -15, 0, -2, 6, 10, -7, -7, -2,
					-- layer=2 filter=132 channel=76
					9, -1, -1, -9, -9, -9, 8, 4, 10,
					-- layer=2 filter=132 channel=77
					-7, -2, 0, -3, -5, -9, -5, -9, -12,
					-- layer=2 filter=132 channel=78
					-4, -10, 8, -11, 1, -1, -11, 0, -11,
					-- layer=2 filter=132 channel=79
					6, 2, 2, -2, 0, 8, -7, 3, 0,
					-- layer=2 filter=132 channel=80
					-9, 3, -9, -2, -8, -2, -2, 0, -5,
					-- layer=2 filter=132 channel=81
					-10, -7, 0, 0, 5, 1, 7, -11, 4,
					-- layer=2 filter=132 channel=82
					9, -4, 4, 8, 0, 5, 3, -9, 1,
					-- layer=2 filter=132 channel=83
					3, -7, -8, 0, 8, -12, -3, -11, 5,
					-- layer=2 filter=132 channel=84
					2, -1, 7, 0, 6, -7, 2, -6, -3,
					-- layer=2 filter=132 channel=85
					0, 6, -6, 3, 7, -5, 8, -2, 1,
					-- layer=2 filter=132 channel=86
					-1, 2, 0, 10, -10, 3, -6, -6, 1,
					-- layer=2 filter=132 channel=87
					3, 0, 6, 7, -5, -14, 7, -9, 1,
					-- layer=2 filter=132 channel=88
					-9, -10, 1, 0, -6, 9, -1, -6, 1,
					-- layer=2 filter=132 channel=89
					-11, 1, -12, -2, -11, -6, 1, 2, 9,
					-- layer=2 filter=132 channel=90
					0, -9, -6, 7, -6, 5, 4, -8, 9,
					-- layer=2 filter=132 channel=91
					-9, -9, 1, 4, -14, 0, 1, -9, -7,
					-- layer=2 filter=132 channel=92
					9, -10, 1, 0, 4, -10, -5, -5, -2,
					-- layer=2 filter=132 channel=93
					-7, -6, 4, -10, 6, -10, 1, 0, 8,
					-- layer=2 filter=132 channel=94
					-8, -4, 0, 1, -7, 4, -15, -7, -3,
					-- layer=2 filter=132 channel=95
					2, 0, -11, -10, 0, 3, 4, -6, -9,
					-- layer=2 filter=132 channel=96
					-8, 4, 0, 5, 0, -10, 3, -2, 0,
					-- layer=2 filter=132 channel=97
					-7, 7, 3, -3, 3, -9, 0, -3, 2,
					-- layer=2 filter=132 channel=98
					-3, -14, 0, -11, -5, -1, -13, -9, -7,
					-- layer=2 filter=132 channel=99
					9, 5, 9, 2, -7, -6, -7, 5, 10,
					-- layer=2 filter=132 channel=100
					-11, 0, -11, -4, -4, 5, 6, -4, -10,
					-- layer=2 filter=132 channel=101
					8, 0, 4, 8, -2, 4, 0, 0, -7,
					-- layer=2 filter=132 channel=102
					2, 0, -10, 0, -10, 1, -9, 1, -5,
					-- layer=2 filter=132 channel=103
					7, 8, -6, -1, 1, 7, -5, -4, 2,
					-- layer=2 filter=132 channel=104
					-6, -7, -6, 6, -4, 4, 1, 5, 6,
					-- layer=2 filter=132 channel=105
					3, 2, 3, -11, -11, 3, 0, -2, -9,
					-- layer=2 filter=132 channel=106
					-4, -7, -2, 2, -15, -2, 0, 6, -3,
					-- layer=2 filter=132 channel=107
					0, 2, 9, 8, 1, 7, -1, 0, -5,
					-- layer=2 filter=132 channel=108
					-3, -10, 1, -2, -12, -11, -12, 1, -5,
					-- layer=2 filter=132 channel=109
					-5, -6, -3, 3, 5, -10, 4, 5, -6,
					-- layer=2 filter=132 channel=110
					-9, -2, -6, -8, 0, 0, -1, 4, 0,
					-- layer=2 filter=132 channel=111
					-3, 5, -3, 8, 4, 10, -6, -5, -4,
					-- layer=2 filter=132 channel=112
					-2, -5, -11, 4, -2, 4, 1, -10, -12,
					-- layer=2 filter=132 channel=113
					7, -9, -14, -3, -12, -10, -3, -6, -6,
					-- layer=2 filter=132 channel=114
					3, -1, 3, 7, 5, 5, -3, -4, 1,
					-- layer=2 filter=132 channel=115
					-8, 0, -8, -4, -2, 0, -2, 5, 10,
					-- layer=2 filter=132 channel=116
					2, -5, 0, -3, -1, 2, 6, -3, -2,
					-- layer=2 filter=132 channel=117
					-14, -7, 0, 0, 1, -12, 7, -4, 9,
					-- layer=2 filter=132 channel=118
					-13, -1, 7, -11, 5, 4, -3, 3, -10,
					-- layer=2 filter=132 channel=119
					-11, -9, -7, -9, 3, 0, -5, 2, -6,
					-- layer=2 filter=132 channel=120
					9, -4, 3, -9, -9, -5, -1, -5, -10,
					-- layer=2 filter=132 channel=121
					-7, -11, 4, -1, -7, 8, 0, -7, 6,
					-- layer=2 filter=132 channel=122
					5, -9, 0, -6, -10, -5, 3, -2, 0,
					-- layer=2 filter=132 channel=123
					-4, 1, -4, 5, -3, 0, 2, -4, -5,
					-- layer=2 filter=132 channel=124
					7, 8, 1, 2, -15, -8, -3, -1, -8,
					-- layer=2 filter=132 channel=125
					0, -4, -10, 3, 10, 6, 9, -5, 7,
					-- layer=2 filter=132 channel=126
					-4, 6, -3, 2, -9, -1, 1, -6, -11,
					-- layer=2 filter=132 channel=127
					7, 0, -9, 0, -5, 0, -5, -9, 5,
					-- layer=2 filter=133 channel=0
					-3, -9, -13, -11, 5, -10, -1, -5, -8,
					-- layer=2 filter=133 channel=1
					-1, 2, -7, 4, 2, -3, -17, 0, -1,
					-- layer=2 filter=133 channel=2
					2, 3, -6, 5, 4, 5, -9, 8, 6,
					-- layer=2 filter=133 channel=3
					-18, -4, -7, 5, -5, -15, -1, 0, 2,
					-- layer=2 filter=133 channel=4
					-10, -10, -13, -9, -16, -5, 0, -7, -4,
					-- layer=2 filter=133 channel=5
					0, 2, -15, -17, -5, -11, -18, -2, -9,
					-- layer=2 filter=133 channel=6
					-3, 0, -12, -3, -3, -9, -4, 1, -3,
					-- layer=2 filter=133 channel=7
					-1, -10, -6, -5, -16, 5, -5, 2, -15,
					-- layer=2 filter=133 channel=8
					9, -5, -5, 8, 5, 0, 3, -2, -2,
					-- layer=2 filter=133 channel=9
					7, -4, 1, 2, -1, 2, -7, 8, -7,
					-- layer=2 filter=133 channel=10
					7, -13, 4, -19, -4, -8, -3, -2, -10,
					-- layer=2 filter=133 channel=11
					-13, -1, -17, -1, -17, -11, -6, -12, -8,
					-- layer=2 filter=133 channel=12
					-7, 0, 4, 2, -11, -4, -17, -2, 4,
					-- layer=2 filter=133 channel=13
					-10, -10, 7, -1, -2, 8, -4, -5, -7,
					-- layer=2 filter=133 channel=14
					-13, -13, 1, 3, -7, -7, -8, -6, 0,
					-- layer=2 filter=133 channel=15
					0, 0, 1, -15, 5, 0, -12, -11, -7,
					-- layer=2 filter=133 channel=16
					-8, -8, 7, -14, 0, -4, -16, -2, 3,
					-- layer=2 filter=133 channel=17
					4, 0, -6, 1, 8, 3, -1, -5, -8,
					-- layer=2 filter=133 channel=18
					-11, -10, -13, 1, 1, -12, -9, -15, -2,
					-- layer=2 filter=133 channel=19
					-12, -7, -18, 4, -8, -4, -4, -8, -8,
					-- layer=2 filter=133 channel=20
					0, 5, -2, 7, 0, -10, 6, 7, 3,
					-- layer=2 filter=133 channel=21
					-10, -11, 6, 0, -7, 4, 6, 2, -5,
					-- layer=2 filter=133 channel=22
					4, -6, 7, -11, -6, -2, -7, -2, 11,
					-- layer=2 filter=133 channel=23
					-10, -1, 5, -17, -12, -3, -18, 1, -20,
					-- layer=2 filter=133 channel=24
					-5, -2, 3, 3, -6, -3, -12, 0, -12,
					-- layer=2 filter=133 channel=25
					5, 2, -19, -10, -11, -2, -6, 7, -8,
					-- layer=2 filter=133 channel=26
					-8, 1, 8, 0, -3, -9, -6, -5, 1,
					-- layer=2 filter=133 channel=27
					2, -5, -2, -12, -10, 1, -7, -3, 3,
					-- layer=2 filter=133 channel=28
					14, 0, 0, 10, 14, 0, 2, -9, -2,
					-- layer=2 filter=133 channel=29
					-8, 0, -8, -5, 0, -4, 7, -3, 0,
					-- layer=2 filter=133 channel=30
					-7, -4, 0, -2, -3, -14, -16, -14, -10,
					-- layer=2 filter=133 channel=31
					-16, 4, -1, -4, -14, -1, -10, -8, -13,
					-- layer=2 filter=133 channel=32
					3, -8, 0, -7, 4, -2, 2, -8, -6,
					-- layer=2 filter=133 channel=33
					-4, 6, 6, -13, 2, -7, 9, 4, 5,
					-- layer=2 filter=133 channel=34
					-1, 1, 0, -10, -12, 2, -2, -11, -8,
					-- layer=2 filter=133 channel=35
					-9, -5, -13, -8, -2, 3, -14, -1, -10,
					-- layer=2 filter=133 channel=36
					-5, -8, -2, 1, -1, 5, -8, 6, -3,
					-- layer=2 filter=133 channel=37
					0, -16, -13, -16, -4, 0, -16, -3, 0,
					-- layer=2 filter=133 channel=38
					-7, -10, -10, 5, -10, -11, -3, 0, 1,
					-- layer=2 filter=133 channel=39
					0, 0, 0, -3, -6, -8, 1, -1, -7,
					-- layer=2 filter=133 channel=40
					15, -12, -14, -6, 9, -17, 15, -9, -11,
					-- layer=2 filter=133 channel=41
					-7, 3, -4, 6, 5, -1, -6, -5, -9,
					-- layer=2 filter=133 channel=42
					0, -5, -5, -18, -5, 0, -10, -5, 4,
					-- layer=2 filter=133 channel=43
					-14, 4, -9, -3, 9, -6, 0, 7, -3,
					-- layer=2 filter=133 channel=44
					10, -10, 0, 0, -4, 1, -8, -4, 1,
					-- layer=2 filter=133 channel=45
					-11, 3, 3, -1, 4, -9, -2, -2, -5,
					-- layer=2 filter=133 channel=46
					3, -2, -6, 0, -7, -4, -4, -8, -9,
					-- layer=2 filter=133 channel=47
					5, -4, 2, -9, 0, 0, 8, -3, -3,
					-- layer=2 filter=133 channel=48
					0, 7, -11, -9, 7, -5, 0, -6, -5,
					-- layer=2 filter=133 channel=49
					-19, -17, -6, -11, -17, 5, -8, -14, -5,
					-- layer=2 filter=133 channel=50
					-1, 5, -2, 7, 2, 5, -1, -2, 6,
					-- layer=2 filter=133 channel=51
					1, -9, -10, -18, -11, -10, -2, -1, -8,
					-- layer=2 filter=133 channel=52
					-11, -10, 2, -5, -15, 0, -5, -3, -10,
					-- layer=2 filter=133 channel=53
					-16, -10, -6, -13, -3, -2, -7, 15, -1,
					-- layer=2 filter=133 channel=54
					3, 6, 5, -15, -11, 3, -9, -14, -17,
					-- layer=2 filter=133 channel=55
					9, 4, -10, -8, -8, 1, 2, 1, 1,
					-- layer=2 filter=133 channel=56
					-7, -14, 0, 2, -14, -11, -13, -1, -4,
					-- layer=2 filter=133 channel=57
					-8, 3, 0, 2, -1, -11, -11, -12, -10,
					-- layer=2 filter=133 channel=58
					-1, -14, 13, 2, -2, 1, -2, -8, 9,
					-- layer=2 filter=133 channel=59
					1, -8, -16, -7, -16, -14, 2, 0, -1,
					-- layer=2 filter=133 channel=60
					-5, 1, -4, 3, 0, -2, -21, -7, -6,
					-- layer=2 filter=133 channel=61
					10, -11, -12, -9, -15, -11, -15, 0, -1,
					-- layer=2 filter=133 channel=62
					12, 5, -11, 0, -14, -15, -16, -5, -16,
					-- layer=2 filter=133 channel=63
					14, -7, -8, -8, -3, -6, -9, -4, 3,
					-- layer=2 filter=133 channel=64
					6, -9, 1, 1, 0, 4, -1, -15, -2,
					-- layer=2 filter=133 channel=65
					0, -11, -10, 11, 6, -8, -13, 0, -4,
					-- layer=2 filter=133 channel=66
					-3, 8, 1, 1, 6, 3, -11, 1, -9,
					-- layer=2 filter=133 channel=67
					-12, -10, -14, 2, -3, -6, -11, -7, -6,
					-- layer=2 filter=133 channel=68
					1, -4, -1, -2, 8, 5, 7, -7, 1,
					-- layer=2 filter=133 channel=69
					5, -11, -1, -12, -3, -15, -4, 2, -11,
					-- layer=2 filter=133 channel=70
					-1, 3, -7, -18, -10, 0, -2, -15, -9,
					-- layer=2 filter=133 channel=71
					-15, -12, -7, -10, -11, -12, -14, -1, 0,
					-- layer=2 filter=133 channel=72
					-9, -7, -17, 5, -5, 10, -12, 5, 2,
					-- layer=2 filter=133 channel=73
					-1, -7, -11, -8, -1, -11, -8, -10, -10,
					-- layer=2 filter=133 channel=74
					5, 6, 0, -7, 0, -6, -5, 0, -1,
					-- layer=2 filter=133 channel=75
					-5, 9, 0, -3, 4, 1, 0, 7, -13,
					-- layer=2 filter=133 channel=76
					7, -4, -13, -9, -2, -7, 15, 6, -2,
					-- layer=2 filter=133 channel=77
					-4, -6, -7, 5, 0, -1, 6, -10, 5,
					-- layer=2 filter=133 channel=78
					-2, -4, -11, 0, -13, -8, 1, 5, -5,
					-- layer=2 filter=133 channel=79
					-11, 0, 7, -9, 2, -6, -1, 9, 7,
					-- layer=2 filter=133 channel=80
					-2, 0, -2, 0, -6, -5, -16, -4, 0,
					-- layer=2 filter=133 channel=81
					-5, 5, 1, 7, -1, 7, -9, 0, 0,
					-- layer=2 filter=133 channel=82
					2, -10, -2, 2, 2, 0, -7, 0, -7,
					-- layer=2 filter=133 channel=83
					-14, 1, 0, 1, 0, -17, -10, -8, -11,
					-- layer=2 filter=133 channel=84
					3, -7, -3, 7, 7, 1, -10, -9, 7,
					-- layer=2 filter=133 channel=85
					-8, -5, -5, -6, 2, -5, 7, 0, -8,
					-- layer=2 filter=133 channel=86
					9, 1, 0, -10, 1, 4, -2, -5, 4,
					-- layer=2 filter=133 channel=87
					2, 1, 0, -8, -5, -6, -8, -10, -17,
					-- layer=2 filter=133 channel=88
					6, -10, -15, 2, 0, -15, 8, -8, -9,
					-- layer=2 filter=133 channel=89
					-2, -3, -13, 7, -7, 3, -4, -9, -7,
					-- layer=2 filter=133 channel=90
					1, -2, -2, -4, -4, -3, -9, 5, -8,
					-- layer=2 filter=133 channel=91
					-12, 5, 7, 6, 1, -11, -7, -14, -11,
					-- layer=2 filter=133 channel=92
					-3, -1, -9, 8, -1, 5, -18, -17, -10,
					-- layer=2 filter=133 channel=93
					-13, 2, 1, 18, 6, -16, -16, 2, -5,
					-- layer=2 filter=133 channel=94
					10, 20, -6, -4, -17, -19, 3, -10, -2,
					-- layer=2 filter=133 channel=95
					4, -3, -7, 6, 0, 0, 8, 8, -3,
					-- layer=2 filter=133 channel=96
					-6, -6, -22, -14, -18, 4, 6, -15, -4,
					-- layer=2 filter=133 channel=97
					-4, -2, -2, -6, -1, -4, 8, 2, -8,
					-- layer=2 filter=133 channel=98
					-9, -6, -17, -18, -4, 16, -11, -18, -2,
					-- layer=2 filter=133 channel=99
					-17, -3, -5, -9, -17, 4, -15, -17, -13,
					-- layer=2 filter=133 channel=100
					4, 5, -5, 16, -1, -12, -8, 6, -10,
					-- layer=2 filter=133 channel=101
					1, -6, -21, 3, -4, -7, -12, -2, -8,
					-- layer=2 filter=133 channel=102
					5, -17, 0, 4, -17, 9, -2, -5, 0,
					-- layer=2 filter=133 channel=103
					-10, 8, 2, -3, 0, 0, -4, 1, -11,
					-- layer=2 filter=133 channel=104
					1, -16, -11, -16, -5, 0, -19, -3, -9,
					-- layer=2 filter=133 channel=105
					-8, -3, -6, 2, -17, 9, 4, -15, -12,
					-- layer=2 filter=133 channel=106
					-13, -8, 0, -6, -14, -18, -17, -7, -3,
					-- layer=2 filter=133 channel=107
					0, 4, -11, 2, 5, -8, 6, -7, 2,
					-- layer=2 filter=133 channel=108
					1, -11, -2, 2, -13, -11, 2, 0, -9,
					-- layer=2 filter=133 channel=109
					6, 1, -9, 0, -11, -10, -4, -5, -2,
					-- layer=2 filter=133 channel=110
					0, -10, -11, -1, -7, -4, 2, -1, -10,
					-- layer=2 filter=133 channel=111
					5, -10, -9, -7, 6, -11, 4, -10, 6,
					-- layer=2 filter=133 channel=112
					-6, -12, -12, -2, -13, -2, -18, -13, 1,
					-- layer=2 filter=133 channel=113
					14, -1, 1, -13, -6, -7, -4, -3, -4,
					-- layer=2 filter=133 channel=114
					8, -6, -8, 7, -4, 2, 2, -3, -9,
					-- layer=2 filter=133 channel=115
					-10, 3, -1, 2, 5, 2, -3, 5, 7,
					-- layer=2 filter=133 channel=116
					-4, -1, -17, -5, 0, 2, 4, -18, -7,
					-- layer=2 filter=133 channel=117
					-13, -16, -25, -17, -2, 6, -7, -7, 3,
					-- layer=2 filter=133 channel=118
					3, 1, -9, -17, 2, -7, 6, -7, 0,
					-- layer=2 filter=133 channel=119
					4, 0, -4, -8, -8, 3, -4, 2, -16,
					-- layer=2 filter=133 channel=120
					6, -1, 0, -1, -2, 5, 7, 6, -1,
					-- layer=2 filter=133 channel=121
					-7, -11, 8, 3, 8, -7, -3, -10, -3,
					-- layer=2 filter=133 channel=122
					0, -2, 0, -6, 6, 2, -9, 6, -9,
					-- layer=2 filter=133 channel=123
					-6, -10, -13, 5, -1, 0, -3, -5, -18,
					-- layer=2 filter=133 channel=124
					-17, -14, -16, -14, -8, -21, -8, -12, -7,
					-- layer=2 filter=133 channel=125
					-4, -3, -8, 3, -6, -2, -10, 2, 0,
					-- layer=2 filter=133 channel=126
					11, -3, -12, 0, 1, -8, 3, -3, 2,
					-- layer=2 filter=133 channel=127
					-12, -9, -1, 2, -11, -3, -2, 0, 1,
					-- layer=2 filter=134 channel=0
					-26, -28, -3, -26, -8, 4, -5, -21, -15,
					-- layer=2 filter=134 channel=1
					28, -3, 5, -2, 25, 12, -13, 9, 14,
					-- layer=2 filter=134 channel=2
					5, 5, 4, -4, 8, -4, 2, 3, -6,
					-- layer=2 filter=134 channel=3
					-9, -38, -20, 13, 0, -19, 11, -16, 5,
					-- layer=2 filter=134 channel=4
					8, 16, 18, -11, 5, 43, 25, 15, -3,
					-- layer=2 filter=134 channel=5
					-7, -12, 1, -17, -12, -3, -6, -11, -21,
					-- layer=2 filter=134 channel=6
					-1, -14, 40, -28, -34, 15, -31, -54, 2,
					-- layer=2 filter=134 channel=7
					-25, 17, 20, 10, 31, -16, 13, -84, -62,
					-- layer=2 filter=134 channel=8
					9, -7, -2, 10, -5, -5, -9, -2, -4,
					-- layer=2 filter=134 channel=9
					-38, -10, 6, -4, -38, -41, 3, 17, 0,
					-- layer=2 filter=134 channel=10
					-52, -45, -21, -15, -14, -2, 3, -13, 0,
					-- layer=2 filter=134 channel=11
					15, 16, 10, 0, 4, -8, -15, -34, -31,
					-- layer=2 filter=134 channel=12
					-7, 18, 52, 25, 31, 1, -28, -5, 43,
					-- layer=2 filter=134 channel=13
					2, -2, -2, -3, 8, 0, 1, 2, 2,
					-- layer=2 filter=134 channel=14
					12, 15, 31, 0, 6, 14, -44, -18, 21,
					-- layer=2 filter=134 channel=15
					-34, 23, 25, -22, -16, -36, 0, 7, -8,
					-- layer=2 filter=134 channel=16
					-18, -7, -42, 39, 45, -18, 40, 49, 7,
					-- layer=2 filter=134 channel=17
					7, 0, 7, 0, 5, -8, -9, -8, -7,
					-- layer=2 filter=134 channel=18
					32, 3, 27, 31, 25, 28, 13, 10, 11,
					-- layer=2 filter=134 channel=19
					24, 10, -11, 8, -16, -9, -15, -4, 23,
					-- layer=2 filter=134 channel=20
					11, 5, -1, -5, -4, -6, -4, -8, -5,
					-- layer=2 filter=134 channel=21
					-5, 16, 5, 9, 7, -1, 8, 0, -6,
					-- layer=2 filter=134 channel=22
					8, 3, 5, 6, -9, -5, -3, -4, -2,
					-- layer=2 filter=134 channel=23
					16, 14, 27, -2, -6, 23, 4, -21, 11,
					-- layer=2 filter=134 channel=24
					-12, 1, -29, -2, -16, 2, 66, -15, 16,
					-- layer=2 filter=134 channel=25
					-17, 15, -13, 18, -7, -28, 12, -7, -23,
					-- layer=2 filter=134 channel=26
					-9, -1, -6, -3, 10, 9, -9, 7, 6,
					-- layer=2 filter=134 channel=27
					16, 23, 0, 16, 15, -25, -15, -2, -29,
					-- layer=2 filter=134 channel=28
					8, 5, 19, -28, 22, 17, -21, 13, 24,
					-- layer=2 filter=134 channel=29
					0, 5, 0, 4, 9, 6, -8, 4, -5,
					-- layer=2 filter=134 channel=30
					-27, -28, -8, -2, -16, 13, 13, 17, 6,
					-- layer=2 filter=134 channel=31
					-63, 14, -14, -16, 20, 33, 23, 26, -48,
					-- layer=2 filter=134 channel=32
					1, 2, -4, -3, 1, -7, 8, 4, 0,
					-- layer=2 filter=134 channel=33
					5, 4, -43, 0, 24, 6, -7, -43, -32,
					-- layer=2 filter=134 channel=34
					-19, 23, 42, -55, 12, 29, 56, 58, 4,
					-- layer=2 filter=134 channel=35
					33, 19, 48, 2, 24, 15, 2, 18, -11,
					-- layer=2 filter=134 channel=36
					6, 9, 17, -3, 13, 3, -11, -7, 3,
					-- layer=2 filter=134 channel=37
					14, 7, -17, -6, 1, -5, -18, -12, -12,
					-- layer=2 filter=134 channel=38
					24, 7, -12, -10, -19, 16, -33, 0, 18,
					-- layer=2 filter=134 channel=39
					-59, -6, 0, -1, 0, -2, 15, 4, 0,
					-- layer=2 filter=134 channel=40
					9, 8, -49, -63, -49, 11, 0, 82, -56,
					-- layer=2 filter=134 channel=41
					-1, 3, -3, 4, -8, -4, 1, 3, 9,
					-- layer=2 filter=134 channel=42
					12, 5, -21, 37, 3, -21, 15, -1, 6,
					-- layer=2 filter=134 channel=43
					-23, -13, -29, -7, 9, -37, 14, 15, -12,
					-- layer=2 filter=134 channel=44
					-3, 8, -10, -5, -1, -7, -1, 0, 2,
					-- layer=2 filter=134 channel=45
					29, 46, -18, -21, 23, 12, 21, 2, -53,
					-- layer=2 filter=134 channel=46
					-64, -31, -6, 17, -4, 10, -13, 0, 18,
					-- layer=2 filter=134 channel=47
					-26, -11, -51, -18, 9, 31, -16, -18, -9,
					-- layer=2 filter=134 channel=48
					6, -2, 3, -8, 7, -2, -5, 4, -9,
					-- layer=2 filter=134 channel=49
					-13, -7, 8, 33, 17, 9, 10, -23, -25,
					-- layer=2 filter=134 channel=50
					-1, -9, 2, 7, 5, 4, -10, 0, 11,
					-- layer=2 filter=134 channel=51
					16, 12, 8, -14, 4, 0, -11, -8, -22,
					-- layer=2 filter=134 channel=52
					-25, -52, -28, -40, -6, 16, -50, -40, -15,
					-- layer=2 filter=134 channel=53
					-35, 20, -46, -18, -19, -44, -53, 5, -25,
					-- layer=2 filter=134 channel=54
					27, 25, 21, -9, -5, 2, 7, -10, -14,
					-- layer=2 filter=134 channel=55
					7, -1, 3, 0, 0, -3, 9, 1, 12,
					-- layer=2 filter=134 channel=56
					-17, 5, 13, 1, 12, -11, -33, -30, -28,
					-- layer=2 filter=134 channel=57
					6, -10, -13, -1, -10, 7, -5, -7, -2,
					-- layer=2 filter=134 channel=58
					0, 6, 42, 5, 39, 11, -34, -10, 21,
					-- layer=2 filter=134 channel=59
					5, -26, -12, -3, 32, 35, -17, -11, 44,
					-- layer=2 filter=134 channel=60
					25, 30, -4, 34, -56, 11, -45, 29, 38,
					-- layer=2 filter=134 channel=61
					7, -1, 13, 27, -30, -17, -1, -73, -44,
					-- layer=2 filter=134 channel=62
					12, 15, 47, 19, -16, 3, 35, -19, -17,
					-- layer=2 filter=134 channel=63
					-33, -36, -12, -5, -3, 1, -19, -4, -3,
					-- layer=2 filter=134 channel=64
					10, 18, 19, 8, 8, 16, 20, 19, -9,
					-- layer=2 filter=134 channel=65
					16, -24, -5, -3, -1, 36, -49, -87, -10,
					-- layer=2 filter=134 channel=66
					-29, 21, 6, 69, 12, 16, 13, -17, -7,
					-- layer=2 filter=134 channel=67
					-71, -44, 3, -15, -69, -6, 5, 7, 17,
					-- layer=2 filter=134 channel=68
					-10, 8, -1, 2, 5, 0, 8, 4, -6,
					-- layer=2 filter=134 channel=69
					0, -4, 19, 24, 16, 4, 26, 39, -22,
					-- layer=2 filter=134 channel=70
					23, 27, 25, -1, 5, -7, -14, 8, -9,
					-- layer=2 filter=134 channel=71
					40, 54, 12, 32, 12, -28, -24, 14, -25,
					-- layer=2 filter=134 channel=72
					-16, 1, 43, 20, 24, 23, 0, -11, 13,
					-- layer=2 filter=134 channel=73
					0, 42, -17, -7, -12, -10, 33, 25, 8,
					-- layer=2 filter=134 channel=74
					-56, -34, -31, -26, -31, 28, -13, 4, 18,
					-- layer=2 filter=134 channel=75
					22, 3, -21, 0, 28, 3, -28, -30, 9,
					-- layer=2 filter=134 channel=76
					-16, 61, 11, -15, -1, -39, -20, 15, -78,
					-- layer=2 filter=134 channel=77
					1, 6, -8, 0, -1, 0, -4, 6, 11,
					-- layer=2 filter=134 channel=78
					12, 11, 21, 0, 22, 27, 8, -9, 0,
					-- layer=2 filter=134 channel=79
					-8, -6, 10, 1, -1, 0, -8, 2, 5,
					-- layer=2 filter=134 channel=80
					-54, -19, -21, 15, -23, -21, 7, 5, 12,
					-- layer=2 filter=134 channel=81
					-5, -7, -4, 3, 5, 9, 9, -5, -1,
					-- layer=2 filter=134 channel=82
					-1, 0, 5, 7, -6, 6, 10, -3, -9,
					-- layer=2 filter=134 channel=83
					20, 2, -1, 6, 11, -9, -6, 6, 35,
					-- layer=2 filter=134 channel=84
					-8, 3, 3, -9, 6, 0, -2, -3, -4,
					-- layer=2 filter=134 channel=85
					14, 3, 0, 4, -1, 15, 5, -9, -1,
					-- layer=2 filter=134 channel=86
					7, -4, -6, 8, 6, -7, 6, 6, -7,
					-- layer=2 filter=134 channel=87
					48, -3, 47, 45, 22, -2, 69, 44, 17,
					-- layer=2 filter=134 channel=88
					1, -11, -5, -19, -13, 6, 5, 27, -24,
					-- layer=2 filter=134 channel=89
					-24, -12, 36, 28, 14, 3, -31, 3, 55,
					-- layer=2 filter=134 channel=90
					-6, -10, -5, -8, 7, -4, 9, 8, -5,
					-- layer=2 filter=134 channel=91
					-10, 1, 11, -2, 32, 0, -28, 26, 41,
					-- layer=2 filter=134 channel=92
					14, -9, 34, 20, 27, -1, -32, 15, 43,
					-- layer=2 filter=134 channel=93
					21, 13, 9, -13, -13, 10, -6, -10, -4,
					-- layer=2 filter=134 channel=94
					-48, -4, 7, 16, -13, -37, -38, -81, -17,
					-- layer=2 filter=134 channel=95
					-6, -13, -6, 1, 0, -5, -8, -9, -7,
					-- layer=2 filter=134 channel=96
					-11, -8, -36, -22, -58, -6, -57, -24, 34,
					-- layer=2 filter=134 channel=97
					-19, -34, -38, 9, -2, 6, 20, -9, -12,
					-- layer=2 filter=134 channel=98
					6, 14, 6, -33, 12, 8, -10, -30, 11,
					-- layer=2 filter=134 channel=99
					-6, -25, -15, -37, 1, -34, -12, -62, -27,
					-- layer=2 filter=134 channel=100
					4, 18, -8, 33, 11, -1, -31, 34, 31,
					-- layer=2 filter=134 channel=101
					-10, 25, -8, -24, -15, -26, -25, -13, -24,
					-- layer=2 filter=134 channel=102
					19, 7, 28, 24, 17, 23, -16, -10, 46,
					-- layer=2 filter=134 channel=103
					-5, -50, 0, -14, 22, 15, 11, 93, 8,
					-- layer=2 filter=134 channel=104
					-18, -11, 8, 15, 9, 2, -11, -7, -22,
					-- layer=2 filter=134 channel=105
					-15, 4, -6, 26, 35, -11, -12, 5, -14,
					-- layer=2 filter=134 channel=106
					-43, 14, 8, -9, -17, -12, -20, -14, -3,
					-- layer=2 filter=134 channel=107
					-9, -23, -18, 50, -13, -23, 9, 26, 18,
					-- layer=2 filter=134 channel=108
					13, 8, -5, -4, 7, -42, -16, -24, 7,
					-- layer=2 filter=134 channel=109
					7, -6, 5, 0, 8, -10, -4, 4, 1,
					-- layer=2 filter=134 channel=110
					4, -18, -31, 13, 22, -20, 35, 23, -3,
					-- layer=2 filter=134 channel=111
					-4, -6, 5, 9, 1, -5, 2, 4, -5,
					-- layer=2 filter=134 channel=112
					16, 11, 10, -29, -20, -11, 8, -29, -44,
					-- layer=2 filter=134 channel=113
					-24, 3, 9, -29, 12, 15, -9, -11, 8,
					-- layer=2 filter=134 channel=114
					-6, 0, -8, -8, 11, 0, -9, 18, -6,
					-- layer=2 filter=134 channel=115
					-5, 7, -5, -1, -4, 6, 3, -8, 10,
					-- layer=2 filter=134 channel=116
					2, -9, 30, 11, -11, -18, 40, 36, 18,
					-- layer=2 filter=134 channel=117
					-5, 22, 6, -44, -34, -9, 2, 0, -23,
					-- layer=2 filter=134 channel=118
					-29, -20, -22, -6, -6, -10, 20, 17, -13,
					-- layer=2 filter=134 channel=119
					2, -1, -4, 12, 41, 8, 37, 34, -23,
					-- layer=2 filter=134 channel=120
					0, 5, -1, 6, 8, 8, 4, 8, 6,
					-- layer=2 filter=134 channel=121
					10, -4, 0, 1, -4, -11, -10, 0, -9,
					-- layer=2 filter=134 channel=122
					11, -17, -13, 8, -15, 6, -5, 4, -5,
					-- layer=2 filter=134 channel=123
					0, -34, 1, 18, 24, 7, 6, -41, -8,
					-- layer=2 filter=134 channel=124
					-1, 24, 10, -10, 15, -58, 38, 23, 43,
					-- layer=2 filter=134 channel=125
					2, 11, -2, 1, -8, 6, 9, -12, 5,
					-- layer=2 filter=134 channel=126
					0, 28, -58, 31, -107, 9, 22, 26, 33,
					-- layer=2 filter=134 channel=127
					8, -11, 19, -9, 7, 50, 0, 14, 25,
					-- layer=2 filter=135 channel=0
					-3, -7, -3, 1, -6, 2, 8, 5, -6,
					-- layer=2 filter=135 channel=1
					-8, 3, -5, 1, -6, -12, 0, 9, -8,
					-- layer=2 filter=135 channel=2
					6, 2, 1, 1, 2, 3, -5, 7, -10,
					-- layer=2 filter=135 channel=3
					-8, -4, 8, -8, 1, 2, 0, -7, 0,
					-- layer=2 filter=135 channel=4
					9, 7, 6, 3, 8, -6, 1, 3, 10,
					-- layer=2 filter=135 channel=5
					2, -11, 3, -4, -13, -2, -7, 4, 3,
					-- layer=2 filter=135 channel=6
					4, -5, -8, -7, -5, -3, -2, 3, -3,
					-- layer=2 filter=135 channel=7
					-2, -8, 0, 0, 1, -6, -8, -1, -8,
					-- layer=2 filter=135 channel=8
					-1, 9, 4, -9, -9, -7, 1, -3, 6,
					-- layer=2 filter=135 channel=9
					-6, 5, 1, -3, -11, 0, 5, -6, 3,
					-- layer=2 filter=135 channel=10
					-13, -5, -1, -12, -3, -1, -14, 1, -4,
					-- layer=2 filter=135 channel=11
					-5, 1, 10, -8, 2, -10, -3, 6, -5,
					-- layer=2 filter=135 channel=12
					-11, 2, 0, -2, 4, -5, -3, 0, -3,
					-- layer=2 filter=135 channel=13
					-5, 7, 4, 6, 2, -1, -6, -9, -8,
					-- layer=2 filter=135 channel=14
					-4, -5, 3, 3, -3, -12, 3, -5, -8,
					-- layer=2 filter=135 channel=15
					-8, 2, 3, -8, 2, 1, -1, 6, -6,
					-- layer=2 filter=135 channel=16
					-5, -11, -4, 1, -10, -3, -9, 1, -7,
					-- layer=2 filter=135 channel=17
					-4, -5, -2, 4, 4, 8, 5, -8, 8,
					-- layer=2 filter=135 channel=18
					-1, -5, 10, -14, 5, 9, -13, -6, -6,
					-- layer=2 filter=135 channel=19
					-7, -2, 11, 5, 8, -1, -2, -8, -9,
					-- layer=2 filter=135 channel=20
					-7, -4, -11, -3, 4, 0, -8, 5, 5,
					-- layer=2 filter=135 channel=21
					0, 0, 4, 3, 8, -2, 1, 7, 5,
					-- layer=2 filter=135 channel=22
					0, -4, -3, 0, -7, 8, -1, 3, -5,
					-- layer=2 filter=135 channel=23
					-4, -8, -5, -5, -3, -12, 0, 0, 6,
					-- layer=2 filter=135 channel=24
					-2, 0, -4, -1, -12, 3, 6, -12, -8,
					-- layer=2 filter=135 channel=25
					2, -7, -9, -4, 8, 9, -7, -10, 0,
					-- layer=2 filter=135 channel=26
					-3, -6, 7, 0, 0, 7, -6, 10, -8,
					-- layer=2 filter=135 channel=27
					-15, 0, -10, 3, -8, -7, -10, -10, -13,
					-- layer=2 filter=135 channel=28
					0, -6, 2, -6, -16, -8, 6, -10, 0,
					-- layer=2 filter=135 channel=29
					8, -9, -4, -3, -3, 1, 2, 8, 5,
					-- layer=2 filter=135 channel=30
					-6, 0, 4, -7, -2, -5, -14, 2, 6,
					-- layer=2 filter=135 channel=31
					-1, -1, -7, 3, -8, -7, -6, 8, 4,
					-- layer=2 filter=135 channel=32
					-5, 0, 8, -11, -8, -10, -6, 0, -7,
					-- layer=2 filter=135 channel=33
					3, 1, -4, -1, 3, 5, 4, -9, -8,
					-- layer=2 filter=135 channel=34
					-8, -2, 0, 0, 0, -1, -7, -7, -10,
					-- layer=2 filter=135 channel=35
					-18, -9, -7, -3, -14, -8, 0, 6, 9,
					-- layer=2 filter=135 channel=36
					0, 1, -10, 3, 3, -8, 2, 3, -3,
					-- layer=2 filter=135 channel=37
					-3, -7, -3, 0, -12, 5, 6, 5, -8,
					-- layer=2 filter=135 channel=38
					-4, 0, 5, -6, -6, 2, 0, -6, -8,
					-- layer=2 filter=135 channel=39
					2, -2, -2, -9, -9, -3, -2, -2, -13,
					-- layer=2 filter=135 channel=40
					5, -7, 9, 1, 0, -8, 4, 2, -1,
					-- layer=2 filter=135 channel=41
					-1, -5, -5, -5, -9, -5, -1, 7, 1,
					-- layer=2 filter=135 channel=42
					1, -2, 8, -6, 5, 1, -9, -5, -3,
					-- layer=2 filter=135 channel=43
					-8, -12, -5, 2, 5, -4, -1, -5, 0,
					-- layer=2 filter=135 channel=44
					4, 6, 6, 4, -3, -6, 2, -5, -9,
					-- layer=2 filter=135 channel=45
					-6, 5, -2, -2, -8, 9, -8, 5, 0,
					-- layer=2 filter=135 channel=46
					3, -14, -2, 6, -13, -7, 0, 2, -12,
					-- layer=2 filter=135 channel=47
					2, -4, -2, -13, 3, 0, -6, 1, -1,
					-- layer=2 filter=135 channel=48
					-3, -1, 8, -2, -9, 2, -5, -8, 5,
					-- layer=2 filter=135 channel=49
					-2, -18, -3, -10, 2, 6, -9, -3, 9,
					-- layer=2 filter=135 channel=50
					3, -6, 11, -3, 0, 0, 2, 0, -8,
					-- layer=2 filter=135 channel=51
					6, 3, 5, -4, 0, 4, -2, -4, -11,
					-- layer=2 filter=135 channel=52
					-6, -4, 4, 5, -9, -4, 5, -5, -6,
					-- layer=2 filter=135 channel=53
					-3, -8, -9, 11, 1, 6, -12, 0, -3,
					-- layer=2 filter=135 channel=54
					-5, -2, 2, 3, 1, -11, -9, -7, -1,
					-- layer=2 filter=135 channel=55
					-2, 0, 4, -1, 4, -7, 7, 3, 8,
					-- layer=2 filter=135 channel=56
					6, -13, 4, -12, 5, 0, -4, 8, 3,
					-- layer=2 filter=135 channel=57
					-4, 8, 2, -3, 0, 7, -1, 0, 10,
					-- layer=2 filter=135 channel=58
					-11, -2, -6, 9, 2, -11, 1, 0, 7,
					-- layer=2 filter=135 channel=59
					-6, 0, -9, -3, -2, -5, 1, -8, -2,
					-- layer=2 filter=135 channel=60
					0, -6, -14, 5, 6, -5, -6, -4, -3,
					-- layer=2 filter=135 channel=61
					8, -10, 0, -1, 0, -5, -11, -2, -6,
					-- layer=2 filter=135 channel=62
					1, -11, -8, 3, 1, -5, 9, 1, -3,
					-- layer=2 filter=135 channel=63
					2, -8, 3, -7, -8, -17, -6, -8, -9,
					-- layer=2 filter=135 channel=64
					-5, 4, -2, -9, -5, -9, -1, 2, 7,
					-- layer=2 filter=135 channel=65
					-8, -4, -7, 4, 1, -13, -4, 4, 1,
					-- layer=2 filter=135 channel=66
					7, -10, 7, -7, -8, -12, 6, 1, 1,
					-- layer=2 filter=135 channel=67
					-12, -11, -2, -5, -4, 5, 5, -3, 8,
					-- layer=2 filter=135 channel=68
					0, -7, -2, -3, 8, -9, -6, 7, -8,
					-- layer=2 filter=135 channel=69
					-10, 9, 6, -2, 3, -9, -10, -7, -6,
					-- layer=2 filter=135 channel=70
					-8, -12, -13, -6, -11, 9, -9, -16, -12,
					-- layer=2 filter=135 channel=71
					1, -8, 4, -1, -3, 7, 2, 5, 9,
					-- layer=2 filter=135 channel=72
					-11, -9, 2, -13, -15, -13, -14, -11, 0,
					-- layer=2 filter=135 channel=73
					-2, 2, 6, -8, 2, -1, -2, 3, -17,
					-- layer=2 filter=135 channel=74
					4, 1, 0, -8, 6, -4, 0, -2, -6,
					-- layer=2 filter=135 channel=75
					-6, 0, -7, 4, -3, -1, 7, -11, 2,
					-- layer=2 filter=135 channel=76
					-9, -6, -6, 5, 7, -11, 1, 8, 3,
					-- layer=2 filter=135 channel=77
					8, 0, 4, 4, 5, 0, -7, 4, 0,
					-- layer=2 filter=135 channel=78
					8, 1, 5, 0, 5, 4, -10, 7, -11,
					-- layer=2 filter=135 channel=79
					5, -10, -11, 9, -1, -7, 8, 3, 0,
					-- layer=2 filter=135 channel=80
					-6, 6, 6, 5, 2, -4, -11, 1, 7,
					-- layer=2 filter=135 channel=81
					6, -10, -4, -9, -2, 7, -5, 5, -1,
					-- layer=2 filter=135 channel=82
					0, -5, 2, 0, 7, -1, -9, 0, -3,
					-- layer=2 filter=135 channel=83
					3, 8, -10, -7, -2, -10, -6, 7, 7,
					-- layer=2 filter=135 channel=84
					0, -4, -7, 4, -3, 6, -9, 0, 1,
					-- layer=2 filter=135 channel=85
					-7, 1, 4, -11, -7, -8, -6, 0, 2,
					-- layer=2 filter=135 channel=86
					6, 1, -7, 3, -4, 8, -5, 0, 4,
					-- layer=2 filter=135 channel=87
					-9, -4, -11, 3, -11, -1, -10, -11, -9,
					-- layer=2 filter=135 channel=88
					0, -13, -14, -6, 5, 2, 2, -4, 1,
					-- layer=2 filter=135 channel=89
					-5, 6, 0, -6, 1, -1, -12, 3, -9,
					-- layer=2 filter=135 channel=90
					0, 1, -9, -5, -10, 5, -6, -9, -9,
					-- layer=2 filter=135 channel=91
					-4, -9, 2, 4, -7, -8, 1, -4, -10,
					-- layer=2 filter=135 channel=92
					2, -8, 3, -8, 0, -19, 0, 2, -3,
					-- layer=2 filter=135 channel=93
					6, -4, -10, -7, -7, -9, -11, -7, -7,
					-- layer=2 filter=135 channel=94
					-6, -10, -2, 7, -1, -3, -5, -5, 2,
					-- layer=2 filter=135 channel=95
					-8, -2, 5, -11, 0, 0, 0, -5, -8,
					-- layer=2 filter=135 channel=96
					2, -9, -10, 3, -1, 6, -5, -2, -3,
					-- layer=2 filter=135 channel=97
					4, -7, -2, 7, -4, -7, 2, -10, -9,
					-- layer=2 filter=135 channel=98
					-10, 6, 0, -15, -15, -8, 0, -4, -5,
					-- layer=2 filter=135 channel=99
					-2, -7, -11, 5, 4, 0, 6, -1, -1,
					-- layer=2 filter=135 channel=100
					1, -1, 0, -5, -12, 2, -3, -4, 0,
					-- layer=2 filter=135 channel=101
					7, -11, 7, 1, -8, -2, -6, 6, 6,
					-- layer=2 filter=135 channel=102
					-2, -2, -6, -4, -3, 5, 0, 5, -4,
					-- layer=2 filter=135 channel=103
					-10, 1, -9, -3, -2, -1, 4, -8, 8,
					-- layer=2 filter=135 channel=104
					-8, 7, -7, -1, -8, -6, 0, 2, 9,
					-- layer=2 filter=135 channel=105
					-3, 5, 7, -1, -4, 5, -4, 2, -3,
					-- layer=2 filter=135 channel=106
					-1, -10, -2, 3, -5, 3, -2, 2, 2,
					-- layer=2 filter=135 channel=107
					-11, 1, -3, -5, 6, 4, -7, 0, 1,
					-- layer=2 filter=135 channel=108
					-2, 3, -5, 3, -6, 0, -6, 3, -3,
					-- layer=2 filter=135 channel=109
					-11, -11, 8, -1, 5, -3, 0, 0, -2,
					-- layer=2 filter=135 channel=110
					-8, 0, 4, -8, 3, -12, -2, -5, -14,
					-- layer=2 filter=135 channel=111
					-2, -9, 4, 1, -5, 2, 5, -5, 3,
					-- layer=2 filter=135 channel=112
					-11, 0, 5, -11, 0, 0, -10, -1, 0,
					-- layer=2 filter=135 channel=113
					-11, -7, 0, 9, -8, -9, -4, -5, -6,
					-- layer=2 filter=135 channel=114
					5, 10, -7, 0, -6, -3, -11, -6, -10,
					-- layer=2 filter=135 channel=115
					0, 0, 8, 6, -3, -6, -7, 1, 7,
					-- layer=2 filter=135 channel=116
					6, 3, 6, -9, -6, 1, -3, 4, 5,
					-- layer=2 filter=135 channel=117
					5, -10, 10, 9, -7, -6, 4, -9, -8,
					-- layer=2 filter=135 channel=118
					0, -12, -8, -11, -6, 1, -3, 0, -10,
					-- layer=2 filter=135 channel=119
					3, -8, -2, -9, -3, 7, -11, 0, -3,
					-- layer=2 filter=135 channel=120
					-3, -3, -5, 6, 3, 9, -9, -6, 3,
					-- layer=2 filter=135 channel=121
					-9, -5, -8, -3, 2, -3, -5, 8, 0,
					-- layer=2 filter=135 channel=122
					-4, 7, -6, -3, 8, -6, 8, 5, -7,
					-- layer=2 filter=135 channel=123
					-3, -6, -6, -13, 2, 1, 10, -5, -12,
					-- layer=2 filter=135 channel=124
					-8, 5, 0, -11, -10, 2, 6, 7, 1,
					-- layer=2 filter=135 channel=125
					0, 1, -5, -2, -8, 5, 6, 8, 6,
					-- layer=2 filter=135 channel=126
					6, -9, -10, -5, -5, -1, -7, -10, 0,
					-- layer=2 filter=135 channel=127
					-6, -9, 2, -1, 0, -8, -7, 9, 3,
					-- layer=2 filter=136 channel=0
					17, 27, 14, 22, -18, -18, -23, -17, 0,
					-- layer=2 filter=136 channel=1
					-19, -16, -48, 13, -8, -10, 16, -2, 17,
					-- layer=2 filter=136 channel=2
					4, -3, -1, -1, -2, -2, -2, -1, -9,
					-- layer=2 filter=136 channel=3
					-1, 9, -2, -21, -52, -15, 2, 33, 44,
					-- layer=2 filter=136 channel=4
					2, -1, -30, 6, 1, -56, -15, -9, -23,
					-- layer=2 filter=136 channel=5
					3, -10, 1, 31, 12, -24, -31, -6, 8,
					-- layer=2 filter=136 channel=6
					20, -3, 37, -7, -2, 7, -34, -22, -45,
					-- layer=2 filter=136 channel=7
					-34, -49, -25, -80, -50, -6, -23, -41, -53,
					-- layer=2 filter=136 channel=8
					5, 8, 10, 1, 4, -7, 6, 11, -10,
					-- layer=2 filter=136 channel=9
					6, -25, -13, -35, 3, -47, -25, -89, 25,
					-- layer=2 filter=136 channel=10
					12, 39, 16, -12, -5, -45, -2, 16, 40,
					-- layer=2 filter=136 channel=11
					-5, 4, -13, 7, 24, 17, 2, -3, -6,
					-- layer=2 filter=136 channel=12
					-37, -28, -37, 1, -3, -53, 7, 1, -11,
					-- layer=2 filter=136 channel=13
					7, 0, 4, 8, -8, -3, 8, -1, -2,
					-- layer=2 filter=136 channel=14
					-25, -46, -48, 10, 9, -24, 43, 16, -10,
					-- layer=2 filter=136 channel=15
					-38, 27, 9, 3, -5, 62, 16, 18, 27,
					-- layer=2 filter=136 channel=16
					44, 16, 14, 7, 13, -31, -17, -13, -18,
					-- layer=2 filter=136 channel=17
					8, 3, 8, -1, 5, -4, -1, -9, 0,
					-- layer=2 filter=136 channel=18
					-18, -18, -39, -38, -27, -9, -25, 13, 13,
					-- layer=2 filter=136 channel=19
					-3, 3, -3, -9, 37, 3, 45, -5, 20,
					-- layer=2 filter=136 channel=20
					7, 0, 0, 8, 0, 7, 3, -8, 1,
					-- layer=2 filter=136 channel=21
					13, 10, 7, 6, 0, -6, 0, 12, -11,
					-- layer=2 filter=136 channel=22
					2, 1, -3, -2, -8, -3, 7, -8, -4,
					-- layer=2 filter=136 channel=23
					19, 11, 21, 1, 4, -13, -24, -24, -21,
					-- layer=2 filter=136 channel=24
					26, 43, 5, -4, -17, -40, -15, 23, 18,
					-- layer=2 filter=136 channel=25
					24, 43, 4, 8, 4, -26, 9, 30, 3,
					-- layer=2 filter=136 channel=26
					10, 2, -11, 0, 8, 7, -11, -7, -1,
					-- layer=2 filter=136 channel=27
					-19, -11, -24, 47, 6, -8, 32, -24, -4,
					-- layer=2 filter=136 channel=28
					-13, 34, -11, -19, -21, -19, 17, 22, -23,
					-- layer=2 filter=136 channel=29
					-7, 9, 4, 2, 9, 8, 8, -4, -9,
					-- layer=2 filter=136 channel=30
					-3, -26, -8, 25, -12, -24, 0, -31, 2,
					-- layer=2 filter=136 channel=31
					15, -35, -54, -3, -27, -6, -19, 9, -35,
					-- layer=2 filter=136 channel=32
					-8, 0, -4, -6, -4, -7, -1, 6, -7,
					-- layer=2 filter=136 channel=33
					-33, -24, 33, 3, 4, 57, -19, 31, 0,
					-- layer=2 filter=136 channel=34
					6, 11, 67, 38, 58, 54, 36, 59, 22,
					-- layer=2 filter=136 channel=35
					-45, -23, -1, -47, -28, 30, 41, 20, 1,
					-- layer=2 filter=136 channel=36
					-10, -8, -1, 5, -11, 5, 6, -12, 19,
					-- layer=2 filter=136 channel=37
					-3, -5, -8, 7, 8, -1, -5, -4, 1,
					-- layer=2 filter=136 channel=38
					-30, -9, 15, 25, 16, 36, 15, -16, 1,
					-- layer=2 filter=136 channel=39
					26, 56, 51, 8, 19, 20, -42, -38, 8,
					-- layer=2 filter=136 channel=40
					-1, 46, -31, -22, -12, -3, 0, 33, 2,
					-- layer=2 filter=136 channel=41
					-9, 9, -11, -4, -2, 8, -4, 5, 3,
					-- layer=2 filter=136 channel=42
					25, 15, 1, -3, -13, -11, 12, -13, 21,
					-- layer=2 filter=136 channel=43
					-26, 54, 4, -12, -74, -3, -35, 2, 62,
					-- layer=2 filter=136 channel=44
					0, 0, 3, 1, -2, 4, -3, -9, 2,
					-- layer=2 filter=136 channel=45
					12, 28, -18, 23, -51, -51, 27, -40, -31,
					-- layer=2 filter=136 channel=46
					-7, 17, -1, 33, -8, 3, -9, -39, 17,
					-- layer=2 filter=136 channel=47
					19, 47, 25, -2, -74, -25, -42, -32, -43,
					-- layer=2 filter=136 channel=48
					-5, -4, 9, -7, 8, 4, -3, 8, 5,
					-- layer=2 filter=136 channel=49
					-24, -23, -48, -54, -9, -27, -10, -28, -24,
					-- layer=2 filter=136 channel=50
					3, 6, -11, 19, -6, -4, 1, -3, 0,
					-- layer=2 filter=136 channel=51
					22, 11, 13, 12, -11, 10, 6, -1, -12,
					-- layer=2 filter=136 channel=52
					-1, 9, -25, 17, 12, 54, -17, -10, 22,
					-- layer=2 filter=136 channel=53
					-32, -60, -82, 2, 43, -56, -22, -44, -49,
					-- layer=2 filter=136 channel=54
					-33, 10, -28, -13, 13, 50, 8, 16, 23,
					-- layer=2 filter=136 channel=55
					12, -2, -2, -4, 4, 2, 9, 4, 6,
					-- layer=2 filter=136 channel=56
					15, 9, 1, 18, 14, 5, -39, -23, -4,
					-- layer=2 filter=136 channel=57
					-16, 11, 15, -6, 3, -10, 0, 6, -7,
					-- layer=2 filter=136 channel=58
					-4, -13, -3, 26, 47, -32, 20, 40, 36,
					-- layer=2 filter=136 channel=59
					-21, 13, 41, 33, 43, 66, 75, 48, 31,
					-- layer=2 filter=136 channel=60
					17, 20, 22, 11, 50, 30, 46, 67, -32,
					-- layer=2 filter=136 channel=61
					3, -31, -39, -46, -13, -45, -50, -34, -58,
					-- layer=2 filter=136 channel=62
					2, -33, 5, 12, 7, 22, 22, 9, -7,
					-- layer=2 filter=136 channel=63
					19, 19, 0, -25, 24, -3, -49, -36, -15,
					-- layer=2 filter=136 channel=64
					57, 38, 14, -29, 20, -44, 2, -7, -4,
					-- layer=2 filter=136 channel=65
					20, -25, 0, -12, -22, 10, -1, -54, -72,
					-- layer=2 filter=136 channel=66
					32, -12, 8, 34, -29, 15, 34, 25, 36,
					-- layer=2 filter=136 channel=67
					-5, -3, -34, 5, -1, -55, 1, -39, 19,
					-- layer=2 filter=136 channel=68
					2, -8, 8, 10, 7, 0, 0, -3, 11,
					-- layer=2 filter=136 channel=69
					42, 24, 7, 10, 0, -21, 14, 3, -8,
					-- layer=2 filter=136 channel=70
					-17, -7, 12, -5, -8, 32, 5, -9, -5,
					-- layer=2 filter=136 channel=71
					-47, -19, -22, 36, 25, -3, 13, 9, 10,
					-- layer=2 filter=136 channel=72
					-40, -42, -25, -35, -44, 18, 29, 11, -20,
					-- layer=2 filter=136 channel=73
					-75, -13, 17, -69, -7, 17, 19, 14, 0,
					-- layer=2 filter=136 channel=74
					-11, 14, -13, 3, 15, -5, 4, 29, 0,
					-- layer=2 filter=136 channel=75
					-29, -31, -34, -20, -14, -103, 55, -10, -77,
					-- layer=2 filter=136 channel=76
					-15, -61, -70, -32, 3, -28, -60, -60, 10,
					-- layer=2 filter=136 channel=77
					-6, 3, 7, -6, -2, 1, 7, -4, 4,
					-- layer=2 filter=136 channel=78
					-17, 6, -17, -24, -13, 12, -14, -23, -8,
					-- layer=2 filter=136 channel=79
					9, 4, 10, 9, -8, -2, -11, 7, 0,
					-- layer=2 filter=136 channel=80
					21, 29, 9, 5, 14, -19, -2, 19, 21,
					-- layer=2 filter=136 channel=81
					6, -8, 11, 13, -2, 2, 4, -12, -6,
					-- layer=2 filter=136 channel=82
					3, -11, 2, -4, -8, 8, -7, 0, 7,
					-- layer=2 filter=136 channel=83
					14, 40, -12, 37, 28, -28, -17, 20, -37,
					-- layer=2 filter=136 channel=84
					7, 9, 9, 8, 7, 1, -3, 0, -11,
					-- layer=2 filter=136 channel=85
					15, -2, 22, 1, 17, 3, 15, 1, -5,
					-- layer=2 filter=136 channel=86
					-14, -18, -7, -1, -2, 0, 6, 1, 3,
					-- layer=2 filter=136 channel=87
					-34, 51, 22, 28, 46, 65, 51, 33, 45,
					-- layer=2 filter=136 channel=88
					19, 17, -6, 8, 14, -13, -2, 2, -48,
					-- layer=2 filter=136 channel=89
					-30, -13, 2, 11, 34, -28, 57, 35, 3,
					-- layer=2 filter=136 channel=90
					0, 2, 0, -5, 5, 9, 6, -6, 12,
					-- layer=2 filter=136 channel=91
					-35, -41, -18, 4, 15, -21, 45, 31, -18,
					-- layer=2 filter=136 channel=92
					-11, -28, -20, 10, -9, -1, 17, -10, 27,
					-- layer=2 filter=136 channel=93
					15, -27, 5, -6, 46, 8, -23, -6, -20,
					-- layer=2 filter=136 channel=94
					-43, -21, -39, -19, -22, -15, -16, -19, -11,
					-- layer=2 filter=136 channel=95
					4, 0, 5, 12, -9, -12, -12, -9, -4,
					-- layer=2 filter=136 channel=96
					38, 10, -19, 35, 44, 18, 13, -24, -9,
					-- layer=2 filter=136 channel=97
					-14, 0, -18, -2, 10, -30, -21, -27, 8,
					-- layer=2 filter=136 channel=98
					-20, 3, -18, -47, -35, -2, -7, -9, -10,
					-- layer=2 filter=136 channel=99
					-26, -21, 4, 19, 33, 3, 37, -1, 43,
					-- layer=2 filter=136 channel=100
					-69, -17, 21, 1, 37, 2, 36, 59, 49,
					-- layer=2 filter=136 channel=101
					-8, -30, -32, 8, 5, -3, 4, -3, 48,
					-- layer=2 filter=136 channel=102
					39, 0, -36, 7, -2, -5, 15, -35, -13,
					-- layer=2 filter=136 channel=103
					-27, 3, -32, -20, -13, -45, -20, -45, -32,
					-- layer=2 filter=136 channel=104
					-84, -20, -52, -13, -12, -18, -20, -10, 8,
					-- layer=2 filter=136 channel=105
					5, -34, -33, 2, -16, -4, 21, 16, -43,
					-- layer=2 filter=136 channel=106
					35, 34, -19, 49, 28, -23, 20, 20, -6,
					-- layer=2 filter=136 channel=107
					-69, -13, 10, -58, 11, -12, 13, 0, -83,
					-- layer=2 filter=136 channel=108
					15, -11, -47, 34, 35, -7, 25, -57, -31,
					-- layer=2 filter=136 channel=109
					12, 8, -7, 2, 12, 6, 1, 10, -1,
					-- layer=2 filter=136 channel=110
					15, 55, 23, -38, 15, -33, -18, 6, -9,
					-- layer=2 filter=136 channel=111
					0, -8, -3, -8, -4, -9, 9, 10, 0,
					-- layer=2 filter=136 channel=112
					15, -14, -23, -24, -33, -44, -4, -57, -48,
					-- layer=2 filter=136 channel=113
					-5, -20, -13, -3, -7, -32, -45, -58, -8,
					-- layer=2 filter=136 channel=114
					5, -11, 5, -5, 10, -2, -8, 3, 9,
					-- layer=2 filter=136 channel=115
					0, 6, 8, 5, 3, -4, 6, -10, 10,
					-- layer=2 filter=136 channel=116
					20, 14, 3, 34, -6, 36, 40, 21, 31,
					-- layer=2 filter=136 channel=117
					-32, -56, -54, -62, -66, -43, 3, -34, -43,
					-- layer=2 filter=136 channel=118
					6, 29, -1, -17, -39, 14, -45, 4, 50,
					-- layer=2 filter=136 channel=119
					2, -13, -6, 50, -43, 1, 26, 26, -18,
					-- layer=2 filter=136 channel=120
					-9, 8, 5, 0, -1, 5, -2, 10, 7,
					-- layer=2 filter=136 channel=121
					-1, 9, 0, 3, 2, -3, 8, 2, 6,
					-- layer=2 filter=136 channel=122
					2, 2, 0, 1, -8, -4, -1, 1, -1,
					-- layer=2 filter=136 channel=123
					-35, 0, 32, -48, -22, 25, 3, -13, -1,
					-- layer=2 filter=136 channel=124
					-69, 11, 23, 33, -33, 49, 33, 40, 66,
					-- layer=2 filter=136 channel=125
					3, -2, 5, 0, 4, 2, -1, 1, -7,
					-- layer=2 filter=136 channel=126
					-27, 30, -35, 22, 4, 9, -1, -13, 64,
					-- layer=2 filter=136 channel=127
					7, -19, -33, 17, -8, 0, 2, 2, -9,
					-- layer=2 filter=137 channel=0
					-5, 24, 1, -6, 0, 16, -5, -2, 22,
					-- layer=2 filter=137 channel=1
					18, -20, -24, -1, -42, -63, 20, 23, -10,
					-- layer=2 filter=137 channel=2
					7, 5, -2, 6, 10, 11, -4, 8, 10,
					-- layer=2 filter=137 channel=3
					-25, -5, 13, -33, 7, -2, -71, -45, -24,
					-- layer=2 filter=137 channel=4
					11, -1, -3, -16, -4, -35, 1, 20, 3,
					-- layer=2 filter=137 channel=5
					4, 12, 20, 6, 16, 10, 7, 3, 32,
					-- layer=2 filter=137 channel=6
					-13, -46, 27, -45, -14, -10, 19, 11, 3,
					-- layer=2 filter=137 channel=7
					-5, 25, 22, 4, -28, -55, -33, -16, -15,
					-- layer=2 filter=137 channel=8
					6, 1, 3, 6, 3, -3, -6, -2, 8,
					-- layer=2 filter=137 channel=9
					41, 4, -15, -32, -22, -15, -67, -82, -31,
					-- layer=2 filter=137 channel=10
					-20, -4, -5, 2, 8, 3, -38, -17, 8,
					-- layer=2 filter=137 channel=11
					15, 29, 14, 23, 25, 27, -7, 27, 25,
					-- layer=2 filter=137 channel=12
					26, 19, 25, 8, -16, -45, 29, -33, -30,
					-- layer=2 filter=137 channel=13
					-8, 0, -8, 7, -8, -5, 2, -5, -5,
					-- layer=2 filter=137 channel=14
					33, 20, 17, 8, 0, -32, 31, 10, -20,
					-- layer=2 filter=137 channel=15
					-22, 35, -18, 15, -27, -9, 41, 37, -34,
					-- layer=2 filter=137 channel=16
					-24, 17, 3, 14, 24, 27, -23, 8, 39,
					-- layer=2 filter=137 channel=17
					6, -2, -8, 2, -8, 8, -6, 7, 4,
					-- layer=2 filter=137 channel=18
					19, -3, 16, 18, 25, -8, 38, 56, -17,
					-- layer=2 filter=137 channel=19
					-8, -34, -23, -4, -18, -52, 5, -10, -42,
					-- layer=2 filter=137 channel=20
					2, 5, 0, 6, -11, -3, -10, -8, 9,
					-- layer=2 filter=137 channel=21
					18, 17, 23, -5, 8, 15, 8, 0, 4,
					-- layer=2 filter=137 channel=22
					3, -4, 2, 8, -8, 1, 0, 10, 7,
					-- layer=2 filter=137 channel=23
					-23, 0, 29, -7, -18, -7, -31, -8, 30,
					-- layer=2 filter=137 channel=24
					-9, 19, 0, -10, 24, 43, -46, -27, -27,
					-- layer=2 filter=137 channel=25
					9, 32, 24, 7, 44, 27, -44, -19, 4,
					-- layer=2 filter=137 channel=26
					-8, 0, 0, -4, 2, -5, 0, 5, 8,
					-- layer=2 filter=137 channel=27
					8, -20, 3, -8, -20, 3, -35, -7, 13,
					-- layer=2 filter=137 channel=28
					-16, 10, 33, 15, -33, -34, 28, -17, -1,
					-- layer=2 filter=137 channel=29
					-7, -2, -7, -2, -2, 9, 3, -3, -1,
					-- layer=2 filter=137 channel=30
					4, 18, -24, 7, 5, -36, -13, -29, -15,
					-- layer=2 filter=137 channel=31
					-49, -56, -54, -28, 22, -29, 10, -39, -30,
					-- layer=2 filter=137 channel=32
					-5, -9, -1, 7, 9, -9, 1, -5, -8,
					-- layer=2 filter=137 channel=33
					-12, 23, 21, -33, -73, -12, -3, -1, -52,
					-- layer=2 filter=137 channel=34
					-5, -23, -3, 55, 17, 0, 28, 33, 17,
					-- layer=2 filter=137 channel=35
					-38, 36, 19, 56, -21, -6, 5, -11, 11,
					-- layer=2 filter=137 channel=36
					11, 9, 14, 1, -9, 13, -6, -14, -3,
					-- layer=2 filter=137 channel=37
					-3, 4, 29, 13, 6, 29, -3, 11, 23,
					-- layer=2 filter=137 channel=38
					-10, -44, -38, -3, -25, -42, 7, -22, -27,
					-- layer=2 filter=137 channel=39
					-28, 16, 0, -18, -16, -4, -22, 6, 80,
					-- layer=2 filter=137 channel=40
					7, -5, -3, -7, -13, -50, -8, 9, -4,
					-- layer=2 filter=137 channel=41
					6, -7, 2, 10, 12, -1, -7, -1, -7,
					-- layer=2 filter=137 channel=42
					-22, 40, -4, -19, -43, -21, -25, -41, 1,
					-- layer=2 filter=137 channel=43
					-10, 0, -4, -9, -37, -7, -57, -5, 25,
					-- layer=2 filter=137 channel=44
					-10, -5, 6, 6, -6, -9, 6, 4, 10,
					-- layer=2 filter=137 channel=45
					-36, -69, -13, -56, -52, -43, -47, -95, -73,
					-- layer=2 filter=137 channel=46
					3, -8, -37, -1, -28, -27, -6, 17, 21,
					-- layer=2 filter=137 channel=47
					29, 19, -5, -9, -13, -25, -25, 0, 6,
					-- layer=2 filter=137 channel=48
					3, 5, -12, -9, -2, 8, 6, 1, -6,
					-- layer=2 filter=137 channel=49
					34, 4, 15, 39, 30, -28, 18, 20, 26,
					-- layer=2 filter=137 channel=50
					-8, -20, -2, 22, 6, 4, 28, -6, 12,
					-- layer=2 filter=137 channel=51
					0, 21, 19, 20, 23, 6, -10, 23, 26,
					-- layer=2 filter=137 channel=52
					-20, 29, -2, 12, -20, 45, 3, 37, 13,
					-- layer=2 filter=137 channel=53
					-38, -51, 25, -36, -5, -51, 10, -61, -54,
					-- layer=2 filter=137 channel=54
					15, 16, 33, 31, 14, -31, 30, 37, 11,
					-- layer=2 filter=137 channel=55
					1, 7, 4, -5, -1, 0, -1, 6, -1,
					-- layer=2 filter=137 channel=56
					2, 6, 32, -9, 3, 6, 0, 26, 10,
					-- layer=2 filter=137 channel=57
					8, -6, -8, 9, -3, 5, -8, 2, -7,
					-- layer=2 filter=137 channel=58
					-7, 28, 3, 36, -10, -10, 43, -16, -43,
					-- layer=2 filter=137 channel=59
					11, -17, 5, -17, -54, -8, 26, 26, -63,
					-- layer=2 filter=137 channel=60
					-2, -27, -3, 36, 15, -29, 28, -16, -26,
					-- layer=2 filter=137 channel=61
					24, 5, 32, 7, 26, -3, -1, 41, -34,
					-- layer=2 filter=137 channel=62
					19, -36, 8, 38, 12, 34, 20, 28, 20,
					-- layer=2 filter=137 channel=63
					8, 8, -3, 5, -28, 40, 7, -5, 50,
					-- layer=2 filter=137 channel=64
					-23, -38, -2, -8, -19, 9, -12, -13, -8,
					-- layer=2 filter=137 channel=65
					10, -8, 50, 21, 3, 10, 6, 20, -14,
					-- layer=2 filter=137 channel=66
					32, 17, 9, 24, 7, -9, 0, 26, 18,
					-- layer=2 filter=137 channel=67
					41, -41, -7, -47, -68, -34, -23, -22, -33,
					-- layer=2 filter=137 channel=68
					-7, 1, 0, -8, 4, 0, 3, 10, -1,
					-- layer=2 filter=137 channel=69
					-28, -17, 14, -31, -6, 28, -33, -13, 12,
					-- layer=2 filter=137 channel=70
					-2, 22, 20, 23, 12, -10, 32, -2, 17,
					-- layer=2 filter=137 channel=71
					-4, -17, 5, 0, -36, 28, -15, -34, 7,
					-- layer=2 filter=137 channel=72
					34, 24, 28, 11, -20, -6, 27, 30, -44,
					-- layer=2 filter=137 channel=73
					-34, -63, -19, 42, 41, -22, 36, -30, -37,
					-- layer=2 filter=137 channel=74
					-11, 15, -17, 23, -60, 11, 29, -6, -14,
					-- layer=2 filter=137 channel=75
					-60, -27, -4, -22, -31, -10, -19, 1, 29,
					-- layer=2 filter=137 channel=76
					-6, -65, -12, -7, 17, -2, 40, 5, -5,
					-- layer=2 filter=137 channel=77
					4, 0, 4, 8, -8, -9, 4, 7, 7,
					-- layer=2 filter=137 channel=78
					0, 21, 29, 3, 16, 41, -5, 13, 17,
					-- layer=2 filter=137 channel=79
					-5, 3, 6, -7, -3, 0, 9, 1, -6,
					-- layer=2 filter=137 channel=80
					-23, -30, -50, 2, 19, 16, -45, 16, 35,
					-- layer=2 filter=137 channel=81
					-4, 2, 3, 0, -7, -3, 4, 1, 2,
					-- layer=2 filter=137 channel=82
					0, -3, -1, -6, -4, -6, 6, -5, -3,
					-- layer=2 filter=137 channel=83
					-37, 16, 58, -4, 24, 19, -15, -9, 11,
					-- layer=2 filter=137 channel=84
					-8, -4, -1, -10, 8, 5, 6, 3, -1,
					-- layer=2 filter=137 channel=85
					9, 6, 12, 6, 1, 4, -10, -1, -2,
					-- layer=2 filter=137 channel=86
					5, -16, 1, 10, -1, 7, -4, -19, 7,
					-- layer=2 filter=137 channel=87
					26, 6, 16, -23, -22, -11, 39, 25, -10,
					-- layer=2 filter=137 channel=88
					17, -18, 0, -1, -17, -14, -2, -26, -31,
					-- layer=2 filter=137 channel=89
					7, 2, 29, 1, -5, -46, 32, 3, -37,
					-- layer=2 filter=137 channel=90
					10, -3, 2, -6, -5, -5, 2, -10, -1,
					-- layer=2 filter=137 channel=91
					10, 5, -4, -25, -74, -76, 4, -95, -43,
					-- layer=2 filter=137 channel=92
					29, 0, 0, -5, -44, -32, 10, 2, -8,
					-- layer=2 filter=137 channel=93
					18, 0, 15, -5, 0, 9, -23, -62, -25,
					-- layer=2 filter=137 channel=94
					-25, 0, 20, -73, -15, -11, 3, 21, -2,
					-- layer=2 filter=137 channel=95
					-2, -6, -10, -7, -14, -7, -3, -13, 5,
					-- layer=2 filter=137 channel=96
					0, -15, -5, -48, 8, 11, 17, 6, -24,
					-- layer=2 filter=137 channel=97
					-18, -31, -32, -9, 47, 3, -51, -18, 7,
					-- layer=2 filter=137 channel=98
					17, 28, 6, 17, -3, -3, 26, 13, 34,
					-- layer=2 filter=137 channel=99
					-52, -9, -7, -18, 37, 21, -18, 14, 13,
					-- layer=2 filter=137 channel=100
					-44, 0, 4, 15, -19, 22, -35, -20, 9,
					-- layer=2 filter=137 channel=101
					-19, 9, 12, 18, -14, 7, -13, -40, 15,
					-- layer=2 filter=137 channel=102
					3, -1, -11, -9, 25, -30, 11, 8, -1,
					-- layer=2 filter=137 channel=103
					-2, -27, -15, -18, 58, 11, 26, 59, 67,
					-- layer=2 filter=137 channel=104
					30, -12, 14, 0, -6, -30, 20, 30, 12,
					-- layer=2 filter=137 channel=105
					0, -7, 43, -32, 45, -48, -36, -16, -12,
					-- layer=2 filter=137 channel=106
					-2, 4, -1, -6, 14, -18, 2, -40, -22,
					-- layer=2 filter=137 channel=107
					-48, -25, -17, -11, -23, 7, -56, 50, -1,
					-- layer=2 filter=137 channel=108
					-9, -31, -14, -26, -5, -29, -19, -24, -26,
					-- layer=2 filter=137 channel=109
					-5, 7, -8, -11, 2, 14, 2, -13, 10,
					-- layer=2 filter=137 channel=110
					15, -7, 22, -14, -33, -32, -29, -40, -52,
					-- layer=2 filter=137 channel=111
					6, -8, 1, -1, 9, 10, 2, 7, 2,
					-- layer=2 filter=137 channel=112
					-6, 11, -13, -18, 22, -3, -47, -32, -19,
					-- layer=2 filter=137 channel=113
					5, 33, 3, 15, 12, 16, 27, -7, 8,
					-- layer=2 filter=137 channel=114
					-16, 6, 4, -12, 0, -6, -6, 4, -1,
					-- layer=2 filter=137 channel=115
					-1, 3, -10, 11, 2, -5, 3, 6, 1,
					-- layer=2 filter=137 channel=116
					-4, -19, 21, -44, -32, -18, 29, 16, -12,
					-- layer=2 filter=137 channel=117
					-12, 16, -7, -19, -16, -47, -13, 1, -70,
					-- layer=2 filter=137 channel=118
					-13, -31, 15, 16, 1, 22, -32, 10, 19,
					-- layer=2 filter=137 channel=119
					-3, 31, -28, -6, 28, -17, -7, 18, 1,
					-- layer=2 filter=137 channel=120
					2, 8, -2, 9, 2, 9, -7, 5, 4,
					-- layer=2 filter=137 channel=121
					6, -7, 1, 11, -6, 9, 5, 9, -6,
					-- layer=2 filter=137 channel=122
					-8, 8, 3, 0, -5, -7, 3, 3, -7,
					-- layer=2 filter=137 channel=123
					-3, 26, 12, -14, -34, -25, 15, -10, -17,
					-- layer=2 filter=137 channel=124
					2, 37, -10, 20, -7, -57, 33, -10, -32,
					-- layer=2 filter=137 channel=125
					13, 5, -6, 11, -8, 7, 5, 10, -4,
					-- layer=2 filter=137 channel=126
					-23, -33, -19, 12, 8, -27, 7, 14, -31,
					-- layer=2 filter=137 channel=127
					-44, -4, 16, -25, 13, 4, 8, 24, -8,
					-- layer=2 filter=138 channel=0
					-10, -13, -10, -19, -16, -13, 0, -16, -6,
					-- layer=2 filter=138 channel=1
					-5, 4, -7, 0, -13, -21, 1, 15, 3,
					-- layer=2 filter=138 channel=2
					-5, -7, -2, 10, 2, 0, 10, -3, -7,
					-- layer=2 filter=138 channel=3
					-3, -10, -10, -2, 2, 1, 0, 2, -3,
					-- layer=2 filter=138 channel=4
					-1, -3, -4, 5, -7, -16, 0, -9, -17,
					-- layer=2 filter=138 channel=5
					-10, -6, -10, -10, -9, -4, -1, -16, -2,
					-- layer=2 filter=138 channel=6
					0, -1, -3, -6, -11, -16, 4, -5, -7,
					-- layer=2 filter=138 channel=7
					-4, -5, 2, -9, -6, -4, -14, -16, 2,
					-- layer=2 filter=138 channel=8
					-7, -1, -6, -2, -4, 0, 0, -6, -9,
					-- layer=2 filter=138 channel=9
					0, 3, 1, -4, -13, -6, -10, -6, 0,
					-- layer=2 filter=138 channel=10
					-14, -9, -10, -12, -11, -1, -3, -9, -8,
					-- layer=2 filter=138 channel=11
					-2, -15, -2, -7, -13, 3, -3, -5, 3,
					-- layer=2 filter=138 channel=12
					-8, 4, -3, 4, -6, 3, 9, 3, -5,
					-- layer=2 filter=138 channel=13
					6, 8, 7, 4, 4, 2, 6, -5, 8,
					-- layer=2 filter=138 channel=14
					-7, 1, -2, -12, -13, -5, -4, 3, -14,
					-- layer=2 filter=138 channel=15
					4, -8, -1, -5, 6, 9, -10, -7, 0,
					-- layer=2 filter=138 channel=16
					-4, -11, -12, -12, -6, -7, 3, -3, 2,
					-- layer=2 filter=138 channel=17
					1, 0, -7, 3, 6, -6, 2, -7, -6,
					-- layer=2 filter=138 channel=18
					5, 8, 14, 0, -8, 1, 0, -23, -19,
					-- layer=2 filter=138 channel=19
					-5, -1, -13, -4, -17, -18, -12, 0, -13,
					-- layer=2 filter=138 channel=20
					8, 0, 10, 0, -2, -5, -1, 0, -9,
					-- layer=2 filter=138 channel=21
					7, -1, 7, 0, -1, -2, -8, -4, -4,
					-- layer=2 filter=138 channel=22
					8, -2, 7, 5, 9, 7, -1, -2, -9,
					-- layer=2 filter=138 channel=23
					-4, 10, 0, -26, 1, -22, -18, 0, -7,
					-- layer=2 filter=138 channel=24
					-6, -10, -7, -3, 3, 5, 4, -5, 0,
					-- layer=2 filter=138 channel=25
					1, 2, -3, 1, -14, 0, -3, 11, -8,
					-- layer=2 filter=138 channel=26
					10, 4, 6, -3, 4, -10, -1, -8, -9,
					-- layer=2 filter=138 channel=27
					-10, -21, -9, -1, -3, -14, -1, -7, -15,
					-- layer=2 filter=138 channel=28
					-14, -4, -10, 9, 6, -11, -8, -1, 8,
					-- layer=2 filter=138 channel=29
					-7, -2, -11, 0, 1, -6, 0, -10, -8,
					-- layer=2 filter=138 channel=30
					-9, 0, 3, 0, 3, -2, -9, -7, -9,
					-- layer=2 filter=138 channel=31
					16, -4, 8, -11, 2, 5, 5, -5, 8,
					-- layer=2 filter=138 channel=32
					-7, -2, 0, 7, 0, -5, -9, 3, -4,
					-- layer=2 filter=138 channel=33
					-16, -1, 8, -28, 3, 1, -14, 16, -10,
					-- layer=2 filter=138 channel=34
					-5, -14, -5, -6, -2, -2, -10, -4, -1,
					-- layer=2 filter=138 channel=35
					1, -15, -18, 7, -7, 1, -4, -5, 1,
					-- layer=2 filter=138 channel=36
					-11, -11, 9, -7, 0, -1, -2, -6, -11,
					-- layer=2 filter=138 channel=37
					-18, -12, -14, -7, 1, -13, -5, -17, -14,
					-- layer=2 filter=138 channel=38
					-10, -1, -12, 0, -7, -13, -10, -19, -7,
					-- layer=2 filter=138 channel=39
					-7, -2, 2, -8, -11, -5, 0, 4, 2,
					-- layer=2 filter=138 channel=40
					10, -14, -10, -3, 6, 5, -4, 0, 3,
					-- layer=2 filter=138 channel=41
					0, 5, -7, 7, -9, 9, 3, -1, -3,
					-- layer=2 filter=138 channel=42
					0, -5, -9, 4, -7, -6, 1, -2, -9,
					-- layer=2 filter=138 channel=43
					5, 0, -17, -5, -15, -4, -17, 1, 11,
					-- layer=2 filter=138 channel=44
					0, -8, -4, -8, -10, 0, 4, 8, 2,
					-- layer=2 filter=138 channel=45
					2, 2, -11, -18, -2, -1, -14, -15, -13,
					-- layer=2 filter=138 channel=46
					7, -14, -10, -1, -11, 1, -14, -9, -8,
					-- layer=2 filter=138 channel=47
					-11, -6, 6, -15, -1, -13, -4, -9, -10,
					-- layer=2 filter=138 channel=48
					-2, 7, -8, 4, 3, 3, -1, 6, -3,
					-- layer=2 filter=138 channel=49
					7, 7, 1, -2, -21, -3, -10, -10, -4,
					-- layer=2 filter=138 channel=50
					-4, 4, -3, 5, 3, 11, -10, -4, -7,
					-- layer=2 filter=138 channel=51
					2, -8, -1, 0, -3, -8, -16, 2, 1,
					-- layer=2 filter=138 channel=52
					-2, -11, 0, -7, -12, -11, -1, -1, -16,
					-- layer=2 filter=138 channel=53
					13, -15, -19, -3, 2, -5, -4, 0, -17,
					-- layer=2 filter=138 channel=54
					-12, -7, -14, -1, -21, -10, -1, -8, -4,
					-- layer=2 filter=138 channel=55
					9, -6, -5, -6, -10, 3, 3, 5, -7,
					-- layer=2 filter=138 channel=56
					-15, -16, -12, -7, -11, -15, 0, -14, 1,
					-- layer=2 filter=138 channel=57
					-3, 6, 4, -2, -6, 2, -4, 0, 4,
					-- layer=2 filter=138 channel=58
					-9, -5, 7, -6, -11, -14, 10, -5, -1,
					-- layer=2 filter=138 channel=59
					-6, -19, -20, -8, -17, -17, 9, 10, -2,
					-- layer=2 filter=138 channel=60
					-10, -16, -4, -6, -2, -22, -7, -12, 4,
					-- layer=2 filter=138 channel=61
					-23, -11, -6, -6, -2, -1, -8, -6, -14,
					-- layer=2 filter=138 channel=62
					18, -14, -3, 6, 0, -6, -14, -19, -18,
					-- layer=2 filter=138 channel=63
					-10, -2, 0, -9, -3, -3, -17, 0, -10,
					-- layer=2 filter=138 channel=64
					2, 6, -12, -2, -10, -11, -10, 3, -16,
					-- layer=2 filter=138 channel=65
					-9, -5, -9, -7, -3, 0, -13, 0, 1,
					-- layer=2 filter=138 channel=66
					2, 0, -1, 10, 4, -5, 2, 2, 8,
					-- layer=2 filter=138 channel=67
					-9, -14, 0, -13, 5, -10, -10, -18, -4,
					-- layer=2 filter=138 channel=68
					2, -11, -6, -9, -2, 6, 0, 3, -4,
					-- layer=2 filter=138 channel=69
					6, 9, -5, 7, -1, -7, 13, -2, -8,
					-- layer=2 filter=138 channel=70
					-7, -21, -5, -24, -7, -14, -26, -24, -2,
					-- layer=2 filter=138 channel=71
					-5, -13, 13, 2, -10, 3, 0, 1, 9,
					-- layer=2 filter=138 channel=72
					-15, -24, 4, -4, 1, -7, -7, -5, 11,
					-- layer=2 filter=138 channel=73
					10, -14, -14, -1, -5, -14, 0, -4, -12,
					-- layer=2 filter=138 channel=74
					-12, -9, -4, -11, -4, 5, -17, 0, -3,
					-- layer=2 filter=138 channel=75
					3, 0, 1, -2, -5, -12, 6, 8, 2,
					-- layer=2 filter=138 channel=76
					-13, -8, -7, 16, -24, -18, 0, 3, 4,
					-- layer=2 filter=138 channel=77
					-6, 11, 4, 2, -8, -9, -2, -1, -8,
					-- layer=2 filter=138 channel=78
					-14, -9, -12, -16, -6, -2, -13, 1, -18,
					-- layer=2 filter=138 channel=79
					5, -9, 7, -2, 2, 4, -4, 0, -3,
					-- layer=2 filter=138 channel=80
					2, -10, -3, -6, -3, 1, -8, -13, -3,
					-- layer=2 filter=138 channel=81
					5, -6, -11, -9, 8, -3, -2, -5, 2,
					-- layer=2 filter=138 channel=82
					-4, 2, -5, -6, -10, -10, 5, -10, -2,
					-- layer=2 filter=138 channel=83
					-12, -3, 1, -5, -1, 2, -22, -3, -14,
					-- layer=2 filter=138 channel=84
					4, 8, 0, 5, -7, -4, 2, -4, 0,
					-- layer=2 filter=138 channel=85
					0, -2, -10, 5, -9, 7, -2, -9, -10,
					-- layer=2 filter=138 channel=86
					9, -2, -10, 0, 4, 1, -8, -2, -7,
					-- layer=2 filter=138 channel=87
					-5, -6, 3, -10, -18, -3, -18, -7, -11,
					-- layer=2 filter=138 channel=88
					1, -10, -1, -1, -6, -11, -13, 3, 4,
					-- layer=2 filter=138 channel=89
					-3, -13, -12, -18, -20, -7, 7, 11, -2,
					-- layer=2 filter=138 channel=90
					4, -8, 5, -6, 0, -8, -10, 8, 6,
					-- layer=2 filter=138 channel=91
					-11, -14, -5, 1, 0, -2, 5, 3, -6,
					-- layer=2 filter=138 channel=92
					-15, 4, -10, 8, 0, -2, 10, 0, 0,
					-- layer=2 filter=138 channel=93
					11, 6, -10, 1, -3, -2, 3, -2, -18,
					-- layer=2 filter=138 channel=94
					-27, -4, -12, -16, -1, -11, 1, -14, -7,
					-- layer=2 filter=138 channel=95
					4, -5, -1, -6, -2, 7, -3, -7, 2,
					-- layer=2 filter=138 channel=96
					-11, -8, -7, -9, -17, -2, -21, -8, -9,
					-- layer=2 filter=138 channel=97
					-4, 2, -15, -9, -9, -13, -4, -11, 6,
					-- layer=2 filter=138 channel=98
					3, -2, -14, -8, -4, -9, 0, 0, 1,
					-- layer=2 filter=138 channel=99
					-3, -18, -18, 2, -4, -19, -9, -10, -13,
					-- layer=2 filter=138 channel=100
					0, -4, -5, -7, -19, -9, -6, -10, -22,
					-- layer=2 filter=138 channel=101
					-6, -9, -3, -11, 5, -9, -6, 2, 9,
					-- layer=2 filter=138 channel=102
					3, 4, -2, -8, -2, 0, -3, -23, -9,
					-- layer=2 filter=138 channel=103
					3, -4, -8, 1, 1, -1, 0, 4, -5,
					-- layer=2 filter=138 channel=104
					13, -2, -2, -13, -16, -1, -14, 7, -8,
					-- layer=2 filter=138 channel=105
					-5, 6, -19, 6, -8, -17, 0, 10, -5,
					-- layer=2 filter=138 channel=106
					-10, -3, -6, -6, -11, 2, -14, 5, -8,
					-- layer=2 filter=138 channel=107
					4, 0, -2, 9, 2, 7, 9, 3, 6,
					-- layer=2 filter=138 channel=108
					-6, -8, -9, -13, -10, -9, -1, -17, -6,
					-- layer=2 filter=138 channel=109
					-4, -1, 3, 5, 10, -4, 2, 3, 8,
					-- layer=2 filter=138 channel=110
					-2, -13, 5, 4, 6, 7, -6, -4, -5,
					-- layer=2 filter=138 channel=111
					-7, 1, 8, 1, 5, -6, -3, 7, 11,
					-- layer=2 filter=138 channel=112
					-15, -8, -3, -11, -3, -7, -2, -10, -3,
					-- layer=2 filter=138 channel=113
					-6, 0, -4, -10, -12, -18, -20, -8, -23,
					-- layer=2 filter=138 channel=114
					-4, -1, 7, -9, 4, -1, 5, -5, -1,
					-- layer=2 filter=138 channel=115
					2, -8, 1, -3, 6, 9, -7, 8, -10,
					-- layer=2 filter=138 channel=116
					-7, -11, 8, -10, 15, -17, 0, 0, -15,
					-- layer=2 filter=138 channel=117
					-1, -6, 0, -5, -1, -12, -10, -3, 5,
					-- layer=2 filter=138 channel=118
					0, -6, -8, -14, -19, -4, -13, -12, -16,
					-- layer=2 filter=138 channel=119
					5, -17, 2, 11, -1, -13, 9, -12, -13,
					-- layer=2 filter=138 channel=120
					8, 0, -6, 6, 2, 7, -3, -5, 0,
					-- layer=2 filter=138 channel=121
					-10, -4, -5, -3, 0, -2, 2, -10, 10,
					-- layer=2 filter=138 channel=122
					0, -4, -3, 6, 5, -1, -4, 4, 7,
					-- layer=2 filter=138 channel=123
					-5, -19, -9, -2, -2, -2, -8, -11, 7,
					-- layer=2 filter=138 channel=124
					5, 5, -1, 8, -5, 12, 12, -6, 0,
					-- layer=2 filter=138 channel=125
					-3, -7, 4, 9, 6, 2, 4, 6, 9,
					-- layer=2 filter=138 channel=126
					-15, -10, 2, -11, 0, -9, -15, -10, 0,
					-- layer=2 filter=138 channel=127
					-18, 2, 1, -10, 0, -9, -5, 0, 0,
					-- layer=2 filter=139 channel=0
					6, -8, -6, -2, -9, -5, -2, 0, -7,
					-- layer=2 filter=139 channel=1
					7, -9, 1, -11, -5, -12, -6, -12, -8,
					-- layer=2 filter=139 channel=2
					0, -1, 0, -9, 7, -8, 8, 0, -8,
					-- layer=2 filter=139 channel=3
					8, -3, 3, -12, -12, 8, -9, -1, -7,
					-- layer=2 filter=139 channel=4
					-3, -9, 0, -11, -6, 5, -10, 3, 3,
					-- layer=2 filter=139 channel=5
					4, -6, 8, -9, -5, 7, 3, -4, -11,
					-- layer=2 filter=139 channel=6
					-10, -13, -5, 2, -10, -10, -5, -11, -9,
					-- layer=2 filter=139 channel=7
					0, -7, -6, -5, 8, 5, 4, 10, -12,
					-- layer=2 filter=139 channel=8
					-4, -3, -1, -4, -4, 0, -4, 4, 0,
					-- layer=2 filter=139 channel=9
					-4, -4, 6, 0, -11, 0, 2, 8, -10,
					-- layer=2 filter=139 channel=10
					4, 4, -12, -7, 6, 8, -7, -8, -4,
					-- layer=2 filter=139 channel=11
					-6, -3, 0, 1, -1, -3, 11, -3, -11,
					-- layer=2 filter=139 channel=12
					3, 4, -4, -11, -3, -7, 0, -3, -1,
					-- layer=2 filter=139 channel=13
					3, -8, -8, 0, -2, 7, 5, 1, -6,
					-- layer=2 filter=139 channel=14
					8, -9, -6, 8, -1, -6, -6, -11, -6,
					-- layer=2 filter=139 channel=15
					-8, 2, -5, 0, -6, -1, -2, -9, 4,
					-- layer=2 filter=139 channel=16
					5, -8, -8, 3, 6, 5, -11, -12, 5,
					-- layer=2 filter=139 channel=17
					10, 6, -6, -3, -2, -4, -2, -3, -5,
					-- layer=2 filter=139 channel=18
					-1, -1, 5, -8, -2, -11, -2, 6, -11,
					-- layer=2 filter=139 channel=19
					-7, -2, -6, -13, -11, -1, -15, 0, -1,
					-- layer=2 filter=139 channel=20
					0, -8, -3, -8, -11, -4, 1, 1, -3,
					-- layer=2 filter=139 channel=21
					-11, -5, -2, 2, -5, 6, 3, -5, -7,
					-- layer=2 filter=139 channel=22
					0, 2, 4, 3, 4, 6, 2, -7, 1,
					-- layer=2 filter=139 channel=23
					-5, 3, -4, -3, -10, 4, 0, 5, 6,
					-- layer=2 filter=139 channel=24
					-9, 4, -12, 0, 0, 4, 5, 3, -13,
					-- layer=2 filter=139 channel=25
					0, 4, -16, 1, 8, -3, -1, 0, -4,
					-- layer=2 filter=139 channel=26
					-10, 5, -6, 7, -1, -2, 10, 8, -3,
					-- layer=2 filter=139 channel=27
					-11, -2, 2, 1, 4, 8, -9, -8, 0,
					-- layer=2 filter=139 channel=28
					-14, -4, -7, -2, -8, -10, -7, -1, -1,
					-- layer=2 filter=139 channel=29
					-5, -7, -12, 7, -4, -8, 4, -4, 8,
					-- layer=2 filter=139 channel=30
					-5, -3, -4, 0, 6, 5, 0, -9, 8,
					-- layer=2 filter=139 channel=31
					8, 7, 0, 2, 8, -7, 8, 1, -1,
					-- layer=2 filter=139 channel=32
					1, 7, -4, -2, 5, -9, -2, 2, 5,
					-- layer=2 filter=139 channel=33
					2, 7, 0, -9, -7, 7, -14, 2, 2,
					-- layer=2 filter=139 channel=34
					-1, -2, -3, 5, 1, 0, -2, -6, 3,
					-- layer=2 filter=139 channel=35
					-4, 2, -6, 0, 5, 3, -4, 8, -6,
					-- layer=2 filter=139 channel=36
					-4, -1, 5, -9, 6, -10, 7, -3, -10,
					-- layer=2 filter=139 channel=37
					-6, -6, 2, 7, -10, 0, 5, 0, -11,
					-- layer=2 filter=139 channel=38
					-1, 1, -11, -3, -8, 0, 1, -2, 2,
					-- layer=2 filter=139 channel=39
					-9, 0, 8, -3, -9, -6, -11, -9, -6,
					-- layer=2 filter=139 channel=40
					-6, 6, 6, 2, 8, -4, 2, 4, 6,
					-- layer=2 filter=139 channel=41
					10, -2, 10, -1, 7, -7, 0, 8, 8,
					-- layer=2 filter=139 channel=42
					1, -6, 3, -3, 0, -8, 4, 0, 3,
					-- layer=2 filter=139 channel=43
					-1, -3, 5, 0, 1, 7, 7, -10, -5,
					-- layer=2 filter=139 channel=44
					0, -8, 5, 6, -4, 8, -7, -10, 4,
					-- layer=2 filter=139 channel=45
					8, 0, 0, 1, 2, -1, -12, -12, -3,
					-- layer=2 filter=139 channel=46
					-2, 0, -8, 6, -1, -2, 5, -2, 3,
					-- layer=2 filter=139 channel=47
					-10, 3, -2, 3, -8, -2, -8, 3, 4,
					-- layer=2 filter=139 channel=48
					-2, -4, 5, -7, 10, 1, 4, 4, 2,
					-- layer=2 filter=139 channel=49
					-5, -4, -7, 1, -10, -13, 8, -10, 1,
					-- layer=2 filter=139 channel=50
					-2, 2, 8, -6, 3, -4, -8, 4, 11,
					-- layer=2 filter=139 channel=51
					-11, -14, 1, -6, -11, -13, -5, -2, 2,
					-- layer=2 filter=139 channel=52
					-11, -8, 7, -7, -1, -6, 0, -6, -13,
					-- layer=2 filter=139 channel=53
					-11, 0, 1, -5, -6, 5, -9, 2, -7,
					-- layer=2 filter=139 channel=54
					1, 8, 0, -1, 1, 5, -3, 7, 2,
					-- layer=2 filter=139 channel=55
					7, -3, 7, 1, 6, -10, -2, 0, -2,
					-- layer=2 filter=139 channel=56
					6, -11, -1, -7, -8, 5, -5, -3, -5,
					-- layer=2 filter=139 channel=57
					7, 2, 3, 8, 5, -10, 0, -7, -9,
					-- layer=2 filter=139 channel=58
					7, -5, -11, -13, -1, 7, -2, -4, 7,
					-- layer=2 filter=139 channel=59
					0, -15, -8, 4, 0, 0, -1, 1, 7,
					-- layer=2 filter=139 channel=60
					-1, -3, 0, -5, -2, -9, 0, 2, -5,
					-- layer=2 filter=139 channel=61
					-6, -1, -1, 2, -1, -7, 8, -1, -12,
					-- layer=2 filter=139 channel=62
					-2, -5, -7, 0, -1, 4, -2, -15, 2,
					-- layer=2 filter=139 channel=63
					1, -6, -3, 4, 1, -10, -1, -11, 2,
					-- layer=2 filter=139 channel=64
					8, -5, 0, -5, -6, -9, -6, -1, -2,
					-- layer=2 filter=139 channel=65
					-2, -5, -10, 0, 1, -10, -7, 0, -4,
					-- layer=2 filter=139 channel=66
					-10, 7, -5, -5, -5, 4, -1, 3, -9,
					-- layer=2 filter=139 channel=67
					-1, -1, -7, -9, 3, 3, 6, 8, 7,
					-- layer=2 filter=139 channel=68
					-11, -4, 6, -2, -12, 2, -1, -3, -3,
					-- layer=2 filter=139 channel=69
					9, -7, -5, -1, -9, 8, -11, -9, -9,
					-- layer=2 filter=139 channel=70
					0, 3, -10, -10, -5, -7, 6, 7, -2,
					-- layer=2 filter=139 channel=71
					1, -2, -1, 3, 0, -2, 2, 6, -9,
					-- layer=2 filter=139 channel=72
					-2, 0, 6, -9, -12, -8, -4, -4, -12,
					-- layer=2 filter=139 channel=73
					6, -11, -15, -2, -3, 0, 0, -6, -4,
					-- layer=2 filter=139 channel=74
					7, 1, 7, -11, 1, -3, -10, 8, 5,
					-- layer=2 filter=139 channel=75
					0, -1, -6, -10, 1, -12, -11, -7, -4,
					-- layer=2 filter=139 channel=76
					3, 2, -12, 0, -4, 6, 1, 5, 0,
					-- layer=2 filter=139 channel=77
					-6, -9, 1, 6, 6, 4, -9, 1, -4,
					-- layer=2 filter=139 channel=78
					7, -10, -3, 7, -1, 5, -10, 6, 2,
					-- layer=2 filter=139 channel=79
					4, -3, 2, -11, -6, 0, 8, 8, 7,
					-- layer=2 filter=139 channel=80
					0, -1, 1, -5, -8, -10, 3, -4, -2,
					-- layer=2 filter=139 channel=81
					-11, 0, -7, 0, 1, 0, -4, 7, 0,
					-- layer=2 filter=139 channel=82
					-2, 2, 1, -6, 8, -6, -1, -2, -7,
					-- layer=2 filter=139 channel=83
					-9, 1, 5, 5, 3, 0, 7, -7, -11,
					-- layer=2 filter=139 channel=84
					1, 4, -1, 4, 9, -4, 6, -8, -9,
					-- layer=2 filter=139 channel=85
					2, 8, 0, 9, 0, 4, 6, -4, -6,
					-- layer=2 filter=139 channel=86
					3, 0, -5, -4, -5, 0, -1, 3, -4,
					-- layer=2 filter=139 channel=87
					-2, 8, 0, 0, -3, -5, 0, 2, 4,
					-- layer=2 filter=139 channel=88
					-5, 1, -6, 4, 4, -10, -12, 2, 3,
					-- layer=2 filter=139 channel=89
					0, -5, 7, -6, -15, -13, -10, -14, 6,
					-- layer=2 filter=139 channel=90
					-7, 2, -4, -6, -5, -7, 0, 10, 8,
					-- layer=2 filter=139 channel=91
					10, -9, -7, 4, -7, -5, 2, -15, -2,
					-- layer=2 filter=139 channel=92
					4, -13, 2, -4, -4, -4, -6, 0, -9,
					-- layer=2 filter=139 channel=93
					-1, -3, 0, 0, -5, 2, 0, 1, 1,
					-- layer=2 filter=139 channel=94
					-6, -5, -8, 0, -1, -3, -3, 1, 4,
					-- layer=2 filter=139 channel=95
					-8, -1, 6, -1, 5, -7, 8, -7, -5,
					-- layer=2 filter=139 channel=96
					-1, 5, -2, 0, 4, -11, 2, 1, 7,
					-- layer=2 filter=139 channel=97
					6, 6, -1, 0, -1, -3, 5, -8, -7,
					-- layer=2 filter=139 channel=98
					-11, -9, -2, -15, -6, 2, 0, -7, -13,
					-- layer=2 filter=139 channel=99
					-5, 3, 4, -6, 0, -6, 1, -12, -9,
					-- layer=2 filter=139 channel=100
					0, -6, -4, -6, 5, -5, -7, -3, -2,
					-- layer=2 filter=139 channel=101
					4, -5, -12, 2, 3, 3, -4, 0, -12,
					-- layer=2 filter=139 channel=102
					3, -2, -5, -4, -8, -7, 6, -1, 5,
					-- layer=2 filter=139 channel=103
					-3, 7, 7, 2, -3, -10, -2, 7, 2,
					-- layer=2 filter=139 channel=104
					0, -11, -9, -10, 6, 8, -2, -2, 2,
					-- layer=2 filter=139 channel=105
					2, -1, 9, -9, -4, 8, 0, 0, -5,
					-- layer=2 filter=139 channel=106
					4, 3, 7, -3, -9, -12, 4, -9, 1,
					-- layer=2 filter=139 channel=107
					-5, -7, 6, 0, 0, -6, 6, -7, -11,
					-- layer=2 filter=139 channel=108
					3, 4, -10, -3, 0, 2, -10, -2, -10,
					-- layer=2 filter=139 channel=109
					8, -1, 0, 0, -4, 7, -5, -9, 8,
					-- layer=2 filter=139 channel=110
					-6, -3, -10, -5, 6, 4, 2, 5, -11,
					-- layer=2 filter=139 channel=111
					-3, 4, 5, -4, 8, -3, -3, -4, -8,
					-- layer=2 filter=139 channel=112
					-11, -12, -10, 6, 7, -1, 0, 1, -1,
					-- layer=2 filter=139 channel=113
					-5, 0, 7, -4, -2, 0, 2, 4, -8,
					-- layer=2 filter=139 channel=114
					5, 5, -9, 5, -4, -1, 9, 0, 4,
					-- layer=2 filter=139 channel=115
					-4, -4, -10, 0, -1, -6, 10, -4, 0,
					-- layer=2 filter=139 channel=116
					4, -9, 4, 2, -10, 5, 5, 5, -6,
					-- layer=2 filter=139 channel=117
					-1, 5, -6, -9, 8, 2, -14, -5, 5,
					-- layer=2 filter=139 channel=118
					-6, -2, -4, -10, -3, 0, -8, -4, 6,
					-- layer=2 filter=139 channel=119
					-1, -11, 6, -5, -9, -1, -2, -5, -3,
					-- layer=2 filter=139 channel=120
					7, -4, 9, 1, 5, 8, 2, 0, 7,
					-- layer=2 filter=139 channel=121
					-9, -4, 5, -10, -4, 0, 5, 1, -11,
					-- layer=2 filter=139 channel=122
					-6, -11, -8, 3, 6, -6, 0, -5, 3,
					-- layer=2 filter=139 channel=123
					-1, 0, 8, 4, -5, -11, -6, -12, 0,
					-- layer=2 filter=139 channel=124
					-3, 6, 3, -4, -6, -12, -9, -1, 3,
					-- layer=2 filter=139 channel=125
					-2, -10, 5, 12, -4, -1, 8, 5, -4,
					-- layer=2 filter=139 channel=126
					-2, 1, 0, -2, -3, 5, 0, 7, 7,
					-- layer=2 filter=139 channel=127
					-10, -11, 6, 3, 7, 0, 6, -4, 4,
					-- layer=2 filter=140 channel=0
					-6, -8, 6, -7, -3, 2, -3, -8, 0,
					-- layer=2 filter=140 channel=1
					4, -5, -3, 4, -8, -11, -4, -9, -9,
					-- layer=2 filter=140 channel=2
					-10, -6, 9, -9, -1, 0, 0, -5, -11,
					-- layer=2 filter=140 channel=3
					4, 0, 0, 1, 0, 7, 5, 0, 10,
					-- layer=2 filter=140 channel=4
					-7, -10, 0, -6, 3, -9, -2, 6, -10,
					-- layer=2 filter=140 channel=5
					-6, -6, -1, 3, -3, -10, -10, 7, 4,
					-- layer=2 filter=140 channel=6
					3, -8, 0, 0, 1, -3, -8, 2, -5,
					-- layer=2 filter=140 channel=7
					0, 0, 7, 6, 11, 8, 0, -2, 3,
					-- layer=2 filter=140 channel=8
					3, 1, -8, 8, -2, 8, -2, -5, 0,
					-- layer=2 filter=140 channel=9
					-11, 5, 7, -6, 5, 3, 7, -6, 4,
					-- layer=2 filter=140 channel=10
					1, 0, -5, -5, 10, -2, 1, -3, -1,
					-- layer=2 filter=140 channel=11
					0, 9, 2, -9, -1, 0, -10, -2, 1,
					-- layer=2 filter=140 channel=12
					-12, 0, -9, -11, -3, -8, 2, -8, 0,
					-- layer=2 filter=140 channel=13
					-7, 9, 8, 1, 7, 1, -6, 7, 5,
					-- layer=2 filter=140 channel=14
					-8, 4, -3, -2, 9, 4, 1, -10, -11,
					-- layer=2 filter=140 channel=15
					-12, -8, 0, -7, -3, -9, 3, -2, 4,
					-- layer=2 filter=140 channel=16
					-8, 2, -15, 2, -5, -9, -2, -1, 8,
					-- layer=2 filter=140 channel=17
					6, 3, 9, 6, 0, 8, -6, -1, 3,
					-- layer=2 filter=140 channel=18
					1, -11, 4, 2, 3, 4, 12, -8, -2,
					-- layer=2 filter=140 channel=19
					0, -6, 4, -2, 0, 0, -1, 2, 9,
					-- layer=2 filter=140 channel=20
					8, 8, -8, 0, -6, 2, -9, -6, -11,
					-- layer=2 filter=140 channel=21
					-3, 7, 3, -1, 0, -8, 4, -3, -2,
					-- layer=2 filter=140 channel=22
					6, -1, -10, 10, -1, 10, 1, -5, -8,
					-- layer=2 filter=140 channel=23
					-2, -9, 0, -5, -10, 0, 7, 9, -4,
					-- layer=2 filter=140 channel=24
					2, -7, -4, -9, -3, -5, -2, 2, 1,
					-- layer=2 filter=140 channel=25
					4, -10, -7, 5, 6, -2, -7, 2, -4,
					-- layer=2 filter=140 channel=26
					1, -5, -2, 9, -3, 9, 0, 5, -5,
					-- layer=2 filter=140 channel=27
					-13, -4, -7, -5, 1, -6, -6, 2, 7,
					-- layer=2 filter=140 channel=28
					-3, 7, -5, -8, -2, -2, 5, 10, -10,
					-- layer=2 filter=140 channel=29
					6, -1, 7, 6, 6, -4, -4, -7, -2,
					-- layer=2 filter=140 channel=30
					6, -3, -1, 0, -12, 0, -9, -5, -4,
					-- layer=2 filter=140 channel=31
					2, 6, 7, 4, 4, 5, -4, 8, -4,
					-- layer=2 filter=140 channel=32
					10, -11, -8, 1, -4, -5, 0, -2, -6,
					-- layer=2 filter=140 channel=33
					-8, 8, -8, -3, 10, -9, 1, -2, -12,
					-- layer=2 filter=140 channel=34
					-11, -2, 6, -8, -1, 9, 0, -8, 1,
					-- layer=2 filter=140 channel=35
					-12, -5, 9, -14, -13, -11, -5, 0, -3,
					-- layer=2 filter=140 channel=36
					0, 1, 7, -7, 9, 0, -3, -8, 7,
					-- layer=2 filter=140 channel=37
					-10, 8, 10, -10, -9, 4, 8, -9, -6,
					-- layer=2 filter=140 channel=38
					1, -2, 1, 0, -3, -6, 4, 0, -7,
					-- layer=2 filter=140 channel=39
					2, -1, -8, -7, 0, 0, 7, 5, -11,
					-- layer=2 filter=140 channel=40
					-6, -9, -3, -14, 9, 6, -7, -10, 1,
					-- layer=2 filter=140 channel=41
					-10, -10, 2, -4, -1, -7, -4, 7, -5,
					-- layer=2 filter=140 channel=42
					-3, -7, 0, -4, 6, 10, 6, 5, -4,
					-- layer=2 filter=140 channel=43
					-3, -10, 3, -2, -6, 8, -12, -7, -3,
					-- layer=2 filter=140 channel=44
					0, -6, 1, 2, -6, 0, 0, 0, 5,
					-- layer=2 filter=140 channel=45
					4, 0, -11, -1, -5, -10, 8, -11, -3,
					-- layer=2 filter=140 channel=46
					7, -9, -11, 1, 5, -1, 5, 7, -9,
					-- layer=2 filter=140 channel=47
					1, 2, -16, -8, -9, -3, 5, -2, 9,
					-- layer=2 filter=140 channel=48
					-3, -8, 2, -2, 1, 2, 2, 0, -7,
					-- layer=2 filter=140 channel=49
					-9, 0, 1, -1, 10, -2, 0, -5, -5,
					-- layer=2 filter=140 channel=50
					1, -6, -1, -9, -9, -4, -1, 10, 6,
					-- layer=2 filter=140 channel=51
					-2, -7, 0, 0, 5, 7, 7, 5, -6,
					-- layer=2 filter=140 channel=52
					-3, 11, 4, 3, 1, -1, 10, 9, 4,
					-- layer=2 filter=140 channel=53
					-1, -3, -3, 1, -1, -5, -10, 0, 4,
					-- layer=2 filter=140 channel=54
					0, -1, -15, -11, -12, -9, -9, 0, -5,
					-- layer=2 filter=140 channel=55
					4, 9, -8, 2, 9, -9, -6, 1, 0,
					-- layer=2 filter=140 channel=56
					-9, 0, -6, 0, -11, -10, 0, 2, 6,
					-- layer=2 filter=140 channel=57
					1, -7, 8, -11, -8, -4, -2, -8, 6,
					-- layer=2 filter=140 channel=58
					-7, 1, -2, -4, -9, -10, 0, -5, -11,
					-- layer=2 filter=140 channel=59
					-7, -4, 1, 0, 5, -7, 3, 4, -1,
					-- layer=2 filter=140 channel=60
					-8, 0, 5, -10, -3, 1, -5, 9, -7,
					-- layer=2 filter=140 channel=61
					0, 2, -4, -5, 3, -8, 5, -12, -7,
					-- layer=2 filter=140 channel=62
					-9, -10, -7, -4, -9, 8, 4, -2, 1,
					-- layer=2 filter=140 channel=63
					7, 2, -4, 3, -9, 9, -4, -11, 2,
					-- layer=2 filter=140 channel=64
					-2, -7, 2, 6, 0, 1, 3, -8, 4,
					-- layer=2 filter=140 channel=65
					0, -5, -7, 1, -8, -10, 3, -1, -9,
					-- layer=2 filter=140 channel=66
					7, 0, -6, 9, -4, 5, -1, 2, -9,
					-- layer=2 filter=140 channel=67
					-5, -6, -3, 4, 0, -1, 0, 7, -9,
					-- layer=2 filter=140 channel=68
					-6, -9, 5, -3, 7, 3, 5, 1, 5,
					-- layer=2 filter=140 channel=69
					8, 1, 5, 0, -6, -4, 0, 0, 1,
					-- layer=2 filter=140 channel=70
					6, -7, 9, -3, -2, 2, -11, 2, -5,
					-- layer=2 filter=140 channel=71
					-7, 3, -3, -2, -1, 4, 1, 5, 6,
					-- layer=2 filter=140 channel=72
					3, 0, 0, -14, 6, 1, -9, 1, -7,
					-- layer=2 filter=140 channel=73
					-8, -3, 7, 7, -7, -2, -4, 4, -2,
					-- layer=2 filter=140 channel=74
					-4, -10, -3, -5, 0, 6, -5, -12, -7,
					-- layer=2 filter=140 channel=75
					1, -13, -11, 2, -5, 10, 7, 2, 7,
					-- layer=2 filter=140 channel=76
					-6, 5, 5, -6, 0, 4, -2, -7, 9,
					-- layer=2 filter=140 channel=77
					-10, -5, -3, -9, -4, -9, -6, 6, 0,
					-- layer=2 filter=140 channel=78
					-4, 1, 0, 7, 0, 5, 3, 0, 4,
					-- layer=2 filter=140 channel=79
					-2, -5, -7, -11, 3, -1, 2, 3, 7,
					-- layer=2 filter=140 channel=80
					-12, 2, -13, -4, -6, 5, 1, -1, -10,
					-- layer=2 filter=140 channel=81
					-9, -7, 0, -3, -10, 5, 4, -6, 3,
					-- layer=2 filter=140 channel=82
					-6, 4, 4, -3, -5, 0, -8, -2, 6,
					-- layer=2 filter=140 channel=83
					1, -7, -8, -2, -12, -4, -12, -7, -10,
					-- layer=2 filter=140 channel=84
					-11, -4, 1, -4, 5, 10, 3, 7, -1,
					-- layer=2 filter=140 channel=85
					10, -6, -6, 0, -6, 3, 5, 2, 0,
					-- layer=2 filter=140 channel=86
					1, -2, 6, -4, -1, 4, 5, 6, -3,
					-- layer=2 filter=140 channel=87
					2, 1, -1, -11, 7, -1, -7, 3, -7,
					-- layer=2 filter=140 channel=88
					-7, -5, 2, -11, -9, 1, 0, -12, -6,
					-- layer=2 filter=140 channel=89
					-1, -8, -7, 10, -4, -5, -3, -9, -4,
					-- layer=2 filter=140 channel=90
					3, -1, 10, 2, 4, 4, 0, -1, -1,
					-- layer=2 filter=140 channel=91
					-9, -11, -2, 7, -12, -9, 2, -8, -8,
					-- layer=2 filter=140 channel=92
					7, -6, -7, 2, 8, 0, 1, -5, -9,
					-- layer=2 filter=140 channel=93
					0, -4, -5, -6, -2, 8, -8, 6, 0,
					-- layer=2 filter=140 channel=94
					4, -11, -12, -9, -6, 6, 5, 5, 5,
					-- layer=2 filter=140 channel=95
					-5, -5, 1, 3, -7, 8, -7, -5, 4,
					-- layer=2 filter=140 channel=96
					0, 1, -4, 5, -2, -4, -4, -10, 4,
					-- layer=2 filter=140 channel=97
					4, -8, 2, 6, 2, -9, -7, -7, -3,
					-- layer=2 filter=140 channel=98
					-12, 0, -4, -12, -6, 7, -8, -1, 0,
					-- layer=2 filter=140 channel=99
					6, -9, 12, 8, 0, -4, -2, -2, 0,
					-- layer=2 filter=140 channel=100
					-5, 0, -4, -7, -4, 10, -3, -1, -9,
					-- layer=2 filter=140 channel=101
					9, 1, -8, 3, -9, -10, -10, -8, 3,
					-- layer=2 filter=140 channel=102
					-8, 3, 3, 2, 6, 4, 0, -10, -10,
					-- layer=2 filter=140 channel=103
					-3, -6, -3, -2, 6, 8, -1, 0, 0,
					-- layer=2 filter=140 channel=104
					-2, -9, -10, 2, -4, 6, -9, 2, -2,
					-- layer=2 filter=140 channel=105
					-11, 2, 1, 10, 2, 4, 4, -7, -4,
					-- layer=2 filter=140 channel=106
					-8, -1, 7, -10, -1, 8, 2, -2, 10,
					-- layer=2 filter=140 channel=107
					0, -1, -8, 4, 11, -1, -8, 6, -5,
					-- layer=2 filter=140 channel=108
					4, 4, 6, -2, 1, 5, -12, -9, -6,
					-- layer=2 filter=140 channel=109
					-8, -7, -2, -1, -4, 1, -6, 3, -5,
					-- layer=2 filter=140 channel=110
					-11, 5, -11, 3, -2, -7, -6, 0, 0,
					-- layer=2 filter=140 channel=111
					1, -1, 0, 3, -4, -1, 0, 0, 3,
					-- layer=2 filter=140 channel=112
					-5, 7, -7, 9, -7, 8, -4, 0, 1,
					-- layer=2 filter=140 channel=113
					4, 0, -12, 10, 5, 0, 1, -4, -3,
					-- layer=2 filter=140 channel=114
					-10, 0, 12, -12, -9, 7, 0, -7, 7,
					-- layer=2 filter=140 channel=115
					0, 10, 0, 1, 7, 0, -1, -9, 8,
					-- layer=2 filter=140 channel=116
					-10, -7, -2, 9, -1, 10, -4, 0, -9,
					-- layer=2 filter=140 channel=117
					-9, -3, -3, -18, -6, -12, -5, 2, -3,
					-- layer=2 filter=140 channel=118
					-5, 6, -3, 6, 0, -6, 5, -9, -10,
					-- layer=2 filter=140 channel=119
					-10, -13, -7, 1, -4, -2, -11, -11, -10,
					-- layer=2 filter=140 channel=120
					3, 6, -6, -8, -6, -7, 2, 4, -8,
					-- layer=2 filter=140 channel=121
					-7, -1, -2, -8, -11, -8, -1, 0, 10,
					-- layer=2 filter=140 channel=122
					-7, 8, 3, 3, -3, 1, 2, 6, -9,
					-- layer=2 filter=140 channel=123
					0, 0, 4, -8, -8, -4, -13, 0, -2,
					-- layer=2 filter=140 channel=124
					2, 7, 1, -11, -2, 4, 1, -8, 8,
					-- layer=2 filter=140 channel=125
					-7, 6, 1, -3, 10, 5, 4, -7, 8,
					-- layer=2 filter=140 channel=126
					-9, -6, 0, -3, -8, -11, 7, -1, 8,
					-- layer=2 filter=140 channel=127
					6, 1, -4, 1, -5, -1, 0, -5, -12,
					-- layer=2 filter=141 channel=0
					0, -2, 10, 12, -9, -3, -6, -11, 3,
					-- layer=2 filter=141 channel=1
					-5, 6, 66, 6, -12, 17, -16, 12, -38,
					-- layer=2 filter=141 channel=2
					-5, 3, 3, -2, 10, 0, -8, -8, 7,
					-- layer=2 filter=141 channel=3
					25, -8, -23, -25, 9, -22, -14, -15, 25,
					-- layer=2 filter=141 channel=4
					19, -11, 7, -5, -25, 0, -16, 0, 6,
					-- layer=2 filter=141 channel=5
					-2, 3, -6, 6, -13, 20, 10, 12, 23,
					-- layer=2 filter=141 channel=6
					0, 40, 27, 3, 24, -28, 23, 20, -50,
					-- layer=2 filter=141 channel=7
					7, -18, -15, 37, 72, 35, 19, 10, -19,
					-- layer=2 filter=141 channel=8
					-9, 6, 0, -2, 7, -1, 4, 5, 0,
					-- layer=2 filter=141 channel=9
					0, -33, -17, -7, -63, -8, 1, 16, 34,
					-- layer=2 filter=141 channel=10
					14, -9, -23, 9, -9, -15, 16, -2, 26,
					-- layer=2 filter=141 channel=11
					-3, 6, -14, -1, 4, 12, -13, -19, 14,
					-- layer=2 filter=141 channel=12
					-2, 31, 7, 26, 15, 17, 10, 19, 5,
					-- layer=2 filter=141 channel=13
					2, 6, -6, -1, -6, 4, 6, 5, 6,
					-- layer=2 filter=141 channel=14
					-6, 11, 27, 24, 10, 3, 4, -8, -13,
					-- layer=2 filter=141 channel=15
					0, -7, -11, -4, 14, -20, -20, -28, 9,
					-- layer=2 filter=141 channel=16
					-15, 19, -23, -31, -11, -36, -43, -16, -51,
					-- layer=2 filter=141 channel=17
					5, 3, -3, 0, 8, 9, 5, -5, -4,
					-- layer=2 filter=141 channel=18
					-16, -18, -14, -15, 3, 16, 17, 8, 7,
					-- layer=2 filter=141 channel=19
					-29, 8, 36, -21, 23, 25, 7, 35, -10,
					-- layer=2 filter=141 channel=20
					-5, 9, 5, 0, -7, 0, -7, -3, 4,
					-- layer=2 filter=141 channel=21
					7, -19, 4, -19, -19, -5, -14, 12, -8,
					-- layer=2 filter=141 channel=22
					-3, 2, 4, -1, -1, 3, -4, -4, -7,
					-- layer=2 filter=141 channel=23
					7, 12, 4, -9, -9, -18, -37, -29, -7,
					-- layer=2 filter=141 channel=24
					21, 0, -30, -4, -22, -1, -7, -55, -23,
					-- layer=2 filter=141 channel=25
					11, 7, -23, 6, 9, -13, -32, -70, -28,
					-- layer=2 filter=141 channel=26
					-1, -7, 4, -3, 5, 3, -8, -6, -1,
					-- layer=2 filter=141 channel=27
					-37, -14, 0, -29, 3, -8, 1, -20, -10,
					-- layer=2 filter=141 channel=28
					8, 24, 10, -21, 35, 11, 44, -2, 28,
					-- layer=2 filter=141 channel=29
					-5, 1, 5, 3, -10, 0, -4, 0, 1,
					-- layer=2 filter=141 channel=30
					15, 2, -2, 3, -27, 22, 31, -8, 5,
					-- layer=2 filter=141 channel=31
					36, 62, -67, 23, 7, -90, 61, 22, -38,
					-- layer=2 filter=141 channel=32
					2, -9, -10, -1, 6, -2, -4, -4, -2,
					-- layer=2 filter=141 channel=33
					-11, -5, -1, 9, -9, -12, -23, -35, -20,
					-- layer=2 filter=141 channel=34
					-14, 17, -4, -38, -18, -26, -22, 29, -18,
					-- layer=2 filter=141 channel=35
					1, 18, 26, -3, 17, -2, 4, 7, -4,
					-- layer=2 filter=141 channel=36
					10, 0, 0, 7, 3, -8, 0, 4, -6,
					-- layer=2 filter=141 channel=37
					-7, -10, -12, -11, 16, 24, -4, -11, 7,
					-- layer=2 filter=141 channel=38
					0, -5, -22, 4, -18, 6, 36, 16, -2,
					-- layer=2 filter=141 channel=39
					-1, -7, -21, -13, 9, -16, -56, -4, 18,
					-- layer=2 filter=141 channel=40
					23, -9, -26, -28, -15, -64, -2, 19, -6,
					-- layer=2 filter=141 channel=41
					4, 0, -4, -6, 1, 1, -7, -3, 7,
					-- layer=2 filter=141 channel=42
					12, 20, -15, 0, 13, -8, -30, -22, -30,
					-- layer=2 filter=141 channel=43
					8, -34, -8, -59, -21, 9, -17, -9, 5,
					-- layer=2 filter=141 channel=44
					10, -8, -5, 11, 8, 3, -7, 6, 6,
					-- layer=2 filter=141 channel=45
					-8, -6, -27, -50, -52, 13, 3, -76, -106,
					-- layer=2 filter=141 channel=46
					22, -1, 3, 36, -26, -6, 18, -6, 6,
					-- layer=2 filter=141 channel=47
					7, 24, -39, 17, 56, -32, 0, -2, -28,
					-- layer=2 filter=141 channel=48
					-3, -3, -4, 6, 0, -6, 3, 1, -3,
					-- layer=2 filter=141 channel=49
					9, -15, -31, -8, -36, -41, 6, -28, -15,
					-- layer=2 filter=141 channel=50
					-9, -3, 4, -4, 17, 1, 0, 4, 9,
					-- layer=2 filter=141 channel=51
					-18, 4, -1, -8, -13, 6, 7, 5, -3,
					-- layer=2 filter=141 channel=52
					-38, -20, 15, -9, -9, 40, -28, 3, 16,
					-- layer=2 filter=141 channel=53
					-30, -57, -20, -20, 62, 31, 2, -16, -21,
					-- layer=2 filter=141 channel=54
					60, 30, 28, 26, 19, 13, 0, -8, -31,
					-- layer=2 filter=141 channel=55
					2, 12, 0, 5, 14, 5, 0, -2, 2,
					-- layer=2 filter=141 channel=56
					-1, -17, -4, -21, 6, 7, -4, -5, 24,
					-- layer=2 filter=141 channel=57
					-7, 1, 8, 7, 3, -2, -5, 6, 4,
					-- layer=2 filter=141 channel=58
					14, 33, 9, 32, 29, 30, -20, 31, 27,
					-- layer=2 filter=141 channel=59
					-20, -35, 20, -13, 47, -12, -13, 4, -4,
					-- layer=2 filter=141 channel=60
					11, 5, -9, -5, 31, -16, -33, -2, -25,
					-- layer=2 filter=141 channel=61
					-23, -16, 7, -11, 29, -64, -27, 6, -27,
					-- layer=2 filter=141 channel=62
					-8, 9, 18, 15, 1, 10, 36, 0, -26,
					-- layer=2 filter=141 channel=63
					27, 12, 2, -11, -2, -33, -18, 7, -11,
					-- layer=2 filter=141 channel=64
					-5, 1, 1, 10, -15, -21, -31, -31, -18,
					-- layer=2 filter=141 channel=65
					-3, -13, 58, 9, 3, -49, -4, -9, -57,
					-- layer=2 filter=141 channel=66
					32, 17, -6, 5, -5, 39, 36, -28, 2,
					-- layer=2 filter=141 channel=67
					-10, -4, -16, 6, -14, -13, -15, 23, 51,
					-- layer=2 filter=141 channel=68
					-7, -2, -8, 10, 1, -3, -7, 0, -4,
					-- layer=2 filter=141 channel=69
					8, 23, 9, 1, -12, -8, -30, -2, -1,
					-- layer=2 filter=141 channel=70
					-2, -3, 17, 0, 21, 0, 6, -11, -12,
					-- layer=2 filter=141 channel=71
					-17, -13, -4, -31, 24, 15, -8, -24, -8,
					-- layer=2 filter=141 channel=72
					-3, 1, 17, -12, 54, 10, 14, 16, -6,
					-- layer=2 filter=141 channel=73
					-29, -47, -93, 0, -30, -24, 15, -29, -23,
					-- layer=2 filter=141 channel=74
					9, -6, -25, 21, -16, -19, -12, 4, 37,
					-- layer=2 filter=141 channel=75
					-9, -21, -8, -8, 46, -28, 0, -34, 1,
					-- layer=2 filter=141 channel=76
					-52, -51, -47, -9, 6, -18, 26, -20, -12,
					-- layer=2 filter=141 channel=77
					10, -8, 3, -9, 7, 4, 5, -8, -13,
					-- layer=2 filter=141 channel=78
					-1, -9, 0, -41, -15, 16, -13, -18, 28,
					-- layer=2 filter=141 channel=79
					-2, 1, -2, 8, 7, -9, -3, 4, -10,
					-- layer=2 filter=141 channel=80
					7, 3, -22, 10, 0, -13, -25, -13, 43,
					-- layer=2 filter=141 channel=81
					-6, -6, 6, -7, 0, 6, -18, -16, -3,
					-- layer=2 filter=141 channel=82
					5, -6, -3, -7, 2, 3, -7, 6, -8,
					-- layer=2 filter=141 channel=83
					-1, 14, 33, -26, 10, 9, -27, -27, 3,
					-- layer=2 filter=141 channel=84
					4, 4, -2, -9, 5, 10, 1, -3, -4,
					-- layer=2 filter=141 channel=85
					4, 0, -3, -1, 13, 10, 4, 9, 3,
					-- layer=2 filter=141 channel=86
					-1, 12, 16, 9, 0, 26, -2, 2, -3,
					-- layer=2 filter=141 channel=87
					-2, 0, 3, -3, 6, -19, 3, 16, 7,
					-- layer=2 filter=141 channel=88
					0, 19, 6, 2, -17, -9, -9, -8, -21,
					-- layer=2 filter=141 channel=89
					-39, -17, 20, 15, -3, -19, -14, 3, -20,
					-- layer=2 filter=141 channel=90
					4, 5, -7, 6, -6, -8, 10, 0, -1,
					-- layer=2 filter=141 channel=91
					-19, 5, 1, -6, 0, -20, -40, -25, -16,
					-- layer=2 filter=141 channel=92
					-8, 11, 41, 26, 20, 10, -16, 33, -40,
					-- layer=2 filter=141 channel=93
					28, 45, 25, -13, -21, -13, -13, -3, -16,
					-- layer=2 filter=141 channel=94
					-7, 21, 28, -16, -1, 36, -14, 5, 8,
					-- layer=2 filter=141 channel=95
					5, -6, 20, -3, 2, 0, 0, 0, -12,
					-- layer=2 filter=141 channel=96
					8, -47, 17, 30, 0, 0, -48, -1, 5,
					-- layer=2 filter=141 channel=97
					16, 0, -8, 23, 21, 10, -35, -18, 27,
					-- layer=2 filter=141 channel=98
					21, 9, -1, -7, 32, -20, 14, 11, -7,
					-- layer=2 filter=141 channel=99
					-50, -18, 2, 0, 17, -6, -43, 13, -9,
					-- layer=2 filter=141 channel=100
					-13, 4, -10, -32, 1, 26, -26, 0, 38,
					-- layer=2 filter=141 channel=101
					-27, 35, 4, -27, 0, -20, -40, -49, -19,
					-- layer=2 filter=141 channel=102
					-12, -15, 48, 22, -39, 2, 1, 16, 13,
					-- layer=2 filter=141 channel=103
					5, -34, 1, -50, -66, -29, 49, -15, -28,
					-- layer=2 filter=141 channel=104
					-23, -20, -8, -50, 11, 26, 3, -13, -4,
					-- layer=2 filter=141 channel=105
					-13, -31, 44, 34, 18, 17, -17, -3, 5,
					-- layer=2 filter=141 channel=106
					0, 1, -22, 4, 12, -25, -17, -26, -8,
					-- layer=2 filter=141 channel=107
					8, -8, -26, -41, 12, -19, 46, -20, -62,
					-- layer=2 filter=141 channel=108
					-27, -21, 21, 8, -33, 24, 12, -27, 11,
					-- layer=2 filter=141 channel=109
					-3, 3, 2, -1, -2, -17, 5, 6, 7,
					-- layer=2 filter=141 channel=110
					-6, -5, 2, -1, -4, -37, -33, -25, -86,
					-- layer=2 filter=141 channel=111
					-10, -9, 1, -6, 10, 0, -3, 4, -2,
					-- layer=2 filter=141 channel=112
					11, -18, 17, 31, 6, -16, 13, 3, 0,
					-- layer=2 filter=141 channel=113
					4, -8, 33, 24, -26, -15, 16, -15, -14,
					-- layer=2 filter=141 channel=114
					-1, 17, -13, 0, 3, -10, 15, 14, 4,
					-- layer=2 filter=141 channel=115
					0, -3, 7, 0, -5, 8, 1, 7, -2,
					-- layer=2 filter=141 channel=116
					5, -17, -2, 17, -1, 12, -20, 27, 25,
					-- layer=2 filter=141 channel=117
					7, -26, -10, -8, 8, -22, -8, -21, -69,
					-- layer=2 filter=141 channel=118
					3, -25, -16, -53, -26, -3, -20, 5, 28,
					-- layer=2 filter=141 channel=119
					-11, 52, -3, 12, 0, 25, 33, -5, 19,
					-- layer=2 filter=141 channel=120
					-2, 1, -4, -2, -4, 8, 7, -10, -5,
					-- layer=2 filter=141 channel=121
					-6, 6, -5, -6, 10, 4, 6, 5, 6,
					-- layer=2 filter=141 channel=122
					8, -9, -9, 9, 9, 7, 9, -4, 0,
					-- layer=2 filter=141 channel=123
					19, -7, 6, 0, 57, -15, 5, -3, -18,
					-- layer=2 filter=141 channel=124
					-5, 15, 12, 6, -3, 11, 10, 12, -11,
					-- layer=2 filter=141 channel=125
					2, -2, 6, 6, -4, 1, -1, -5, 6,
					-- layer=2 filter=141 channel=126
					-13, -68, 21, 45, 8, 3, -47, -30, -7,
					-- layer=2 filter=141 channel=127
					0, 9, 37, 24, -8, 12, -9, -8, -28,
					-- layer=2 filter=142 channel=0
					30, 15, 3, 36, 4, 12, 14, 18, 4,
					-- layer=2 filter=142 channel=1
					-17, -11, 14, -34, -38, -45, 9, -38, -47,
					-- layer=2 filter=142 channel=2
					3, 5, 0, -2, 8, -6, -6, 1, 4,
					-- layer=2 filter=142 channel=3
					21, 9, 4, 2, -10, -7, -25, -26, -29,
					-- layer=2 filter=142 channel=4
					28, 19, 3, 6, -5, -28, 1, 6, 6,
					-- layer=2 filter=142 channel=5
					2, 11, 9, 0, 5, -5, -14, 12, -16,
					-- layer=2 filter=142 channel=6
					12, 36, 29, 45, 15, 33, 63, 41, 25,
					-- layer=2 filter=142 channel=7
					20, 14, -13, -15, -72, -27, 18, -20, -6,
					-- layer=2 filter=142 channel=8
					7, 4, -3, -7, 2, 6, -5, -8, -6,
					-- layer=2 filter=142 channel=9
					-8, 4, 0, -6, 21, -8, -7, -24, -11,
					-- layer=2 filter=142 channel=10
					21, 17, -7, 25, 42, 8, 2, -13, -5,
					-- layer=2 filter=142 channel=11
					9, -1, -4, 19, -11, -8, 30, 14, -6,
					-- layer=2 filter=142 channel=12
					-6, -17, 30, -19, -45, -2, 7, -66, -59,
					-- layer=2 filter=142 channel=13
					-8, 3, -2, 7, 11, 5, -1, 2, 5,
					-- layer=2 filter=142 channel=14
					-1, 18, 12, -8, -38, -62, 25, -22, -15,
					-- layer=2 filter=142 channel=15
					31, -7, 3, 40, -32, 45, 13, 56, -9,
					-- layer=2 filter=142 channel=16
					33, -13, 11, 31, -21, -4, -21, -62, 3,
					-- layer=2 filter=142 channel=17
					9, -1, 4, -1, -3, 5, -8, 3, -10,
					-- layer=2 filter=142 channel=18
					-11, -29, -17, -32, -44, -5, -27, 3, 15,
					-- layer=2 filter=142 channel=19
					-32, -41, -1, 7, -1, 20, -35, -53, -29,
					-- layer=2 filter=142 channel=20
					-3, 4, 7, -2, 7, 0, 0, 1, 1,
					-- layer=2 filter=142 channel=21
					-5, -2, -11, 3, -7, -5, -4, -1, -13,
					-- layer=2 filter=142 channel=22
					0, 4, 2, 1, -7, 7, -9, 6, 8,
					-- layer=2 filter=142 channel=23
					10, 18, -10, 4, 23, 0, -21, -26, -10,
					-- layer=2 filter=142 channel=24
					19, 6, -34, -12, -21, -37, -48, -28, -25,
					-- layer=2 filter=142 channel=25
					1, 9, -40, -3, -13, -12, -16, 0, 21,
					-- layer=2 filter=142 channel=26
					3, -4, 2, 5, 6, -8, 9, -3, -9,
					-- layer=2 filter=142 channel=27
					-21, -8, 38, 13, 12, 20, 0, -12, 3,
					-- layer=2 filter=142 channel=28
					-30, 24, -32, 11, 1, -4, 20, -16, -1,
					-- layer=2 filter=142 channel=29
					-6, 4, -5, -3, 0, -3, -1, -2, 6,
					-- layer=2 filter=142 channel=30
					9, 5, -13, 8, 25, -25, -5, 10, -3,
					-- layer=2 filter=142 channel=31
					-15, 51, -8, 6, 80, 29, -22, 76, -4,
					-- layer=2 filter=142 channel=32
					6, -4, -1, -1, -3, 8, -6, 1, -1,
					-- layer=2 filter=142 channel=33
					37, -11, -9, 28, -54, -32, 18, 12, 27,
					-- layer=2 filter=142 channel=34
					-65, 9, 15, -28, 44, 24, 11, 16, 72,
					-- layer=2 filter=142 channel=35
					-31, -11, -23, 1, 11, 38, 28, -1, 13,
					-- layer=2 filter=142 channel=36
					11, -2, 0, -1, 3, -14, 9, -11, 10,
					-- layer=2 filter=142 channel=37
					-11, -15, 1, -1, 6, 0, -9, -4, -15,
					-- layer=2 filter=142 channel=38
					-17, -25, 16, 28, 12, -10, 37, 22, 21,
					-- layer=2 filter=142 channel=39
					23, -16, -5, -8, -38, -32, -19, -62, -8,
					-- layer=2 filter=142 channel=40
					14, -10, 43, 29, -21, -10, -49, -7, 67,
					-- layer=2 filter=142 channel=41
					2, -6, 2, -4, -3, 0, -6, -5, 0,
					-- layer=2 filter=142 channel=42
					29, -20, 32, -17, -21, 18, -15, -58, -10,
					-- layer=2 filter=142 channel=43
					-3, 10, 3, 14, 24, -14, 12, 3, 8,
					-- layer=2 filter=142 channel=44
					6, -8, 11, 7, 6, 8, 8, -7, 4,
					-- layer=2 filter=142 channel=45
					-45, -20, 1, -48, -37, -7, -7, 5, 31,
					-- layer=2 filter=142 channel=46
					4, 2, -5, 6, 16, -10, 3, 17, -8,
					-- layer=2 filter=142 channel=47
					6, 36, -2, 51, 0, -36, 25, 0, 11,
					-- layer=2 filter=142 channel=48
					7, 2, 7, 3, 6, -7, -7, 6, 4,
					-- layer=2 filter=142 channel=49
					13, 17, -11, -18, 1, 17, -34, -4, 47,
					-- layer=2 filter=142 channel=50
					-14, -18, -17, -6, -11, -8, -7, -8, -10,
					-- layer=2 filter=142 channel=51
					20, 5, -9, -3, 11, -18, 31, 36, 10,
					-- layer=2 filter=142 channel=52
					12, -11, 17, -3, -32, 1, 10, 0, -2,
					-- layer=2 filter=142 channel=53
					40, 6, -34, 3, -34, -18, 20, -19, -18,
					-- layer=2 filter=142 channel=54
					-19, -26, -16, 5, -13, 8, 27, -2, -19,
					-- layer=2 filter=142 channel=55
					-7, -7, 9, 0, -5, -2, 3, -5, -3,
					-- layer=2 filter=142 channel=56
					20, 19, 5, 24, 2, -18, 0, 0, -8,
					-- layer=2 filter=142 channel=57
					12, 6, 11, -3, 0, -5, -6, 7, 3,
					-- layer=2 filter=142 channel=58
					-29, -15, 8, 16, -4, -14, 17, -46, -63,
					-- layer=2 filter=142 channel=59
					-8, -20, 39, 28, -9, -7, -13, -6, -4,
					-- layer=2 filter=142 channel=60
					-30, -16, 9, 0, -34, 14, 5, -14, 3,
					-- layer=2 filter=142 channel=61
					-30, 5, 17, -7, -16, 23, -32, 0, 30,
					-- layer=2 filter=142 channel=62
					-30, -5, 8, -5, -27, -4, 0, 12, 41,
					-- layer=2 filter=142 channel=63
					25, 29, 25, 20, -27, 3, -2, -1, 43,
					-- layer=2 filter=142 channel=64
					13, 19, -16, 10, 0, -34, -15, -6, -14,
					-- layer=2 filter=142 channel=65
					-31, 5, 30, 3, 10, 39, -18, 24, 12,
					-- layer=2 filter=142 channel=66
					22, -3, -14, 15, -18, -3, -19, 8, -34,
					-- layer=2 filter=142 channel=67
					25, -9, -24, 14, 18, -32, 24, 16, -22,
					-- layer=2 filter=142 channel=68
					0, -6, -1, -2, 0, 10, 10, -8, 5,
					-- layer=2 filter=142 channel=69
					23, 14, 13, 0, -26, -30, 10, -40, -12,
					-- layer=2 filter=142 channel=70
					-26, -15, -16, 17, 15, 23, 7, -8, 15,
					-- layer=2 filter=142 channel=71
					-27, -12, -28, 32, 0, 3, 28, 10, 15,
					-- layer=2 filter=142 channel=72
					37, 2, 3, 15, 0, -12, -22, -61, -46,
					-- layer=2 filter=142 channel=73
					30, 67, 77, 44, 33, 8, 39, 6, -6,
					-- layer=2 filter=142 channel=74
					25, 6, 1, 17, 20, -22, 33, 4, 12,
					-- layer=2 filter=142 channel=75
					16, 29, 3, -2, 0, -22, 6, -24, 41,
					-- layer=2 filter=142 channel=76
					-17, 30, 14, 20, 17, -3, 6, 35, 3,
					-- layer=2 filter=142 channel=77
					-6, 9, -2, -5, 0, 9, 1, -4, -9,
					-- layer=2 filter=142 channel=78
					-23, -3, -33, 13, -22, -30, -6, 13, -23,
					-- layer=2 filter=142 channel=79
					11, 7, 12, 8, 9, -1, 2, 11, -2,
					-- layer=2 filter=142 channel=80
					6, -4, -3, 31, 19, 2, -30, -11, 5,
					-- layer=2 filter=142 channel=81
					-3, 0, 7, 5, 12, 1, 6, 9, 3,
					-- layer=2 filter=142 channel=82
					2, 0, 2, 6, 5, 0, 9, 9, 1,
					-- layer=2 filter=142 channel=83
					-6, 26, -1, 3, 9, 12, -27, -39, -12,
					-- layer=2 filter=142 channel=84
					9, -6, -9, 1, 10, 3, 0, 10, 0,
					-- layer=2 filter=142 channel=85
					-10, 6, -9, -17, -10, -4, -7, -3, -15,
					-- layer=2 filter=142 channel=86
					8, 2, 2, 11, -11, 0, -8, -18, 8,
					-- layer=2 filter=142 channel=87
					7, -25, -1, 2, -6, 7, 7, 17, 13,
					-- layer=2 filter=142 channel=88
					-4, 23, 2, -18, 21, -5, 15, 36, -5,
					-- layer=2 filter=142 channel=89
					-14, 0, 2, -26, -20, -23, -2, -40, -55,
					-- layer=2 filter=142 channel=90
					-4, -5, 0, 4, 0, 9, -7, -5, 0,
					-- layer=2 filter=142 channel=91
					-2, -11, 15, -1, -28, -23, 17, -65, 2,
					-- layer=2 filter=142 channel=92
					-36, -28, 10, 6, -3, 0, 0, -67, -52,
					-- layer=2 filter=142 channel=93
					-27, 16, -7, 35, -15, 15, 1, -20, -61,
					-- layer=2 filter=142 channel=94
					1, 12, 37, 0, -29, -9, 11, -68, -24,
					-- layer=2 filter=142 channel=95
					7, -2, 4, 9, -5, -9, -11, 7, 3,
					-- layer=2 filter=142 channel=96
					6, 42, 3, 0, 18, 40, 18, 34, 50,
					-- layer=2 filter=142 channel=97
					10, 25, 8, 35, -32, -25, -8, -10, -16,
					-- layer=2 filter=142 channel=98
					-22, 5, -4, 34, 5, 21, 15, -9, -1,
					-- layer=2 filter=142 channel=99
					-2, 5, -24, 25, -67, 6, 37, -11, -49,
					-- layer=2 filter=142 channel=100
					-10, -3, 31, 4, -12, 4, -5, -46, -36,
					-- layer=2 filter=142 channel=101
					14, 17, -15, 38, 13, -2, 4, 17, 14,
					-- layer=2 filter=142 channel=102
					23, 3, -26, 1, 0, 17, -9, -12, -9,
					-- layer=2 filter=142 channel=103
					-7, 75, 2, 35, 64, -17, 59, 43, 47,
					-- layer=2 filter=142 channel=104
					18, 7, -28, -32, -21, 12, -23, 6, -4,
					-- layer=2 filter=142 channel=105
					-21, -2, 8, -10, -11, -15, 7, -28, -19,
					-- layer=2 filter=142 channel=106
					43, 17, -16, 38, 15, -26, 16, 0, 2,
					-- layer=2 filter=142 channel=107
					14, 13, 53, -19, 40, -13, 27, -21, -34,
					-- layer=2 filter=142 channel=108
					-40, -22, -15, -14, -14, 13, -4, 0, 9,
					-- layer=2 filter=142 channel=109
					5, 13, -16, -9, 10, -4, 6, 0, -8,
					-- layer=2 filter=142 channel=110
					-6, 4, -49, -31, -12, -42, -94, -61, -49,
					-- layer=2 filter=142 channel=111
					10, 5, 1, -9, 5, 11, 3, 6, 0,
					-- layer=2 filter=142 channel=112
					26, 9, -19, 8, 22, 0, 13, 20, 26,
					-- layer=2 filter=142 channel=113
					3, 17, -36, 28, 1, -9, 4, 6, -24,
					-- layer=2 filter=142 channel=114
					8, -8, 9, 11, -13, 6, 11, -2, 9,
					-- layer=2 filter=142 channel=115
					1, 4, 0, -1, -8, -3, 4, -10, -9,
					-- layer=2 filter=142 channel=116
					11, 20, -1, -32, -28, -7, -12, 3, 48,
					-- layer=2 filter=142 channel=117
					37, -2, 27, 13, -1, -3, 31, -32, -7,
					-- layer=2 filter=142 channel=118
					-6, -4, 2, 14, 9, -5, -34, 28, 28,
					-- layer=2 filter=142 channel=119
					33, -29, -6, -9, -16, -12, -21, -31, 25,
					-- layer=2 filter=142 channel=120
					10, 10, -9, 0, 10, 0, -8, -5, 4,
					-- layer=2 filter=142 channel=121
					6, 0, 0, -5, 1, 1, 0, 8, -7,
					-- layer=2 filter=142 channel=122
					-3, -3, -2, 0, 4, -3, 8, -1, -16,
					-- layer=2 filter=142 channel=123
					20, 11, -3, 43, -43, 7, 30, -10, -16,
					-- layer=2 filter=142 channel=124
					13, -41, -18, 30, 11, -2, 7, 75, -44,
					-- layer=2 filter=142 channel=125
					1, -12, 8, -2, -1, 13, 4, 0, -9,
					-- layer=2 filter=142 channel=126
					-6, 87, -10, 56, 22, 29, 30, -7, -27,
					-- layer=2 filter=142 channel=127
					-10, 8, 20, -8, 13, -12, -12, -1, 11,
					-- layer=2 filter=143 channel=0
					9, -5, -18, 19, -20, 17, 27, -2, 19,
					-- layer=2 filter=143 channel=1
					-2, 28, 13, -9, -3, 21, 37, 0, 23,
					-- layer=2 filter=143 channel=2
					9, -5, 3, -9, -2, 3, -1, -3, -1,
					-- layer=2 filter=143 channel=3
					-40, -20, -6, 8, -39, -7, -10, -45, -36,
					-- layer=2 filter=143 channel=4
					-33, -4, 8, -6, -17, -6, 4, 21, 10,
					-- layer=2 filter=143 channel=5
					13, 6, -36, 20, -7, -7, 1, 8, -5,
					-- layer=2 filter=143 channel=6
					0, 16, 19, -14, -7, -22, 15, 23, -3,
					-- layer=2 filter=143 channel=7
					-11, -31, 29, -6, 0, 20, -2, 9, -9,
					-- layer=2 filter=143 channel=8
					2, 2, 8, 2, -2, -3, -8, -5, 1,
					-- layer=2 filter=143 channel=9
					-34, -11, -7, -21, -25, -37, -1, 22, 4,
					-- layer=2 filter=143 channel=10
					7, -1, -27, 19, -14, 13, 32, 1, 11,
					-- layer=2 filter=143 channel=11
					-8, 13, 18, 7, 8, -7, 3, 8, 9,
					-- layer=2 filter=143 channel=12
					-23, 11, -3, -43, -7, -6, 2, -12, 7,
					-- layer=2 filter=143 channel=13
					0, -2, 0, 6, -8, -7, -3, 2, -9,
					-- layer=2 filter=143 channel=14
					10, 24, 24, -9, -7, 3, 17, 5, 32,
					-- layer=2 filter=143 channel=15
					24, 22, 38, 0, -17, 17, 27, -7, 0,
					-- layer=2 filter=143 channel=16
					-22, -4, -6, -27, -63, -35, -6, 3, -42,
					-- layer=2 filter=143 channel=17
					0, -3, -1, 7, -4, 7, 11, 11, 7,
					-- layer=2 filter=143 channel=18
					4, 29, 12, 6, 33, 14, 0, 37, 20,
					-- layer=2 filter=143 channel=19
					37, 29, 0, 3, 13, 16, 23, 24, 15,
					-- layer=2 filter=143 channel=20
					-1, 3, -9, -10, -6, 3, -1, -8, -7,
					-- layer=2 filter=143 channel=21
					7, 4, -9, 2, 9, 6, -16, 2, -5,
					-- layer=2 filter=143 channel=22
					-1, -1, -2, -4, 4, -11, 2, 4, 0,
					-- layer=2 filter=143 channel=23
					-33, -41, -40, -35, 2, -26, 12, 0, -29,
					-- layer=2 filter=143 channel=24
					-44, -52, -29, -41, -95, -54, -8, -83, -53,
					-- layer=2 filter=143 channel=25
					-25, -32, 0, -25, -67, -34, -2, -61, -39,
					-- layer=2 filter=143 channel=26
					8, -4, -6, 5, 0, 7, 5, 6, -5,
					-- layer=2 filter=143 channel=27
					0, -4, -11, -1, -25, -17, 0, 1, 19,
					-- layer=2 filter=143 channel=28
					1, 10, -7, 4, 4, 54, -1, 26, 21,
					-- layer=2 filter=143 channel=29
					8, -7, 7, 6, -10, 3, -8, -2, -7,
					-- layer=2 filter=143 channel=30
					9, -22, -34, 6, -7, -21, 10, 10, 11,
					-- layer=2 filter=143 channel=31
					-16, 41, -32, -23, -51, -24, -18, -9, 35,
					-- layer=2 filter=143 channel=32
					7, 6, -1, -4, 5, 9, 0, 8, -4,
					-- layer=2 filter=143 channel=33
					-10, -5, 24, -45, -67, 27, 9, -35, 27,
					-- layer=2 filter=143 channel=34
					-22, 16, 19, -26, 13, 17, -32, 1, 11,
					-- layer=2 filter=143 channel=35
					3, -8, -3, 12, -4, 35, -6, -29, -13,
					-- layer=2 filter=143 channel=36
					-9, -6, 3, -9, 8, 6, -1, 8, -1,
					-- layer=2 filter=143 channel=37
					6, 15, -6, 16, 5, -12, 14, 0, 16,
					-- layer=2 filter=143 channel=38
					-12, -16, -13, -14, -14, 1, 9, 9, 7,
					-- layer=2 filter=143 channel=39
					-51, -74, 1, 22, -7, -61, 16, 2, -18,
					-- layer=2 filter=143 channel=40
					14, 42, 11, -4, 24, 46, -31, -3, 33,
					-- layer=2 filter=143 channel=41
					11, -4, -3, -4, 3, 8, -6, -7, 4,
					-- layer=2 filter=143 channel=42
					-66, -6, -34, -45, -53, -40, -46, -7, -33,
					-- layer=2 filter=143 channel=43
					16, -12, -31, 1, -21, -2, -3, -2, 5,
					-- layer=2 filter=143 channel=44
					-7, -4, 0, 3, -9, -5, -9, 6, -5,
					-- layer=2 filter=143 channel=45
					-25, -32, -40, 7, -81, -15, 2, -23, -11,
					-- layer=2 filter=143 channel=46
					20, 0, -25, 23, -18, -32, 17, 13, 26,
					-- layer=2 filter=143 channel=47
					-33, -14, -8, -33, -37, 15, 0, -4, -4,
					-- layer=2 filter=143 channel=48
					-4, -7, -2, 0, 10, 8, 6, 4, -7,
					-- layer=2 filter=143 channel=49
					-18, 14, 13, 1, 32, -11, -23, -18, -34,
					-- layer=2 filter=143 channel=50
					-11, -12, -3, -1, 16, -2, 9, -19, 1,
					-- layer=2 filter=143 channel=51
					9, -7, -2, 7, 9, 2, 14, 19, 17,
					-- layer=2 filter=143 channel=52
					-4, 4, 8, 13, 5, -4, 0, -5, 3,
					-- layer=2 filter=143 channel=53
					-45, 12, -33, -11, 31, -7, 33, 33, 34,
					-- layer=2 filter=143 channel=54
					0, 29, 2, -8, 13, 30, 0, 2, -2,
					-- layer=2 filter=143 channel=55
					-8, 2, 5, -6, 3, -12, 0, 7, -3,
					-- layer=2 filter=143 channel=56
					-11, 10, 9, -6, 0, -25, 4, 6, 3,
					-- layer=2 filter=143 channel=57
					-7, 5, 14, -4, 13, 8, 2, 1, 3,
					-- layer=2 filter=143 channel=58
					-2, 17, 0, -34, -5, 0, 7, -35, 1,
					-- layer=2 filter=143 channel=59
					5, -2, 7, -7, 34, 5, 27, 1, 22,
					-- layer=2 filter=143 channel=60
					18, 8, 9, -6, 16, 44, 41, -2, 1,
					-- layer=2 filter=143 channel=61
					16, -4, -10, 5, 22, -40, 56, 11, -35,
					-- layer=2 filter=143 channel=62
					-6, -2, 5, -33, -10, -4, 1, 0, -27,
					-- layer=2 filter=143 channel=63
					3, -35, 3, 1, 4, -14, 33, 0, -9,
					-- layer=2 filter=143 channel=64
					-49, -68, -23, -49, -49, -40, -34, -19, -42,
					-- layer=2 filter=143 channel=65
					31, 9, 3, -10, 0, -21, 34, 16, -64,
					-- layer=2 filter=143 channel=66
					8, 10, -23, -36, 43, -29, -2, -2, -22,
					-- layer=2 filter=143 channel=67
					0, 0, -3, 10, -3, -12, 2, -8, 14,
					-- layer=2 filter=143 channel=68
					2, 5, 2, -13, -9, 3, 0, 0, -7,
					-- layer=2 filter=143 channel=69
					-41, -21, 0, -32, -27, -39, -38, -48, -39,
					-- layer=2 filter=143 channel=70
					34, 11, -7, 9, -4, 40, -11, -9, 27,
					-- layer=2 filter=143 channel=71
					-4, 0, -1, -21, -29, 20, -18, 0, 10,
					-- layer=2 filter=143 channel=72
					1, 8, 45, 17, -2, 25, 1, 3, 14,
					-- layer=2 filter=143 channel=73
					-25, -7, 14, -2, 10, 24, 0, -9, -13,
					-- layer=2 filter=143 channel=74
					-7, -5, 27, 24, 5, 11, 29, 0, 57,
					-- layer=2 filter=143 channel=75
					-9, 25, 10, -22, -31, 12, -24, -54, 27,
					-- layer=2 filter=143 channel=76
					-25, -25, -21, -42, 9, -10, -37, -5, 21,
					-- layer=2 filter=143 channel=77
					4, 12, -5, -2, -2, 4, 0, -6, 5,
					-- layer=2 filter=143 channel=78
					-6, 3, 0, 0, -1, -1, 14, 11, -23,
					-- layer=2 filter=143 channel=79
					6, 1, -2, -10, -8, -1, 7, 5, -3,
					-- layer=2 filter=143 channel=80
					-17, -6, -12, -2, -24, -15, 29, 1, 11,
					-- layer=2 filter=143 channel=81
					-16, -7, -4, -3, -9, 0, 0, 0, -1,
					-- layer=2 filter=143 channel=82
					2, 1, -7, -1, 3, -9, 0, 0, 5,
					-- layer=2 filter=143 channel=83
					2, -9, -22, 12, -24, -18, 5, 1, -26,
					-- layer=2 filter=143 channel=84
					6, -3, -8, 0, -9, -10, 2, 7, -2,
					-- layer=2 filter=143 channel=85
					4, 4, 12, -12, 10, -12, 8, 10, 0,
					-- layer=2 filter=143 channel=86
					2, -2, 7, 5, 16, 11, -9, -16, 4,
					-- layer=2 filter=143 channel=87
					9, 23, -33, -27, 30, 7, -6, -13, -39,
					-- layer=2 filter=143 channel=88
					9, -13, 10, 10, -6, -2, 26, -14, 8,
					-- layer=2 filter=143 channel=89
					0, 16, 19, -13, 2, 7, -7, -9, -3,
					-- layer=2 filter=143 channel=90
					-3, 6, -5, -3, 3, 7, 0, 9, 10,
					-- layer=2 filter=143 channel=91
					-20, 20, 16, -35, -30, 2, -24, -32, -33,
					-- layer=2 filter=143 channel=92
					-2, 21, -16, -20, -19, -11, 5, -5, -23,
					-- layer=2 filter=143 channel=93
					37, 9, 16, -21, -63, -4, -28, -34, -8,
					-- layer=2 filter=143 channel=94
					-8, 1, -7, 16, 23, -29, 60, 43, 9,
					-- layer=2 filter=143 channel=95
					-8, -9, -5, 1, 2, 6, 1, -7, 8,
					-- layer=2 filter=143 channel=96
					18, 33, 15, -3, 24, 25, 1, -7, 23,
					-- layer=2 filter=143 channel=97
					-19, -4, 10, -40, -39, -37, -17, -14, -3,
					-- layer=2 filter=143 channel=98
					-7, 10, -3, 12, 3, 24, 8, 5, 19,
					-- layer=2 filter=143 channel=99
					4, 4, 35, -8, 39, 28, 0, 30, 68,
					-- layer=2 filter=143 channel=100
					-5, 9, -56, -5, -27, 7, 23, -3, -12,
					-- layer=2 filter=143 channel=101
					26, 36, 25, -14, -24, 22, -17, -22, 4,
					-- layer=2 filter=143 channel=102
					-23, 9, 50, 0, 9, -1, -27, -15, -21,
					-- layer=2 filter=143 channel=103
					36, -26, 8, -57, -22, -1, 31, 10, 7,
					-- layer=2 filter=143 channel=104
					-30, 19, 10, 28, 40, 16, 23, 7, -8,
					-- layer=2 filter=143 channel=105
					35, 3, -10, 0, -4, -17, 14, -7, 1,
					-- layer=2 filter=143 channel=106
					-36, 13, 44, -35, -29, 14, 19, -40, 25,
					-- layer=2 filter=143 channel=107
					-34, -45, -23, -37, -13, -31, 17, -3, -35,
					-- layer=2 filter=143 channel=108
					-2, -10, 16, -8, -28, 8, 5, 1, 3,
					-- layer=2 filter=143 channel=109
					-6, -1, 3, 0, 3, 5, 4, -1, 3,
					-- layer=2 filter=143 channel=110
					-20, -4, -15, -25, -30, -42, -40, -41, -9,
					-- layer=2 filter=143 channel=111
					-1, -4, -5, 7, 6, 4, 3, 7, 0,
					-- layer=2 filter=143 channel=112
					-21, -15, 8, -2, 5, -11, 11, 6, -29,
					-- layer=2 filter=143 channel=113
					-4, -28, -5, 12, -32, -1, -2, 8, -16,
					-- layer=2 filter=143 channel=114
					5, 2, -5, -10, -11, 5, -10, 0, 3,
					-- layer=2 filter=143 channel=115
					-8, 2, 4, -6, 7, -7, -3, 7, -1,
					-- layer=2 filter=143 channel=116
					2, 38, 5, -20, 24, 31, -6, -10, -30,
					-- layer=2 filter=143 channel=117
					32, 15, 23, 7, 4, 30, -8, 35, 16,
					-- layer=2 filter=143 channel=118
					9, 11, -18, 8, 13, 3, 17, -1, -10,
					-- layer=2 filter=143 channel=119
					-12, 11, -10, -2, 27, 0, -17, 0, 10,
					-- layer=2 filter=143 channel=120
					5, -6, -6, 6, -4, -3, -7, -2, -6,
					-- layer=2 filter=143 channel=121
					-1, -4, 5, -7, 4, 0, 8, -8, -6,
					-- layer=2 filter=143 channel=122
					13, 1, 16, 2, -1, -5, 0, 3, 6,
					-- layer=2 filter=143 channel=123
					34, 7, 42, -4, 19, 26, -9, -2, 42,
					-- layer=2 filter=143 channel=124
					11, 26, 14, -45, -32, -2, -2, 9, 23,
					-- layer=2 filter=143 channel=125
					-9, 0, -10, 7, 6, 6, -2, 1, -7,
					-- layer=2 filter=143 channel=126
					53, -54, -16, -8, -79, 15, 12, -27, -13,
					-- layer=2 filter=143 channel=127
					3, -19, -23, 6, -12, 3, 40, -33, 5,
					-- layer=2 filter=144 channel=0
					-1, -7, 1, 6, -6, 7, 1, 2, 9,
					-- layer=2 filter=144 channel=1
					-8, -13, -1, -2, -7, -10, -13, -11, 0,
					-- layer=2 filter=144 channel=2
					-6, 1, -6, 7, 4, -4, -4, 5, 8,
					-- layer=2 filter=144 channel=3
					3, 8, -4, 6, 6, -3, -5, 7, -1,
					-- layer=2 filter=144 channel=4
					0, -4, 1, 0, -9, 6, 5, -4, -7,
					-- layer=2 filter=144 channel=5
					-9, -9, -7, 6, 5, -8, -7, 4, -3,
					-- layer=2 filter=144 channel=6
					0, -11, -8, -7, 7, 0, -3, 2, 6,
					-- layer=2 filter=144 channel=7
					2, 4, -1, -11, 5, -13, -7, 1, -2,
					-- layer=2 filter=144 channel=8
					8, -4, -4, -7, 4, -2, 6, 3, -5,
					-- layer=2 filter=144 channel=9
					5, 1, 6, -9, -6, 8, -1, -3, -1,
					-- layer=2 filter=144 channel=10
					2, -1, 4, 8, -1, -5, -7, 4, -5,
					-- layer=2 filter=144 channel=11
					-12, 0, 5, 6, -11, -1, -2, -13, -3,
					-- layer=2 filter=144 channel=12
					-5, -9, 3, -2, -6, 1, -13, -12, 0,
					-- layer=2 filter=144 channel=13
					6, 1, 6, -8, 9, 0, 1, 3, 7,
					-- layer=2 filter=144 channel=14
					-9, -2, -10, -7, 7, -8, -6, -4, 6,
					-- layer=2 filter=144 channel=15
					-4, -11, 6, -10, 8, 2, 2, -10, 0,
					-- layer=2 filter=144 channel=16
					5, -3, -5, 5, -9, -6, 0, 1, 1,
					-- layer=2 filter=144 channel=17
					-11, 0, 0, 0, 10, 6, 10, -9, 5,
					-- layer=2 filter=144 channel=18
					-6, -13, -9, 7, -4, 6, 2, 0, -9,
					-- layer=2 filter=144 channel=19
					-9, -5, -14, -3, -1, -10, -4, 4, 0,
					-- layer=2 filter=144 channel=20
					-8, 2, -2, 0, -4, 4, -6, -3, 4,
					-- layer=2 filter=144 channel=21
					-2, 6, -9, 3, -5, -5, -3, -8, 5,
					-- layer=2 filter=144 channel=22
					-1, 4, -2, 3, 5, -8, -5, 1, -3,
					-- layer=2 filter=144 channel=23
					-12, -11, -2, 2, -2, 3, -2, 4, -1,
					-- layer=2 filter=144 channel=24
					-1, -7, 2, -6, 4, 0, -6, 5, -9,
					-- layer=2 filter=144 channel=25
					-4, -10, -2, -14, -2, -11, 5, -5, -1,
					-- layer=2 filter=144 channel=26
					-9, -1, 0, -4, -2, 3, -1, 5, -8,
					-- layer=2 filter=144 channel=27
					-5, 8, -11, -6, -9, 2, -3, -2, 4,
					-- layer=2 filter=144 channel=28
					1, 0, -3, -4, -9, 0, 7, 0, 8,
					-- layer=2 filter=144 channel=29
					8, 1, -5, -9, -6, 4, 0, -7, -7,
					-- layer=2 filter=144 channel=30
					8, -6, -4, -8, 6, 1, 6, 2, 5,
					-- layer=2 filter=144 channel=31
					2, -12, -10, -7, 1, 0, 3, 7, -9,
					-- layer=2 filter=144 channel=32
					3, -3, -4, 9, 0, -7, -9, -2, 9,
					-- layer=2 filter=144 channel=33
					0, -2, 5, -5, -7, -4, 5, 9, 1,
					-- layer=2 filter=144 channel=34
					0, -11, 8, 0, -8, -9, -7, -7, -10,
					-- layer=2 filter=144 channel=35
					0, 3, 5, 0, 5, -3, -11, -14, -11,
					-- layer=2 filter=144 channel=36
					6, 3, -12, -3, 6, -7, 0, -1, 1,
					-- layer=2 filter=144 channel=37
					-9, -4, -4, -6, 1, -12, -9, -12, -2,
					-- layer=2 filter=144 channel=38
					5, -1, 8, -10, 6, -7, 3, 3, -9,
					-- layer=2 filter=144 channel=39
					-7, 7, 0, 6, -5, -7, -8, -4, -3,
					-- layer=2 filter=144 channel=40
					3, -3, 3, 3, -10, -10, -3, -10, 1,
					-- layer=2 filter=144 channel=41
					-2, -8, 4, 6, -7, 9, -4, -5, 1,
					-- layer=2 filter=144 channel=42
					6, -11, -5, 6, 4, 5, -4, 4, 6,
					-- layer=2 filter=144 channel=43
					-10, -8, -1, 5, -6, 6, 6, 7, 2,
					-- layer=2 filter=144 channel=44
					-2, 5, 1, 0, -2, -2, -7, 4, -6,
					-- layer=2 filter=144 channel=45
					-4, -4, 9, -1, 3, 0, -7, -4, -5,
					-- layer=2 filter=144 channel=46
					-5, -8, -2, -3, -6, -11, -9, 6, -9,
					-- layer=2 filter=144 channel=47
					-6, 1, 4, -4, 0, 4, -10, 9, -4,
					-- layer=2 filter=144 channel=48
					0, 10, -1, 11, 8, 1, -2, 4, -5,
					-- layer=2 filter=144 channel=49
					-8, -9, -9, 2, -10, 0, 4, 4, 0,
					-- layer=2 filter=144 channel=50
					9, 2, 9, -9, 9, 11, -7, -3, 3,
					-- layer=2 filter=144 channel=51
					-1, 5, 2, -10, -6, 7, -11, 5, 2,
					-- layer=2 filter=144 channel=52
					-5, -10, -5, 3, -8, 7, -13, -4, -3,
					-- layer=2 filter=144 channel=53
					-5, 1, 1, -9, 5, 0, -5, 4, -4,
					-- layer=2 filter=144 channel=54
					0, -3, -15, -7, 3, -9, 0, 0, -5,
					-- layer=2 filter=144 channel=55
					6, -7, -5, -5, 0, 5, 1, -7, 3,
					-- layer=2 filter=144 channel=56
					-4, -11, -2, -12, -1, -8, 2, -5, 1,
					-- layer=2 filter=144 channel=57
					2, 7, -4, -5, 0, -5, 2, -2, 2,
					-- layer=2 filter=144 channel=58
					-6, -1, -11, -4, 1, -3, -4, 8, 2,
					-- layer=2 filter=144 channel=59
					-15, 8, 6, 1, 3, -12, 5, -7, 0,
					-- layer=2 filter=144 channel=60
					-5, 3, -3, 0, 5, 6, -4, -5, 7,
					-- layer=2 filter=144 channel=61
					0, -9, -10, -4, -2, 2, -12, 7, -5,
					-- layer=2 filter=144 channel=62
					-6, -10, 4, -13, -16, -11, -8, -3, -8,
					-- layer=2 filter=144 channel=63
					-3, 5, -6, -12, 3, 4, -12, -5, 4,
					-- layer=2 filter=144 channel=64
					5, -11, -12, 5, -8, 4, 7, -2, 6,
					-- layer=2 filter=144 channel=65
					0, -2, -6, -3, -9, 4, -1, -5, 5,
					-- layer=2 filter=144 channel=66
					-5, 3, 5, 2, -7, 4, -3, 0, 0,
					-- layer=2 filter=144 channel=67
					-10, 2, 1, 5, 5, 3, -5, 0, 6,
					-- layer=2 filter=144 channel=68
					-8, 1, 3, 7, 4, 1, -8, -8, -9,
					-- layer=2 filter=144 channel=69
					-10, -1, -6, 1, 0, -8, -9, -12, -13,
					-- layer=2 filter=144 channel=70
					-3, 3, -14, -11, 0, 2, -13, 5, -8,
					-- layer=2 filter=144 channel=71
					6, -3, -10, -5, 2, -7, -6, -11, -11,
					-- layer=2 filter=144 channel=72
					5, -7, -6, 6, -11, -8, -5, 1, -3,
					-- layer=2 filter=144 channel=73
					-6, -14, 1, 1, -7, -14, 1, -4, -4,
					-- layer=2 filter=144 channel=74
					0, -8, -7, 9, 3, -11, -4, -7, 1,
					-- layer=2 filter=144 channel=75
					7, 5, -2, 1, 1, -8, 8, 7, 5,
					-- layer=2 filter=144 channel=76
					-9, -1, 0, -12, 5, -8, 8, 0, -3,
					-- layer=2 filter=144 channel=77
					-9, 0, -9, 3, 7, 2, -8, 0, -9,
					-- layer=2 filter=144 channel=78
					6, 0, -9, -6, -4, 0, 8, 1, -9,
					-- layer=2 filter=144 channel=79
					4, -1, -1, 0, -9, -3, -3, 1, 5,
					-- layer=2 filter=144 channel=80
					-2, 9, 4, -1, -11, 0, -3, 6, -9,
					-- layer=2 filter=144 channel=81
					-4, -10, -7, 3, 2, 0, 4, 2, -7,
					-- layer=2 filter=144 channel=82
					-2, 4, 0, 11, 0, -6, -8, -1, 5,
					-- layer=2 filter=144 channel=83
					-9, 2, 3, -10, 2, -11, 0, -3, -3,
					-- layer=2 filter=144 channel=84
					-5, -2, 4, -8, 0, -1, 1, 5, 3,
					-- layer=2 filter=144 channel=85
					-7, 2, -4, -5, 10, 5, 7, -8, 6,
					-- layer=2 filter=144 channel=86
					0, -2, -2, -10, -1, -7, 2, -8, 7,
					-- layer=2 filter=144 channel=87
					1, -1, -2, 0, -9, 2, -1, -8, -1,
					-- layer=2 filter=144 channel=88
					0, -5, -7, 0, -6, 4, -8, 1, 3,
					-- layer=2 filter=144 channel=89
					-10, -2, -10, -7, -1, 0, 6, 6, -10,
					-- layer=2 filter=144 channel=90
					7, 9, -4, -4, 10, -3, -6, 1, 5,
					-- layer=2 filter=144 channel=91
					-16, -9, -12, -10, -13, 6, -5, 0, 2,
					-- layer=2 filter=144 channel=92
					1, 0, 3, -2, -1, 0, -3, 1, -9,
					-- layer=2 filter=144 channel=93
					-8, -3, -13, 1, -6, -11, -3, 6, 3,
					-- layer=2 filter=144 channel=94
					0, -13, -8, -15, -13, -11, -16, 3, -4,
					-- layer=2 filter=144 channel=95
					-9, -2, -3, -11, 0, -2, -7, 2, -9,
					-- layer=2 filter=144 channel=96
					-4, 5, -3, -1, -10, -5, -7, 0, -3,
					-- layer=2 filter=144 channel=97
					-9, 3, -10, 2, -8, 4, -9, -10, -6,
					-- layer=2 filter=144 channel=98
					-3, 2, 2, -9, 3, 3, -10, 3, -11,
					-- layer=2 filter=144 channel=99
					-11, -3, 1, -13, -15, -7, -14, -15, -1,
					-- layer=2 filter=144 channel=100
					1, -6, 12, 4, 1, -7, -7, 3, -1,
					-- layer=2 filter=144 channel=101
					8, 0, -11, -8, 3, -11, 3, -12, 4,
					-- layer=2 filter=144 channel=102
					7, -4, -2, -2, -10, -7, 0, 4, 5,
					-- layer=2 filter=144 channel=103
					-7, 0, -9, -1, 2, 3, 1, 5, -4,
					-- layer=2 filter=144 channel=104
					-7, 3, -10, -3, 6, -9, 3, -9, 3,
					-- layer=2 filter=144 channel=105
					7, -2, 7, -2, 7, 4, -3, -3, -6,
					-- layer=2 filter=144 channel=106
					-9, -6, -13, 10, 2, -1, 4, -4, 1,
					-- layer=2 filter=144 channel=107
					8, -2, 3, 0, -8, -10, -7, 5, -6,
					-- layer=2 filter=144 channel=108
					6, 3, 4, -4, 0, 4, -3, 4, 7,
					-- layer=2 filter=144 channel=109
					4, 3, 11, 5, -3, -8, 10, 7, 9,
					-- layer=2 filter=144 channel=110
					-8, -7, -9, 0, -4, -11, 2, 2, -7,
					-- layer=2 filter=144 channel=111
					2, 6, -3, -1, -7, -9, 1, 0, 6,
					-- layer=2 filter=144 channel=112
					-13, -3, -1, -10, 1, 6, 1, 0, -7,
					-- layer=2 filter=144 channel=113
					-11, 6, -12, 5, 2, 7, 7, 6, -8,
					-- layer=2 filter=144 channel=114
					6, -2, 4, 0, 0, -9, 7, 0, -4,
					-- layer=2 filter=144 channel=115
					2, 1, 7, 2, 9, 6, -2, -3, 5,
					-- layer=2 filter=144 channel=116
					-2, -11, -4, -2, -1, -8, -3, 4, -2,
					-- layer=2 filter=144 channel=117
					4, -1, 4, -5, -3, -13, -1, -13, 2,
					-- layer=2 filter=144 channel=118
					-6, -11, -5, 9, 1, 7, -2, 4, -2,
					-- layer=2 filter=144 channel=119
					-5, -9, 0, -7, -2, -4, 3, -1, -1,
					-- layer=2 filter=144 channel=120
					5, -3, 10, -5, 1, -2, 8, 9, 0,
					-- layer=2 filter=144 channel=121
					3, 5, -11, 4, -3, 0, -7, -10, 3,
					-- layer=2 filter=144 channel=122
					5, -5, 3, 10, 2, 0, 10, -1, -3,
					-- layer=2 filter=144 channel=123
					0, -13, -4, -11, 5, 1, -6, -6, -17,
					-- layer=2 filter=144 channel=124
					-5, -6, -1, 7, -7, 3, -9, 2, 1,
					-- layer=2 filter=144 channel=125
					-2, -7, 11, 3, 2, 6, 8, -11, 6,
					-- layer=2 filter=144 channel=126
					0, -5, 3, 3, 6, 6, 3, 6, 6,
					-- layer=2 filter=144 channel=127
					7, 10, -3, -12, -3, -10, -2, -4, 7,
					-- layer=2 filter=145 channel=0
					0, 21, 7, 2, 9, 41, 0, -1, 12,
					-- layer=2 filter=145 channel=1
					36, -15, -17, 3, 10, 3, 15, 18, 9,
					-- layer=2 filter=145 channel=2
					0, 6, 1, -2, -1, -5, 5, -2, -10,
					-- layer=2 filter=145 channel=3
					9, 12, -7, 2, 23, 3, -11, -4, -15,
					-- layer=2 filter=145 channel=4
					37, 27, -28, 33, -6, -85, 18, -30, -49,
					-- layer=2 filter=145 channel=5
					-19, -7, 41, -30, -1, 44, -27, 13, 39,
					-- layer=2 filter=145 channel=6
					-24, -44, -18, -36, -40, -37, -39, -21, -36,
					-- layer=2 filter=145 channel=7
					7, 0, -12, -18, -28, -43, 0, 23, -24,
					-- layer=2 filter=145 channel=8
					7, 7, -4, -7, -6, -2, 5, -2, 4,
					-- layer=2 filter=145 channel=9
					25, 27, -15, -8, 9, -39, -16, -20, -22,
					-- layer=2 filter=145 channel=10
					24, 22, -6, 18, 16, 24, -15, -11, 12,
					-- layer=2 filter=145 channel=11
					-40, 20, 34, -24, 16, 40, -31, 1, 39,
					-- layer=2 filter=145 channel=12
					7, -5, -6, 8, -12, 1, 19, 38, 1,
					-- layer=2 filter=145 channel=13
					-3, 3, -7, -4, -5, 11, -2, 9, -11,
					-- layer=2 filter=145 channel=14
					-14, -18, 15, -1, 13, 6, 11, 15, 7,
					-- layer=2 filter=145 channel=15
					-34, -35, 16, 15, 34, 77, 13, -16, 20,
					-- layer=2 filter=145 channel=16
					38, 12, -48, 29, -3, -85, 19, -21, -80,
					-- layer=2 filter=145 channel=17
					0, -5, -4, -6, 2, 8, -1, 9, 0,
					-- layer=2 filter=145 channel=18
					0, -19, 2, 4, 10, 12, 50, 30, 40,
					-- layer=2 filter=145 channel=19
					-9, -17, 8, 7, 1, -5, 13, 2, -12,
					-- layer=2 filter=145 channel=20
					11, 6, 2, 2, 4, -6, 1, 8, 6,
					-- layer=2 filter=145 channel=21
					4, 7, 3, 1, 4, -2, 5, 2, -8,
					-- layer=2 filter=145 channel=22
					-4, 0, -5, 2, 1, 10, 0, -8, 6,
					-- layer=2 filter=145 channel=23
					19, 0, -43, 72, -29, -93, 26, -29, -67,
					-- layer=2 filter=145 channel=24
					23, 28, -12, 27, 17, -5, 13, -8, -13,
					-- layer=2 filter=145 channel=25
					-13, 4, 15, -4, 32, 31, -21, 11, 15,
					-- layer=2 filter=145 channel=26
					0, 7, 9, 9, -3, -8, 5, -10, 13,
					-- layer=2 filter=145 channel=27
					-52, 3, 47, -31, 24, 28, -71, 0, 33,
					-- layer=2 filter=145 channel=28
					-37, 1, -27, -59, -15, -1, -7, -7, -3,
					-- layer=2 filter=145 channel=29
					-1, 0, 8, 0, -4, 0, -7, -4, -3,
					-- layer=2 filter=145 channel=30
					10, -5, -8, 47, 6, 15, 7, -1, -29,
					-- layer=2 filter=145 channel=31
					-45, -77, -30, -23, -35, 10, 11, 13, 2,
					-- layer=2 filter=145 channel=32
					5, 11, 10, -4, -3, 7, -4, -5, -7,
					-- layer=2 filter=145 channel=33
					-19, 9, 5, 33, 31, 16, 5, -13, 10,
					-- layer=2 filter=145 channel=34
					-48, -17, -9, -8, -5, -2, 74, 11, -9,
					-- layer=2 filter=145 channel=35
					-8, -3, -8, -16, 20, 9, 4, -7, -20,
					-- layer=2 filter=145 channel=36
					-9, -7, -2, -2, -7, -4, -1, -18, 1,
					-- layer=2 filter=145 channel=37
					-32, -2, 49, -36, 12, 38, -39, 20, 44,
					-- layer=2 filter=145 channel=38
					-43, -32, 12, -25, -7, 30, -39, 2, 0,
					-- layer=2 filter=145 channel=39
					17, 24, -49, 42, -29, -64, 9, -4, -46,
					-- layer=2 filter=145 channel=40
					-24, -22, 15, 14, -9, 43, -4, 24, 23,
					-- layer=2 filter=145 channel=41
					7, 6, 0, 5, -4, 4, -7, 0, 2,
					-- layer=2 filter=145 channel=42
					11, -13, -54, 38, 9, -52, 46, 7, -40,
					-- layer=2 filter=145 channel=43
					2, -9, -34, -15, 5, 17, -35, 28, 26,
					-- layer=2 filter=145 channel=44
					1, 6, 0, 4, 7, 7, -4, 6, -8,
					-- layer=2 filter=145 channel=45
					-24, -5, -11, 53, 21, -34, 7, 51, 15,
					-- layer=2 filter=145 channel=46
					9, -11, -28, 45, 31, -1, 5, -35, -11,
					-- layer=2 filter=145 channel=47
					-35, 23, 8, 5, 12, 3, -28, -43, -22,
					-- layer=2 filter=145 channel=48
					-8, -3, -1, 1, 1, 6, 8, 11, -5,
					-- layer=2 filter=145 channel=49
					24, -33, -1, -16, -29, -5, 21, -5, 11,
					-- layer=2 filter=145 channel=50
					-14, -16, -6, -25, 0, 1, 16, 12, 17,
					-- layer=2 filter=145 channel=51
					-10, 1, 34, -30, 5, 41, -8, 0, 26,
					-- layer=2 filter=145 channel=52
					-32, -19, 31, -9, -1, 21, -25, 2, 13,
					-- layer=2 filter=145 channel=53
					37, -74, 31, -30, -26, -12, -51, -28, -34,
					-- layer=2 filter=145 channel=54
					-32, -23, 14, 4, 3, -3, 17, -6, -27,
					-- layer=2 filter=145 channel=55
					-2, -2, -3, 5, -6, 14, 5, 5, -2,
					-- layer=2 filter=145 channel=56
					-66, 16, 27, -59, 0, 42, -56, 20, 48,
					-- layer=2 filter=145 channel=57
					-1, 6, 6, -3, -3, 3, -7, -15, 7,
					-- layer=2 filter=145 channel=58
					-22, -2, -26, 28, -8, 11, 8, 41, 0,
					-- layer=2 filter=145 channel=59
					-2, -9, 9, 33, -13, 8, -9, 1, -21,
					-- layer=2 filter=145 channel=60
					-4, -26, 19, 15, 14, -15, 1, 6, 18,
					-- layer=2 filter=145 channel=61
					64, 11, 40, 33, 40, 4, -25, 0, 5,
					-- layer=2 filter=145 channel=62
					-21, -38, -1, -36, -34, -35, 23, -11, -12,
					-- layer=2 filter=145 channel=63
					47, -9, -30, 41, -11, -47, 5, -9, -42,
					-- layer=2 filter=145 channel=64
					49, -1, -37, 83, -1, -45, 32, -9, -47,
					-- layer=2 filter=145 channel=65
					53, -4, 35, -6, 4, -8, -28, 12, 0,
					-- layer=2 filter=145 channel=66
					11, -40, 0, -6, -55, -60, 13, -32, 4,
					-- layer=2 filter=145 channel=67
					4, -3, -17, 25, 27, -2, -10, 25, 2,
					-- layer=2 filter=145 channel=68
					-4, 1, 5, 0, -1, -7, 8, -4, 8,
					-- layer=2 filter=145 channel=69
					30, -14, -53, 55, 4, -83, 38, 2, -49,
					-- layer=2 filter=145 channel=70
					-16, -23, -10, -18, -8, 0, 15, -24, 1,
					-- layer=2 filter=145 channel=71
					-34, -2, 20, -49, 11, 32, -49, 4, 4,
					-- layer=2 filter=145 channel=72
					-20, -1, 21, -4, 33, 0, 23, -4, 10,
					-- layer=2 filter=145 channel=73
					1, 0, 8, 3, 18, 15, 16, 20, 1,
					-- layer=2 filter=145 channel=74
					-7, -15, -53, 48, -1, -14, -1, 17, -17,
					-- layer=2 filter=145 channel=75
					5, 33, 7, -11, 32, -9, -21, -7, 12,
					-- layer=2 filter=145 channel=76
					12, 1, 13, -30, -32, -18, 4, 14, -5,
					-- layer=2 filter=145 channel=77
					-1, -2, 1, -9, -5, 12, -9, 2, 3,
					-- layer=2 filter=145 channel=78
					-23, 1, 33, -28, -3, 31, 2, 6, 24,
					-- layer=2 filter=145 channel=79
					-9, -4, 2, 5, 0, 0, 4, -5, 7,
					-- layer=2 filter=145 channel=80
					59, 35, -56, 39, 26, -63, -12, -29, -39,
					-- layer=2 filter=145 channel=81
					-5, 9, 2, -7, 17, 7, 0, 18, 11,
					-- layer=2 filter=145 channel=82
					0, 0, -2, -5, 2, -11, 6, -1, 10,
					-- layer=2 filter=145 channel=83
					60, 15, -19, 57, -2, -13, 36, -28, -24,
					-- layer=2 filter=145 channel=84
					4, -1, -4, 9, 7, 8, -9, 11, 2,
					-- layer=2 filter=145 channel=85
					-9, -3, 0, -14, 9, 8, 0, -7, 9,
					-- layer=2 filter=145 channel=86
					-19, 0, 1, 0, -13, 4, 2, 7, 11,
					-- layer=2 filter=145 channel=87
					5, -20, 6, 33, -12, -16, 9, -19, -20,
					-- layer=2 filter=145 channel=88
					27, 3, 9, 70, -4, 0, 5, 4, -13,
					-- layer=2 filter=145 channel=89
					15, -1, -23, 1, 14, -8, 47, 14, 4,
					-- layer=2 filter=145 channel=90
					-11, 0, -1, 6, 10, -3, -1, -2, 6,
					-- layer=2 filter=145 channel=91
					-4, 6, -33, -17, 5, -8, 13, 43, 30,
					-- layer=2 filter=145 channel=92
					12, -37, 2, 0, 18, 35, 19, 22, 12,
					-- layer=2 filter=145 channel=93
					22, -29, -11, -30, -44, -90, -29, -7, -55,
					-- layer=2 filter=145 channel=94
					8, 5, -1, 9, -17, -51, -19, 1, -20,
					-- layer=2 filter=145 channel=95
					3, -7, 4, 10, -14, 4, -15, 0, 1,
					-- layer=2 filter=145 channel=96
					16, -21, -55, -6, -80, -63, 3, -22, -73,
					-- layer=2 filter=145 channel=97
					13, 0, -3, 19, 28, -25, -23, -45, -31,
					-- layer=2 filter=145 channel=98
					-27, 32, -15, 0, 23, 12, -8, 1, -12,
					-- layer=2 filter=145 channel=99
					-54, -4, 50, 17, -2, 9, -17, 13, 26,
					-- layer=2 filter=145 channel=100
					15, 14, -29, 11, -24, -15, -8, 5, -5,
					-- layer=2 filter=145 channel=101
					-58, 7, 1, -62, 25, 14, -51, 12, 0,
					-- layer=2 filter=145 channel=102
					29, -77, -46, -20, -53, -58, 47, -30, -23,
					-- layer=2 filter=145 channel=103
					41, 5, -5, -10, -2, 20, 0, -7, 30,
					-- layer=2 filter=145 channel=104
					13, 4, 10, -33, -45, 14, 13, -9, -26,
					-- layer=2 filter=145 channel=105
					-25, 39, -53, -34, 5, -65, 52, 20, 41,
					-- layer=2 filter=145 channel=106
					-15, 12, -24, -10, 22, 8, -6, 4, -12,
					-- layer=2 filter=145 channel=107
					25, -11, -39, 0, -13, 46, 48, 39, -12,
					-- layer=2 filter=145 channel=108
					-18, -10, 11, -55, 4, -4, -50, -12, -10,
					-- layer=2 filter=145 channel=109
					6, -13, 3, -5, 23, 14, 0, -1, 4,
					-- layer=2 filter=145 channel=110
					85, 6, -20, 94, 11, -38, 66, 19, -30,
					-- layer=2 filter=145 channel=111
					-8, -11, 5, -5, 0, -1, 3, -9, 2,
					-- layer=2 filter=145 channel=112
					17, 32, 26, -10, 19, 31, -23, -21, 18,
					-- layer=2 filter=145 channel=113
					31, 0, 0, 32, -6, 13, 23, -4, -35,
					-- layer=2 filter=145 channel=114
					2, -5, 0, -3, -5, -9, -3, -10, -7,
					-- layer=2 filter=145 channel=115
					9, -6, -10, 0, 3, -6, -13, -5, -2,
					-- layer=2 filter=145 channel=116
					26, -26, 18, 21, 19, -6, 31, -18, -30,
					-- layer=2 filter=145 channel=117
					-43, 3, 16, 9, 26, 3, 9, 36, -16,
					-- layer=2 filter=145 channel=118
					34, 22, -1, 0, 15, 2, -22, 11, 19,
					-- layer=2 filter=145 channel=119
					-17, 11, -25, 12, -9, -50, 4, -19, -18,
					-- layer=2 filter=145 channel=120
					0, 8, 4, -8, -8, 4, 2, 10, 2,
					-- layer=2 filter=145 channel=121
					4, 0, -1, 7, 8, -4, -12, 5, 6,
					-- layer=2 filter=145 channel=122
					3, 0, -5, 0, -1, -14, 8, -8, -2,
					-- layer=2 filter=145 channel=123
					14, 0, 0, 17, 1, -48, 11, -1, -44,
					-- layer=2 filter=145 channel=124
					5, -51, -26, 58, 12, 1, 83, 38, 26,
					-- layer=2 filter=145 channel=125
					-4, 0, 8, -2, 0, 5, -4, 4, 16,
					-- layer=2 filter=145 channel=126
					13, -19, -25, -24, -11, -2, 9, -13, 20,
					-- layer=2 filter=145 channel=127
					41, -30, -44, 45, 1, -34, 27, 0, 1,
					-- layer=2 filter=146 channel=0
					3, 4, 4, -18, -12, -17, 2, 1, 14,
					-- layer=2 filter=146 channel=1
					-35, 17, 27, -36, -32, -29, -15, -30, -16,
					-- layer=2 filter=146 channel=2
					4, 6, -11, -2, -4, 6, 5, -2, 5,
					-- layer=2 filter=146 channel=3
					-7, 33, 16, 9, 13, 4, 4, 9, 32,
					-- layer=2 filter=146 channel=4
					18, 11, -3, 5, -15, 7, -3, -16, -32,
					-- layer=2 filter=146 channel=5
					14, -7, 4, 9, -2, -12, -31, 1, -36,
					-- layer=2 filter=146 channel=6
					11, -31, 44, 34, 16, 27, 20, 1, 38,
					-- layer=2 filter=146 channel=7
					-63, 9, -15, -22, 40, 44, -16, 34, 51,
					-- layer=2 filter=146 channel=8
					-4, -1, -8, 9, 1, 3, -9, -10, 1,
					-- layer=2 filter=146 channel=9
					-10, 26, 23, -1, 2, 8, -37, -22, -38,
					-- layer=2 filter=146 channel=10
					-1, 6, 11, -4, -3, 14, 1, 15, 25,
					-- layer=2 filter=146 channel=11
					-31, -16, -25, -21, -8, -38, 11, 0, -1,
					-- layer=2 filter=146 channel=12
					-4, 34, 25, -48, -14, 6, -41, -21, 15,
					-- layer=2 filter=146 channel=13
					7, -4, -6, 6, 0, -6, 1, -4, -5,
					-- layer=2 filter=146 channel=14
					-22, 4, 28, -37, -16, -20, -35, -15, 1,
					-- layer=2 filter=146 channel=15
					19, -21, 55, -55, -28, -39, -26, -31, -40,
					-- layer=2 filter=146 channel=16
					6, -12, -19, -19, 6, 4, -27, -9, 3,
					-- layer=2 filter=146 channel=17
					-2, 1, -7, 2, -5, 0, 8, 8, -2,
					-- layer=2 filter=146 channel=18
					-29, -29, -64, -70, -79, -58, -30, -68, -106,
					-- layer=2 filter=146 channel=19
					-4, 25, -7, 13, 6, 15, -1, -6, 0,
					-- layer=2 filter=146 channel=20
					2, 7, 4, -3, 8, -9, -7, -9, 7,
					-- layer=2 filter=146 channel=21
					-6, 11, 6, 14, 10, 5, -9, 8, -4,
					-- layer=2 filter=146 channel=22
					1, 10, 3, -10, 9, -10, 7, 1, -1,
					-- layer=2 filter=146 channel=23
					-8, -11, -10, 0, 3, -12, -13, -9, 29,
					-- layer=2 filter=146 channel=24
					3, 19, -17, -8, 33, 12, 35, 40, 19,
					-- layer=2 filter=146 channel=25
					-23, -8, -30, 5, 33, 7, 17, 29, 28,
					-- layer=2 filter=146 channel=26
					10, -3, -7, -7, -1, 0, -8, -3, 10,
					-- layer=2 filter=146 channel=27
					29, 12, 31, -8, -11, 17, -4, -38, -61,
					-- layer=2 filter=146 channel=28
					-56, 3, 36, -16, -4, -1, -7, 9, 24,
					-- layer=2 filter=146 channel=29
					-9, 1, 6, 2, -6, -2, 3, -7, -7,
					-- layer=2 filter=146 channel=30
					25, -5, 22, 23, -25, -26, -15, 7, -8,
					-- layer=2 filter=146 channel=31
					-18, -35, 30, -20, -31, 23, -42, -16, -36,
					-- layer=2 filter=146 channel=32
					0, 8, 5, 7, 4, 5, 5, -9, -2,
					-- layer=2 filter=146 channel=33
					-103, 2, 54, -76, -5, 7, -28, 13, 15,
					-- layer=2 filter=146 channel=34
					-10, -11, -56, -27, -8, -25, -29, 11, -20,
					-- layer=2 filter=146 channel=35
					-63, 13, 0, -24, 6, 1, -6, 36, 16,
					-- layer=2 filter=146 channel=36
					-3, 12, -4, 1, 10, 2, 9, 3, -8,
					-- layer=2 filter=146 channel=37
					11, -21, -4, -10, -22, -3, -9, -11, -32,
					-- layer=2 filter=146 channel=38
					29, 22, 47, 28, -44, 3, 1, -20, -35,
					-- layer=2 filter=146 channel=39
					-12, -11, -13, -3, 19, 25, -34, -6, 27,
					-- layer=2 filter=146 channel=40
					77, 33, -29, -62, 16, -23, -24, 7, -42,
					-- layer=2 filter=146 channel=41
					-12, -12, 5, 6, 7, 4, -2, -5, 0,
					-- layer=2 filter=146 channel=42
					-14, 7, 15, -21, 6, -13, -22, -3, 7,
					-- layer=2 filter=146 channel=43
					25, 19, 7, 5, 5, 22, 21, 21, -44,
					-- layer=2 filter=146 channel=44
					7, -10, -1, 2, -8, 0, -2, -3, 6,
					-- layer=2 filter=146 channel=45
					-56, -8, 35, -60, -10, 0, -20, 16, 20,
					-- layer=2 filter=146 channel=46
					11, 0, 10, -6, -21, -14, -5, 15, 6,
					-- layer=2 filter=146 channel=47
					-78, -19, 15, -34, -9, 32, -2, 12, 0,
					-- layer=2 filter=146 channel=48
					0, -9, -4, 0, -6, -5, 4, 7, 6,
					-- layer=2 filter=146 channel=49
					-1, -41, -22, -15, -20, 5, -5, -76, -8,
					-- layer=2 filter=146 channel=50
					11, 17, 5, -1, 0, 5, 20, 1, 7,
					-- layer=2 filter=146 channel=51
					-6, -17, -16, 1, -4, -27, -5, 4, 7,
					-- layer=2 filter=146 channel=52
					24, -16, -21, 11, -3, -1, 48, -15, -12,
					-- layer=2 filter=146 channel=53
					-10, -5, 0, -32, 0, 20, -6, 1, -17,
					-- layer=2 filter=146 channel=54
					-82, -1, -20, -36, 3, -19, 25, 5, 46,
					-- layer=2 filter=146 channel=55
					4, 8, -5, -5, -4, -6, -1, 0, -6,
					-- layer=2 filter=146 channel=56
					13, -9, -2, -8, 0, -23, -17, -18, -38,
					-- layer=2 filter=146 channel=57
					-12, -2, 5, -9, -9, -4, -14, 0, 5,
					-- layer=2 filter=146 channel=58
					-31, 39, 24, -72, -35, 13, -18, -23, 25,
					-- layer=2 filter=146 channel=59
					47, 31, -4, -11, -5, -31, 13, -66, 0,
					-- layer=2 filter=146 channel=60
					11, -1, -16, 0, -35, -9, 4, 13, -20,
					-- layer=2 filter=146 channel=61
					7, -45, -24, -5, -42, -12, -2, -19, 4,
					-- layer=2 filter=146 channel=62
					13, -45, 5, 7, -34, -23, 7, 2, -33,
					-- layer=2 filter=146 channel=63
					38, -21, -14, -3, 12, 16, -2, -1, -15,
					-- layer=2 filter=146 channel=64
					2, -4, -24, 12, -5, 5, -19, -11, 0,
					-- layer=2 filter=146 channel=65
					36, -55, 43, 50, -12, 0, 40, 17, -1,
					-- layer=2 filter=146 channel=66
					17, 41, -22, 1, 9, 29, -4, 62, -14,
					-- layer=2 filter=146 channel=67
					48, 4, -5, 8, -14, 3, -9, -25, -62,
					-- layer=2 filter=146 channel=68
					1, 10, 3, 2, 8, -2, -2, 7, 0,
					-- layer=2 filter=146 channel=69
					-10, -24, -20, 4, 13, 0, -25, -18, 6,
					-- layer=2 filter=146 channel=70
					-56, -2, 17, -34, -24, -5, -4, 42, 43,
					-- layer=2 filter=146 channel=71
					23, -4, 28, -16, -6, 28, -10, -64, -53,
					-- layer=2 filter=146 channel=72
					-50, 8, 38, -35, -1, 11, 5, -3, -3,
					-- layer=2 filter=146 channel=73
					8, 31, 2, -41, 51, 71, -10, 42, 67,
					-- layer=2 filter=146 channel=74
					18, 12, -2, -18, -15, 7, -15, -8, 0,
					-- layer=2 filter=146 channel=75
					-63, -5, -19, -48, -28, 0, -14, 57, 51,
					-- layer=2 filter=146 channel=76
					-13, -64, -59, -60, -31, -48, -21, -72, 12,
					-- layer=2 filter=146 channel=77
					0, 0, 12, -4, 6, -2, -9, -2, -6,
					-- layer=2 filter=146 channel=78
					-9, 14, -23, 25, -7, -18, 35, 28, -1,
					-- layer=2 filter=146 channel=79
					4, -7, -7, -4, -11, 3, -3, -6, -5,
					-- layer=2 filter=146 channel=80
					16, 2, 1, 0, 19, 13, -9, 0, 2,
					-- layer=2 filter=146 channel=81
					8, 4, 0, -11, 2, -4, -9, 4, -11,
					-- layer=2 filter=146 channel=82
					-8, -2, 4, -8, 7, -10, -3, -9, 5,
					-- layer=2 filter=146 channel=83
					-3, 11, 17, 9, -16, -1, 19, 2, -8,
					-- layer=2 filter=146 channel=84
					-5, 0, -3, 8, -6, -3, -3, 3, -5,
					-- layer=2 filter=146 channel=85
					15, 11, 12, 13, -3, -9, -3, 4, -7,
					-- layer=2 filter=146 channel=86
					-18, 0, -11, -21, 0, -4, -8, -8, -13,
					-- layer=2 filter=146 channel=87
					14, -15, -15, -19, -52, -90, 30, -16, -40,
					-- layer=2 filter=146 channel=88
					40, 0, 3, 12, -27, -4, -26, -12, -18,
					-- layer=2 filter=146 channel=89
					-18, 16, 12, -34, 2, 1, -41, -3, 22,
					-- layer=2 filter=146 channel=90
					2, -1, -8, 0, -3, -7, -9, -6, 0,
					-- layer=2 filter=146 channel=91
					-16, 31, 35, -37, -1, 34, -16, -2, 11,
					-- layer=2 filter=146 channel=92
					-21, 3, 41, -61, -44, -16, -29, -20, -19,
					-- layer=2 filter=146 channel=93
					21, -41, 33, 52, -27, 38, 27, 25, -19,
					-- layer=2 filter=146 channel=94
					-9, 30, 24, -2, 22, 17, -19, -28, -52,
					-- layer=2 filter=146 channel=95
					11, -5, 10, -9, 5, -3, 8, -4, 4,
					-- layer=2 filter=146 channel=96
					19, 21, -61, 35, 47, -85, 35, 29, -17,
					-- layer=2 filter=146 channel=97
					-4, 7, 1, 20, 16, 19, 19, -5, 5,
					-- layer=2 filter=146 channel=98
					-54, -22, 1, -44, 9, 8, 13, 25, 39,
					-- layer=2 filter=146 channel=99
					18, 0, -10, 2, 2, 4, -24, 8, 2,
					-- layer=2 filter=146 channel=100
					1, 43, 28, 16, -36, -2, 0, 8, -42,
					-- layer=2 filter=146 channel=101
					0, 0, -20, -30, 10, 8, 7, -9, 3,
					-- layer=2 filter=146 channel=102
					-10, 1, -83, 0, 23, -50, 4, -37, -20,
					-- layer=2 filter=146 channel=103
					16, 10, 55, 6, -29, -2, 37, 25, 34,
					-- layer=2 filter=146 channel=104
					-44, 3, -63, -27, 16, -52, 5, -45, -81,
					-- layer=2 filter=146 channel=105
					62, 32, -63, -75, -8, 3, -20, -60, 36,
					-- layer=2 filter=146 channel=106
					-20, 3, -3, -16, -17, 3, -12, 7, 36,
					-- layer=2 filter=146 channel=107
					-4, 9, 61, -8, -4, -40, -13, 30, 38,
					-- layer=2 filter=146 channel=108
					13, 28, 24, 6, -8, -16, -44, -21, -35,
					-- layer=2 filter=146 channel=109
					5, -5, -14, -3, -2, 8, -14, -7, -3,
					-- layer=2 filter=146 channel=110
					-6, 20, -8, 12, 15, 29, -11, 20, -5,
					-- layer=2 filter=146 channel=111
					5, 3, -3, 0, -3, 2, 7, -5, 8,
					-- layer=2 filter=146 channel=112
					5, -65, -12, 12, -24, -2, -17, -4, 17,
					-- layer=2 filter=146 channel=113
					12, -27, 5, 0, -25, 18, -24, -1, -22,
					-- layer=2 filter=146 channel=114
					-14, -2, -6, 7, -23, 2, -18, -5, -2,
					-- layer=2 filter=146 channel=115
					7, -9, 9, 2, 6, 3, -7, -8, 4,
					-- layer=2 filter=146 channel=116
					43, -21, -56, -43, -28, -104, 32, -21, -62,
					-- layer=2 filter=146 channel=117
					-57, 36, 10, -38, 7, 2, 8, 53, 31,
					-- layer=2 filter=146 channel=118
					23, 18, 3, 27, 13, 19, 49, 18, -4,
					-- layer=2 filter=146 channel=119
					-10, -23, -10, 25, -29, -25, 28, -8, -46,
					-- layer=2 filter=146 channel=120
					-1, 9, 3, 1, -5, -9, 7, -10, 3,
					-- layer=2 filter=146 channel=121
					1, -5, 6, -5, -5, -1, 7, 8, 5,
					-- layer=2 filter=146 channel=122
					4, 9, 0, 4, 10, 0, -8, -6, 1,
					-- layer=2 filter=146 channel=123
					-42, -29, -7, -15, 16, 20, 3, 12, 27,
					-- layer=2 filter=146 channel=124
					-41, -40, -7, -96, -89, -14, -64, -16, -30,
					-- layer=2 filter=146 channel=125
					-4, 13, 11, 12, 10, -3, 8, 5, 0,
					-- layer=2 filter=146 channel=126
					-6, 16, -23, -38, 43, 19, -49, -16, 20,
					-- layer=2 filter=146 channel=127
					-15, -15, 14, -10, -26, -18, -14, -28, -59,
					-- layer=2 filter=147 channel=0
					-4, 38, -10, 2, 11, -13, -8, -3, -22,
					-- layer=2 filter=147 channel=1
					11, 8, -20, -6, -1, 27, 11, 7, -13,
					-- layer=2 filter=147 channel=2
					1, -4, 1, 9, -2, 1, 0, 0, 3,
					-- layer=2 filter=147 channel=3
					20, 5, 2, -10, 13, -14, -33, -17, -37,
					-- layer=2 filter=147 channel=4
					-3, 3, -15, -3, -23, -18, -14, -2, 12,
					-- layer=2 filter=147 channel=5
					-11, -8, 9, 22, 40, 5, -2, 16, -1,
					-- layer=2 filter=147 channel=6
					-19, -29, -10, -27, -22, -75, 26, 12, -22,
					-- layer=2 filter=147 channel=7
					41, 16, -33, 4, 12, 51, -35, -24, 10,
					-- layer=2 filter=147 channel=8
					-5, -6, 0, 3, -8, 0, 3, -6, 3,
					-- layer=2 filter=147 channel=9
					14, 28, -15, 35, 0, -31, 9, 0, -15,
					-- layer=2 filter=147 channel=10
					-8, -2, -10, -3, 14, -24, -19, -26, -9,
					-- layer=2 filter=147 channel=11
					-42, -8, 19, 36, 21, 20, 0, 27, 15,
					-- layer=2 filter=147 channel=12
					19, 9, -2, 3, -32, 19, 30, 13, -51,
					-- layer=2 filter=147 channel=13
					-6, -7, -7, 5, 11, 4, -11, 5, -7,
					-- layer=2 filter=147 channel=14
					14, -4, 8, 0, -6, 13, 36, 26, 9,
					-- layer=2 filter=147 channel=15
					-33, 19, 15, 27, 38, -46, -4, 10, -11,
					-- layer=2 filter=147 channel=16
					17, 15, 28, -20, 12, 36, -59, -44, 8,
					-- layer=2 filter=147 channel=17
					-7, -2, 0, -2, 4, 6, 4, -3, -6,
					-- layer=2 filter=147 channel=18
					-43, 1, 35, -16, -56, -26, 5, 30, 11,
					-- layer=2 filter=147 channel=19
					10, -35, -53, -26, -5, 10, 0, 11, 12,
					-- layer=2 filter=147 channel=20
					-6, -5, 7, -7, -5, 2, -7, 4, -2,
					-- layer=2 filter=147 channel=21
					20, 11, 0, -10, 3, 19, -6, 0, 0,
					-- layer=2 filter=147 channel=22
					-2, -8, -7, 8, 0, 3, 2, 0, -2,
					-- layer=2 filter=147 channel=23
					9, -24, 9, 2, -29, 3, 11, 1, -11,
					-- layer=2 filter=147 channel=24
					12, 14, 10, -1, 27, 40, -18, -14, -20,
					-- layer=2 filter=147 channel=25
					-31, -9, -23, -8, 13, -1, -33, -2, -3,
					-- layer=2 filter=147 channel=26
					0, 8, -1, -7, 4, 9, -1, -9, 3,
					-- layer=2 filter=147 channel=27
					-8, -13, -44, -21, 8, 22, 7, 39, 25,
					-- layer=2 filter=147 channel=28
					25, -22, -18, -11, 11, 29, 27, 8, 50,
					-- layer=2 filter=147 channel=29
					7, -8, -9, -2, -3, 2, 2, -7, -2,
					-- layer=2 filter=147 channel=30
					22, 9, 6, 10, 22, -12, 1, -30, 34,
					-- layer=2 filter=147 channel=31
					5, 28, -12, -34, 45, 14, -76, 13, 31,
					-- layer=2 filter=147 channel=32
					9, 0, 10, 4, -4, 9, 1, 11, -2,
					-- layer=2 filter=147 channel=33
					-4, -2, -21, 38, 26, -23, -61, 16, -16,
					-- layer=2 filter=147 channel=34
					-38, -29, -71, 17, 0, -29, 13, 5, 26,
					-- layer=2 filter=147 channel=35
					4, 13, -59, 14, 8, 1, -9, 13, 44,
					-- layer=2 filter=147 channel=36
					4, 3, 0, 0, 12, 20, 10, 8, -1,
					-- layer=2 filter=147 channel=37
					-29, -27, 7, -5, 18, 8, 0, 24, 22,
					-- layer=2 filter=147 channel=38
					-1, -17, -25, 17, 53, 4, -6, 42, 23,
					-- layer=2 filter=147 channel=39
					4, 1, -5, -12, 8, 42, -4, -1, -2,
					-- layer=2 filter=147 channel=40
					-60, -11, 35, 32, -31, -20, 3, -26, 6,
					-- layer=2 filter=147 channel=41
					-4, 4, -10, 4, 0, 11, -4, 7, -2,
					-- layer=2 filter=147 channel=42
					5, -13, -16, 1, 29, 27, 19, -18, -54,
					-- layer=2 filter=147 channel=43
					-1, 9, -19, -9, 5, -49, -26, -7, -27,
					-- layer=2 filter=147 channel=44
					7, -6, 1, -9, -4, 5, -9, 7, 5,
					-- layer=2 filter=147 channel=45
					-12, -54, -59, -49, -1, 0, -82, -12, -14,
					-- layer=2 filter=147 channel=46
					13, -4, -20, 17, 17, -6, -11, -3, -9,
					-- layer=2 filter=147 channel=47
					7, 24, 6, 30, 32, 29, -23, -4, 30,
					-- layer=2 filter=147 channel=48
					0, 3, -7, 3, 2, -2, 4, 0, -2,
					-- layer=2 filter=147 channel=49
					4, 37, 40, -41, 16, 1, 16, 52, 5,
					-- layer=2 filter=147 channel=50
					-26, -1, -12, 3, 0, 21, -3, -10, 3,
					-- layer=2 filter=147 channel=51
					-5, -2, -1, 2, 30, 8, 0, 26, 25,
					-- layer=2 filter=147 channel=52
					-34, 0, -41, -1, -6, 3, -12, 27, 34,
					-- layer=2 filter=147 channel=53
					22, 6, -19, -8, -16, 2, 6, -9, -28,
					-- layer=2 filter=147 channel=54
					-15, 15, -20, -5, 7, 4, -3, -18, -20,
					-- layer=2 filter=147 channel=55
					-8, -8, 7, 7, -10, 0, -1, 6, -11,
					-- layer=2 filter=147 channel=56
					-14, 5, 1, 32, 57, 33, 19, 38, 27,
					-- layer=2 filter=147 channel=57
					10, -6, 8, 0, 5, 3, 1, 3, 9,
					-- layer=2 filter=147 channel=58
					-10, -6, 0, 38, -19, 4, 55, 23, -18,
					-- layer=2 filter=147 channel=59
					-27, 11, -71, 9, 7, 15, 14, 42, 5,
					-- layer=2 filter=147 channel=60
					2, -2, -35, 14, 10, 55, 22, 5, 37,
					-- layer=2 filter=147 channel=61
					17, 35, 9, -1, 12, 49, 2, -11, 54,
					-- layer=2 filter=147 channel=62
					-56, -59, -9, -51, -56, -32, 0, 22, 0,
					-- layer=2 filter=147 channel=63
					-2, 19, 10, 12, 0, 5, -24, -11, 1,
					-- layer=2 filter=147 channel=64
					15, 19, 8, 3, 0, -6, 1, -32, -23,
					-- layer=2 filter=147 channel=65
					12, -6, 12, -2, 11, 38, 18, 0, 70,
					-- layer=2 filter=147 channel=66
					27, 9, -10, -49, -16, -8, 19, 28, 55,
					-- layer=2 filter=147 channel=67
					11, -6, -14, 27, 19, 0, -35, 4, 10,
					-- layer=2 filter=147 channel=68
					5, 0, -2, 10, -2, -1, -5, 5, -2,
					-- layer=2 filter=147 channel=69
					-1, -12, -12, -17, 0, 27, -18, -24, -10,
					-- layer=2 filter=147 channel=70
					4, -6, -20, 12, 1, -23, -4, 2, 39,
					-- layer=2 filter=147 channel=71
					10, -21, -37, 6, -32, 4, 15, 53, -4,
					-- layer=2 filter=147 channel=72
					10, -28, -1, 14, -7, 30, 0, -7, 2,
					-- layer=2 filter=147 channel=73
					34, 16, -31, 26, 42, 16, -58, -6, 7,
					-- layer=2 filter=147 channel=74
					4, -10, -9, 34, -5, -5, -11, 10, 4,
					-- layer=2 filter=147 channel=75
					15, 11, 25, -22, -54, -5, 15, 17, -15,
					-- layer=2 filter=147 channel=76
					-10, 32, -15, -36, 13, 36, -43, -50, 18,
					-- layer=2 filter=147 channel=77
					0, 9, -6, 5, 10, 10, -8, -3, -1,
					-- layer=2 filter=147 channel=78
					-45, -2, 18, 0, 19, -9, -11, 8, -15,
					-- layer=2 filter=147 channel=79
					-1, -1, -9, 5, 4, -7, -3, 3, 0,
					-- layer=2 filter=147 channel=80
					27, -11, 16, 1, 9, -1, 1, 8, 0,
					-- layer=2 filter=147 channel=81
					-7, 0, -9, -16, 6, 0, -11, -14, 5,
					-- layer=2 filter=147 channel=82
					-7, -7, 0, 0, -3, -7, 0, 3, -2,
					-- layer=2 filter=147 channel=83
					15, -1, -2, -33, -44, -30, -7, -2, -13,
					-- layer=2 filter=147 channel=84
					-2, -4, -9, 7, 8, 6, 0, 9, 1,
					-- layer=2 filter=147 channel=85
					2, -2, -2, 9, 1, 15, 8, -11, -9,
					-- layer=2 filter=147 channel=86
					-17, -19, 9, 1, -25, 0, -12, 0, -14,
					-- layer=2 filter=147 channel=87
					-73, -27, -35, -14, -53, -67, 0, 11, 32,
					-- layer=2 filter=147 channel=88
					0, 15, -14, 36, 0, -1, -2, -7, -5,
					-- layer=2 filter=147 channel=89
					-23, -13, -42, -13, -21, 21, 13, 10, -21,
					-- layer=2 filter=147 channel=90
					-7, 1, -2, 1, 2, 0, 8, -12, -1,
					-- layer=2 filter=147 channel=91
					18, -10, -37, -12, -38, 7, 19, -12, -9,
					-- layer=2 filter=147 channel=92
					4, 10, -19, -10, 0, 13, 18, 19, -12,
					-- layer=2 filter=147 channel=93
					11, -20, -56, -9, -26, 27, 7, 10, -4,
					-- layer=2 filter=147 channel=94
					4, 3, 16, -50, 5, 8, -15, -10, -41,
					-- layer=2 filter=147 channel=95
					-6, -4, 5, 2, 10, 16, 20, 8, 11,
					-- layer=2 filter=147 channel=96
					-26, -4, -72, 30, -4, 9, -4, 12, -39,
					-- layer=2 filter=147 channel=97
					15, 5, -16, 43, 15, -4, -19, -35, -59,
					-- layer=2 filter=147 channel=98
					23, -6, -3, 23, 21, 21, 12, 1, 63,
					-- layer=2 filter=147 channel=99
					-2, -47, -37, -3, 8, 46, -25, 0, 25,
					-- layer=2 filter=147 channel=100
					3, 1, -12, 30, 9, -3, 6, 7, -48,
					-- layer=2 filter=147 channel=101
					-6, -4, -6, -7, 5, -1, 0, 11, 13,
					-- layer=2 filter=147 channel=102
					-25, 9, -20, -1, -50, -1, -12, -43, 12,
					-- layer=2 filter=147 channel=103
					-16, -6, -14, 28, -1, 25, 23, -3, 17,
					-- layer=2 filter=147 channel=104
					-43, 4, 4, -14, -5, 10, 6, 56, -35,
					-- layer=2 filter=147 channel=105
					-10, -56, -44, -70, 0, -32, -35, -64, -15,
					-- layer=2 filter=147 channel=106
					-21, -25, -34, -1, 5, -4, 14, 2, -3,
					-- layer=2 filter=147 channel=107
					-28, -22, 6, -13, 64, 2, -3, -46, 18,
					-- layer=2 filter=147 channel=108
					-9, -33, -44, -40, -7, -6, -25, 11, 19,
					-- layer=2 filter=147 channel=109
					41, 8, 11, 9, 9, -23, -2, 4, -5,
					-- layer=2 filter=147 channel=110
					20, 5, 9, -4, -21, 27, 50, -47, 18,
					-- layer=2 filter=147 channel=111
					-7, -3, 0, -3, 12, 3, 2, -7, -7,
					-- layer=2 filter=147 channel=112
					31, 4, -8, -14, 42, 34, -20, -40, 11,
					-- layer=2 filter=147 channel=113
					38, 11, 37, 3, 34, 7, 22, -3, 40,
					-- layer=2 filter=147 channel=114
					2, 16, 6, 17, 10, 9, -19, 5, -5,
					-- layer=2 filter=147 channel=115
					0, 10, -7, -8, 2, -6, 1, -7, -6,
					-- layer=2 filter=147 channel=116
					-54, -25, -34, -15, -63, -66, 8, 5, 29,
					-- layer=2 filter=147 channel=117
					39, 23, -24, -30, 6, 8, -72, -10, -14,
					-- layer=2 filter=147 channel=118
					22, -4, 18, 2, 4, -42, -27, 11, -40,
					-- layer=2 filter=147 channel=119
					-39, 36, -1, -13, -3, 2, -16, 12, -7,
					-- layer=2 filter=147 channel=120
					-2, -4, -6, 0, 1, -1, 8, -5, 0,
					-- layer=2 filter=147 channel=121
					5, -3, 0, 5, -8, -11, -10, 4, 0,
					-- layer=2 filter=147 channel=122
					-5, 5, 1, -4, 2, 5, -8, -5, -16,
					-- layer=2 filter=147 channel=123
					3, -40, -6, -13, 8, 11, -60, -15, 0,
					-- layer=2 filter=147 channel=124
					0, -30, -36, -3, 33, -13, -36, 6, -86,
					-- layer=2 filter=147 channel=125
					-6, -2, 7, 2, -4, -8, 9, -3, 6,
					-- layer=2 filter=147 channel=126
					-24, 47, -30, -23, -31, -5, 15, -10, -63,
					-- layer=2 filter=147 channel=127
					-5, 15, 4, 15, 7, -14, -7, 3, -8,
					-- layer=2 filter=148 channel=0
					17, 9, 32, -8, 10, 6, 0, 6, 14,
					-- layer=2 filter=148 channel=1
					11, 20, 15, 20, 24, 12, -1, 20, -22,
					-- layer=2 filter=148 channel=2
					2, 3, -9, 12, 4, 0, 0, 5, -1,
					-- layer=2 filter=148 channel=3
					-10, 7, -14, -24, -17, -28, -20, 2, -28,
					-- layer=2 filter=148 channel=4
					5, -13, -2, -8, 5, -16, -10, 19, 16,
					-- layer=2 filter=148 channel=5
					2, -6, 6, 19, 8, 4, 9, -11, 8,
					-- layer=2 filter=148 channel=6
					28, 15, 26, 3, -8, 3, 6, 30, -12,
					-- layer=2 filter=148 channel=7
					-15, -16, 25, -22, 10, 32, 3, 21, 8,
					-- layer=2 filter=148 channel=8
					3, -10, 4, -3, -3, 11, 4, -3, 8,
					-- layer=2 filter=148 channel=9
					-7, 11, -41, 5, -28, -32, 23, 6, 6,
					-- layer=2 filter=148 channel=10
					-4, 6, -9, 10, 15, -20, 13, -8, 2,
					-- layer=2 filter=148 channel=11
					29, 17, 13, 15, 5, 5, 2, -27, -11,
					-- layer=2 filter=148 channel=12
					64, 18, 28, 27, 34, 32, 6, 11, 22,
					-- layer=2 filter=148 channel=13
					3, -6, -9, -6, 0, -10, 12, 4, -7,
					-- layer=2 filter=148 channel=14
					40, 30, 22, -7, 11, 5, -26, -11, -16,
					-- layer=2 filter=148 channel=15
					29, 6, 29, 31, -14, -27, 7, -17, -16,
					-- layer=2 filter=148 channel=16
					-28, -25, -28, -31, -31, -10, -22, -9, 0,
					-- layer=2 filter=148 channel=17
					-5, -4, -8, 6, -8, -10, 2, 6, -1,
					-- layer=2 filter=148 channel=18
					9, -47, 7, -36, -3, -32, -38, -12, -3,
					-- layer=2 filter=148 channel=19
					-29, -23, -45, 16, 25, -6, 9, -7, 5,
					-- layer=2 filter=148 channel=20
					-1, 3, 5, 1, 1, 1, 9, 1, -6,
					-- layer=2 filter=148 channel=21
					4, 9, 15, 7, 6, 10, 15, 1, -16,
					-- layer=2 filter=148 channel=22
					-2, 7, -6, 8, 0, 0, 0, 8, 2,
					-- layer=2 filter=148 channel=23
					-23, -34, 8, -34, -5, 28, -22, -18, 13,
					-- layer=2 filter=148 channel=24
					0, 70, 48, -48, -26, -3, -45, -39, -23,
					-- layer=2 filter=148 channel=25
					28, 77, 49, -39, -4, -7, -60, -39, -3,
					-- layer=2 filter=148 channel=26
					12, 5, 4, -5, 4, -3, 6, 8, -11,
					-- layer=2 filter=148 channel=27
					-8, -38, -38, 4, -9, -16, 28, 16, -13,
					-- layer=2 filter=148 channel=28
					2, -1, 1, -11, 7, 22, -50, -38, 3,
					-- layer=2 filter=148 channel=29
					-4, -9, -9, -3, -10, 3, 8, 5, -1,
					-- layer=2 filter=148 channel=30
					-23, 6, -29, 16, -8, 13, 3, 7, -14,
					-- layer=2 filter=148 channel=31
					0, 42, -1, 43, 18, -52, 14, -58, -51,
					-- layer=2 filter=148 channel=32
					-7, -5, 3, -5, 11, -4, -7, 8, 0,
					-- layer=2 filter=148 channel=33
					14, -26, -12, 0, -58, -22, -43, -14, -12,
					-- layer=2 filter=148 channel=34
					6, 38, 0, 15, -11, 37, -67, -46, 36,
					-- layer=2 filter=148 channel=35
					15, 0, -7, -19, 12, 25, -48, -40, -13,
					-- layer=2 filter=148 channel=36
					2, -16, -1, 7, -3, 8, 6, -11, -6,
					-- layer=2 filter=148 channel=37
					16, 6, -20, 21, 6, -11, 3, -2, 17,
					-- layer=2 filter=148 channel=38
					1, -17, -11, 20, -16, 3, 13, -17, -4,
					-- layer=2 filter=148 channel=39
					-14, -18, -10, 16, -1, 25, 1, 27, -7,
					-- layer=2 filter=148 channel=40
					37, 13, 26, 7, -1, -1, -24, -15, 35,
					-- layer=2 filter=148 channel=41
					3, -2, 0, -2, 8, 8, 4, -6, 6,
					-- layer=2 filter=148 channel=42
					5, -5, 3, 4, 17, 3, 10, 9, 6,
					-- layer=2 filter=148 channel=43
					-31, -28, -50, 25, -26, -49, 25, 0, 3,
					-- layer=2 filter=148 channel=44
					1, -1, 0, -1, 8, -5, 3, -7, 11,
					-- layer=2 filter=148 channel=45
					-24, -18, -21, -50, -47, -53, 5, 9, 4,
					-- layer=2 filter=148 channel=46
					8, 12, 14, 27, -5, -32, 35, 8, 16,
					-- layer=2 filter=148 channel=47
					10, 15, 24, -28, -11, 29, -36, 16, 18,
					-- layer=2 filter=148 channel=48
					-4, 1, -10, -10, 1, 8, -5, 4, -11,
					-- layer=2 filter=148 channel=49
					-7, -6, 24, -5, -8, -17, -3, 11, 11,
					-- layer=2 filter=148 channel=50
					-7, -20, -16, 4, -1, -11, -5, 15, -10,
					-- layer=2 filter=148 channel=51
					17, 29, 13, -2, 7, -4, 0, -6, -6,
					-- layer=2 filter=148 channel=52
					-9, 16, -16, 33, 2, 25, 20, 16, 13,
					-- layer=2 filter=148 channel=53
					-64, -14, 21, 34, -5, -21, -59, -68, -11,
					-- layer=2 filter=148 channel=54
					59, 54, 33, -9, 14, 29, -19, 10, 19,
					-- layer=2 filter=148 channel=55
					-1, -7, 6, -1, 11, 1, -6, -6, -2,
					-- layer=2 filter=148 channel=56
					38, -10, -8, 7, -11, -14, 4, -16, 0,
					-- layer=2 filter=148 channel=57
					-2, 1, -5, 4, -9, -8, -3, 1, 4,
					-- layer=2 filter=148 channel=58
					50, 41, -18, 40, 37, 36, 16, 4, 36,
					-- layer=2 filter=148 channel=59
					1, 16, -25, -15, 19, 4, 19, -17, -20,
					-- layer=2 filter=148 channel=60
					24, 23, 22, 25, 26, -5, -13, -35, 0,
					-- layer=2 filter=148 channel=61
					-38, -12, 2, -57, -28, -13, -48, -33, -71,
					-- layer=2 filter=148 channel=62
					22, 17, 33, 16, 6, -15, 4, 22, 10,
					-- layer=2 filter=148 channel=63
					6, -4, 25, -17, -13, 7, -28, -4, -4,
					-- layer=2 filter=148 channel=64
					-36, -6, 6, -19, 4, 19, -23, 16, 1,
					-- layer=2 filter=148 channel=65
					-8, -23, 18, 10, 2, -20, -21, 7, -20,
					-- layer=2 filter=148 channel=66
					55, -11, -6, -9, -5, -28, 7, 16, 28,
					-- layer=2 filter=148 channel=67
					7, -6, -8, 5, -14, -53, 22, 6, 4,
					-- layer=2 filter=148 channel=68
					-1, 8, -1, -2, -7, -11, -9, 10, -1,
					-- layer=2 filter=148 channel=69
					-16, 0, -7, -6, -5, -9, 4, 14, -2,
					-- layer=2 filter=148 channel=70
					39, -15, -23, -4, -1, 26, -21, 9, 32,
					-- layer=2 filter=148 channel=71
					11, -2, -28, -4, 1, 0, 18, -2, -54,
					-- layer=2 filter=148 channel=72
					59, 6, 22, 13, 12, 67, -5, 8, 19,
					-- layer=2 filter=148 channel=73
					-18, 27, 27, 50, 33, -49, 38, -29, -20,
					-- layer=2 filter=148 channel=74
					11, 11, 12, -3, 8, -30, 30, 8, 15,
					-- layer=2 filter=148 channel=75
					-3, 11, -4, 25, 48, -2, -17, -15, 8,
					-- layer=2 filter=148 channel=76
					-45, -27, -4, -2, -20, -62, -11, -49, 18,
					-- layer=2 filter=148 channel=77
					-5, 0, 5, 5, 1, -8, -9, 5, -1,
					-- layer=2 filter=148 channel=78
					14, 27, 48, -20, -5, -9, -12, -3, 2,
					-- layer=2 filter=148 channel=79
					10, -9, -2, 6, 3, -5, -3, -2, 1,
					-- layer=2 filter=148 channel=80
					4, -3, 8, 9, -17, -27, 23, 28, 17,
					-- layer=2 filter=148 channel=81
					3, 15, 11, -12, 7, 13, 12, 2, 11,
					-- layer=2 filter=148 channel=82
					-7, 3, -4, -3, -8, 0, 0, 0, 0,
					-- layer=2 filter=148 channel=83
					-2, -6, -4, -15, 4, 15, -10, 18, 2,
					-- layer=2 filter=148 channel=84
					-3, -5, 2, 5, 0, 0, 6, 0, 7,
					-- layer=2 filter=148 channel=85
					1, 9, -13, 2, 0, -4, 1, 0, 15,
					-- layer=2 filter=148 channel=86
					2, -9, 16, 0, -5, 4, -13, -18, -5,
					-- layer=2 filter=148 channel=87
					38, -6, 47, 23, -22, -67, -10, -18, -18,
					-- layer=2 filter=148 channel=88
					-7, 1, 4, 7, 0, 0, -1, 2, -3,
					-- layer=2 filter=148 channel=89
					21, 31, -14, 2, 15, 23, -28, -8, 6,
					-- layer=2 filter=148 channel=90
					-1, 4, 0, -2, 5, -2, -8, 4, -7,
					-- layer=2 filter=148 channel=91
					37, 17, 4, 23, 12, 36, -25, 0, 32,
					-- layer=2 filter=148 channel=92
					19, 18, 16, 35, 13, 21, -6, 33, 11,
					-- layer=2 filter=148 channel=93
					15, 44, -39, 8, -7, -42, -14, 32, 18,
					-- layer=2 filter=148 channel=94
					-53, -24, 15, -9, -18, -4, -32, -3, -25,
					-- layer=2 filter=148 channel=95
					-2, 4, 18, 0, 8, 15, 1, 13, 11,
					-- layer=2 filter=148 channel=96
					20, 9, -32, -9, 27, 24, 0, -5, 17,
					-- layer=2 filter=148 channel=97
					12, 18, -3, 20, 0, -24, -17, -24, 20,
					-- layer=2 filter=148 channel=98
					43, -18, 23, -25, -18, 43, -31, 2, 24,
					-- layer=2 filter=148 channel=99
					-2, 16, 14, 29, -12, -5, -7, -14, -21,
					-- layer=2 filter=148 channel=100
					0, -4, 31, 42, 11, 4, 11, 7, 4,
					-- layer=2 filter=148 channel=101
					19, 58, 27, -12, 1, 16, -18, -15, -27,
					-- layer=2 filter=148 channel=102
					1, -14, -30, -38, 24, -6, -13, -15, -42,
					-- layer=2 filter=148 channel=103
					-61, -51, -22, 17, -57, -79, 17, 11, -13,
					-- layer=2 filter=148 channel=104
					6, -61, 23, -19, -9, -3, -7, -6, 29,
					-- layer=2 filter=148 channel=105
					-33, -5, -23, -9, -54, -90, 0, -9, -28,
					-- layer=2 filter=148 channel=106
					8, 36, 11, -32, -6, -14, -32, -48, -6,
					-- layer=2 filter=148 channel=107
					-9, -4, 9, -31, 24, -18, 0, -4, -11,
					-- layer=2 filter=148 channel=108
					-43, 13, -27, 10, 24, 12, 41, 6, -16,
					-- layer=2 filter=148 channel=109
					3, 5, -16, 0, -10, -8, 2, 7, -14,
					-- layer=2 filter=148 channel=110
					5, -12, 18, -52, 5, 11, -19, 10, 14,
					-- layer=2 filter=148 channel=111
					-1, 8, 3, -5, 2, -3, -6, -6, 3,
					-- layer=2 filter=148 channel=112
					1, 4, 11, -7, 14, -8, -6, -22, -18,
					-- layer=2 filter=148 channel=113
					21, -17, 5, 15, -7, 1, -25, -17, -1,
					-- layer=2 filter=148 channel=114
					11, 5, 13, 22, 19, 1, 12, 15, 8,
					-- layer=2 filter=148 channel=115
					-3, 7, -2, 7, 5, 8, 4, -5, 1,
					-- layer=2 filter=148 channel=116
					28, -34, 8, 14, -4, -47, 6, -9, -13,
					-- layer=2 filter=148 channel=117
					-16, 0, 33, 1, -49, -19, 3, -31, -10,
					-- layer=2 filter=148 channel=118
					-4, -21, 2, 8, -3, -18, 34, 43, 30,
					-- layer=2 filter=148 channel=119
					-12, -3, 7, -19, 8, -8, -4, -14, -15,
					-- layer=2 filter=148 channel=120
					3, 6, 6, -7, 7, 7, -5, 0, -1,
					-- layer=2 filter=148 channel=121
					9, -2, -6, 5, -3, -8, 0, 2, -7,
					-- layer=2 filter=148 channel=122
					-12, 2, -4, -11, -2, 17, -16, -7, -3,
					-- layer=2 filter=148 channel=123
					13, -27, 5, -24, -19, 59, 0, 9, 46,
					-- layer=2 filter=148 channel=124
					-23, 7, -36, 0, -41, -67, 2, 1, -5,
					-- layer=2 filter=148 channel=125
					-4, 5, -5, -4, -6, -5, 7, 4, 7,
					-- layer=2 filter=148 channel=126
					-25, 23, 8, -23, -64, -8, -39, -60, -80,
					-- layer=2 filter=148 channel=127
					4, 40, 11, 35, 20, 5, -12, -10, 0,
					-- layer=2 filter=149 channel=0
					-3, -6, -4, 5, -6, -13, 2, -9, 6,
					-- layer=2 filter=149 channel=1
					14, -18, 1, -4, -4, -13, -17, -19, -8,
					-- layer=2 filter=149 channel=2
					-1, 0, 9, -6, 0, 6, -4, -6, 10,
					-- layer=2 filter=149 channel=3
					-13, -4, -7, -4, -13, 0, -7, -4, -8,
					-- layer=2 filter=149 channel=4
					-12, -12, 1, 13, 5, -5, 5, -13, -5,
					-- layer=2 filter=149 channel=5
					-10, 5, 2, -1, -13, -11, 7, 11, 0,
					-- layer=2 filter=149 channel=6
					11, 18, 11, -5, -7, -11, -5, -9, -7,
					-- layer=2 filter=149 channel=7
					-8, -21, -7, 10, 17, -1, 1, -16, -17,
					-- layer=2 filter=149 channel=8
					-6, 5, 3, 11, -8, -10, -5, 2, 0,
					-- layer=2 filter=149 channel=9
					-17, 3, -15, -2, 2, -3, -4, -8, 0,
					-- layer=2 filter=149 channel=10
					-4, -3, -5, -13, -9, 0, 5, -6, -9,
					-- layer=2 filter=149 channel=11
					-3, -9, 0, 2, 3, -11, 5, 3, 0,
					-- layer=2 filter=149 channel=12
					-11, 0, -6, -8, 0, 2, 4, -4, -9,
					-- layer=2 filter=149 channel=13
					5, 11, 8, -7, 3, 6, 1, 6, 3,
					-- layer=2 filter=149 channel=14
					3, -7, -10, -17, 5, 0, -7, -6, -13,
					-- layer=2 filter=149 channel=15
					1, -5, -11, -27, -13, -5, -7, -8, -8,
					-- layer=2 filter=149 channel=16
					-4, 10, -5, -10, 10, -9, -8, -5, -9,
					-- layer=2 filter=149 channel=17
					2, 0, 6, -7, -6, 0, -6, 3, -1,
					-- layer=2 filter=149 channel=18
					8, -5, -10, 0, -22, -4, -20, -9, -10,
					-- layer=2 filter=149 channel=19
					1, -5, 4, 3, -5, -8, -6, -11, 0,
					-- layer=2 filter=149 channel=20
					0, 5, 3, 10, -8, 1, -7, 7, 0,
					-- layer=2 filter=149 channel=21
					0, 5, -8, -4, -10, -7, 8, 8, -6,
					-- layer=2 filter=149 channel=22
					-8, 7, 2, -5, -2, 1, -1, -6, 3,
					-- layer=2 filter=149 channel=23
					7, -4, -5, 0, -2, -4, -16, -10, -13,
					-- layer=2 filter=149 channel=24
					-4, -4, -16, -11, 1, -12, 4, -3, 0,
					-- layer=2 filter=149 channel=25
					-15, 0, -5, -16, -14, -9, 7, -7, -2,
					-- layer=2 filter=149 channel=26
					-5, 0, -8, -10, 10, -3, -7, 0, -6,
					-- layer=2 filter=149 channel=27
					-22, -28, -28, -12, -5, -18, -11, -6, -12,
					-- layer=2 filter=149 channel=28
					-19, -1, -12, 1, -15, -24, -7, -8, 0,
					-- layer=2 filter=149 channel=29
					-10, -5, 6, -4, -3, 3, 6, -7, 5,
					-- layer=2 filter=149 channel=30
					12, 5, 5, 0, -11, 4, 7, -1, -10,
					-- layer=2 filter=149 channel=31
					6, 0, -8, -2, -5, -5, 0, 4, -12,
					-- layer=2 filter=149 channel=32
					-2, -9, 3, 6, 1, -4, 2, -8, 0,
					-- layer=2 filter=149 channel=33
					-11, -10, 0, -2, 12, 0, 3, 6, -7,
					-- layer=2 filter=149 channel=34
					20, -15, 7, -17, -10, -9, -22, 4, -23,
					-- layer=2 filter=149 channel=35
					9, -7, -16, -2, -5, -23, 0, -1, 9,
					-- layer=2 filter=149 channel=36
					6, -5, -3, 6, -5, -11, -7, -10, 0,
					-- layer=2 filter=149 channel=37
					0, -8, -6, 0, -5, -11, -8, -3, 1,
					-- layer=2 filter=149 channel=38
					-11, -8, -1, -1, -4, -14, -8, -1, -12,
					-- layer=2 filter=149 channel=39
					-8, -10, -7, -17, 16, 5, -9, 5, -4,
					-- layer=2 filter=149 channel=40
					-12, -9, 6, -7, -14, -6, 1, 8, -4,
					-- layer=2 filter=149 channel=41
					0, -1, 2, -6, -4, -6, 2, 3, 11,
					-- layer=2 filter=149 channel=42
					-1, 6, -16, -9, -6, -6, -14, -15, -15,
					-- layer=2 filter=149 channel=43
					-7, 3, -6, 3, 2, -12, -9, -2, 4,
					-- layer=2 filter=149 channel=44
					10, -9, 6, -6, 1, -7, -7, 0, -11,
					-- layer=2 filter=149 channel=45
					-12, -4, -12, 9, 16, -2, 10, 6, -5,
					-- layer=2 filter=149 channel=46
					4, -9, 6, 3, -5, -2, -8, -4, -6,
					-- layer=2 filter=149 channel=47
					-11, -14, -14, 3, -11, -14, -12, -7, -10,
					-- layer=2 filter=149 channel=48
					9, -3, -2, 0, -3, 8, 4, -8, -5,
					-- layer=2 filter=149 channel=49
					11, -7, -30, -12, -17, -9, -28, -14, -9,
					-- layer=2 filter=149 channel=50
					10, 1, 1, 9, 9, 0, -2, -2, 0,
					-- layer=2 filter=149 channel=51
					-12, -4, 1, -5, -12, -17, -6, -4, -1,
					-- layer=2 filter=149 channel=52
					-2, -11, -9, 2, -14, -1, -6, 0, -12,
					-- layer=2 filter=149 channel=53
					-2, 0, -5, -10, -7, -8, 3, 7, 13,
					-- layer=2 filter=149 channel=54
					13, 11, -7, 9, 15, 0, -4, -6, -3,
					-- layer=2 filter=149 channel=55
					-10, -7, 2, -6, -3, -6, 1, 8, -6,
					-- layer=2 filter=149 channel=56
					-11, -5, -1, 5, 7, -7, 7, 1, -3,
					-- layer=2 filter=149 channel=57
					-9, 1, -10, -9, 2, -1, 4, 0, -8,
					-- layer=2 filter=149 channel=58
					-12, -11, -7, -19, 8, -17, 12, 7, 12,
					-- layer=2 filter=149 channel=59
					1, -18, -3, -6, 9, 6, -11, 0, -3,
					-- layer=2 filter=149 channel=60
					-16, -24, 21, -16, -6, -8, -17, -13, -20,
					-- layer=2 filter=149 channel=61
					-13, -2, -3, -24, -15, -5, -9, -5, -6,
					-- layer=2 filter=149 channel=62
					6, 1, 7, -15, -24, -21, -15, 1, -12,
					-- layer=2 filter=149 channel=63
					-4, 1, -2, 0, 0, -12, 5, 0, 2,
					-- layer=2 filter=149 channel=64
					2, 8, -6, -3, -5, 3, 3, 2, 1,
					-- layer=2 filter=149 channel=65
					-8, 12, 10, -6, -5, 5, -8, -10, -11,
					-- layer=2 filter=149 channel=66
					-13, -10, 6, -5, 0, 9, 0, -14, -5,
					-- layer=2 filter=149 channel=67
					0, 0, -6, 3, 4, -13, -6, -9, -10,
					-- layer=2 filter=149 channel=68
					-7, -5, -7, 5, 7, -8, -2, -8, 3,
					-- layer=2 filter=149 channel=69
					12, -8, -5, 0, 1, -12, 0, -12, -1,
					-- layer=2 filter=149 channel=70
					-3, 5, -14, 0, -3, 6, 1, 8, 3,
					-- layer=2 filter=149 channel=71
					-15, -6, -13, 5, 2, -4, 3, -15, 3,
					-- layer=2 filter=149 channel=72
					-8, -18, -15, 4, -1, -4, 0, -21, -26,
					-- layer=2 filter=149 channel=73
					0, -20, -6, 0, -25, -12, 0, -4, 4,
					-- layer=2 filter=149 channel=74
					-9, -2, -16, -4, -9, -7, 1, -1, -8,
					-- layer=2 filter=149 channel=75
					-22, -1, -1, -3, -3, 2, -9, -10, -13,
					-- layer=2 filter=149 channel=76
					0, -7, -1, -17, -20, 2, -9, 3, -9,
					-- layer=2 filter=149 channel=77
					-2, 4, 2, 1, -5, -3, 0, 0, 0,
					-- layer=2 filter=149 channel=78
					7, -4, -4, 0, -4, 1, -5, 0, -1,
					-- layer=2 filter=149 channel=79
					7, 9, -6, 0, -1, -12, 1, 7, -2,
					-- layer=2 filter=149 channel=80
					-8, 0, -3, 2, -10, 2, -2, -2, 0,
					-- layer=2 filter=149 channel=81
					-10, -9, 1, -5, 4, -8, 8, 2, -9,
					-- layer=2 filter=149 channel=82
					-10, 6, 12, -8, -2, 6, -2, 3, 7,
					-- layer=2 filter=149 channel=83
					-21, -2, 1, -11, -16, -13, -17, -12, -4,
					-- layer=2 filter=149 channel=84
					4, -5, 10, 3, 3, 5, 9, 8, -7,
					-- layer=2 filter=149 channel=85
					-7, 11, -7, -10, -7, 0, 8, 0, 5,
					-- layer=2 filter=149 channel=86
					8, 11, 0, 2, -11, 0, 6, -10, -2,
					-- layer=2 filter=149 channel=87
					-11, -6, -18, -10, -18, -9, -21, -23, -22,
					-- layer=2 filter=149 channel=88
					-7, 1, 2, -4, 0, -1, -4, -8, -5,
					-- layer=2 filter=149 channel=89
					-9, -7, -7, -18, -4, -12, -7, -13, -16,
					-- layer=2 filter=149 channel=90
					9, -8, -7, 8, -8, 0, -6, 0, -8,
					-- layer=2 filter=149 channel=91
					-20, -21, -12, -8, -9, -30, -10, -13, -21,
					-- layer=2 filter=149 channel=92
					9, -2, -7, 0, 6, -15, -2, -7, -3,
					-- layer=2 filter=149 channel=93
					7, 4, 28, -9, -4, 17, -2, -1, -7,
					-- layer=2 filter=149 channel=94
					-12, 9, -5, 0, -16, -2, -11, -11, 2,
					-- layer=2 filter=149 channel=95
					3, 7, -5, -10, 0, 7, -7, 10, -5,
					-- layer=2 filter=149 channel=96
					-34, -21, -23, 0, -23, -9, -26, -2, 1,
					-- layer=2 filter=149 channel=97
					-16, -4, 4, -5, 0, 0, -11, -9, -10,
					-- layer=2 filter=149 channel=98
					-25, 0, -22, 1, -17, -2, -25, -2, 0,
					-- layer=2 filter=149 channel=99
					-11, -18, -10, -12, -17, 2, -2, 0, -11,
					-- layer=2 filter=149 channel=100
					-28, -24, -14, 1, -11, -11, -9, -8, -3,
					-- layer=2 filter=149 channel=101
					-14, 0, -12, 5, -8, -15, 8, 15, 5,
					-- layer=2 filter=149 channel=102
					3, -15, -20, -2, -4, 2, -5, -15, 8,
					-- layer=2 filter=149 channel=103
					-4, -8, 9, 11, 0, 0, 6, 7, 1,
					-- layer=2 filter=149 channel=104
					-8, -12, -16, -15, -3, -6, -7, -12, -3,
					-- layer=2 filter=149 channel=105
					-19, -17, 4, -5, -16, -12, 6, 5, 3,
					-- layer=2 filter=149 channel=106
					-15, -11, -5, -8, -13, -11, 12, -9, -8,
					-- layer=2 filter=149 channel=107
					-3, 3, -9, 1, -13, -19, 9, -4, 1,
					-- layer=2 filter=149 channel=108
					-13, -1, -1, -1, -6, 0, -8, 2, 0,
					-- layer=2 filter=149 channel=109
					-6, -8, -8, -6, 10, -7, -5, -6, 0,
					-- layer=2 filter=149 channel=110
					5, -4, 8, -19, -1, 11, -4, -2, -10,
					-- layer=2 filter=149 channel=111
					-4, 4, 8, -4, -3, 1, -8, 10, -3,
					-- layer=2 filter=149 channel=112
					-2, -9, -10, 6, -2, -1, -11, -10, -8,
					-- layer=2 filter=149 channel=113
					7, -3, 3, -6, -6, 5, -15, 2, -3,
					-- layer=2 filter=149 channel=114
					10, 11, -10, -4, 0, 5, 4, -9, 0,
					-- layer=2 filter=149 channel=115
					4, 7, -3, 1, 5, 0, 0, -8, -6,
					-- layer=2 filter=149 channel=116
					9, -5, -11, -10, -21, -21, -16, -8, 0,
					-- layer=2 filter=149 channel=117
					8, -16, -17, 16, 15, 10, -10, -5, -3,
					-- layer=2 filter=149 channel=118
					0, 0, -9, 2, -17, -18, -7, 1, -15,
					-- layer=2 filter=149 channel=119
					14, -9, -10, 9, -3, -7, -13, -1, -14,
					-- layer=2 filter=149 channel=120
					7, -1, 0, -10, -9, -2, -8, -1, 6,
					-- layer=2 filter=149 channel=121
					7, -6, 7, 7, 0, 12, -8, 4, 0,
					-- layer=2 filter=149 channel=122
					-10, 8, 0, -2, -4, -5, -8, -8, 9,
					-- layer=2 filter=149 channel=123
					-9, -1, 4, 6, 4, -4, -9, -18, -20,
					-- layer=2 filter=149 channel=124
					5, -21, -18, -1, 27, 1, -3, -24, -7,
					-- layer=2 filter=149 channel=125
					1, -3, -8, -8, 8, 1, -5, 0, -4,
					-- layer=2 filter=149 channel=126
					-5, 3, -7, -4, 7, -5, 4, 3, -4,
					-- layer=2 filter=149 channel=127
					4, -16, -1, 0, -11, -3, -7, -3, -6,
					-- layer=2 filter=150 channel=0
					-22, -6, -21, -16, 0, 23, -8, 10, 13,
					-- layer=2 filter=150 channel=1
					5, -21, 0, -25, 2, -1, -27, -25, 12,
					-- layer=2 filter=150 channel=2
					-2, 6, 5, 0, 8, 3, 0, -4, -6,
					-- layer=2 filter=150 channel=3
					9, 16, 0, 0, 25, -4, 13, 11, 34,
					-- layer=2 filter=150 channel=4
					9, -100, -35, -89, -57, -32, 1, -47, -20,
					-- layer=2 filter=150 channel=5
					9, 20, 20, 15, 22, -3, -21, -29, -5,
					-- layer=2 filter=150 channel=6
					24, 25, -17, 52, 21, -22, 30, -17, 8,
					-- layer=2 filter=150 channel=7
					2, 10, -51, -89, -30, 27, -24, 37, 57,
					-- layer=2 filter=150 channel=8
					3, 7, 6, -2, 0, 6, 3, -1, -11,
					-- layer=2 filter=150 channel=9
					39, 54, 52, -25, 4, -7, -32, -25, -24,
					-- layer=2 filter=150 channel=10
					-27, -17, -5, -17, -8, -19, 4, -1, 1,
					-- layer=2 filter=150 channel=11
					12, 4, 2, 5, 0, 1, -20, -20, -1,
					-- layer=2 filter=150 channel=12
					7, -4, -8, -20, -18, 6, -39, -12, 45,
					-- layer=2 filter=150 channel=13
					2, -9, -8, -10, 6, 12, 8, 3, 2,
					-- layer=2 filter=150 channel=14
					45, 16, -4, -15, -14, -19, -62, -33, -28,
					-- layer=2 filter=150 channel=15
					20, 15, 25, -3, -3, 36, 1, 45, 50,
					-- layer=2 filter=150 channel=16
					5, 23, -20, -23, -42, 20, -16, -6, -13,
					-- layer=2 filter=150 channel=17
					-9, 5, -2, 2, 8, -6, -1, 9, -8,
					-- layer=2 filter=150 channel=18
					41, -3, -15, -31, -12, 0, 22, 3, 13,
					-- layer=2 filter=150 channel=19
					-24, -22, -36, 14, 20, 25, 25, 3, 17,
					-- layer=2 filter=150 channel=20
					0, 1, -10, -3, -1, -4, 10, -9, -5,
					-- layer=2 filter=150 channel=21
					8, 6, -7, -9, -8, -5, -7, 10, 14,
					-- layer=2 filter=150 channel=22
					4, 1, -7, -8, 0, -4, -7, -7, -2,
					-- layer=2 filter=150 channel=23
					-51, -4, -16, -50, -26, -9, 40, -10, 1,
					-- layer=2 filter=150 channel=24
					26, 34, 14, 0, -12, 13, -20, -11, 8,
					-- layer=2 filter=150 channel=25
					20, 17, 17, -3, -3, -10, -12, -14, 19,
					-- layer=2 filter=150 channel=26
					-12, 5, -5, 1, 5, 2, 10, -5, -6,
					-- layer=2 filter=150 channel=27
					14, 6, 25, -8, 21, 35, -55, -45, -38,
					-- layer=2 filter=150 channel=28
					-62, -30, 0, -65, -49, -34, -7, -7, 11,
					-- layer=2 filter=150 channel=29
					-6, 6, -5, -7, 0, 6, -2, 1, 0,
					-- layer=2 filter=150 channel=30
					12, -36, -22, -17, -10, -24, -2, -19, 19,
					-- layer=2 filter=150 channel=31
					-29, -83, -21, -63, -44, 33, -40, 3, 31,
					-- layer=2 filter=150 channel=32
					-5, 7, -6, 5, -6, -1, 2, -3, -3,
					-- layer=2 filter=150 channel=33
					28, 43, 7, -108, -32, -39, -66, -3, 35,
					-- layer=2 filter=150 channel=34
					-30, 3, -19, -27, 1, 11, -81, 47, 9,
					-- layer=2 filter=150 channel=35
					-51, -73, -75, -115, -80, -35, -52, 4, 41,
					-- layer=2 filter=150 channel=36
					5, 4, -9, 4, -1, -1, 0, -1, -15,
					-- layer=2 filter=150 channel=37
					8, 22, 21, 21, 9, 12, -7, -18, -8,
					-- layer=2 filter=150 channel=38
					47, 27, 22, 4, -5, -1, -55, -71, -39,
					-- layer=2 filter=150 channel=39
					19, -18, -44, -59, -10, -22, 2, -40, -21,
					-- layer=2 filter=150 channel=40
					41, 18, -19, -58, -4, -1, -35, 56, 51,
					-- layer=2 filter=150 channel=41
					4, -1, -7, -4, 2, -9, 9, 5, -9,
					-- layer=2 filter=150 channel=42
					-1, -5, -3, 2, -24, -13, 58, 27, 46,
					-- layer=2 filter=150 channel=43
					-10, -28, 1, -29, 18, -21, -30, -25, 15,
					-- layer=2 filter=150 channel=44
					3, -7, 1, 0, -6, -5, 4, -6, 6,
					-- layer=2 filter=150 channel=45
					1, 0, 37, -25, -14, 28, -77, 5, 54,
					-- layer=2 filter=150 channel=46
					-2, -55, -24, -7, 15, -18, -58, 10, -34,
					-- layer=2 filter=150 channel=47
					-34, -18, 23, -69, -10, -29, -13, 12, 8,
					-- layer=2 filter=150 channel=48
					9, 1, -5, -1, -7, -1, 0, 2, -1,
					-- layer=2 filter=150 channel=49
					13, -52, -15, -2, -5, 32, 6, 11, 5,
					-- layer=2 filter=150 channel=50
					2, 28, 7, 14, -3, 23, 10, -8, 6,
					-- layer=2 filter=150 channel=51
					24, 6, 6, 12, -11, -8, -5, -9, 10,
					-- layer=2 filter=150 channel=52
					-34, -28, -21, -48, 3, -22, 0, 10, 3,
					-- layer=2 filter=150 channel=53
					10, -26, -14, 50, 29, 38, 38, -16, 45,
					-- layer=2 filter=150 channel=54
					-31, -60, -73, -40, -37, -18, -31, 34, 45,
					-- layer=2 filter=150 channel=55
					6, -2, 0, -6, 2, 2, 6, 0, -9,
					-- layer=2 filter=150 channel=56
					14, 6, 23, 27, -12, 1, -25, -15, 4,
					-- layer=2 filter=150 channel=57
					11, -5, 11, 11, -1, -9, 4, -5, -8,
					-- layer=2 filter=150 channel=58
					20, -8, -6, -2, 19, 3, -41, -26, 80,
					-- layer=2 filter=150 channel=59
					31, 0, -33, -21, 34, 12, -1, -3, 14,
					-- layer=2 filter=150 channel=60
					9, -2, -24, 36, 10, 16, 27, -16, -30,
					-- layer=2 filter=150 channel=61
					-17, -24, -36, 23, -22, 27, 35, -9, -7,
					-- layer=2 filter=150 channel=62
					26, -31, -48, 38, -20, 12, 9, -10, 13,
					-- layer=2 filter=150 channel=63
					11, -15, -31, -35, -18, -22, 15, 14, -10,
					-- layer=2 filter=150 channel=64
					-8, -12, -30, -23, -6, -5, 18, -17, 2,
					-- layer=2 filter=150 channel=65
					4, 5, 21, 29, -41, -8, 23, -46, -28,
					-- layer=2 filter=150 channel=66
					20, 18, -38, 49, 19, 49, -5, -22, 16,
					-- layer=2 filter=150 channel=67
					29, -24, 3, 0, -11, -7, -23, -42, -34,
					-- layer=2 filter=150 channel=68
					9, -7, 6, 8, -7, 7, 1, 11, -9,
					-- layer=2 filter=150 channel=69
					13, -1, -8, -41, -19, -17, 31, -35, -10,
					-- layer=2 filter=150 channel=70
					-78, -42, -47, -72, -54, -27, -72, 10, 36,
					-- layer=2 filter=150 channel=71
					28, -5, 13, 1, 16, 50, -57, -30, -40,
					-- layer=2 filter=150 channel=72
					36, 68, 27, -23, 2, -17, 18, 31, 2,
					-- layer=2 filter=150 channel=73
					-46, -48, -18, 5, 12, -14, 7, 1, 40,
					-- layer=2 filter=150 channel=74
					16, -29, -60, -30, -52, -29, -11, 8, -13,
					-- layer=2 filter=150 channel=75
					6, -6, -11, -1, 8, -9, -105, 18, 27,
					-- layer=2 filter=150 channel=76
					-37, -35, -12, 19, 7, 19, 59, -19, 57,
					-- layer=2 filter=150 channel=77
					-6, 6, 6, 6, -8, -3, 6, 0, 3,
					-- layer=2 filter=150 channel=78
					27, 19, 3, 7, 0, 2, -4, 2, 14,
					-- layer=2 filter=150 channel=79
					3, 11, 11, 9, -4, 0, 0, -1, 5,
					-- layer=2 filter=150 channel=80
					-103, -61, -62, -63, -18, -53, 11, -29, -15,
					-- layer=2 filter=150 channel=81
					5, -4, 1, -7, 8, -10, 6, 3, -2,
					-- layer=2 filter=150 channel=82
					0, 2, -5, -6, 8, -4, -9, -3, 2,
					-- layer=2 filter=150 channel=83
					-23, -19, 14, -22, -25, 19, 10, 7, 0,
					-- layer=2 filter=150 channel=84
					-8, 2, -3, -1, 7, -3, 11, 6, -3,
					-- layer=2 filter=150 channel=85
					-4, 0, 5, -14, 7, -6, -17, 10, 0,
					-- layer=2 filter=150 channel=86
					0, 10, -4, 10, -11, 0, 0, 8, 0,
					-- layer=2 filter=150 channel=87
					30, -19, 11, 16, -14, -23, -23, 8, 4,
					-- layer=2 filter=150 channel=88
					8, -1, 0, -29, -73, -67, -10, -8, 12,
					-- layer=2 filter=150 channel=89
					13, 22, -14, 3, 12, 2, -16, 1, 3,
					-- layer=2 filter=150 channel=90
					1, 7, 3, -4, 3, -9, 1, 8, 3,
					-- layer=2 filter=150 channel=91
					23, 40, 18, 8, -3, 1, -10, 13, 56,
					-- layer=2 filter=150 channel=92
					37, 1, 0, -26, 10, 5, -12, -13, 13,
					-- layer=2 filter=150 channel=93
					-12, -66, 44, 8, -32, 46, 8, -47, 24,
					-- layer=2 filter=150 channel=94
					-8, -52, -66, 26, 17, -16, 51, -25, -3,
					-- layer=2 filter=150 channel=95
					-1, 8, -4, 3, 5, 2, 8, 12, -4,
					-- layer=2 filter=150 channel=96
					-19, -23, 1, -1, 31, 24, 37, 40, 15,
					-- layer=2 filter=150 channel=97
					29, 59, 32, -38, 34, 17, -26, 26, 7,
					-- layer=2 filter=150 channel=98
					-109, -60, -32, -95, -53, -14, -26, 12, 20,
					-- layer=2 filter=150 channel=99
					-33, -32, -68, 30, 27, 23, 66, 18, -15,
					-- layer=2 filter=150 channel=100
					-9, -25, 5, -9, -29, -12, -31, -65, -44,
					-- layer=2 filter=150 channel=101
					5, -15, -16, 24, 8, 39, -73, 1, 7,
					-- layer=2 filter=150 channel=102
					-17, -31, 12, -28, 3, -1, 31, 50, -9,
					-- layer=2 filter=150 channel=103
					-35, 8, -16, -6, 33, 21, 6, 17, 43,
					-- layer=2 filter=150 channel=104
					21, -60, -20, 12, -20, 14, 13, 14, 35,
					-- layer=2 filter=150 channel=105
					-18, 18, -20, -24, -17, -13, 28, -37, -33,
					-- layer=2 filter=150 channel=106
					48, 48, 4, -3, 0, 12, -47, -30, 23,
					-- layer=2 filter=150 channel=107
					-36, -39, -22, 61, -24, 3, 5, 9, -7,
					-- layer=2 filter=150 channel=108
					25, -16, 23, -11, 10, 16, -13, -13, -51,
					-- layer=2 filter=150 channel=109
					5, 12, -6, 15, 9, -3, -3, -12, -1,
					-- layer=2 filter=150 channel=110
					-13, 10, -29, -19, -1, -34, 39, 28, 14,
					-- layer=2 filter=150 channel=111
					4, -11, 0, 0, 7, 0, 0, 10, 4,
					-- layer=2 filter=150 channel=112
					5, -17, -9, 21, -20, 78, -32, -12, 15,
					-- layer=2 filter=150 channel=113
					-10, -46, -9, -3, -69, 0, -8, -5, 50,
					-- layer=2 filter=150 channel=114
					12, -9, 9, -1, -7, -8, 4, -15, -2,
					-- layer=2 filter=150 channel=115
					0, -5, 5, -6, 7, -9, -8, 2, 1,
					-- layer=2 filter=150 channel=116
					69, 22, 30, -7, 11, -7, -14, 44, 18,
					-- layer=2 filter=150 channel=117
					-61, -74, -64, -45, -42, 34, -8, 46, 52,
					-- layer=2 filter=150 channel=118
					-33, 2, -10, -35, 20, -21, -1, 2, 19,
					-- layer=2 filter=150 channel=119
					40, -35, 3, -37, -61, -32, 22, 3, 15,
					-- layer=2 filter=150 channel=120
					9, -1, 6, -9, 8, -7, 0, -2, -3,
					-- layer=2 filter=150 channel=121
					-7, -8, -6, 8, 6, -1, 10, -8, 7,
					-- layer=2 filter=150 channel=122
					-4, 6, -10, -2, 0, -1, -1, 3, 3,
					-- layer=2 filter=150 channel=123
					-1, 18, -27, -79, -10, 0, -2, 45, 34,
					-- layer=2 filter=150 channel=124
					-6, -16, -28, -1, -1, 3, 29, 41, 49,
					-- layer=2 filter=150 channel=125
					1, 4, -7, 1, -4, -11, -7, -12, 9,
					-- layer=2 filter=150 channel=126
					-12, -20, -12, 22, 49, 18, 7, 5, 26,
					-- layer=2 filter=150 channel=127
					13, -10, -3, -68, -52, -71, -12, -12, 23,
					-- layer=2 filter=151 channel=0
					-5, 6, -8, 4, 0, -7, 0, 6, -2,
					-- layer=2 filter=151 channel=1
					-14, -10, -4, -4, -4, 7, -1, -16, -9,
					-- layer=2 filter=151 channel=2
					-2, -6, 1, -3, 3, 2, 4, -9, -2,
					-- layer=2 filter=151 channel=3
					-2, 3, -11, -11, 6, -5, 6, 7, 5,
					-- layer=2 filter=151 channel=4
					1, -10, 6, 0, -6, -6, -5, 0, 6,
					-- layer=2 filter=151 channel=5
					-1, -7, 7, 3, -8, -8, 3, -4, 1,
					-- layer=2 filter=151 channel=6
					-5, 7, -2, -4, 3, 1, -7, 0, 0,
					-- layer=2 filter=151 channel=7
					0, -6, 5, 6, -4, -4, -2, -5, -6,
					-- layer=2 filter=151 channel=8
					-5, -3, -6, 6, 3, 3, 0, 0, -5,
					-- layer=2 filter=151 channel=9
					-4, -5, -5, 5, -6, -1, -5, 1, -6,
					-- layer=2 filter=151 channel=10
					0, -9, 5, -12, 1, -12, -8, 0, -6,
					-- layer=2 filter=151 channel=11
					-1, 3, -4, -4, 4, -2, -11, -11, -5,
					-- layer=2 filter=151 channel=12
					7, 0, -9, -8, -8, -7, 2, 3, -13,
					-- layer=2 filter=151 channel=13
					-2, 2, -1, 7, 1, 8, 9, 0, 0,
					-- layer=2 filter=151 channel=14
					-6, -2, -8, -2, -2, -14, 4, 0, 5,
					-- layer=2 filter=151 channel=15
					-9, -5, 3, -5, -5, 4, -11, -9, 1,
					-- layer=2 filter=151 channel=16
					4, -8, 1, 1, -7, 0, 5, 7, -1,
					-- layer=2 filter=151 channel=17
					-6, 4, -8, -2, -9, 0, 10, 6, -11,
					-- layer=2 filter=151 channel=18
					8, 9, -11, 2, -11, 0, 1, 8, -4,
					-- layer=2 filter=151 channel=19
					-15, -4, -2, 4, 3, -7, 6, -7, 6,
					-- layer=2 filter=151 channel=20
					-5, -7, -4, 0, -2, 9, 4, 6, 9,
					-- layer=2 filter=151 channel=21
					5, 1, -5, 1, -2, 9, -10, 5, -6,
					-- layer=2 filter=151 channel=22
					-6, -3, -5, 2, 2, -5, 0, 1, 5,
					-- layer=2 filter=151 channel=23
					0, 2, 2, 1, 5, 8, -6, 0, 4,
					-- layer=2 filter=151 channel=24
					-6, -9, -5, 7, -10, 6, 9, -11, -8,
					-- layer=2 filter=151 channel=25
					-4, 4, -3, -3, 3, -8, 3, 0, 4,
					-- layer=2 filter=151 channel=26
					-10, -8, 7, -1, -6, -3, 1, -1, 9,
					-- layer=2 filter=151 channel=27
					-6, 0, -2, 6, -5, 3, -8, 6, -1,
					-- layer=2 filter=151 channel=28
					0, 8, -10, -10, 6, -1, 4, -7, -11,
					-- layer=2 filter=151 channel=29
					2, -11, 0, -11, 4, -2, 7, -8, -1,
					-- layer=2 filter=151 channel=30
					7, 4, 4, -10, -9, 5, 5, -7, -8,
					-- layer=2 filter=151 channel=31
					-3, 5, 0, 4, -4, 4, 0, 8, -4,
					-- layer=2 filter=151 channel=32
					-2, -4, -2, -7, 3, 10, 10, 2, -7,
					-- layer=2 filter=151 channel=33
					1, -8, 4, 5, -7, -7, 8, -10, -1,
					-- layer=2 filter=151 channel=34
					-6, -12, -3, 1, 8, -2, -7, 3, -9,
					-- layer=2 filter=151 channel=35
					2, -7, -14, 3, -10, 3, -3, 4, -12,
					-- layer=2 filter=151 channel=36
					5, 8, -8, -4, -9, -7, 9, -10, -10,
					-- layer=2 filter=151 channel=37
					-12, 5, -8, 0, 4, -2, -5, 5, 7,
					-- layer=2 filter=151 channel=38
					0, 1, -10, 0, 5, 2, -4, -5, 3,
					-- layer=2 filter=151 channel=39
					2, -7, 6, -3, 2, -10, 2, -6, 0,
					-- layer=2 filter=151 channel=40
					3, -9, -1, 7, -7, 3, 4, 0, 1,
					-- layer=2 filter=151 channel=41
					-7, -6, -9, -12, 9, 8, -2, 2, -4,
					-- layer=2 filter=151 channel=42
					0, -10, -11, 3, -7, 0, 1, -6, -2,
					-- layer=2 filter=151 channel=43
					-6, -11, -8, 2, -8, -8, -2, -4, 8,
					-- layer=2 filter=151 channel=44
					8, 6, -6, 2, -7, 6, 7, -9, 2,
					-- layer=2 filter=151 channel=45
					0, -7, -3, 4, 3, -10, -8, -5, 1,
					-- layer=2 filter=151 channel=46
					4, 6, 3, -11, -9, -9, 5, 0, -5,
					-- layer=2 filter=151 channel=47
					8, -8, -2, 4, -2, -8, -4, -5, -7,
					-- layer=2 filter=151 channel=48
					1, -8, 11, -6, -7, -11, -6, 4, -10,
					-- layer=2 filter=151 channel=49
					-3, 2, 1, 0, 0, 1, 2, -9, -7,
					-- layer=2 filter=151 channel=50
					4, -7, -8, -7, -1, 1, 2, 3, 2,
					-- layer=2 filter=151 channel=51
					-4, -1, 1, -5, -1, -8, -3, -9, 6,
					-- layer=2 filter=151 channel=52
					-9, -9, -9, -12, -9, -4, -11, 0, 3,
					-- layer=2 filter=151 channel=53
					2, 5, 5, -5, 8, -1, -1, -8, 0,
					-- layer=2 filter=151 channel=54
					4, 5, 0, -14, -12, -9, 6, 7, 7,
					-- layer=2 filter=151 channel=55
					5, -1, -8, -1, -9, 8, 4, -2, 4,
					-- layer=2 filter=151 channel=56
					-9, -2, -4, -11, -5, -7, -3, -10, -7,
					-- layer=2 filter=151 channel=57
					8, 1, 9, -5, -7, 8, -5, -7, 7,
					-- layer=2 filter=151 channel=58
					6, 3, 4, 0, 4, 4, -8, -5, 1,
					-- layer=2 filter=151 channel=59
					-10, 8, 1, -2, 10, 2, 0, -13, -8,
					-- layer=2 filter=151 channel=60
					7, 1, 2, 8, 3, -3, -6, -8, -7,
					-- layer=2 filter=151 channel=61
					-2, -16, -18, 1, -7, 1, -13, -2, 0,
					-- layer=2 filter=151 channel=62
					-7, 9, 4, 6, 8, -1, -11, 4, -9,
					-- layer=2 filter=151 channel=63
					2, 1, 4, -3, 0, 1, -11, -11, 5,
					-- layer=2 filter=151 channel=64
					-10, 2, -8, 2, -1, 2, 0, 1, 3,
					-- layer=2 filter=151 channel=65
					0, 5, -5, -6, 4, -2, 9, 1, 1,
					-- layer=2 filter=151 channel=66
					10, 0, 7, -5, 9, 3, -2, 7, 7,
					-- layer=2 filter=151 channel=67
					-11, -2, -5, -9, 8, 8, 5, 0, -5,
					-- layer=2 filter=151 channel=68
					1, -9, 6, 8, 5, 7, 7, 5, -10,
					-- layer=2 filter=151 channel=69
					-10, -4, 0, 4, -4, -3, -1, 6, -3,
					-- layer=2 filter=151 channel=70
					0, 6, -1, -4, -12, 1, 2, 9, -10,
					-- layer=2 filter=151 channel=71
					-8, -8, -13, 5, -9, 2, -2, -5, 3,
					-- layer=2 filter=151 channel=72
					-13, 5, 7, -12, -7, 4, -6, -11, -6,
					-- layer=2 filter=151 channel=73
					-9, -13, -12, 2, -15, -9, -1, -5, 0,
					-- layer=2 filter=151 channel=74
					-6, 3, 5, 0, -11, 4, 0, -11, 2,
					-- layer=2 filter=151 channel=75
					4, 7, -6, 4, -1, 0, 5, -7, 3,
					-- layer=2 filter=151 channel=76
					0, 8, -14, 2, -6, 1, 3, -6, -14,
					-- layer=2 filter=151 channel=77
					1, 4, 1, 6, -5, 6, 4, 3, -11,
					-- layer=2 filter=151 channel=78
					-2, -12, -12, -10, 2, -4, -3, 0, -11,
					-- layer=2 filter=151 channel=79
					-1, 4, -8, -8, -10, 2, 12, -4, 10,
					-- layer=2 filter=151 channel=80
					-5, -2, -11, 2, -1, 0, -10, 7, -4,
					-- layer=2 filter=151 channel=81
					-10, -7, -10, 1, -10, 1, 3, -7, 8,
					-- layer=2 filter=151 channel=82
					3, -2, -9, -2, -1, -6, 10, 0, 7,
					-- layer=2 filter=151 channel=83
					3, 6, -6, -8, 5, -9, 0, 0, -6,
					-- layer=2 filter=151 channel=84
					5, -5, -7, -4, 0, -8, 6, 8, -1,
					-- layer=2 filter=151 channel=85
					2, 7, -3, -8, 9, 2, 3, 9, 8,
					-- layer=2 filter=151 channel=86
					-3, -8, 6, -7, -4, 0, -3, 3, -6,
					-- layer=2 filter=151 channel=87
					1, 3, -1, 0, -1, -9, -9, -9, -6,
					-- layer=2 filter=151 channel=88
					0, -5, -9, 7, -6, -13, 9, -2, 1,
					-- layer=2 filter=151 channel=89
					1, -11, 2, -7, 0, -6, 0, -6, -2,
					-- layer=2 filter=151 channel=90
					-5, 3, -6, -1, -10, -3, -6, -3, 6,
					-- layer=2 filter=151 channel=91
					-8, -8, -7, 1, 2, -5, -3, 4, -2,
					-- layer=2 filter=151 channel=92
					-3, -2, -5, 8, -6, -7, -4, -3, -14,
					-- layer=2 filter=151 channel=93
					5, 0, 0, -3, -4, 2, -3, -4, -9,
					-- layer=2 filter=151 channel=94
					3, 0, -5, 7, -11, -7, -2, 5, -16,
					-- layer=2 filter=151 channel=95
					1, -6, 4, -2, -7, -6, 0, 1, -9,
					-- layer=2 filter=151 channel=96
					-8, -8, 5, -9, 2, -2, -5, 6, 4,
					-- layer=2 filter=151 channel=97
					-10, 1, -10, 3, 3, 3, 0, -12, 5,
					-- layer=2 filter=151 channel=98
					4, -11, 3, -4, 8, -6, -12, 2, 1,
					-- layer=2 filter=151 channel=99
					-12, -12, -10, -14, -6, 2, 0, -5, -21,
					-- layer=2 filter=151 channel=100
					1, -8, -11, 0, 6, -6, -8, -3, 2,
					-- layer=2 filter=151 channel=101
					-11, 0, 0, 2, 0, 6, 0, -7, 6,
					-- layer=2 filter=151 channel=102
					-10, 1, -6, -10, 8, -4, -5, -3, 7,
					-- layer=2 filter=151 channel=103
					-5, 5, -5, -1, 2, -11, -2, -8, -9,
					-- layer=2 filter=151 channel=104
					0, 2, -1, -9, 0, -7, 0, 1, 2,
					-- layer=2 filter=151 channel=105
					-8, -4, -9, -2, -5, -4, 4, -9, 4,
					-- layer=2 filter=151 channel=106
					-2, 0, -4, 9, 2, -1, -12, -3, -2,
					-- layer=2 filter=151 channel=107
					1, 0, 0, 1, 0, 6, -13, 3, -11,
					-- layer=2 filter=151 channel=108
					4, -2, 3, -2, 4, -4, -3, 0, -6,
					-- layer=2 filter=151 channel=109
					1, 8, 9, -7, 4, 6, 1, 2, -2,
					-- layer=2 filter=151 channel=110
					-10, -5, -2, -3, -12, -7, -1, 6, -9,
					-- layer=2 filter=151 channel=111
					-1, -5, 2, -8, 8, 1, -4, 6, 1,
					-- layer=2 filter=151 channel=112
					0, -4, -4, -3, -8, 5, 3, 2, 8,
					-- layer=2 filter=151 channel=113
					7, 5, -11, 5, 0, 4, -9, 4, -9,
					-- layer=2 filter=151 channel=114
					-4, 2, 2, 6, 4, -6, 5, 9, -10,
					-- layer=2 filter=151 channel=115
					3, -9, -10, -2, -9, 1, -7, -5, -10,
					-- layer=2 filter=151 channel=116
					3, 4, -6, 4, 1, -2, -11, -12, -13,
					-- layer=2 filter=151 channel=117
					0, -4, -16, 0, -10, -4, -3, 0, 0,
					-- layer=2 filter=151 channel=118
					5, -7, -4, 7, 1, -10, 0, -3, -11,
					-- layer=2 filter=151 channel=119
					6, 1, 2, 2, 0, 4, -8, 7, 0,
					-- layer=2 filter=151 channel=120
					6, 4, 5, -7, 8, -1, 2, 4, 10,
					-- layer=2 filter=151 channel=121
					-7, 7, -3, 0, -10, 2, -8, 10, -2,
					-- layer=2 filter=151 channel=122
					-8, 2, -10, -9, -2, 8, -1, -11, 10,
					-- layer=2 filter=151 channel=123
					-4, 8, 5, -1, 3, 0, 2, -5, -10,
					-- layer=2 filter=151 channel=124
					2, -9, -9, -13, -11, -12, -8, -14, -1,
					-- layer=2 filter=151 channel=125
					0, 1, 0, 0, 0, 1, -2, 8, 10,
					-- layer=2 filter=151 channel=126
					-8, 2, -6, 9, -1, -12, -6, 7, 2,
					-- layer=2 filter=151 channel=127
					0, -11, 0, -7, -8, 6, -12, -12, 7,
					-- layer=2 filter=152 channel=0
					-19, -27, -16, -13, -26, -17, -14, -7, -22,
					-- layer=2 filter=152 channel=1
					-1, -1, -2, -7, 2, -18, -7, -2, -20,
					-- layer=2 filter=152 channel=2
					-6, -6, 5, 9, 0, -6, 11, -4, -7,
					-- layer=2 filter=152 channel=3
					0, 0, -8, -4, -2, -1, -6, -14, -12,
					-- layer=2 filter=152 channel=4
					-10, -11, -5, -4, -10, -6, 4, -19, -2,
					-- layer=2 filter=152 channel=5
					-22, -2, -20, -16, -9, -24, -25, -9, -12,
					-- layer=2 filter=152 channel=6
					-11, -20, 1, -2, 10, -11, 0, 2, 5,
					-- layer=2 filter=152 channel=7
					-27, -5, 0, -11, -11, -20, -10, -16, -5,
					-- layer=2 filter=152 channel=8
					2, -6, 0, -5, 0, -8, 8, -10, -8,
					-- layer=2 filter=152 channel=9
					-13, -3, -19, -6, -9, -12, -19, -8, -11,
					-- layer=2 filter=152 channel=10
					-16, -23, -4, -18, -16, -13, -17, -21, -5,
					-- layer=2 filter=152 channel=11
					-20, -10, -15, -17, -12, -4, -11, -21, -11,
					-- layer=2 filter=152 channel=12
					-9, 11, -7, -14, -2, -13, 9, 8, -3,
					-- layer=2 filter=152 channel=13
					3, 0, 10, 6, 1, 8, 8, 1, -4,
					-- layer=2 filter=152 channel=14
					0, 1, -7, -10, -10, -26, -4, 3, -20,
					-- layer=2 filter=152 channel=15
					1, -2, -5, 0, -5, -3, -2, -9, 0,
					-- layer=2 filter=152 channel=16
					19, 4, -6, -2, 8, 2, -6, -1, -7,
					-- layer=2 filter=152 channel=17
					4, 9, 4, 10, 5, -2, 3, 8, -6,
					-- layer=2 filter=152 channel=18
					-9, -18, -7, -37, 0, -6, -5, -8, -18,
					-- layer=2 filter=152 channel=19
					-18, -16, -4, -24, 7, -5, 0, -6, -12,
					-- layer=2 filter=152 channel=20
					-10, 2, -6, 2, -2, 10, 1, 6, 5,
					-- layer=2 filter=152 channel=21
					9, 11, -8, -6, 0, 8, 5, -3, 7,
					-- layer=2 filter=152 channel=22
					-3, -6, -7, -10, 2, 7, -6, 0, 0,
					-- layer=2 filter=152 channel=23
					1, -3, -2, 9, 7, -9, 5, -9, -3,
					-- layer=2 filter=152 channel=24
					-1, -3, 1, -1, -12, -16, -11, -1, -14,
					-- layer=2 filter=152 channel=25
					-15, -13, -3, 7, -16, -14, -7, -16, 2,
					-- layer=2 filter=152 channel=26
					3, 6, 7, 9, -10, 3, -2, 10, 2,
					-- layer=2 filter=152 channel=27
					-30, -5, -6, -21, -7, -5, -20, -11, -12,
					-- layer=2 filter=152 channel=28
					-23, -24, -24, -5, 0, -19, 12, 0, -21,
					-- layer=2 filter=152 channel=29
					-4, 4, -2, -3, 11, 11, -6, 0, 11,
					-- layer=2 filter=152 channel=30
					2, 5, -21, -13, -11, -7, -12, -9, -13,
					-- layer=2 filter=152 channel=31
					4, -6, -12, -4, -9, 14, 1, 4, -4,
					-- layer=2 filter=152 channel=32
					1, -4, 11, 0, 7, 10, 4, -2, -1,
					-- layer=2 filter=152 channel=33
					-12, 12, 2, -8, 0, -14, -15, -35, -14,
					-- layer=2 filter=152 channel=34
					6, -7, -5, -19, -8, -4, 6, -18, -8,
					-- layer=2 filter=152 channel=35
					-9, -26, -15, -13, -11, -2, 2, -18, -8,
					-- layer=2 filter=152 channel=36
					5, 0, -6, -2, 4, -4, -8, -1, 2,
					-- layer=2 filter=152 channel=37
					-14, -7, -21, -20, -14, -12, -14, -17, -17,
					-- layer=2 filter=152 channel=38
					-18, -8, -11, -27, -13, -9, -25, -7, -5,
					-- layer=2 filter=152 channel=39
					16, 9, 9, 2, -4, -5, 7, -12, -8,
					-- layer=2 filter=152 channel=40
					-15, -4, -22, -8, -7, 18, 3, -4, -7,
					-- layer=2 filter=152 channel=41
					1, 2, 7, 4, 6, -5, -1, -4, 9,
					-- layer=2 filter=152 channel=42
					4, -5, -7, 8, -3, -7, -6, -1, -22,
					-- layer=2 filter=152 channel=43
					-15, -8, -17, -10, -14, -9, -1, -3, -17,
					-- layer=2 filter=152 channel=44
					0, -7, -1, -8, -2, -10, 2, 2, 2,
					-- layer=2 filter=152 channel=45
					-22, -7, 1, -6, -5, -4, -7, -18, 0,
					-- layer=2 filter=152 channel=46
					-16, -8, -19, -1, -12, -5, -6, -12, 3,
					-- layer=2 filter=152 channel=47
					-8, -2, -6, -8, -2, 0, -9, -23, -8,
					-- layer=2 filter=152 channel=48
					-8, 0, -8, 0, 1, 5, 7, -9, -5,
					-- layer=2 filter=152 channel=49
					-2, -16, -9, -21, -5, -23, -9, 5, -20,
					-- layer=2 filter=152 channel=50
					8, 4, 3, 7, -9, 0, -5, -2, -9,
					-- layer=2 filter=152 channel=51
					-23, -6, -22, -15, -9, 0, -11, -12, -14,
					-- layer=2 filter=152 channel=52
					-26, -24, -18, -23, -13, -20, -11, -20, -1,
					-- layer=2 filter=152 channel=53
					-12, -5, 14, -14, -10, -6, -21, 15, 0,
					-- layer=2 filter=152 channel=54
					-13, -21, -1, -16, -18, -17, -7, -6, -9,
					-- layer=2 filter=152 channel=55
					0, -3, 0, 0, -6, 6, 0, 4, -7,
					-- layer=2 filter=152 channel=56
					0, -6, -11, -13, 2, -3, 0, -17, -11,
					-- layer=2 filter=152 channel=57
					-3, -7, 1, 0, 4, 5, 0, -6, 5,
					-- layer=2 filter=152 channel=58
					2, 5, 3, -10, -2, -5, -7, -11, -18,
					-- layer=2 filter=152 channel=59
					-10, -9, 6, -26, 15, -20, -3, 5, 6,
					-- layer=2 filter=152 channel=60
					-18, 6, -12, -18, 9, -27, 5, -4, 7,
					-- layer=2 filter=152 channel=61
					-17, 8, 17, 0, -1, -8, 0, -3, 4,
					-- layer=2 filter=152 channel=62
					-8, -29, 2, -16, -7, -22, -11, -2, -17,
					-- layer=2 filter=152 channel=63
					2, 4, -3, -3, -2, -11, 7, 5, -20,
					-- layer=2 filter=152 channel=64
					-4, -9, 0, 1, -5, -3, 9, 3, -1,
					-- layer=2 filter=152 channel=65
					-11, 6, -1, -17, 12, 0, -6, -9, -1,
					-- layer=2 filter=152 channel=66
					0, -6, 2, 5, -6, 9, -4, -3, 5,
					-- layer=2 filter=152 channel=67
					-9, 1, -10, -20, -23, -2, -12, -12, 6,
					-- layer=2 filter=152 channel=68
					9, -6, -2, -6, 10, 4, 0, -6, 8,
					-- layer=2 filter=152 channel=69
					6, -8, 0, 0, -4, -16, 5, 7, -11,
					-- layer=2 filter=152 channel=70
					-12, -11, -22, -9, -3, -14, -4, -19, -8,
					-- layer=2 filter=152 channel=71
					-31, -20, -28, -17, -29, -4, -16, -18, -1,
					-- layer=2 filter=152 channel=72
					-3, -1, -5, -28, -5, -33, 11, -7, -24,
					-- layer=2 filter=152 channel=73
					-11, -10, -6, 0, -7, 3, -27, 0, 0,
					-- layer=2 filter=152 channel=74
					0, -12, -15, -14, -12, -12, -11, -12, -16,
					-- layer=2 filter=152 channel=75
					-7, 9, -13, 8, 0, -6, 1, 14, -2,
					-- layer=2 filter=152 channel=76
					-22, -13, -8, -1, -9, -11, -7, 5, 8,
					-- layer=2 filter=152 channel=77
					0, 2, 2, -10, 5, 6, 11, 4, 5,
					-- layer=2 filter=152 channel=78
					-3, -24, -21, -15, -3, -15, -3, -12, -3,
					-- layer=2 filter=152 channel=79
					-9, 9, 5, -11, 9, 5, -2, 5, 12,
					-- layer=2 filter=152 channel=80
					-12, 0, -8, -9, 1, -14, -9, -7, -7,
					-- layer=2 filter=152 channel=81
					0, 7, 6, 0, 3, -1, 1, 5, 4,
					-- layer=2 filter=152 channel=82
					-4, -5, 9, 0, 0, -10, -2, 3, -8,
					-- layer=2 filter=152 channel=83
					2, 8, -17, -10, -10, -4, -4, -7, 4,
					-- layer=2 filter=152 channel=84
					-4, 4, -9, 2, -4, 3, -6, 3, -10,
					-- layer=2 filter=152 channel=85
					1, -2, -11, 0, 6, -5, -6, 0, -11,
					-- layer=2 filter=152 channel=86
					-7, 11, 7, 1, -3, -5, 1, 2, 0,
					-- layer=2 filter=152 channel=87
					-15, -18, -19, -20, 3, -6, -5, 8, -14,
					-- layer=2 filter=152 channel=88
					-14, -2, -16, -9, -17, -19, -2, -5, -9,
					-- layer=2 filter=152 channel=89
					-9, -5, 1, -8, 0, -21, 8, 9, -16,
					-- layer=2 filter=152 channel=90
					2, -7, -1, -9, -5, -1, -9, 7, 4,
					-- layer=2 filter=152 channel=91
					-6, 1, -14, -13, -2, -23, 7, 17, -2,
					-- layer=2 filter=152 channel=92
					-2, 0, 3, -7, -8, -22, 11, 0, -19,
					-- layer=2 filter=152 channel=93
					-10, -21, -15, -10, 21, -2, -11, 1, 3,
					-- layer=2 filter=152 channel=94
					-10, 2, 11, -15, -1, -15, -6, -2, 1,
					-- layer=2 filter=152 channel=95
					0, -6, -9, -8, 10, -4, -5, 6, -1,
					-- layer=2 filter=152 channel=96
					4, -20, 9, -10, -16, -14, 27, 23, 4,
					-- layer=2 filter=152 channel=97
					-9, 0, -13, 0, -1, -10, -2, -4, 3,
					-- layer=2 filter=152 channel=98
					-20, -12, -23, -19, -16, 5, 14, -17, -25,
					-- layer=2 filter=152 channel=99
					-26, -11, -18, -17, 1, -10, -4, -6, 12,
					-- layer=2 filter=152 channel=100
					-10, 2, -4, -16, -7, -24, -28, -10, -21,
					-- layer=2 filter=152 channel=101
					-2, -20, -21, 0, -22, -28, -2, -21, -13,
					-- layer=2 filter=152 channel=102
					2, 2, -16, -15, 8, -35, 2, 2, -26,
					-- layer=2 filter=152 channel=103
					-8, -9, -6, 0, 3, -4, -3, 0, 7,
					-- layer=2 filter=152 channel=104
					-2, -6, 8, -12, -5, -25, -15, -3, -3,
					-- layer=2 filter=152 channel=105
					-8, -7, -7, -13, 8, -5, -10, 15, -10,
					-- layer=2 filter=152 channel=106
					-6, 0, -14, -1, -2, -12, 8, 6, -13,
					-- layer=2 filter=152 channel=107
					0, -7, 0, 2, 1, -3, -2, 5, -3,
					-- layer=2 filter=152 channel=108
					4, -17, -17, -17, 2, -22, 5, -10, -11,
					-- layer=2 filter=152 channel=109
					-1, -1, -7, 7, -7, 6, -4, -5, 4,
					-- layer=2 filter=152 channel=110
					9, 12, 8, 10, -4, -8, 13, -2, -6,
					-- layer=2 filter=152 channel=111
					9, 5, -3, 3, 4, 13, -8, 6, 5,
					-- layer=2 filter=152 channel=112
					-26, -5, 9, -22, -16, 6, -8, -6, -6,
					-- layer=2 filter=152 channel=113
					-10, 3, -17, -12, -16, -5, 0, 0, -14,
					-- layer=2 filter=152 channel=114
					-3, -2, 0, -3, 3, -3, 10, -8, -12,
					-- layer=2 filter=152 channel=115
					-3, 2, -4, 0, 3, -1, -5, -1, 9,
					-- layer=2 filter=152 channel=116
					-13, -4, 0, -16, -3, -11, 9, -3, -26,
					-- layer=2 filter=152 channel=117
					-15, -10, -5, -9, -18, -5, -9, -17, -14,
					-- layer=2 filter=152 channel=118
					-13, -9, -20, 1, -1, -11, -1, 2, 1,
					-- layer=2 filter=152 channel=119
					-3, -10, -25, -6, -22, -16, -10, -2, -26,
					-- layer=2 filter=152 channel=120
					7, 3, -2, -5, -10, 5, -5, -10, 0,
					-- layer=2 filter=152 channel=121
					8, 4, 3, -9, 2, -1, 0, 3, 8,
					-- layer=2 filter=152 channel=122
					0, 5, 7, 7, -1, -10, 8, -3, 6,
					-- layer=2 filter=152 channel=123
					-7, -13, -6, -17, -4, -14, -15, -12, -11,
					-- layer=2 filter=152 channel=124
					-5, 2, -14, 3, -13, -20, -20, -16, -14,
					-- layer=2 filter=152 channel=125
					-7, 5, -10, -5, 6, 2, 10, 6, 5,
					-- layer=2 filter=152 channel=126
					9, -6, 27, 2, -9, -10, 5, 3, 11,
					-- layer=2 filter=152 channel=127
					-12, 1, 3, -4, -17, -25, 0, -12, -28,
					-- layer=2 filter=153 channel=0
					-27, -11, -3, -11, -4, -18, -6, -39, -35,
					-- layer=2 filter=153 channel=1
					0, -1, 8, -18, 1, 19, 13, -9, 0,
					-- layer=2 filter=153 channel=2
					4, 2, 2, -3, 8, 0, -6, 9, -6,
					-- layer=2 filter=153 channel=3
					4, -14, -37, 5, 12, -53, 11, 29, -9,
					-- layer=2 filter=153 channel=4
					-16, 40, 49, -6, 12, 34, -58, -42, -35,
					-- layer=2 filter=153 channel=5
					12, 10, -3, -37, 12, -39, -17, 6, -44,
					-- layer=2 filter=153 channel=6
					-15, -38, 27, 0, -19, 31, 5, -17, -9,
					-- layer=2 filter=153 channel=7
					-16, 25, -33, -12, -14, -1, -55, -58, -11,
					-- layer=2 filter=153 channel=8
					-3, 2, 5, -5, -12, 5, -2, -7, -3,
					-- layer=2 filter=153 channel=9
					-14, -9, -12, -26, -22, -7, -17, 4, -9,
					-- layer=2 filter=153 channel=10
					-20, -9, -2, -6, 3, -34, -15, -9, -21,
					-- layer=2 filter=153 channel=11
					22, 24, -6, 3, 10, -7, 10, -3, -17,
					-- layer=2 filter=153 channel=12
					0, -3, 10, -3, 18, 35, -28, 2, 22,
					-- layer=2 filter=153 channel=13
					0, -3, -6, -3, 1, -6, -3, 6, -8,
					-- layer=2 filter=153 channel=14
					-12, 11, 23, -16, 11, 19, 11, 17, 18,
					-- layer=2 filter=153 channel=15
					-3, 69, 29, 22, -18, 25, 14, -8, 9,
					-- layer=2 filter=153 channel=16
					23, 21, 2, 41, 10, -14, 6, -14, -4,
					-- layer=2 filter=153 channel=17
					-7, 4, 7, 3, -9, 8, -7, -1, 0,
					-- layer=2 filter=153 channel=18
					30, 49, 44, 20, 55, 55, 31, 10, 22,
					-- layer=2 filter=153 channel=19
					16, -6, 13, -1, -2, 18, 21, -32, -13,
					-- layer=2 filter=153 channel=20
					-5, -8, -9, 6, -6, -5, -4, -5, 10,
					-- layer=2 filter=153 channel=21
					9, -3, -3, -10, 2, 2, 0, 18, 0,
					-- layer=2 filter=153 channel=22
					2, -2, -4, 9, -6, -6, -6, -9, -10,
					-- layer=2 filter=153 channel=23
					8, 5, 14, 27, 24, 40, -8, -18, -6,
					-- layer=2 filter=153 channel=24
					-5, -8, -33, 10, -14, -36, 23, 17, 5,
					-- layer=2 filter=153 channel=25
					14, -27, -47, 11, 10, -16, 1, 6, 0,
					-- layer=2 filter=153 channel=26
					-2, -7, 5, 0, 9, 6, -6, -7, 0,
					-- layer=2 filter=153 channel=27
					26, 14, 20, -27, -42, -1, -33, -25, 0,
					-- layer=2 filter=153 channel=28
					-32, -23, 1, -24, -14, 17, -33, -6, -29,
					-- layer=2 filter=153 channel=29
					6, 9, 1, 2, -9, -6, -1, -6, 9,
					-- layer=2 filter=153 channel=30
					-17, -28, 15, 23, -30, -41, 3, -20, -25,
					-- layer=2 filter=153 channel=31
					-28, 40, 13, 3, -1, -1, 11, -27, 28,
					-- layer=2 filter=153 channel=32
					8, -2, -2, 4, 9, -5, 4, 8, -7,
					-- layer=2 filter=153 channel=33
					-18, 28, -4, -16, -33, 13, -66, -21, 0,
					-- layer=2 filter=153 channel=34
					15, 23, -9, 31, 10, -5, 46, -33, -26,
					-- layer=2 filter=153 channel=35
					-30, 8, 26, -1, -3, 8, -74, -84, -58,
					-- layer=2 filter=153 channel=36
					12, 4, -8, 5, -6, 9, -4, -11, 1,
					-- layer=2 filter=153 channel=37
					34, 12, 3, 10, 0, -32, -8, 0, -16,
					-- layer=2 filter=153 channel=38
					-28, -33, 12, -39, -18, -5, -25, 0, -5,
					-- layer=2 filter=153 channel=39
					-60, 7, -20, 24, -29, -33, -38, -34, 13,
					-- layer=2 filter=153 channel=40
					6, -29, 42, 44, 5, 40, 31, 3, 35,
					-- layer=2 filter=153 channel=41
					8, 1, -4, -1, -8, -1, 3, 0, 0,
					-- layer=2 filter=153 channel=42
					5, 3, 7, 14, 12, -6, -18, 11, 39,
					-- layer=2 filter=153 channel=43
					17, 5, 33, 36, 1, -24, -20, 17, 15,
					-- layer=2 filter=153 channel=44
					-5, 7, -1, -8, 2, -7, 4, 6, 4,
					-- layer=2 filter=153 channel=45
					35, 53, 35, -56, -45, 25, -61, -23, 42,
					-- layer=2 filter=153 channel=46
					-78, -11, 20, -28, -22, 17, -5, -62, -43,
					-- layer=2 filter=153 channel=47
					-12, 18, 8, -15, -16, -57, -39, -60, -11,
					-- layer=2 filter=153 channel=48
					6, 9, -1, 1, -7, -2, -6, -6, -8,
					-- layer=2 filter=153 channel=49
					35, 39, 77, 12, 30, 73, 51, 32, 47,
					-- layer=2 filter=153 channel=50
					18, -4, -2, -24, -11, -18, -16, -9, 5,
					-- layer=2 filter=153 channel=51
					7, 22, -7, 12, 9, -47, -2, 3, -19,
					-- layer=2 filter=153 channel=52
					-28, 43, 19, 28, -16, -25, 0, -35, -23,
					-- layer=2 filter=153 channel=53
					-30, 2, 0, -2, -35, -7, -19, 6, 2,
					-- layer=2 filter=153 channel=54
					12, 19, 18, -6, 44, 35, -12, -20, 15,
					-- layer=2 filter=153 channel=55
					0, -1, -3, -9, 2, 2, 8, -3, 0,
					-- layer=2 filter=153 channel=56
					39, 30, -18, 0, 25, -22, 5, 10, 6,
					-- layer=2 filter=153 channel=57
					0, 4, 5, -3, -12, 7, -12, 3, 12,
					-- layer=2 filter=153 channel=58
					-10, -14, 15, -34, 3, 15, -14, -7, 37,
					-- layer=2 filter=153 channel=59
					-16, -43, 11, -79, -34, 50, 13, -30, 18,
					-- layer=2 filter=153 channel=60
					-11, -39, -22, -50, 12, 0, 14, -7, 20,
					-- layer=2 filter=153 channel=61
					-11, -62, 3, -33, -23, -6, 21, -14, -27,
					-- layer=2 filter=153 channel=62
					30, 0, 37, 5, 0, 53, 46, -5, 7,
					-- layer=2 filter=153 channel=63
					-22, -13, -18, -23, -27, -6, -21, -51, 9,
					-- layer=2 filter=153 channel=64
					-21, -37, -9, 29, 29, 13, 14, 7, 22,
					-- layer=2 filter=153 channel=65
					-15, -57, -41, -18, -8, 22, -4, -39, -27,
					-- layer=2 filter=153 channel=66
					-31, 43, -26, 15, 14, 12, 5, 39, 4,
					-- layer=2 filter=153 channel=67
					-24, -5, -13, -44, -6, -41, 0, -6, -38,
					-- layer=2 filter=153 channel=68
					11, -7, -2, -2, -2, -3, -8, -1, -4,
					-- layer=2 filter=153 channel=69
					-28, -23, 29, 24, -2, -10, 16, -8, 11,
					-- layer=2 filter=153 channel=70
					-16, 2, 14, -29, 6, -25, -76, -41, -35,
					-- layer=2 filter=153 channel=71
					44, -6, 8, 1, -28, 8, 12, 9, 32,
					-- layer=2 filter=153 channel=72
					37, 10, 8, -14, 5, 31, -47, -4, 30,
					-- layer=2 filter=153 channel=73
					65, 23, 8, 53, 19, -14, 42, 49, 46,
					-- layer=2 filter=153 channel=74
					-78, 5, -2, -40, -11, 28, -34, -21, -41,
					-- layer=2 filter=153 channel=75
					-6, -3, -4, 42, 20, 11, 92, 50, -2,
					-- layer=2 filter=153 channel=76
					-27, 23, 38, 10, -16, -2, -5, 4, 8,
					-- layer=2 filter=153 channel=77
					9, 2, -4, 2, 2, -4, 5, -2, 6,
					-- layer=2 filter=153 channel=78
					18, 8, -9, 23, 19, -7, 33, 4, -24,
					-- layer=2 filter=153 channel=79
					3, 9, -9, 0, -1, 3, -10, -1, 5,
					-- layer=2 filter=153 channel=80
					0, -1, 14, 3, -1, -25, -21, -11, -39,
					-- layer=2 filter=153 channel=81
					16, 1, 6, 12, -2, 1, -2, 1, 7,
					-- layer=2 filter=153 channel=82
					-2, 0, 13, 1, 8, -3, -1, -3, 9,
					-- layer=2 filter=153 channel=83
					28, 21, 39, 7, -12, 12, -25, 4, -17,
					-- layer=2 filter=153 channel=84
					-6, 7, -6, -2, 4, 1, -6, 3, -3,
					-- layer=2 filter=153 channel=85
					2, -4, 16, 3, 1, 18, 0, 1, 10,
					-- layer=2 filter=153 channel=86
					-6, 8, -6, 1, -12, -13, 20, 5, 12,
					-- layer=2 filter=153 channel=87
					-3, 15, 64, 1, -15, 48, -32, -20, 24,
					-- layer=2 filter=153 channel=88
					-54, -11, 1, -17, -34, -41, -44, -28, 7,
					-- layer=2 filter=153 channel=89
					-9, -25, 27, -19, -20, 14, -26, -18, 0,
					-- layer=2 filter=153 channel=90
					-6, -11, -3, -5, 6, 2, 1, 5, -2,
					-- layer=2 filter=153 channel=91
					11, -4, 7, -11, -18, 24, -21, 0, 21,
					-- layer=2 filter=153 channel=92
					-10, -3, 8, -13, -1, 29, -16, -5, 24,
					-- layer=2 filter=153 channel=93
					22, -46, 0, 57, 32, 14, 13, -29, -35,
					-- layer=2 filter=153 channel=94
					-30, -18, 27, -4, -34, -15, 0, -20, -32,
					-- layer=2 filter=153 channel=95
					10, 20, 7, 22, 13, 11, 12, 8, 7,
					-- layer=2 filter=153 channel=96
					-26, -32, -1, -14, -16, -16, 9, 39, 4,
					-- layer=2 filter=153 channel=97
					-16, -18, 48, 2, 2, -3, 0, 16, 0,
					-- layer=2 filter=153 channel=98
					2, -2, 17, -9, 3, 8, -43, -20, -21,
					-- layer=2 filter=153 channel=99
					13, -18, 57, -8, -6, 7, 3, -18, -21,
					-- layer=2 filter=153 channel=100
					-7, -18, 16, -52, 4, 5, -21, -38, 13,
					-- layer=2 filter=153 channel=101
					25, 33, -19, 24, 16, 18, 12, 4, 29,
					-- layer=2 filter=153 channel=102
					27, 53, 33, -8, 31, 31, 37, 9, 22,
					-- layer=2 filter=153 channel=103
					-47, 2, -7, -1, 36, -39, -34, -11, -20,
					-- layer=2 filter=153 channel=104
					27, 67, 50, -1, 32, 36, 6, -4, 10,
					-- layer=2 filter=153 channel=105
					44, 6, -5, 25, 32, -40, 0, -37, -60,
					-- layer=2 filter=153 channel=106
					-11, -6, -26, -23, -28, -20, -6, 13, -6,
					-- layer=2 filter=153 channel=107
					-44, 4, -13, 36, 32, -4, -6, -23, 33,
					-- layer=2 filter=153 channel=108
					2, 0, 11, -35, -7, 13, 16, 32, -13,
					-- layer=2 filter=153 channel=109
					1, -14, 22, 14, -4, 13, 7, 12, -9,
					-- layer=2 filter=153 channel=110
					0, -4, -55, 24, 12, -13, 14, 19, 7,
					-- layer=2 filter=153 channel=111
					6, -11, 2, -1, 0, -1, 7, 6, -3,
					-- layer=2 filter=153 channel=112
					-24, 45, -9, -41, -13, -29, -37, -44, -9,
					-- layer=2 filter=153 channel=113
					-35, -20, 11, -39, 10, -23, -23, -22, -15,
					-- layer=2 filter=153 channel=114
					-11, -2, 0, -7, -3, -5, -4, -6, -23,
					-- layer=2 filter=153 channel=115
					-1, 0, 8, 1, 4, -9, -4, 4, -2,
					-- layer=2 filter=153 channel=116
					9, 35, 35, -19, -1, 24, -15, 31, 8,
					-- layer=2 filter=153 channel=117
					32, 41, -30, 0, 3, 15, -33, -25, -7,
					-- layer=2 filter=153 channel=118
					25, 4, 27, 31, 24, 19, 19, 17, -18,
					-- layer=2 filter=153 channel=119
					1, 31, 61, -42, 4, 29, -13, 0, 11,
					-- layer=2 filter=153 channel=120
					0, 6, -3, 5, -6, -1, -1, -3, -10,
					-- layer=2 filter=153 channel=121
					-8, 9, 9, -9, 9, -6, -5, -6, 7,
					-- layer=2 filter=153 channel=122
					-8, -8, -1, 0, 0, 0, 0, -3, 2,
					-- layer=2 filter=153 channel=123
					-4, -13, 7, 6, -25, 26, -33, -38, -15,
					-- layer=2 filter=153 channel=124
					-28, -4, 29, 36, 0, 16, 1, 10, 18,
					-- layer=2 filter=153 channel=125
					9, -1, 1, -11, 2, 5, -1, 5, 8,
					-- layer=2 filter=153 channel=126
					-9, -56, -26, 13, -69, 15, 60, 19, 36,
					-- layer=2 filter=153 channel=127
					-34, 9, 28, -59, 1, 8, -37, 0, 20,
					-- layer=2 filter=154 channel=0
					-2, -6, -7, -8, 6, 1, -4, 0, 6,
					-- layer=2 filter=154 channel=1
					-10, -8, 8, -16, -8, -1, -12, -17, -13,
					-- layer=2 filter=154 channel=2
					5, 1, 7, 0, 4, 8, -1, 8, -7,
					-- layer=2 filter=154 channel=3
					-6, 7, -8, 0, 6, -10, 1, -6, 5,
					-- layer=2 filter=154 channel=4
					-12, 0, 0, -5, 8, -6, -4, 5, 1,
					-- layer=2 filter=154 channel=5
					-6, -2, -4, -6, -8, -7, -9, -5, 7,
					-- layer=2 filter=154 channel=6
					-2, -10, -13, -1, -7, 3, -18, -4, -3,
					-- layer=2 filter=154 channel=7
					5, -5, -4, 4, -1, -3, -10, -5, -15,
					-- layer=2 filter=154 channel=8
					2, 1, 8, -1, -1, 9, 6, 9, -2,
					-- layer=2 filter=154 channel=9
					8, 2, -4, -6, -9, -6, 6, -4, 0,
					-- layer=2 filter=154 channel=10
					4, -13, 0, -5, -8, 0, 3, -6, 8,
					-- layer=2 filter=154 channel=11
					4, -13, 4, 6, -13, -13, -15, -6, -17,
					-- layer=2 filter=154 channel=12
					6, -8, 1, 6, -2, -11, -3, -9, -7,
					-- layer=2 filter=154 channel=13
					0, 5, 0, -2, 1, -1, -10, -1, 0,
					-- layer=2 filter=154 channel=14
					5, 7, -2, 2, 4, 1, -11, -5, 2,
					-- layer=2 filter=154 channel=15
					-1, -8, 5, -11, -4, -1, -14, 5, 5,
					-- layer=2 filter=154 channel=16
					-1, 3, -4, 3, -11, -5, 1, 8, -3,
					-- layer=2 filter=154 channel=17
					-8, -4, 10, -4, -6, -6, 8, 11, 0,
					-- layer=2 filter=154 channel=18
					-15, 1, -2, -7, -5, -18, -7, -3, -1,
					-- layer=2 filter=154 channel=19
					-5, 3, 4, -2, 8, -1, -22, 0, -2,
					-- layer=2 filter=154 channel=20
					1, -9, -4, 9, 0, 6, 10, -8, -8,
					-- layer=2 filter=154 channel=21
					7, 0, 5, 5, -3, 3, 0, 0, 0,
					-- layer=2 filter=154 channel=22
					3, 8, 5, -6, -9, -11, -6, 4, 2,
					-- layer=2 filter=154 channel=23
					5, -5, 5, -4, 1, -13, 8, 6, -10,
					-- layer=2 filter=154 channel=24
					-1, 4, -2, 2, -8, -2, 0, 3, -3,
					-- layer=2 filter=154 channel=25
					-5, -12, -13, -1, -17, -5, -11, -16, -1,
					-- layer=2 filter=154 channel=26
					8, -6, -3, 2, 6, 6, -8, 1, -2,
					-- layer=2 filter=154 channel=27
					-7, 2, 0, 7, 8, 0, -5, 7, -3,
					-- layer=2 filter=154 channel=28
					-2, 10, 6, -3, -5, 0, 0, -5, -6,
					-- layer=2 filter=154 channel=29
					-11, -9, 4, 1, 0, 6, -8, -9, -3,
					-- layer=2 filter=154 channel=30
					4, 8, 4, 9, -10, -3, 7, 4, -11,
					-- layer=2 filter=154 channel=31
					0, 1, 1, 5, -4, -5, -1, 1, 7,
					-- layer=2 filter=154 channel=32
					0, 3, 5, 12, 5, 9, -6, 0, 11,
					-- layer=2 filter=154 channel=33
					-7, -8, -2, -3, -6, -4, 3, -11, 2,
					-- layer=2 filter=154 channel=34
					5, -11, -3, -13, -5, -13, -12, 8, -1,
					-- layer=2 filter=154 channel=35
					-13, 3, 6, -2, 9, -12, 5, 2, -14,
					-- layer=2 filter=154 channel=36
					-8, -5, 1, -6, 0, 1, 0, 4, 0,
					-- layer=2 filter=154 channel=37
					-11, -14, -15, -7, -15, -12, -6, -2, 0,
					-- layer=2 filter=154 channel=38
					-8, 0, 1, -4, -8, 2, -6, 2, -1,
					-- layer=2 filter=154 channel=39
					2, -4, -6, -9, -5, 0, -8, -9, -10,
					-- layer=2 filter=154 channel=40
					-5, -4, -2, 1, -7, -12, -3, 7, -1,
					-- layer=2 filter=154 channel=41
					2, -1, 8, 1, -2, 3, 5, -4, -3,
					-- layer=2 filter=154 channel=42
					-6, 8, -3, -8, -10, -4, 1, 7, 3,
					-- layer=2 filter=154 channel=43
					-2, 6, -14, -3, -5, -2, -6, 6, -9,
					-- layer=2 filter=154 channel=44
					3, -6, -8, 8, 4, 7, 3, -9, -4,
					-- layer=2 filter=154 channel=45
					-12, 9, -2, -4, 1, -16, 4, -5, 0,
					-- layer=2 filter=154 channel=46
					-7, -4, -7, -10, 1, 0, 3, -8, -4,
					-- layer=2 filter=154 channel=47
					-4, 0, -8, -4, 0, -8, 3, 5, -13,
					-- layer=2 filter=154 channel=48
					4, -12, 1, -7, 1, -3, 3, 8, 2,
					-- layer=2 filter=154 channel=49
					5, -11, -12, -8, -1, -11, -9, -16, -8,
					-- layer=2 filter=154 channel=50
					0, -10, -7, -5, 0, 11, 10, 1, -3,
					-- layer=2 filter=154 channel=51
					-8, -10, 4, -2, 6, -5, -1, -2, -12,
					-- layer=2 filter=154 channel=52
					-15, 0, -14, 4, -14, -9, -5, -1, -11,
					-- layer=2 filter=154 channel=53
					4, 10, -6, 8, -4, -1, -9, 0, 4,
					-- layer=2 filter=154 channel=54
					-10, -4, 0, 11, -7, -5, -7, 4, -14,
					-- layer=2 filter=154 channel=55
					0, 10, 1, -8, 10, -9, 9, -3, 7,
					-- layer=2 filter=154 channel=56
					1, -4, -2, -1, -8, -10, 0, -7, -5,
					-- layer=2 filter=154 channel=57
					5, -7, 1, -5, -1, 10, -3, 2, 4,
					-- layer=2 filter=154 channel=58
					-8, 5, -6, -3, 5, -9, -4, -4, -8,
					-- layer=2 filter=154 channel=59
					-6, -10, 3, 0, -8, -11, -3, -4, -6,
					-- layer=2 filter=154 channel=60
					2, 3, -9, -6, 4, 2, -5, 6, 0,
					-- layer=2 filter=154 channel=61
					-5, -6, 2, 5, 4, -1, 0, 13, 5,
					-- layer=2 filter=154 channel=62
					-4, -13, 2, -3, -9, -18, -4, -6, -18,
					-- layer=2 filter=154 channel=63
					-10, -9, -12, -3, -8, -7, -2, -9, 0,
					-- layer=2 filter=154 channel=64
					-6, 6, 4, -5, -6, -2, 1, 3, 1,
					-- layer=2 filter=154 channel=65
					1, 1, -6, -6, 5, 2, 9, -4, 2,
					-- layer=2 filter=154 channel=66
					1, -8, -2, 6, -9, 8, 5, 9, -3,
					-- layer=2 filter=154 channel=67
					-2, -9, -8, 1, 4, -8, 7, -1, 7,
					-- layer=2 filter=154 channel=68
					6, -2, 8, 3, 7, -6, -12, -2, 5,
					-- layer=2 filter=154 channel=69
					5, -4, 8, 0, -10, -11, -5, -4, 7,
					-- layer=2 filter=154 channel=70
					3, 0, -12, -3, 10, 3, -5, 0, -17,
					-- layer=2 filter=154 channel=71
					0, -9, -4, -3, -8, 7, 1, -10, -3,
					-- layer=2 filter=154 channel=72
					-11, 11, -9, -4, -1, -5, -14, 6, -20,
					-- layer=2 filter=154 channel=73
					-4, 4, -13, 6, 0, -5, -16, -3, -5,
					-- layer=2 filter=154 channel=74
					-4, 2, -2, 0, 0, 0, -9, 6, -9,
					-- layer=2 filter=154 channel=75
					1, 9, 8, 9, -3, 4, -9, 2, -5,
					-- layer=2 filter=154 channel=76
					-9, -2, 0, -1, -18, -6, -14, -2, -16,
					-- layer=2 filter=154 channel=77
					-8, -1, 10, 2, 1, 7, 0, 3, 0,
					-- layer=2 filter=154 channel=78
					-7, 8, -13, -5, 4, -4, 0, 1, 6,
					-- layer=2 filter=154 channel=79
					3, 4, 8, 0, -2, -5, 5, 2, 7,
					-- layer=2 filter=154 channel=80
					6, 8, -9, -9, 5, -11, -7, -10, -11,
					-- layer=2 filter=154 channel=81
					8, 3, 8, -6, 8, 0, -1, 5, 4,
					-- layer=2 filter=154 channel=82
					8, 0, 3, -5, 0, 0, 4, -3, -3,
					-- layer=2 filter=154 channel=83
					0, 4, 8, -10, 3, 5, 0, 0, 0,
					-- layer=2 filter=154 channel=84
					4, 5, 10, -1, -3, -9, -10, 3, 3,
					-- layer=2 filter=154 channel=85
					-7, 7, 4, -3, -10, -6, -5, -2, 4,
					-- layer=2 filter=154 channel=86
					-4, 5, 5, -8, 1, -6, -5, -8, 7,
					-- layer=2 filter=154 channel=87
					-9, 2, -8, -2, -5, 1, -11, -2, 3,
					-- layer=2 filter=154 channel=88
					-8, -4, -3, -4, 6, 1, 0, -12, -5,
					-- layer=2 filter=154 channel=89
					-3, -10, 0, 5, -11, -1, 5, -3, 6,
					-- layer=2 filter=154 channel=90
					0, -1, 4, 10, 10, -3, 8, -7, 5,
					-- layer=2 filter=154 channel=91
					0, -16, 4, -13, 0, -14, -5, 0, -4,
					-- layer=2 filter=154 channel=92
					-10, -11, -1, 0, 1, -4, -5, -15, -17,
					-- layer=2 filter=154 channel=93
					-14, -16, -8, -2, 5, 2, 8, -6, -10,
					-- layer=2 filter=154 channel=94
					0, 0, -1, -3, 0, -5, -10, -2, -11,
					-- layer=2 filter=154 channel=95
					0, 5, 0, -9, 5, -10, -6, 5, -11,
					-- layer=2 filter=154 channel=96
					-6, 5, -1, -7, 3, 2, -2, -6, 9,
					-- layer=2 filter=154 channel=97
					2, -9, 5, 4, 7, 0, -6, -5, 0,
					-- layer=2 filter=154 channel=98
					-8, -11, -11, 4, -7, 2, 5, 3, -15,
					-- layer=2 filter=154 channel=99
					3, 4, -7, 2, -3, 4, -6, -5, -8,
					-- layer=2 filter=154 channel=100
					7, -3, -4, -6, -2, 0, 0, -6, 0,
					-- layer=2 filter=154 channel=101
					-11, -3, -11, -8, -2, -7, -21, -18, -13,
					-- layer=2 filter=154 channel=102
					3, -3, 0, -12, -4, -5, -12, -2, -9,
					-- layer=2 filter=154 channel=103
					-9, -3, 4, -3, -4, -10, -4, -3, 5,
					-- layer=2 filter=154 channel=104
					4, 0, -7, 7, 0, 0, -4, -9, -13,
					-- layer=2 filter=154 channel=105
					-5, 6, 9, 2, -12, -6, -5, 8, 7,
					-- layer=2 filter=154 channel=106
					-3, -7, -7, 1, 0, -3, 6, -3, -3,
					-- layer=2 filter=154 channel=107
					-4, -5, -3, 7, 0, 2, 5, 2, -6,
					-- layer=2 filter=154 channel=108
					5, -9, -5, -2, -6, -9, -11, 4, -8,
					-- layer=2 filter=154 channel=109
					0, -8, -4, 5, 3, 5, 4, 1, -3,
					-- layer=2 filter=154 channel=110
					-10, 1, -7, -6, 1, -10, -4, 5, 6,
					-- layer=2 filter=154 channel=111
					-2, 0, -5, 9, -9, 1, 2, 7, 9,
					-- layer=2 filter=154 channel=112
					-13, -12, -3, -2, -2, -11, 0, 8, -6,
					-- layer=2 filter=154 channel=113
					-8, -11, 6, -6, 4, -2, 7, 5, 0,
					-- layer=2 filter=154 channel=114
					6, -10, 5, -11, 4, 3, 2, -5, -5,
					-- layer=2 filter=154 channel=115
					-3, 0, -5, -1, -8, -4, 8, -5, -5,
					-- layer=2 filter=154 channel=116
					-10, -10, 1, 4, 0, 2, 1, -4, -9,
					-- layer=2 filter=154 channel=117
					3, -6, 2, 9, -12, 1, -8, 3, -9,
					-- layer=2 filter=154 channel=118
					-7, -7, 0, -12, -10, -13, -5, 2, 6,
					-- layer=2 filter=154 channel=119
					1, -4, 9, -3, 7, -4, -14, -10, 6,
					-- layer=2 filter=154 channel=120
					-5, -1, 10, 6, 5, -4, 2, 1, -6,
					-- layer=2 filter=154 channel=121
					0, -4, 9, -4, 12, -1, 0, -9, 0,
					-- layer=2 filter=154 channel=122
					4, -1, 3, 5, 3, 6, 4, -8, -6,
					-- layer=2 filter=154 channel=123
					1, -5, 2, 0, -9, -3, -1, -14, -17,
					-- layer=2 filter=154 channel=124
					0, -7, 6, -15, -9, -9, -7, -4, -19,
					-- layer=2 filter=154 channel=125
					6, -8, -7, 0, -4, 8, 11, -3, 1,
					-- layer=2 filter=154 channel=126
					0, -2, -9, -3, 0, 7, 3, -9, 10,
					-- layer=2 filter=154 channel=127
					-11, -5, 10, 7, 9, -1, 0, 1, -7,
					-- layer=2 filter=155 channel=0
					-2, -6, -11, -6, -8, -12, 4, -4, 0,
					-- layer=2 filter=155 channel=1
					-10, -6, -10, 7, 7, -8, 4, -14, -11,
					-- layer=2 filter=155 channel=2
					-5, -6, 9, -4, 2, 6, 6, -5, 10,
					-- layer=2 filter=155 channel=3
					-2, -5, 8, -12, 4, -10, -7, -7, 0,
					-- layer=2 filter=155 channel=4
					-8, -1, -8, 1, -12, -5, 0, 0, -3,
					-- layer=2 filter=155 channel=5
					2, 1, -12, -6, 6, 5, -1, 6, 6,
					-- layer=2 filter=155 channel=6
					0, -2, 3, -4, 0, -7, -4, -5, -8,
					-- layer=2 filter=155 channel=7
					-8, -13, -5, 0, -6, -10, 0, -5, -15,
					-- layer=2 filter=155 channel=8
					5, -3, -5, -6, -2, 4, 2, -6, 2,
					-- layer=2 filter=155 channel=9
					0, 1, 3, 4, -9, -8, -9, 6, 3,
					-- layer=2 filter=155 channel=10
					3, 6, -8, 0, -4, -3, 5, 0, -13,
					-- layer=2 filter=155 channel=11
					-15, 3, -9, -4, -12, 3, -9, -4, 3,
					-- layer=2 filter=155 channel=12
					-7, -9, 1, 9, -8, 8, -4, 0, -11,
					-- layer=2 filter=155 channel=13
					-10, 7, -4, 0, 0, -4, 2, 0, 8,
					-- layer=2 filter=155 channel=14
					5, 0, -8, 0, 5, -5, -3, 5, 0,
					-- layer=2 filter=155 channel=15
					-9, 3, -7, -8, 4, 2, -1, -8, 4,
					-- layer=2 filter=155 channel=16
					3, -2, 6, -7, 5, 6, -4, -8, -6,
					-- layer=2 filter=155 channel=17
					-1, 7, 0, 4, -1, -1, 9, -9, -6,
					-- layer=2 filter=155 channel=18
					-15, 3, 6, -12, -16, 6, -3, -1, -3,
					-- layer=2 filter=155 channel=19
					-7, 4, -9, 0, -4, 7, -6, -12, 6,
					-- layer=2 filter=155 channel=20
					-11, 5, 7, -7, -1, 6, -7, -5, 6,
					-- layer=2 filter=155 channel=21
					3, 7, -3, 1, 0, -12, -3, 0, -10,
					-- layer=2 filter=155 channel=22
					6, 7, -1, 4, -3, 6, -5, 8, -3,
					-- layer=2 filter=155 channel=23
					-3, 7, 7, -9, 6, -4, -4, 2, -6,
					-- layer=2 filter=155 channel=24
					4, -4, -3, -3, 0, -9, 0, -10, -10,
					-- layer=2 filter=155 channel=25
					-11, -7, 9, -12, 9, -9, 2, -9, 4,
					-- layer=2 filter=155 channel=26
					4, 2, -1, 0, -1, 2, 6, 9, -2,
					-- layer=2 filter=155 channel=27
					-1, -11, 2, -11, -6, -15, -9, -8, -3,
					-- layer=2 filter=155 channel=28
					-10, 2, -1, 0, 0, 2, 4, -5, -12,
					-- layer=2 filter=155 channel=29
					6, 11, -5, 7, 0, -4, -4, -7, -1,
					-- layer=2 filter=155 channel=30
					2, -1, -10, -8, 6, 8, -3, -9, -8,
					-- layer=2 filter=155 channel=31
					-2, 6, 5, 5, -10, -4, 0, 2, -6,
					-- layer=2 filter=155 channel=32
					5, 7, 2, -4, 5, 4, 7, -5, 6,
					-- layer=2 filter=155 channel=33
					-8, -6, -11, -13, -6, -8, -3, -13, -7,
					-- layer=2 filter=155 channel=34
					-2, 3, 5, -2, -4, -14, 9, 5, 8,
					-- layer=2 filter=155 channel=35
					-10, -5, -11, 3, 1, -3, -6, 5, 9,
					-- layer=2 filter=155 channel=36
					0, 5, 2, 5, -7, 8, -4, -2, 8,
					-- layer=2 filter=155 channel=37
					2, 3, -1, 0, 0, -6, -3, -11, -7,
					-- layer=2 filter=155 channel=38
					-5, -11, -5, -6, -14, 1, 0, 2, 2,
					-- layer=2 filter=155 channel=39
					-3, -10, -5, -7, -5, 8, -3, -2, 9,
					-- layer=2 filter=155 channel=40
					-8, -13, -13, 0, -2, -5, 0, -2, 7,
					-- layer=2 filter=155 channel=41
					-2, 3, 6, 9, -8, -8, 5, 7, -4,
					-- layer=2 filter=155 channel=42
					0, -9, 3, 3, 9, -7, -1, 0, 3,
					-- layer=2 filter=155 channel=43
					-14, -7, 0, 3, 5, -5, 5, 0, -4,
					-- layer=2 filter=155 channel=44
					-3, -5, -5, 5, -10, -8, 2, -8, -7,
					-- layer=2 filter=155 channel=45
					-2, -8, -6, -8, 6, 0, 5, 9, 2,
					-- layer=2 filter=155 channel=46
					0, -8, -10, -3, 0, 6, -1, -7, -5,
					-- layer=2 filter=155 channel=47
					3, 5, 1, 2, 3, -2, 8, -6, -1,
					-- layer=2 filter=155 channel=48
					6, 5, 10, 5, -3, 5, -1, -5, 1,
					-- layer=2 filter=155 channel=49
					0, -11, -14, -17, -19, 10, -12, -15, -2,
					-- layer=2 filter=155 channel=50
					7, 4, 5, 0, -2, -2, 7, -6, 3,
					-- layer=2 filter=155 channel=51
					-2, -12, 3, 2, -7, -4, -9, -7, -2,
					-- layer=2 filter=155 channel=52
					-11, 0, -6, -14, -12, -11, -2, 0, -9,
					-- layer=2 filter=155 channel=53
					8, 5, -8, -7, -4, 10, 3, 1, 0,
					-- layer=2 filter=155 channel=54
					-5, -3, -12, -1, 2, -9, -11, -3, -6,
					-- layer=2 filter=155 channel=55
					8, -8, -6, 10, 3, -4, -2, -11, 2,
					-- layer=2 filter=155 channel=56
					-8, 6, 4, 1, 3, -1, -7, -13, -3,
					-- layer=2 filter=155 channel=57
					6, -9, -2, 7, -8, -1, 9, 11, -1,
					-- layer=2 filter=155 channel=58
					0, -2, 2, -6, -7, 0, -2, -4, -2,
					-- layer=2 filter=155 channel=59
					8, 4, 5, 0, 0, -9, -9, 0, -12,
					-- layer=2 filter=155 channel=60
					-4, 0, -10, 0, 4, -6, -4, 2, -11,
					-- layer=2 filter=155 channel=61
					-13, -5, -13, -7, 0, -13, -10, 1, -10,
					-- layer=2 filter=155 channel=62
					-4, 0, -1, 6, 2, -2, -12, -9, -3,
					-- layer=2 filter=155 channel=63
					2, 8, -6, 1, 1, 1, 0, 6, 0,
					-- layer=2 filter=155 channel=64
					8, -1, 6, -1, 9, 2, 2, -10, -5,
					-- layer=2 filter=155 channel=65
					-8, -10, 9, -2, 3, 10, -3, -8, 0,
					-- layer=2 filter=155 channel=66
					11, 7, 2, 0, -3, 9, 5, 9, -5,
					-- layer=2 filter=155 channel=67
					-8, -6, 6, -2, 0, -7, 4, -1, 0,
					-- layer=2 filter=155 channel=68
					9, 11, 1, 0, -4, -4, 10, -4, -8,
					-- layer=2 filter=155 channel=69
					5, 0, -1, -5, 4, -8, -10, -10, 6,
					-- layer=2 filter=155 channel=70
					-6, 1, -12, -8, -7, -8, 5, 2, -11,
					-- layer=2 filter=155 channel=71
					2, 4, -3, 1, 2, -6, -6, -1, 8,
					-- layer=2 filter=155 channel=72
					5, 5, 1, -4, -14, -15, -11, -4, 0,
					-- layer=2 filter=155 channel=73
					-15, -3, -6, -12, -8, -9, -16, 1, -8,
					-- layer=2 filter=155 channel=74
					-11, -10, 4, -1, -5, -7, 1, 2, 5,
					-- layer=2 filter=155 channel=75
					3, -12, 0, 9, 8, 6, 3, 0, -3,
					-- layer=2 filter=155 channel=76
					-9, -1, 3, 1, -15, -7, -6, -6, 2,
					-- layer=2 filter=155 channel=77
					-3, -1, 0, 0, 1, 4, 7, -2, 2,
					-- layer=2 filter=155 channel=78
					0, 6, -11, -11, 4, -9, 9, 6, -8,
					-- layer=2 filter=155 channel=79
					-3, 10, -2, 1, -2, 7, 10, -2, 3,
					-- layer=2 filter=155 channel=80
					1, 5, 2, 1, 3, 0, -7, 1, -4,
					-- layer=2 filter=155 channel=81
					-9, 11, 0, 4, -5, 5, 5, 3, 1,
					-- layer=2 filter=155 channel=82
					-3, -7, 6, 10, -8, 10, 9, 9, 6,
					-- layer=2 filter=155 channel=83
					-10, -4, 6, -6, -7, -6, 9, -1, -6,
					-- layer=2 filter=155 channel=84
					2, -11, -9, -3, 0, -1, -6, 4, 5,
					-- layer=2 filter=155 channel=85
					6, 8, 5, 5, 7, 5, -8, 1, 5,
					-- layer=2 filter=155 channel=86
					5, 8, -6, 7, -6, -7, -1, 2, 2,
					-- layer=2 filter=155 channel=87
					5, -4, -10, 0, -7, -11, -4, 1, -3,
					-- layer=2 filter=155 channel=88
					-6, -3, 3, 6, -4, -5, -5, 1, -7,
					-- layer=2 filter=155 channel=89
					1, 0, -1, -6, -10, -2, -5, 0, 1,
					-- layer=2 filter=155 channel=90
					4, -3, 2, 10, -5, 7, -3, 9, -10,
					-- layer=2 filter=155 channel=91
					-6, -6, 1, -13, 0, -12, -4, 4, 2,
					-- layer=2 filter=155 channel=92
					-14, 5, -3, 0, 11, 0, -4, -18, -9,
					-- layer=2 filter=155 channel=93
					-10, 2, -1, 1, -6, 1, -6, -5, -7,
					-- layer=2 filter=155 channel=94
					-6, -21, -3, -17, -9, -6, -18, 0, -6,
					-- layer=2 filter=155 channel=95
					2, -10, 5, 1, 6, -4, -4, -10, 4,
					-- layer=2 filter=155 channel=96
					-13, -4, 0, -3, -3, 6, -3, -3, -10,
					-- layer=2 filter=155 channel=97
					8, -1, -11, -4, -2, 7, -7, -11, 1,
					-- layer=2 filter=155 channel=98
					-4, -4, -12, -4, -18, -7, -3, -8, -18,
					-- layer=2 filter=155 channel=99
					6, -6, 3, -2, -2, 3, -11, 3, -1,
					-- layer=2 filter=155 channel=100
					2, -3, 6, -7, 10, 6, 1, 0, -3,
					-- layer=2 filter=155 channel=101
					0, 3, -7, 5, -13, 7, -1, 5, -10,
					-- layer=2 filter=155 channel=102
					-8, -9, -7, 0, 2, 0, -6, -6, 5,
					-- layer=2 filter=155 channel=103
					3, -9, 0, 9, 5, 5, 2, 5, -5,
					-- layer=2 filter=155 channel=104
					-1, -2, -9, 2, -16, 7, -10, 2, 4,
					-- layer=2 filter=155 channel=105
					0, -6, -6, -8, 7, 0, -2, 0, 1,
					-- layer=2 filter=155 channel=106
					-10, 2, 2, 1, -3, 6, -1, 4, -5,
					-- layer=2 filter=155 channel=107
					-3, -2, 5, -5, 3, 0, 5, 1, -8,
					-- layer=2 filter=155 channel=108
					1, -1, -3, 0, -4, -8, -4, 1, 4,
					-- layer=2 filter=155 channel=109
					8, 11, -1, 10, 0, 0, -1, 1, 10,
					-- layer=2 filter=155 channel=110
					-8, 7, -6, -11, -9, -7, 1, -5, -3,
					-- layer=2 filter=155 channel=111
					0, 2, -6, 0, 7, 3, 9, 0, -9,
					-- layer=2 filter=155 channel=112
					7, 6, 8, -7, -9, 0, -7, -9, 7,
					-- layer=2 filter=155 channel=113
					-6, 7, 5, -10, 4, 0, -9, 7, 5,
					-- layer=2 filter=155 channel=114
					-1, 6, -7, -7, 2, -7, 0, -1, -3,
					-- layer=2 filter=155 channel=115
					-4, -1, 6, 9, 5, 1, 1, -2, -9,
					-- layer=2 filter=155 channel=116
					-6, -2, 5, -6, -13, -6, 6, -7, 6,
					-- layer=2 filter=155 channel=117
					-10, -14, -10, -6, -3, 2, -10, 1, 5,
					-- layer=2 filter=155 channel=118
					4, 1, 0, 0, 3, -12, 1, -5, -10,
					-- layer=2 filter=155 channel=119
					6, 0, -13, 2, 6, -8, -6, 4, -8,
					-- layer=2 filter=155 channel=120
					-10, -3, -7, 7, -3, 0, 0, 2, 2,
					-- layer=2 filter=155 channel=121
					8, 0, -12, 7, 9, -7, 4, 1, 8,
					-- layer=2 filter=155 channel=122
					-3, 1, 11, -3, -4, 5, 5, 6, 9,
					-- layer=2 filter=155 channel=123
					-14, 7, -9, 3, -11, 2, -10, -6, -14,
					-- layer=2 filter=155 channel=124
					-14, 0, -17, -11, 0, -7, 1, 1, -6,
					-- layer=2 filter=155 channel=125
					-7, 7, 7, 8, 0, 2, 5, -4, 5,
					-- layer=2 filter=155 channel=126
					9, 10, -5, 3, 0, 9, -2, -2, 10,
					-- layer=2 filter=155 channel=127
					7, -12, -13, -7, -3, 7, -4, -11, -9,
					-- layer=2 filter=156 channel=0
					1, 9, 5, -11, 3, -37, 16, 21, 21,
					-- layer=2 filter=156 channel=1
					-36, -18, -13, 39, 2, -26, 2, -38, -14,
					-- layer=2 filter=156 channel=2
					-4, -7, 9, 9, -10, -5, 7, 7, 5,
					-- layer=2 filter=156 channel=3
					0, -3, -9, -4, -9, 18, 17, 9, -17,
					-- layer=2 filter=156 channel=4
					-5, -16, 0, -3, 8, -14, 19, 17, 8,
					-- layer=2 filter=156 channel=5
					19, -16, -18, -10, -2, -35, -31, 4, -4,
					-- layer=2 filter=156 channel=6
					-37, 12, 17, -27, 21, 24, -38, -44, 44,
					-- layer=2 filter=156 channel=7
					-7, -12, -39, 41, -22, -68, -18, -41, -12,
					-- layer=2 filter=156 channel=8
					-3, -6, 1, -1, -8, -3, 2, -9, -1,
					-- layer=2 filter=156 channel=9
					-28, -8, 11, -8, 17, -1, -30, -28, 1,
					-- layer=2 filter=156 channel=10
					12, 16, 14, 26, -6, 5, 30, 24, 27,
					-- layer=2 filter=156 channel=11
					23, 14, 20, -15, 4, -4, -16, 20, 0,
					-- layer=2 filter=156 channel=12
					-8, 5, -16, 40, -3, -12, 8, -17, -31,
					-- layer=2 filter=156 channel=13
					-9, 8, -8, 9, -4, 4, -6, 8, -1,
					-- layer=2 filter=156 channel=14
					14, 8, 13, 54, 19, 2, 40, -11, -50,
					-- layer=2 filter=156 channel=15
					0, 25, -32, 49, 30, -28, 17, 72, -18,
					-- layer=2 filter=156 channel=16
					-31, 14, -2, -4, 1, -4, -4, 3, -2,
					-- layer=2 filter=156 channel=17
					7, -1, 8, 4, -3, -10, -6, 2, -5,
					-- layer=2 filter=156 channel=18
					49, 15, 13, 10, 30, -3, 14, 30, 14,
					-- layer=2 filter=156 channel=19
					-37, -22, -35, 7, -31, -17, -7, -41, -31,
					-- layer=2 filter=156 channel=20
					-10, 1, 8, -4, 0, 2, 4, 1, -1,
					-- layer=2 filter=156 channel=21
					7, 13, 25, 0, 5, 5, 6, 10, 0,
					-- layer=2 filter=156 channel=22
					9, 8, -7, -3, 0, -3, 9, -12, 2,
					-- layer=2 filter=156 channel=23
					-2, -1, 15, -5, -1, 6, -48, -2, -26,
					-- layer=2 filter=156 channel=24
					24, 15, 48, -34, -14, 16, -19, 3, 15,
					-- layer=2 filter=156 channel=25
					31, 31, 18, -14, 0, 12, 5, 11, 24,
					-- layer=2 filter=156 channel=26
					0, -3, -1, 5, -10, 0, -7, 3, 7,
					-- layer=2 filter=156 channel=27
					-8, -26, -15, 13, 8, 24, 24, -11, 16,
					-- layer=2 filter=156 channel=28
					47, -25, -41, 55, -34, -56, 50, 13, -40,
					-- layer=2 filter=156 channel=29
					10, 7, -4, -10, -2, 7, 0, 0, -8,
					-- layer=2 filter=156 channel=30
					20, -2, 11, 15, 6, 8, 15, 46, -8,
					-- layer=2 filter=156 channel=31
					39, -4, -28, 9, -9, -30, -50, 77, -22,
					-- layer=2 filter=156 channel=32
					-1, 12, -2, -7, -11, 9, 1, -9, -8,
					-- layer=2 filter=156 channel=33
					47, 14, -26, 65, 2, 1, 66, 14, -19,
					-- layer=2 filter=156 channel=34
					-30, -7, 6, 19, 33, 9, -2, 0, 15,
					-- layer=2 filter=156 channel=35
					-3, 1, -49, 102, 30, -49, 55, 6, 12,
					-- layer=2 filter=156 channel=36
					5, -5, 10, -9, 0, 3, 3, -6, 3,
					-- layer=2 filter=156 channel=37
					19, -9, -11, -6, 7, 4, -24, 8, 2,
					-- layer=2 filter=156 channel=38
					-7, 2, -5, 33, 24, 36, 3, -25, -11,
					-- layer=2 filter=156 channel=39
					36, 21, 23, 8, 22, 39, 32, -29, -22,
					-- layer=2 filter=156 channel=40
					-7, -17, -26, -32, 11, 3, -17, 50, 1,
					-- layer=2 filter=156 channel=41
					-7, -8, 4, 6, 7, 3, 1, 0, -11,
					-- layer=2 filter=156 channel=42
					3, 31, 8, 34, 30, -13, -1, 20, 21,
					-- layer=2 filter=156 channel=43
					54, -11, -65, -21, 0, -19, 16, 36, 1,
					-- layer=2 filter=156 channel=44
					2, -3, 3, 5, 8, -8, 11, 1, -1,
					-- layer=2 filter=156 channel=45
					22, 9, -8, 35, -37, -10, 35, 0, -3,
					-- layer=2 filter=156 channel=46
					16, -1, -27, -5, -17, -26, 55, 31, 8,
					-- layer=2 filter=156 channel=47
					48, 2, -34, 26, -13, -31, 62, 1, -42,
					-- layer=2 filter=156 channel=48
					-12, -8, -1, 3, -8, -4, -3, 2, -7,
					-- layer=2 filter=156 channel=49
					46, 23, 51, 14, 17, 6, -23, 13, 50,
					-- layer=2 filter=156 channel=50
					8, -6, 2, -5, 5, -7, -8, 17, -2,
					-- layer=2 filter=156 channel=51
					0, 9, 22, -16, 11, 0, 0, 19, -2,
					-- layer=2 filter=156 channel=52
					-20, 24, 0, -7, 8, -1, -47, -19, -31,
					-- layer=2 filter=156 channel=53
					50, 23, 6, -31, -14, 27, -24, -1, 12,
					-- layer=2 filter=156 channel=54
					16, 17, -7, 12, -9, -30, -12, -3, 12,
					-- layer=2 filter=156 channel=55
					12, 5, -1, 5, 10, -7, -13, 13, -4,
					-- layer=2 filter=156 channel=56
					29, -3, -11, -15, 8, 2, -2, 4, -2,
					-- layer=2 filter=156 channel=57
					8, 12, 5, 0, 0, 7, 6, -5, 8,
					-- layer=2 filter=156 channel=58
					-10, 6, -3, 59, 3, 11, -8, -7, -72,
					-- layer=2 filter=156 channel=59
					-6, 10, -23, 2, 11, 32, 26, 21, -31,
					-- layer=2 filter=156 channel=60
					-51, 0, -14, 4, 16, 17, -8, -32, -3,
					-- layer=2 filter=156 channel=61
					-27, -11, 20, -34, 6, -5, -22, 10, 28,
					-- layer=2 filter=156 channel=62
					-7, 0, 18, 12, -2, -9, -41, -19, 31,
					-- layer=2 filter=156 channel=63
					-11, -2, 10, -5, -3, 16, -15, -15, 11,
					-- layer=2 filter=156 channel=64
					-14, 0, 58, -7, 1, 37, -45, 9, 26,
					-- layer=2 filter=156 channel=65
					-44, -23, 14, -57, -10, -7, -41, -38, 27,
					-- layer=2 filter=156 channel=66
					1, -5, -15, 9, -15, -38, 8, -2, -58,
					-- layer=2 filter=156 channel=67
					-12, -16, -29, -26, -56, -16, -14, -15, 2,
					-- layer=2 filter=156 channel=68
					1, -5, 10, 4, -1, -9, -4, 4, 8,
					-- layer=2 filter=156 channel=69
					-30, -5, 18, 21, 22, 18, -10, 25, 21,
					-- layer=2 filter=156 channel=70
					16, 5, -45, 52, -7, -48, 37, 9, -23,
					-- layer=2 filter=156 channel=71
					-12, -17, 9, -5, 28, 54, 13, -4, -7,
					-- layer=2 filter=156 channel=72
					-22, -26, -19, 11, -4, -3, 42, -14, -49,
					-- layer=2 filter=156 channel=73
					3, 23, -47, 32, -11, -32, 49, 26, 0,
					-- layer=2 filter=156 channel=74
					-3, -15, -15, 43, -27, -26, 36, 24, 14,
					-- layer=2 filter=156 channel=75
					24, -20, 50, 12, -9, 12, -27, -10, -38,
					-- layer=2 filter=156 channel=76
					1, 14, -99, -18, 6, -60, -72, 17, -61,
					-- layer=2 filter=156 channel=77
					0, -3, 9, 1, 11, 0, 6, 11, 0,
					-- layer=2 filter=156 channel=78
					29, 34, 22, -11, -7, 17, -76, -13, 10,
					-- layer=2 filter=156 channel=79
					3, 11, -2, 6, -6, -6, 0, -2, -1,
					-- layer=2 filter=156 channel=80
					1, -6, -3, 24, -5, 14, 34, 11, 9,
					-- layer=2 filter=156 channel=81
					-13, -9, 0, 15, -7, -6, 6, 5, 4,
					-- layer=2 filter=156 channel=82
					5, 3, -11, -7, -5, 8, 3, 1, 7,
					-- layer=2 filter=156 channel=83
					34, -3, -3, 25, 3, 2, -14, -3, 5,
					-- layer=2 filter=156 channel=84
					1, 7, 4, 5, -8, -5, -11, 8, 7,
					-- layer=2 filter=156 channel=85
					11, -9, -11, 10, 8, -5, 5, -3, -13,
					-- layer=2 filter=156 channel=86
					10, -5, -3, 0, -17, 0, 21, -6, 1,
					-- layer=2 filter=156 channel=87
					-1, 12, -35, -19, 46, -4, -17, 34, 13,
					-- layer=2 filter=156 channel=88
					1, -33, -15, 40, 4, 3, 28, 12, 0,
					-- layer=2 filter=156 channel=89
					-18, 2, -29, 62, 16, 9, 64, 1, -57,
					-- layer=2 filter=156 channel=90
					-1, -7, -3, -1, -7, -5, 5, -2, 0,
					-- layer=2 filter=156 channel=91
					0, 0, -23, 64, -7, -11, 15, -9, -12,
					-- layer=2 filter=156 channel=92
					-18, -14, -31, 60, 8, -2, 44, -15, -4,
					-- layer=2 filter=156 channel=93
					35, 20, -29, 43, -6, -26, 12, -21, 35,
					-- layer=2 filter=156 channel=94
					-76, -31, 1, -103, 22, 15, -25, -38, -2,
					-- layer=2 filter=156 channel=95
					9, 16, 25, 3, 17, 3, -17, 5, -5,
					-- layer=2 filter=156 channel=96
					-89, 5, -4, -96, 6, 60, -65, -35, 11,
					-- layer=2 filter=156 channel=97
					-6, -12, 20, 13, 62, 69, -7, -7, 35,
					-- layer=2 filter=156 channel=98
					13, -15, -53, 58, -27, -50, 48, -11, -26,
					-- layer=2 filter=156 channel=99
					-17, 2, -47, -5, 4, -58, -35, -19, 12,
					-- layer=2 filter=156 channel=100
					13, 8, -16, 14, -3, 24, -31, 9, 17,
					-- layer=2 filter=156 channel=101
					32, 19, -39, 29, 32, 24, 18, 15, 6,
					-- layer=2 filter=156 channel=102
					-63, 17, 11, -18, 27, 10, -22, -27, -17,
					-- layer=2 filter=156 channel=103
					14, -4, 25, 11, -43, -11, -33, 4, 66,
					-- layer=2 filter=156 channel=104
					27, -17, 0, -3, 7, 2, -52, 5, -5,
					-- layer=2 filter=156 channel=105
					-47, -70, -58, -23, 20, -36, -33, 11, 21,
					-- layer=2 filter=156 channel=106
					0, -4, -11, 7, 15, 0, 16, 33, -23,
					-- layer=2 filter=156 channel=107
					9, 40, -28, -4, 15, -2, 8, -14, 20,
					-- layer=2 filter=156 channel=108
					-24, -1, 3, 9, 3, 25, -11, -49, -28,
					-- layer=2 filter=156 channel=109
					-6, -13, -1, 5, -5, -7, 8, 8, 20,
					-- layer=2 filter=156 channel=110
					3, -13, 61, -4, -22, 15, -15, -18, 3,
					-- layer=2 filter=156 channel=111
					3, -10, -8, 12, 8, 8, 3, -8, -7,
					-- layer=2 filter=156 channel=112
					-18, -10, 0, -1, 27, -12, 0, -1, 7,
					-- layer=2 filter=156 channel=113
					18, -6, 50, 5, -26, 7, -21, 8, -20,
					-- layer=2 filter=156 channel=114
					3, -5, 10, -11, 11, 8, 1, -14, -12,
					-- layer=2 filter=156 channel=115
					4, -6, -4, 0, -3, -3, 0, -1, 11,
					-- layer=2 filter=156 channel=116
					-19, -9, -25, 2, 46, -10, -61, -5, -12,
					-- layer=2 filter=156 channel=117
					-38, 61, -15, 21, -22, -33, 17, -43, -2,
					-- layer=2 filter=156 channel=118
					11, -8, -10, -14, -2, 14, -3, 27, 28,
					-- layer=2 filter=156 channel=119
					30, -7, -16, 22, -7, -16, 31, 15, -19,
					-- layer=2 filter=156 channel=120
					-9, -2, 7, -9, 8, -6, 7, 8, 4,
					-- layer=2 filter=156 channel=121
					-2, 4, -3, -7, -2, -7, -2, 5, -9,
					-- layer=2 filter=156 channel=122
					1, 9, -6, 1, 0, 3, -7, 10, 16,
					-- layer=2 filter=156 channel=123
					-35, -30, -12, -19, -23, -58, -3, -19, -49,
					-- layer=2 filter=156 channel=124
					17, 12, 13, 57, 13, -74, -11, 64, 26,
					-- layer=2 filter=156 channel=125
					-7, -5, -4, 5, 0, 0, 6, 4, -3,
					-- layer=2 filter=156 channel=126
					-72, 7, 22, -24, 50, -11, 80, 13, 29,
					-- layer=2 filter=156 channel=127
					-26, -27, 7, 1, -16, 5, -29, -39, -34,
					-- layer=2 filter=157 channel=0
					-7, -3, 3, -5, -4, -10, -7, 1, -5,
					-- layer=2 filter=157 channel=1
					-3, -2, -7, -6, 0, -9, 0, -4, 2,
					-- layer=2 filter=157 channel=2
					-2, 6, -4, 0, -6, -2, 4, -10, 1,
					-- layer=2 filter=157 channel=3
					0, -1, -12, -1, -9, 4, -4, 7, -2,
					-- layer=2 filter=157 channel=4
					2, -12, -5, -6, -8, -10, -11, -1, -5,
					-- layer=2 filter=157 channel=5
					-9, 3, 0, -7, -2, 5, -3, 1, 4,
					-- layer=2 filter=157 channel=6
					-1, -9, -5, 4, -5, 8, -2, 3, -7,
					-- layer=2 filter=157 channel=7
					-7, 2, 2, -6, 7, 0, 1, -13, 10,
					-- layer=2 filter=157 channel=8
					1, 9, 0, 10, 11, -6, 7, 5, 6,
					-- layer=2 filter=157 channel=9
					0, 0, 8, -8, 0, -7, -10, 8, -10,
					-- layer=2 filter=157 channel=10
					-10, -11, -5, -10, -2, -6, -7, -3, 0,
					-- layer=2 filter=157 channel=11
					-5, -5, 5, 2, -12, 0, 1, -16, 7,
					-- layer=2 filter=157 channel=12
					-9, -16, -9, 2, -11, -9, -6, -3, 0,
					-- layer=2 filter=157 channel=13
					3, 8, -9, -7, 7, 7, 0, 2, -2,
					-- layer=2 filter=157 channel=14
					-8, 4, -4, 0, -3, -12, -3, -6, -6,
					-- layer=2 filter=157 channel=15
					8, -1, 5, 5, -4, -10, -5, -4, -7,
					-- layer=2 filter=157 channel=16
					-11, -1, 4, -2, -11, -8, -2, -11, 9,
					-- layer=2 filter=157 channel=17
					-2, -3, 9, 5, -7, -1, 3, -6, -9,
					-- layer=2 filter=157 channel=18
					-8, -4, 5, 3, 5, -12, -9, 1, 0,
					-- layer=2 filter=157 channel=19
					-6, -15, 6, 0, 3, -6, -12, -10, 2,
					-- layer=2 filter=157 channel=20
					3, -7, 4, -9, 0, -4, -11, -3, -11,
					-- layer=2 filter=157 channel=21
					-2, -7, -7, 4, -5, -9, -4, 11, -4,
					-- layer=2 filter=157 channel=22
					2, -3, -6, -11, -6, 0, -9, -7, -3,
					-- layer=2 filter=157 channel=23
					-12, -6, -6, 5, 3, 0, 2, -2, 5,
					-- layer=2 filter=157 channel=24
					-11, 6, -7, 7, -9, -7, -12, 6, -10,
					-- layer=2 filter=157 channel=25
					-2, -1, -10, -12, 1, -10, -5, -12, -8,
					-- layer=2 filter=157 channel=26
					-4, -4, 5, 3, -9, -7, 8, -4, 4,
					-- layer=2 filter=157 channel=27
					6, 2, 0, -6, -4, -2, -8, 6, 1,
					-- layer=2 filter=157 channel=28
					1, 0, 6, -15, 2, 2, -7, 10, -4,
					-- layer=2 filter=157 channel=29
					-6, 1, -7, -8, -7, 6, -1, -1, 5,
					-- layer=2 filter=157 channel=30
					-10, 9, -2, -1, 3, -11, -4, -6, -3,
					-- layer=2 filter=157 channel=31
					3, -9, -11, 8, -2, 1, -1, -2, 4,
					-- layer=2 filter=157 channel=32
					-1, 5, 6, 0, -5, 0, 0, 6, 8,
					-- layer=2 filter=157 channel=33
					-4, -6, -2, -8, -8, 3, -4, 3, 12,
					-- layer=2 filter=157 channel=34
					6, -9, 8, -7, -9, 3, -5, 0, -9,
					-- layer=2 filter=157 channel=35
					-9, 0, -12, 0, -7, 6, -10, -18, -7,
					-- layer=2 filter=157 channel=36
					5, 2, -11, 11, 5, -2, -2, 6, -11,
					-- layer=2 filter=157 channel=37
					-5, -6, 3, -8, -9, -8, 4, 4, 0,
					-- layer=2 filter=157 channel=38
					-8, 0, -11, 0, -6, 1, -9, -4, -8,
					-- layer=2 filter=157 channel=39
					3, 0, 2, -3, 4, 5, -8, 0, 7,
					-- layer=2 filter=157 channel=40
					0, -9, 8, 7, -10, 0, 10, -5, 0,
					-- layer=2 filter=157 channel=41
					-9, -10, -3, -5, 9, 2, 2, -4, 9,
					-- layer=2 filter=157 channel=42
					8, 7, -2, 0, -14, -15, -4, 0, -1,
					-- layer=2 filter=157 channel=43
					0, 0, 3, -7, 0, -3, -10, -11, 3,
					-- layer=2 filter=157 channel=44
					-3, -3, -9, -6, 9, -1, 7, 0, 6,
					-- layer=2 filter=157 channel=45
					7, -10, -10, 0, -2, -6, 7, -6, -5,
					-- layer=2 filter=157 channel=46
					2, 0, -1, 8, -1, -10, 5, 6, -4,
					-- layer=2 filter=157 channel=47
					-5, 1, 9, 5, -7, 5, -2, -5, 3,
					-- layer=2 filter=157 channel=48
					9, -6, 0, -3, 9, -4, 5, -8, 3,
					-- layer=2 filter=157 channel=49
					-11, 6, -5, 4, 1, 6, 6, 2, 0,
					-- layer=2 filter=157 channel=50
					4, 2, 1, -6, 4, -5, -4, 7, -5,
					-- layer=2 filter=157 channel=51
					-14, -5, -6, -1, -13, -1, 1, -14, -15,
					-- layer=2 filter=157 channel=52
					-15, -5, -7, 3, -12, -6, -12, 5, -2,
					-- layer=2 filter=157 channel=53
					1, 3, 7, -5, 11, -8, 4, -4, 4,
					-- layer=2 filter=157 channel=54
					-12, -10, 6, -14, -4, -2, -12, -16, -14,
					-- layer=2 filter=157 channel=55
					-1, 8, 8, -7, 6, -6, 9, 7, -11,
					-- layer=2 filter=157 channel=56
					0, -13, -5, -6, -4, 3, -5, -7, -14,
					-- layer=2 filter=157 channel=57
					9, 10, 10, -7, 11, -1, 10, -4, 3,
					-- layer=2 filter=157 channel=58
					5, -7, -9, -9, -6, -16, 0, 5, -7,
					-- layer=2 filter=157 channel=59
					-4, 2, 5, -5, -1, -5, -3, 1, 10,
					-- layer=2 filter=157 channel=60
					-7, -6, -11, 0, 0, -1, -4, -13, -6,
					-- layer=2 filter=157 channel=61
					-13, 3, 3, -11, -6, -1, 3, 4, -4,
					-- layer=2 filter=157 channel=62
					6, 5, -7, -10, 1, -5, 1, -11, -8,
					-- layer=2 filter=157 channel=63
					-14, -4, 7, -12, -7, -1, 1, -10, -10,
					-- layer=2 filter=157 channel=64
					-1, -4, -1, -12, -5, 1, 2, -5, 1,
					-- layer=2 filter=157 channel=65
					-2, -7, 4, -2, 6, -1, -6, 4, -1,
					-- layer=2 filter=157 channel=66
					-7, 5, 4, 1, 6, 0, -6, 6, -8,
					-- layer=2 filter=157 channel=67
					-7, -10, 1, -4, -5, -1, -3, -11, -5,
					-- layer=2 filter=157 channel=68
					7, 0, 6, 8, -10, -11, -5, 6, 4,
					-- layer=2 filter=157 channel=69
					-10, 0, -5, -8, 5, 2, 11, 0, -2,
					-- layer=2 filter=157 channel=70
					-6, 5, -6, -6, 0, -15, -5, -19, -7,
					-- layer=2 filter=157 channel=71
					-8, 0, 0, 5, -2, 6, 3, 0, -2,
					-- layer=2 filter=157 channel=72
					-5, -7, 3, -7, -11, -5, 3, -3, 13,
					-- layer=2 filter=157 channel=73
					-3, -8, 3, -5, -9, 7, 5, 2, -11,
					-- layer=2 filter=157 channel=74
					7, 7, -4, 7, 8, 4, -6, 0, -2,
					-- layer=2 filter=157 channel=75
					-6, 2, 5, 8, 7, 7, -5, 6, 1,
					-- layer=2 filter=157 channel=76
					8, 7, 8, 0, -7, 1, 4, -6, 0,
					-- layer=2 filter=157 channel=77
					2, -5, -2, 0, 0, 3, 0, 1, -2,
					-- layer=2 filter=157 channel=78
					8, 3, 6, 0, 8, 7, -4, -6, 5,
					-- layer=2 filter=157 channel=79
					6, 0, 2, 0, -1, -5, 0, -12, -8,
					-- layer=2 filter=157 channel=80
					-10, -3, -4, -7, 3, -2, -3, -3, 7,
					-- layer=2 filter=157 channel=81
					3, 0, -7, 1, -8, -9, -11, -5, 0,
					-- layer=2 filter=157 channel=82
					-11, -2, -10, -6, -10, 1, -8, -9, 10,
					-- layer=2 filter=157 channel=83
					7, 5, -4, 9, -10, -11, -7, 8, -7,
					-- layer=2 filter=157 channel=84
					4, -9, 1, 9, -4, -4, -8, 4, 3,
					-- layer=2 filter=157 channel=85
					10, 2, -5, -2, 0, 7, 4, -7, -7,
					-- layer=2 filter=157 channel=86
					-7, 5, -8, 7, 10, 2, 9, 9, -4,
					-- layer=2 filter=157 channel=87
					-1, 2, -7, -9, 0, -1, -10, -10, 0,
					-- layer=2 filter=157 channel=88
					-2, 3, -15, -6, 0, 2, -9, -8, -5,
					-- layer=2 filter=157 channel=89
					-8, -11, -1, -15, -18, -1, -8, -6, -7,
					-- layer=2 filter=157 channel=90
					3, -3, 8, 5, 6, 2, -1, 0, 4,
					-- layer=2 filter=157 channel=91
					-15, -12, 0, -13, -4, -11, 6, 5, -5,
					-- layer=2 filter=157 channel=92
					-3, -10, 4, -2, -9, -4, -1, -12, 0,
					-- layer=2 filter=157 channel=93
					4, -3, -3, 7, -9, -11, -6, 2, 5,
					-- layer=2 filter=157 channel=94
					-4, -12, 1, -3, -3, 9, 2, -1, -13,
					-- layer=2 filter=157 channel=95
					-9, -5, -10, 0, -5, 0, -6, -10, -6,
					-- layer=2 filter=157 channel=96
					3, 3, 6, -3, -3, -4, -1, 7, -5,
					-- layer=2 filter=157 channel=97
					4, -10, 7, 1, 0, 3, 2, 7, -7,
					-- layer=2 filter=157 channel=98
					4, 1, 0, -15, -4, -13, -15, -12, -4,
					-- layer=2 filter=157 channel=99
					-4, 3, -15, -7, -6, 2, -7, -5, -5,
					-- layer=2 filter=157 channel=100
					-5, -9, 1, -3, 2, -10, -10, -3, -7,
					-- layer=2 filter=157 channel=101
					-5, 5, -12, 0, 0, -6, -7, -2, -11,
					-- layer=2 filter=157 channel=102
					-13, 0, -1, 7, 6, 0, -9, -8, -2,
					-- layer=2 filter=157 channel=103
					-10, -4, -10, 1, 0, 3, 6, -9, -4,
					-- layer=2 filter=157 channel=104
					0, 0, 6, 4, -12, 7, -8, 1, 2,
					-- layer=2 filter=157 channel=105
					-6, -9, -8, -9, -7, 0, -9, 1, 6,
					-- layer=2 filter=157 channel=106
					4, 3, -7, -11, -3, -19, 8, -13, 1,
					-- layer=2 filter=157 channel=107
					-5, 8, -1, 0, -1, 0, 7, 1, -6,
					-- layer=2 filter=157 channel=108
					-2, -2, 5, -11, 7, 5, 2, -6, 1,
					-- layer=2 filter=157 channel=109
					-9, 0, 2, 4, -3, -1, -7, 1, -7,
					-- layer=2 filter=157 channel=110
					-8, -10, -9, 6, 1, -6, -7, 7, 0,
					-- layer=2 filter=157 channel=111
					-8, -8, 0, 3, -2, -8, 9, 0, 0,
					-- layer=2 filter=157 channel=112
					-11, -6, -1, 0, 4, -1, -12, -16, -7,
					-- layer=2 filter=157 channel=113
					0, -1, -9, -4, 7, -7, -12, -2, -7,
					-- layer=2 filter=157 channel=114
					4, 0, -8, 6, 0, -8, -3, -10, -4,
					-- layer=2 filter=157 channel=115
					5, 7, 4, 4, 3, 10, 9, 2, -3,
					-- layer=2 filter=157 channel=116
					7, -4, 12, -4, -8, -14, 7, -14, 0,
					-- layer=2 filter=157 channel=117
					7, -2, 4, -19, 3, 3, -12, 1, 2,
					-- layer=2 filter=157 channel=118
					0, -10, 3, 1, -4, 5, -9, -5, -1,
					-- layer=2 filter=157 channel=119
					-4, 6, -5, -5, -7, 7, -4, -7, 0,
					-- layer=2 filter=157 channel=120
					-7, 1, -1, 3, -8, -3, -3, 5, -2,
					-- layer=2 filter=157 channel=121
					-3, -1, -1, -11, 5, 8, 7, 9, 4,
					-- layer=2 filter=157 channel=122
					-5, -2, -2, -7, -1, 2, -9, 7, 0,
					-- layer=2 filter=157 channel=123
					4, -3, 4, 1, -7, -7, 1, -8, 6,
					-- layer=2 filter=157 channel=124
					0, 5, -5, 0, 7, -11, 11, 9, 12,
					-- layer=2 filter=157 channel=125
					-4, 9, -5, -4, -6, 0, 1, -5, -1,
					-- layer=2 filter=157 channel=126
					0, 1, 4, 3, -11, -5, 0, 8, -5,
					-- layer=2 filter=157 channel=127
					-3, 1, -6, -11, 3, 0, 1, -4, -3,
					-- layer=2 filter=158 channel=0
					15, 39, 14, 6, -33, -21, 33, 31, 27,
					-- layer=2 filter=158 channel=1
					38, -20, 6, 21, 44, 37, -3, -31, -31,
					-- layer=2 filter=158 channel=2
					-2, -2, 6, 0, -5, -6, -6, -4, 10,
					-- layer=2 filter=158 channel=3
					11, -23, -5, -3, -26, -33, 57, 22, 6,
					-- layer=2 filter=158 channel=4
					29, 3, 16, 0, -24, -9, -22, 3, -12,
					-- layer=2 filter=158 channel=5
					30, 36, 0, 14, -21, -43, 28, 10, -21,
					-- layer=2 filter=158 channel=6
					-10, -1, -3, -74, -62, -2, -72, 2, -31,
					-- layer=2 filter=158 channel=7
					19, 6, 39, 42, 66, 17, 21, -27, -37,
					-- layer=2 filter=158 channel=8
					4, 1, -1, 7, -5, -6, -4, 1, 6,
					-- layer=2 filter=158 channel=9
					-23, -27, 5, -73, -39, -49, 8, -13, -26,
					-- layer=2 filter=158 channel=10
					16, -10, 9, 6, -32, -59, 40, 32, 28,
					-- layer=2 filter=158 channel=11
					37, 11, 0, 7, 0, -22, -5, 17, -7,
					-- layer=2 filter=158 channel=12
					32, 1, 12, 51, 62, 63, -15, -99, -91,
					-- layer=2 filter=158 channel=13
					-5, -1, 2, -9, 7, 6, 0, -2, 4,
					-- layer=2 filter=158 channel=14
					27, 8, -3, 12, 33, 36, -19, -48, -72,
					-- layer=2 filter=158 channel=15
					15, -4, -43, 15, 37, 19, 23, 33, 25,
					-- layer=2 filter=158 channel=16
					24, 18, 8, 12, 5, -13, 0, 1, 9,
					-- layer=2 filter=158 channel=17
					-8, 10, -4, -3, -7, -4, 1, -3, 2,
					-- layer=2 filter=158 channel=18
					36, -13, -33, -23, -3, 0, -48, 48, 22,
					-- layer=2 filter=158 channel=19
					18, 22, 29, -8, -11, -7, 20, 15, -20,
					-- layer=2 filter=158 channel=20
					4, 0, 4, -8, -7, 0, 0, 1, 4,
					-- layer=2 filter=158 channel=21
					17, 2, 1, 8, 3, 9, 14, 10, 17,
					-- layer=2 filter=158 channel=22
					-9, -6, 1, -1, -10, 8, -7, -2, 0,
					-- layer=2 filter=158 channel=23
					-15, 4, -3, -7, -12, -13, -44, -20, -15,
					-- layer=2 filter=158 channel=24
					-3, -6, -19, -11, -37, -31, 16, -10, -28,
					-- layer=2 filter=158 channel=25
					12, 21, -23, 17, -1, -25, 9, -6, -38,
					-- layer=2 filter=158 channel=26
					-5, 6, 1, -6, -7, -9, 0, 10, -8,
					-- layer=2 filter=158 channel=27
					11, 17, 7, -5, 0, -6, 25, -9, -26,
					-- layer=2 filter=158 channel=28
					-3, 24, 9, -4, -1, -16, -3, -8, 13,
					-- layer=2 filter=158 channel=29
					-1, -10, 7, 6, -6, 0, 1, 3, 3,
					-- layer=2 filter=158 channel=30
					-1, -28, -52, -17, -26, -16, -5, 2, 14,
					-- layer=2 filter=158 channel=31
					48, -4, -17, 82, 74, 102, 13, 11, -35,
					-- layer=2 filter=158 channel=32
					3, -1, 1, -3, -1, -5, -1, 3, -7,
					-- layer=2 filter=158 channel=33
					40, 20, 6, 47, 55, 18, 27, -2, -26,
					-- layer=2 filter=158 channel=34
					-12, -38, 18, -42, -45, -40, -77, -46, 18,
					-- layer=2 filter=158 channel=35
					-23, 26, 0, 3, -19, -57, -14, 15, 0,
					-- layer=2 filter=158 channel=36
					5, -4, 7, -12, -1, -2, -11, -3, -1,
					-- layer=2 filter=158 channel=37
					6, 11, -8, -10, -11, -9, -6, 9, 9,
					-- layer=2 filter=158 channel=38
					-6, 0, -10, 25, -7, -4, -7, 1, -21,
					-- layer=2 filter=158 channel=39
					4, 37, 23, -7, 21, 27, 30, 24, -25,
					-- layer=2 filter=158 channel=40
					-18, 24, -11, 22, 2, -32, -1, 7, 0,
					-- layer=2 filter=158 channel=41
					-3, 6, -2, 8, 8, -7, -2, -6, 8,
					-- layer=2 filter=158 channel=42
					-28, 9, 8, 8, 39, 25, 14, -47, -16,
					-- layer=2 filter=158 channel=43
					1, -1, -33, 12, -78, -30, 78, 57, 36,
					-- layer=2 filter=158 channel=44
					6, 0, 6, 10, -4, -4, 4, -7, 3,
					-- layer=2 filter=158 channel=45
					13, 5, -15, 8, 0, -14, 40, 11, -19,
					-- layer=2 filter=158 channel=46
					-10, -28, 11, -30, -16, -46, 38, 32, 34,
					-- layer=2 filter=158 channel=47
					-2, 13, 34, -1, 10, -60, 3, 1, 2,
					-- layer=2 filter=158 channel=48
					-8, 7, 6, 1, 2, -8, 8, -11, 6,
					-- layer=2 filter=158 channel=49
					1, -65, -34, -27, -20, -3, -47, 69, 54,
					-- layer=2 filter=158 channel=50
					17, 0, 21, 12, 1, -4, -11, 5, -3,
					-- layer=2 filter=158 channel=51
					42, 22, 1, -8, -30, -43, 14, 22, 0,
					-- layer=2 filter=158 channel=52
					11, -18, 9, -41, -58, -3, -10, -5, 27,
					-- layer=2 filter=158 channel=53
					25, -32, 47, -19, -8, -48, 42, 81, -1,
					-- layer=2 filter=158 channel=54
					37, 8, 6, 45, 29, 6, -24, -17, -27,
					-- layer=2 filter=158 channel=55
					-6, -4, -7, 1, 9, 2, -9, 10, 8,
					-- layer=2 filter=158 channel=56
					6, 19, 8, 19, -2, 3, 8, 4, -12,
					-- layer=2 filter=158 channel=57
					0, 8, -2, -11, -11, -3, -1, -8, -3,
					-- layer=2 filter=158 channel=58
					28, 22, -3, 44, 69, 81, -10, -69, -92,
					-- layer=2 filter=158 channel=59
					1, -8, -4, 26, 0, -1, -21, -27, -85,
					-- layer=2 filter=158 channel=60
					-3, -25, 22, 40, 19, -9, 0, -21, -33,
					-- layer=2 filter=158 channel=61
					1, -5, -13, -24, -80, -110, 7, 12, 7,
					-- layer=2 filter=158 channel=62
					16, 8, 45, -33, -44, 24, -56, 32, 35,
					-- layer=2 filter=158 channel=63
					-13, 12, -1, -23, -12, -39, 15, 0, 13,
					-- layer=2 filter=158 channel=64
					-31, -30, -18, -31, -23, -20, -41, -3, -32,
					-- layer=2 filter=158 channel=65
					-32, -31, -25, -42, -60, -55, -46, 16, -21,
					-- layer=2 filter=158 channel=66
					-12, 6, -33, 35, 24, 35, -38, -7, 7,
					-- layer=2 filter=158 channel=67
					3, -3, -14, -24, -55, -85, 59, 20, 18,
					-- layer=2 filter=158 channel=68
					-6, -1, -7, 7, -2, -2, 9, 7, 2,
					-- layer=2 filter=158 channel=69
					-28, -17, -11, -35, -21, -3, 8, -26, -43,
					-- layer=2 filter=158 channel=70
					2, 25, -5, 20, 11, -11, -15, 4, -24,
					-- layer=2 filter=158 channel=71
					23, -17, -7, -26, -15, -41, 18, -21, -35,
					-- layer=2 filter=158 channel=72
					-2, -7, 21, 17, 57, -1, 16, -3, -9,
					-- layer=2 filter=158 channel=73
					-23, -13, -4, -1, 16, -6, 11, 36, 30,
					-- layer=2 filter=158 channel=74
					-31, -16, -13, -23, -8, -23, 37, 28, 6,
					-- layer=2 filter=158 channel=75
					-1, 18, 20, 62, 50, 64, -33, -27, -38,
					-- layer=2 filter=158 channel=76
					1, -24, -9, -33, -51, -48, -10, 52, 24,
					-- layer=2 filter=158 channel=77
					-1, -7, 5, 1, -5, -6, 6, -12, -10,
					-- layer=2 filter=158 channel=78
					-4, 10, -22, -43, -25, -10, 6, 43, 7,
					-- layer=2 filter=158 channel=79
					-9, -1, -10, 3, 9, -2, -10, 7, 10,
					-- layer=2 filter=158 channel=80
					-35, -32, -10, 33, 18, 8, 1, 30, 18,
					-- layer=2 filter=158 channel=81
					17, 7, 20, 5, -1, 22, 18, 4, 25,
					-- layer=2 filter=158 channel=82
					0, -6, 10, -9, 1, 4, 7, 5, 1,
					-- layer=2 filter=158 channel=83
					-16, -5, 18, -20, 32, 3, -25, -12, -18,
					-- layer=2 filter=158 channel=84
					8, -6, -6, 11, -5, 4, -6, 3, 2,
					-- layer=2 filter=158 channel=85
					2, -6, -11, -2, 6, 3, 16, 4, 7,
					-- layer=2 filter=158 channel=86
					3, 0, 7, 19, -17, -11, -9, -10, 11,
					-- layer=2 filter=158 channel=87
					4, -1, -25, -40, -53, 0, -41, -28, 13,
					-- layer=2 filter=158 channel=88
					-23, -46, -30, -42, -20, 4, -13, 6, -12,
					-- layer=2 filter=158 channel=89
					10, -5, 0, 16, 29, 25, -23, -33, -53,
					-- layer=2 filter=158 channel=90
					-3, 7, 0, -10, 9, 1, 2, 3, -9,
					-- layer=2 filter=158 channel=91
					6, 31, 30, 29, 53, 35, 21, -46, -74,
					-- layer=2 filter=158 channel=92
					39, 0, 4, 15, 59, 40, 3, -53, -56,
					-- layer=2 filter=158 channel=93
					-11, -36, 22, 20, -6, 80, -54, 12, 2,
					-- layer=2 filter=158 channel=94
					-10, -33, -1, -19, -67, -83, -14, 57, -49,
					-- layer=2 filter=158 channel=95
					-11, 3, 0, -3, -9, -13, -8, 8, 3,
					-- layer=2 filter=158 channel=96
					-14, -38, -11, -21, -102, -24, -42, -33, 3,
					-- layer=2 filter=158 channel=97
					-2, -24, 11, -4, -31, -35, 32, 9, -40,
					-- layer=2 filter=158 channel=98
					-5, 33, 32, -22, 0, -42, -15, -9, -9,
					-- layer=2 filter=158 channel=99
					-31, -5, -18, -52, -90, -35, 3, 30, -36,
					-- layer=2 filter=158 channel=100
					-34, 27, -2, 43, 32, 12, -12, -10, -32,
					-- layer=2 filter=158 channel=101
					35, 15, 7, 24, -4, -18, 17, -4, -38,
					-- layer=2 filter=158 channel=102
					30, -33, -53, -24, -42, 9, -52, 28, 32,
					-- layer=2 filter=158 channel=103
					15, 20, -8, 25, 27, -13, -26, -56, -17,
					-- layer=2 filter=158 channel=104
					-14, -46, 20, -21, -22, -15, -47, 84, 33,
					-- layer=2 filter=158 channel=105
					-10, -10, 22, -32, -72, -38, -26, -4, -2,
					-- layer=2 filter=158 channel=106
					16, 40, 14, 28, 44, -6, 14, -37, -56,
					-- layer=2 filter=158 channel=107
					11, -7, -3, -2, -19, -1, -39, -34, 40,
					-- layer=2 filter=158 channel=108
					-24, -11, -46, -25, -3, -28, 13, 13, 29,
					-- layer=2 filter=158 channel=109
					-18, 13, -3, -8, 14, 1, 0, 9, 11,
					-- layer=2 filter=158 channel=110
					0, -15, -42, -6, -12, -40, -39, -30, -45,
					-- layer=2 filter=158 channel=111
					2, 0, 3, 8, -7, -1, -9, -5, 1,
					-- layer=2 filter=158 channel=112
					24, 20, 16, 9, -40, -98, 20, 32, 37,
					-- layer=2 filter=158 channel=113
					-40, 9, -32, -24, -60, -56, -17, 2, -20,
					-- layer=2 filter=158 channel=114
					18, 5, 5, -4, -4, -1, 8, -9, -8,
					-- layer=2 filter=158 channel=115
					9, -3, -7, 8, -6, 9, -9, 10, -5,
					-- layer=2 filter=158 channel=116
					34, -4, -19, -36, -30, 0, -14, 1, 15,
					-- layer=2 filter=158 channel=117
					17, -19, -5, 28, 40, -26, 1, -25, -16,
					-- layer=2 filter=158 channel=118
					-23, -8, -2, -38, -55, -12, 42, 50, 46,
					-- layer=2 filter=158 channel=119
					23, -32, -13, 25, 3, 3, -46, -24, -19,
					-- layer=2 filter=158 channel=120
					-5, -1, 6, 3, 5, -8, 0, -10, 8,
					-- layer=2 filter=158 channel=121
					4, -7, 3, 2, 5, 10, 0, 4, 6,
					-- layer=2 filter=158 channel=122
					2, 5, -7, 4, -6, -5, -7, -1, -11,
					-- layer=2 filter=158 channel=123
					2, -1, 24, -4, 13, -11, 13, -17, 7,
					-- layer=2 filter=158 channel=124
					18, 4, -22, 7, 1, -11, -9, 2, 6,
					-- layer=2 filter=158 channel=125
					-8, -8, -1, -12, 5, -3, 3, -3, -4,
					-- layer=2 filter=158 channel=126
					-38, 9, -18, 6, -4, 11, 43, -3, -68,
					-- layer=2 filter=158 channel=127
					-11, -15, -13, -8, -8, 0, 1, -18, -33,
					-- layer=2 filter=159 channel=0
					-10, 0, 0, -6, -4, -6, -4, -6, -9,
					-- layer=2 filter=159 channel=1
					4, 6, 7, -6, -10, -10, -23, -8, -4,
					-- layer=2 filter=159 channel=2
					5, -10, 0, 1, -1, 1, -9, 8, 7,
					-- layer=2 filter=159 channel=3
					-5, 1, -13, 3, -9, -6, 4, 6, -10,
					-- layer=2 filter=159 channel=4
					-14, -4, -16, 2, 5, -14, -4, -8, -12,
					-- layer=2 filter=159 channel=5
					-13, -7, -4, -3, 7, -4, -4, -5, -2,
					-- layer=2 filter=159 channel=6
					-22, -10, -2, -20, -9, 9, -12, 11, 0,
					-- layer=2 filter=159 channel=7
					6, -13, -15, -15, -20, -11, -12, -3, 0,
					-- layer=2 filter=159 channel=8
					-7, -3, 0, 0, 11, 10, 2, 2, 0,
					-- layer=2 filter=159 channel=9
					-1, -10, -6, -8, 0, -6, -1, -13, 0,
					-- layer=2 filter=159 channel=10
					6, -7, -16, -10, -1, -15, -2, -10, -10,
					-- layer=2 filter=159 channel=11
					-8, 2, 3, 7, 0, -9, -10, 9, 5,
					-- layer=2 filter=159 channel=12
					-9, -16, -9, 0, -7, 1, -23, -8, -2,
					-- layer=2 filter=159 channel=13
					0, -9, 1, -11, -4, 7, 0, -1, 7,
					-- layer=2 filter=159 channel=14
					5, 4, 6, -3, 6, -14, -17, 0, 4,
					-- layer=2 filter=159 channel=15
					0, 4, -1, -7, -10, -3, 3, -1, -7,
					-- layer=2 filter=159 channel=16
					-1, 3, -17, -7, 1, -4, -14, -7, -3,
					-- layer=2 filter=159 channel=17
					10, 4, -9, 0, 5, -5, 4, 1, 7,
					-- layer=2 filter=159 channel=18
					4, -4, -4, -23, 1, 5, -8, -2, 1,
					-- layer=2 filter=159 channel=19
					-11, 0, 11, 2, -3, 1, -18, -7, -5,
					-- layer=2 filter=159 channel=20
					-9, -3, -2, 1, 8, -1, -4, -1, -6,
					-- layer=2 filter=159 channel=21
					-2, -11, 3, -7, -5, 4, -5, 9, 0,
					-- layer=2 filter=159 channel=22
					8, -2, -3, -9, -9, 2, -1, -9, 0,
					-- layer=2 filter=159 channel=23
					-10, -15, -5, -11, 3, -15, -13, -13, -14,
					-- layer=2 filter=159 channel=24
					3, -4, -4, -8, 6, -15, 6, -14, -8,
					-- layer=2 filter=159 channel=25
					13, -4, 2, 0, -2, -13, 8, 6, -5,
					-- layer=2 filter=159 channel=26
					1, 0, 10, -2, -2, 0, 7, 8, -2,
					-- layer=2 filter=159 channel=27
					4, -4, 0, 5, -8, 4, -4, 7, 7,
					-- layer=2 filter=159 channel=28
					-9, -10, -8, -16, 9, -8, -7, -13, -2,
					-- layer=2 filter=159 channel=29
					-5, -1, -9, -5, -1, 5, 3, 0, -2,
					-- layer=2 filter=159 channel=30
					9, -14, -11, -7, -10, -17, 1, 3, 0,
					-- layer=2 filter=159 channel=31
					3, -1, -2, -9, -13, -1, -4, 1, -8,
					-- layer=2 filter=159 channel=32
					8, 2, 9, 2, -1, 5, -1, -4, 5,
					-- layer=2 filter=159 channel=33
					0, -19, -22, -22, -5, 8, -19, -6, -14,
					-- layer=2 filter=159 channel=34
					-1, -8, -12, -4, -8, -8, 6, -3, -2,
					-- layer=2 filter=159 channel=35
					-11, -9, -7, -5, 3, -14, -11, -4, -12,
					-- layer=2 filter=159 channel=36
					4, -5, 5, -8, 4, -9, 6, -6, -8,
					-- layer=2 filter=159 channel=37
					6, 2, 2, -2, 1, -5, -10, -10, -1,
					-- layer=2 filter=159 channel=38
					4, 5, -3, -8, 1, -11, 0, -8, 5,
					-- layer=2 filter=159 channel=39
					-9, -13, -5, -2, -1, -7, -10, -10, -9,
					-- layer=2 filter=159 channel=40
					0, -2, 15, 4, -8, -11, 3, -14, -9,
					-- layer=2 filter=159 channel=41
					-2, -4, 2, -1, 7, -9, -6, -6, -8,
					-- layer=2 filter=159 channel=42
					0, 0, 0, 1, -1, 7, -10, -9, 0,
					-- layer=2 filter=159 channel=43
					-10, -12, 0, 6, -1, -6, 4, -16, 4,
					-- layer=2 filter=159 channel=44
					7, 2, 2, 8, 10, 10, 0, -4, 1,
					-- layer=2 filter=159 channel=45
					3, 0, 2, -3, 5, -1, -12, -9, 2,
					-- layer=2 filter=159 channel=46
					-5, -1, 4, -6, -13, 5, -11, -6, -2,
					-- layer=2 filter=159 channel=47
					-9, -20, -16, -3, -11, -9, 1, -4, -17,
					-- layer=2 filter=159 channel=48
					0, -6, -9, 8, -4, 0, -3, -2, 10,
					-- layer=2 filter=159 channel=49
					-3, -14, 16, -17, -11, 4, -3, 4, 6,
					-- layer=2 filter=159 channel=50
					-3, 6, 5, -10, 10, 10, 5, 5, -9,
					-- layer=2 filter=159 channel=51
					6, -5, -10, 7, -3, 5, 5, -12, -9,
					-- layer=2 filter=159 channel=52
					-5, -5, -5, 2, 1, 0, -14, -6, 12,
					-- layer=2 filter=159 channel=53
					-13, -16, -4, -6, -4, 6, -4, -4, 2,
					-- layer=2 filter=159 channel=54
					-13, -17, -13, -15, -15, -8, -9, -11, 0,
					-- layer=2 filter=159 channel=55
					-8, 10, 8, 1, 1, 4, -4, 0, 11,
					-- layer=2 filter=159 channel=56
					2, 4, 1, -3, 5, -11, -13, -13, -12,
					-- layer=2 filter=159 channel=57
					-3, -2, -4, 4, -4, -4, 8, -6, -6,
					-- layer=2 filter=159 channel=58
					-3, -10, -10, 9, 0, 2, -24, -13, -15,
					-- layer=2 filter=159 channel=59
					-9, 6, 2, -3, -16, 2, -22, 0, 8,
					-- layer=2 filter=159 channel=60
					-12, -8, 8, -6, -18, -4, -17, -3, 0,
					-- layer=2 filter=159 channel=61
					-19, -6, 0, 0, -10, 1, -11, 0, -12,
					-- layer=2 filter=159 channel=62
					-6, 0, -5, -2, -15, 18, -4, 0, 10,
					-- layer=2 filter=159 channel=63
					1, -9, -14, -5, -5, -8, -16, 1, 0,
					-- layer=2 filter=159 channel=64
					1, 5, 1, -12, -7, -3, -2, -2, -1,
					-- layer=2 filter=159 channel=65
					-20, 4, -5, -12, -3, -8, -5, 4, 3,
					-- layer=2 filter=159 channel=66
					-9, -8, 5, -10, 0, -3, -4, 0, 6,
					-- layer=2 filter=159 channel=67
					13, -1, -5, -4, -4, -5, -9, -8, 2,
					-- layer=2 filter=159 channel=68
					-6, -3, -9, 2, -1, -4, -7, -4, -8,
					-- layer=2 filter=159 channel=69
					-8, 3, -6, -8, -1, -3, -1, -12, -4,
					-- layer=2 filter=159 channel=70
					-22, -15, -2, -5, 14, 8, 2, -18, 4,
					-- layer=2 filter=159 channel=71
					9, -5, -10, -9, -3, 1, -7, 8, 2,
					-- layer=2 filter=159 channel=72
					4, 1, -9, -20, -14, -3, -3, -9, -6,
					-- layer=2 filter=159 channel=73
					1, 2, 15, 8, 13, 0, 5, 9, 0,
					-- layer=2 filter=159 channel=74
					0, -3, -7, -10, -2, 0, -7, 7, -6,
					-- layer=2 filter=159 channel=75
					-11, 4, 0, 5, 0, 5, -9, 0, 0,
					-- layer=2 filter=159 channel=76
					0, -16, 8, -7, -5, 2, -14, 2, -2,
					-- layer=2 filter=159 channel=77
					-3, -5, -8, -1, 6, 2, 5, -5, -11,
					-- layer=2 filter=159 channel=78
					-3, 6, -1, -5, -14, -13, -11, -1, -2,
					-- layer=2 filter=159 channel=79
					0, 3, -8, -3, -3, 0, -6, 5, -4,
					-- layer=2 filter=159 channel=80
					0, 1, -10, -2, 5, 4, 2, -3, -11,
					-- layer=2 filter=159 channel=81
					0, 1, 8, -10, -6, -2, 3, 5, 1,
					-- layer=2 filter=159 channel=82
					-8, 6, 0, -4, 8, -5, 0, 7, 6,
					-- layer=2 filter=159 channel=83
					2, -3, -14, 2, -3, 0, 2, -7, -8,
					-- layer=2 filter=159 channel=84
					6, -5, -8, 0, 8, 1, 3, 3, -4,
					-- layer=2 filter=159 channel=85
					11, 9, 1, 2, -11, 9, -3, 3, -4,
					-- layer=2 filter=159 channel=86
					-7, 0, -4, 0, 4, 9, -2, 0, -2,
					-- layer=2 filter=159 channel=87
					-2, -19, 1, -13, -12, 5, -3, -3, -7,
					-- layer=2 filter=159 channel=88
					-6, -4, -6, -9, 6, 1, -11, 7, -7,
					-- layer=2 filter=159 channel=89
					3, -2, 13, 0, -5, 10, -25, 0, 1,
					-- layer=2 filter=159 channel=90
					-5, -8, 0, -9, -5, 5, 4, -3, -9,
					-- layer=2 filter=159 channel=91
					-16, -4, -6, -1, -5, 6, -20, -10, -14,
					-- layer=2 filter=159 channel=92
					-4, -7, 8, 1, -10, -8, -21, -7, -10,
					-- layer=2 filter=159 channel=93
					-10, 8, 3, 3, -9, 11, -2, -2, 11,
					-- layer=2 filter=159 channel=94
					-8, -20, -13, -14, -11, 2, -15, 1, -2,
					-- layer=2 filter=159 channel=95
					-10, 0, 5, 7, 4, 6, -2, -10, 0,
					-- layer=2 filter=159 channel=96
					-19, 2, 6, 9, 0, -10, -13, -22, -7,
					-- layer=2 filter=159 channel=97
					3, -11, -19, -3, -3, -12, 0, 0, -6,
					-- layer=2 filter=159 channel=98
					-20, -20, 5, -13, -1, 0, -12, -6, -15,
					-- layer=2 filter=159 channel=99
					-2, 14, 13, -1, -5, -5, -14, -11, 1,
					-- layer=2 filter=159 channel=100
					-6, -4, 1, 7, 6, -2, 3, -11, -3,
					-- layer=2 filter=159 channel=101
					3, 12, 8, -2, 0, 0, 8, 0, 1,
					-- layer=2 filter=159 channel=102
					-18, 3, -8, -7, 6, 14, -5, -20, -6,
					-- layer=2 filter=159 channel=103
					2, 0, -8, -5, -8, -10, 8, 7, 0,
					-- layer=2 filter=159 channel=104
					-11, 5, -3, -7, -2, -3, -5, 4, -9,
					-- layer=2 filter=159 channel=105
					0, 5, 7, 2, -3, -7, -5, -9, 13,
					-- layer=2 filter=159 channel=106
					1, -9, -9, 5, 0, -15, 0, 8, -4,
					-- layer=2 filter=159 channel=107
					-8, 0, 3, 3, 11, -5, 3, -1, 7,
					-- layer=2 filter=159 channel=108
					2, -2, 2, 3, -10, -8, 4, -10, 9,
					-- layer=2 filter=159 channel=109
					-1, 8, -6, -6, -4, -11, 2, 4, 0,
					-- layer=2 filter=159 channel=110
					0, -11, 0, 0, 1, 0, 4, -7, 3,
					-- layer=2 filter=159 channel=111
					0, 5, 0, -7, -6, -6, 3, 3, -6,
					-- layer=2 filter=159 channel=112
					-3, -10, -10, 2, 5, -13, -12, -8, -9,
					-- layer=2 filter=159 channel=113
					7, -14, -12, -1, -4, -17, -6, -18, -10,
					-- layer=2 filter=159 channel=114
					-10, 2, -2, 1, -8, -9, 3, -3, -1,
					-- layer=2 filter=159 channel=115
					-6, -6, -4, -1, 8, 8, -6, 9, 0,
					-- layer=2 filter=159 channel=116
					-10, 0, 1, -20, 0, 10, -5, -7, 2,
					-- layer=2 filter=159 channel=117
					7, 1, 0, 2, 3, -8, -14, -14, 3,
					-- layer=2 filter=159 channel=118
					-4, -10, -5, -6, -15, -8, -7, -16, 3,
					-- layer=2 filter=159 channel=119
					-14, -9, -1, -5, 2, 0, -4, 0, -3,
					-- layer=2 filter=159 channel=120
					-2, -1, 6, -4, 6, -1, 4, 8, -8,
					-- layer=2 filter=159 channel=121
					-8, -1, -11, -7, -2, 0, -3, -4, 3,
					-- layer=2 filter=159 channel=122
					0, -5, -10, 6, 0, -5, -3, 10, -7,
					-- layer=2 filter=159 channel=123
					0, -10, -3, -19, -7, 7, -13, 6, -10,
					-- layer=2 filter=159 channel=124
					11, 6, -5, -18, -14, 0, -13, 0, -12,
					-- layer=2 filter=159 channel=125
					4, 0, 0, -10, 1, -2, -10, 2, -1,
					-- layer=2 filter=159 channel=126
					-7, -9, -5, 9, 7, -11, -4, 4, 3,
					-- layer=2 filter=159 channel=127
					5, -3, -14, 3, -4, 5, 4, 0, 0,
					-- layer=2 filter=160 channel=0
					-6, 2, -5, 13, 11, 10, 15, 31, 0,
					-- layer=2 filter=160 channel=1
					32, 16, 7, -15, -13, 4, -24, -24, 15,
					-- layer=2 filter=160 channel=2
					-8, -5, -11, -8, -8, 0, -10, -6, -1,
					-- layer=2 filter=160 channel=3
					-44, 1, -20, -2, -33, -13, 17, 8, -17,
					-- layer=2 filter=160 channel=4
					-24, -39, -12, -1, -25, -7, 29, 28, 31,
					-- layer=2 filter=160 channel=5
					-5, 10, -7, 11, 18, 0, 3, 17, 38,
					-- layer=2 filter=160 channel=6
					54, 34, 35, -10, -4, 16, -25, -16, -2,
					-- layer=2 filter=160 channel=7
					8, 3, 11, 0, -14, 5, 47, 14, -14,
					-- layer=2 filter=160 channel=8
					1, 3, -4, 4, 0, -3, 10, 11, -3,
					-- layer=2 filter=160 channel=9
					-2, -1, -23, -65, -76, -57, 5, 5, -17,
					-- layer=2 filter=160 channel=10
					-20, -19, -22, 5, 16, 10, 39, 17, 17,
					-- layer=2 filter=160 channel=11
					10, 14, 4, 19, 12, 1, 11, -3, 3,
					-- layer=2 filter=160 channel=12
					14, 4, 16, -23, -34, -20, -9, -25, 17,
					-- layer=2 filter=160 channel=13
					-5, -3, -1, -1, 2, 3, 2, 3, -4,
					-- layer=2 filter=160 channel=14
					38, 29, 10, -5, -22, 1, -42, -36, 16,
					-- layer=2 filter=160 channel=15
					10, -13, -6, -5, -4, 5, -4, -2, 19,
					-- layer=2 filter=160 channel=16
					-21, 4, -5, -26, -18, -5, -17, -6, -27,
					-- layer=2 filter=160 channel=17
					3, 3, 2, 3, 3, 10, -10, -2, -1,
					-- layer=2 filter=160 channel=18
					38, -8, 12, -3, 3, -25, -24, -4, 7,
					-- layer=2 filter=160 channel=19
					-2, 0, 10, -3, -18, 12, 7, -40, -10,
					-- layer=2 filter=160 channel=20
					9, 0, -1, -11, 2, 4, -11, -12, -8,
					-- layer=2 filter=160 channel=21
					-10, -5, -9, -16, 6, -19, 7, 9, 4,
					-- layer=2 filter=160 channel=22
					-2, -8, 0, 0, -1, 2, 5, 0, -3,
					-- layer=2 filter=160 channel=23
					-19, 5, 2, -13, -11, 21, 12, 36, 19,
					-- layer=2 filter=160 channel=24
					-25, -2, 4, -12, -26, -15, 3, 18, -14,
					-- layer=2 filter=160 channel=25
					11, 19, 19, 7, -9, -12, -6, 12, 9,
					-- layer=2 filter=160 channel=26
					-3, 2, 4, 2, -5, 9, 4, 1, 0,
					-- layer=2 filter=160 channel=27
					7, 15, -1, -10, -14, 10, 21, 30, 24,
					-- layer=2 filter=160 channel=28
					-33, -26, 5, 1, -11, -22, 3, 29, 14,
					-- layer=2 filter=160 channel=29
					-8, -6, -7, -11, -1, -5, -1, -10, 0,
					-- layer=2 filter=160 channel=30
					-21, 9, -11, -20, 6, -13, -11, -15, 6,
					-- layer=2 filter=160 channel=31
					-36, -27, 4, 28, -21, 18, 0, -29, 28,
					-- layer=2 filter=160 channel=32
					0, 4, 5, 2, -6, -13, -4, -11, 10,
					-- layer=2 filter=160 channel=33
					0, -6, -1, -16, -27, -6, -44, -56, -28,
					-- layer=2 filter=160 channel=34
					34, 4, 14, 22, -31, 27, -28, -42, 3,
					-- layer=2 filter=160 channel=35
					35, -16, -16, 15, 8, -5, 13, 8, 21,
					-- layer=2 filter=160 channel=36
					1, 8, -1, -11, 0, 4, 9, 8, 14,
					-- layer=2 filter=160 channel=37
					19, 1, -4, 17, 6, 9, 12, -9, 16,
					-- layer=2 filter=160 channel=38
					17, 10, 18, -9, 13, -6, 0, 0, 23,
					-- layer=2 filter=160 channel=39
					-24, -1, 7, 12, -38, -10, 7, 11, 1,
					-- layer=2 filter=160 channel=40
					15, 7, -6, 9, -14, -27, 23, -13, 22,
					-- layer=2 filter=160 channel=41
					-9, 5, 3, 1, 2, -4, 0, -4, 7,
					-- layer=2 filter=160 channel=42
					12, 28, 7, 0, 5, -23, 20, 12, -4,
					-- layer=2 filter=160 channel=43
					-37, -48, -46, -1, -18, -20, 19, -15, -4,
					-- layer=2 filter=160 channel=44
					-11, 0, 3, -7, 9, -5, -7, -2, -3,
					-- layer=2 filter=160 channel=45
					-68, -39, -48, -55, -66, -79, -54, -39, -67,
					-- layer=2 filter=160 channel=46
					-22, -46, -30, 21, -28, -7, 25, -4, 14,
					-- layer=2 filter=160 channel=47
					-51, -63, -47, -40, -50, -54, -34, -21, -10,
					-- layer=2 filter=160 channel=48
					0, 4, -7, 1, 1, -1, -5, 3, -2,
					-- layer=2 filter=160 channel=49
					17, 18, 28, 23, -3, -4, -60, -1, -16,
					-- layer=2 filter=160 channel=50
					-16, -6, -18, 14, -18, 17, 3, 28, 4,
					-- layer=2 filter=160 channel=51
					-4, 8, 1, 12, -4, 10, 2, 4, -6,
					-- layer=2 filter=160 channel=52
					21, -1, 9, 40, -20, 15, 20, 7, 27,
					-- layer=2 filter=160 channel=53
					-83, -25, -14, -37, -4, -15, -95, -19, 14,
					-- layer=2 filter=160 channel=54
					19, 5, 24, 23, 12, -2, 35, -7, 33,
					-- layer=2 filter=160 channel=55
					-8, -12, 0, 9, -2, -11, 4, -11, -6,
					-- layer=2 filter=160 channel=56
					0, 0, 9, 16, -9, 8, 7, 5, 15,
					-- layer=2 filter=160 channel=57
					-12, -5, 3, 13, -4, 0, 9, 3, 7,
					-- layer=2 filter=160 channel=58
					11, 8, -3, -15, -30, 15, 15, -35, 13,
					-- layer=2 filter=160 channel=59
					-20, 25, 29, -23, -9, 38, 1, -6, 26,
					-- layer=2 filter=160 channel=60
					10, 2, 45, -18, 12, 10, -8, -12, 20,
					-- layer=2 filter=160 channel=61
					-4, -17, 17, -22, -13, -25, 0, 0, -50,
					-- layer=2 filter=160 channel=62
					39, 8, 6, -1, 18, 43, -45, -7, 1,
					-- layer=2 filter=160 channel=63
					-31, -2, 22, -5, -41, 16, 4, 37, 9,
					-- layer=2 filter=160 channel=64
					8, 30, 15, -7, -1, -11, 31, 26, 13,
					-- layer=2 filter=160 channel=65
					-3, -1, 7, -31, 7, 4, -3, -17, -10,
					-- layer=2 filter=160 channel=66
					27, 8, -44, -41, 44, -5, 1, -26, -41,
					-- layer=2 filter=160 channel=67
					-38, -63, -36, -119, -102, -51, -37, -29, -19,
					-- layer=2 filter=160 channel=68
					-1, 6, -4, -9, 5, -5, 0, 0, 5,
					-- layer=2 filter=160 channel=69
					20, 21, 19, 19, 30, 22, 13, 24, -3,
					-- layer=2 filter=160 channel=70
					11, -8, 12, 29, 1, -3, 28, 21, 44,
					-- layer=2 filter=160 channel=71
					30, 17, -24, -12, -8, 8, -26, -24, -25,
					-- layer=2 filter=160 channel=72
					47, 43, 23, 5, 1, -7, 31, 20, -2,
					-- layer=2 filter=160 channel=73
					-7, -4, 5, 8, -10, -17, 25, 1, -56,
					-- layer=2 filter=160 channel=74
					-29, -45, -13, -39, -1, 5, 40, -11, 55,
					-- layer=2 filter=160 channel=75
					-3, -22, -49, -6, -35, -30, -91, -26, -24,
					-- layer=2 filter=160 channel=76
					-47, -33, -13, 16, -12, -24, -51, -43, -11,
					-- layer=2 filter=160 channel=77
					9, -1, 3, 2, -4, -12, 6, -8, -1,
					-- layer=2 filter=160 channel=78
					19, 5, 15, 14, -8, 6, 12, 7, 2,
					-- layer=2 filter=160 channel=79
					-2, -10, 0, -4, -7, 9, -6, 7, 1,
					-- layer=2 filter=160 channel=80
					-40, -2, -19, -8, -2, -11, 14, -5, 5,
					-- layer=2 filter=160 channel=81
					-2, -9, -5, -5, -3, -3, -15, -8, -10,
					-- layer=2 filter=160 channel=82
					0, -2, 5, -4, 1, 5, 2, 0, 6,
					-- layer=2 filter=160 channel=83
					-41, -18, 1, -23, -17, 4, 20, 0, 29,
					-- layer=2 filter=160 channel=84
					6, -5, 7, -3, 2, -7, 11, -6, 2,
					-- layer=2 filter=160 channel=85
					0, -2, 2, 10, 1, 6, -19, -9, 8,
					-- layer=2 filter=160 channel=86
					1, 2, -2, -10, -2, -2, 0, -10, -17,
					-- layer=2 filter=160 channel=87
					-6, 19, 8, 13, 11, -22, -38, 13, -15,
					-- layer=2 filter=160 channel=88
					21, 16, 27, -87, 12, -27, -32, -16, 17,
					-- layer=2 filter=160 channel=89
					46, 38, 4, 9, -21, 29, -38, -11, 26,
					-- layer=2 filter=160 channel=90
					-11, -7, 7, 8, 8, 9, 2, -4, 0,
					-- layer=2 filter=160 channel=91
					12, 5, -13, 3, -21, -3, -29, -37, -4,
					-- layer=2 filter=160 channel=92
					46, 24, 32, -3, -21, 6, -7, -4, 10,
					-- layer=2 filter=160 channel=93
					-18, -31, -28, -35, -24, -37, 21, -7, 0,
					-- layer=2 filter=160 channel=94
					-4, 41, 41, 5, 1, -7, -21, 13, -2,
					-- layer=2 filter=160 channel=95
					-17, -2, -5, -3, 1, 4, 10, 0, 7,
					-- layer=2 filter=160 channel=96
					36, 46, 24, 43, 23, 6, 20, 5, 6,
					-- layer=2 filter=160 channel=97
					0, 6, -11, -49, -28, -36, -6, 2, -7,
					-- layer=2 filter=160 channel=98
					14, 0, -9, 0, 4, 8, 21, 39, 32,
					-- layer=2 filter=160 channel=99
					-2, 14, 1, 2, -14, 25, 8, -35, 11,
					-- layer=2 filter=160 channel=100
					11, -12, -10, 12, 21, 1, 23, 0, 59,
					-- layer=2 filter=160 channel=101
					18, 15, -12, 0, -7, 4, -29, -10, -44,
					-- layer=2 filter=160 channel=102
					27, 3, 27, -12, 9, -32, 34, -14, -49,
					-- layer=2 filter=160 channel=103
					-3, -31, 5, -31, 19, 13, -8, -26, -16,
					-- layer=2 filter=160 channel=104
					-15, -9, 21, 8, -8, -8, -48, 20, 16,
					-- layer=2 filter=160 channel=105
					-73, -46, -15, -19, -23, -49, -21, 7, -66,
					-- layer=2 filter=160 channel=106
					12, 2, 1, -25, -18, -23, -46, -23, -16,
					-- layer=2 filter=160 channel=107
					29, 9, 19, 0, 27, 17, -1, -20, -41,
					-- layer=2 filter=160 channel=108
					28, 25, 32, 9, 16, 0, -13, -14, 16,
					-- layer=2 filter=160 channel=109
					-4, 1, -15, 6, -22, -1, 6, -2, -8,
					-- layer=2 filter=160 channel=110
					8, 16, -7, 2, 2, -16, 17, 18, 14,
					-- layer=2 filter=160 channel=111
					0, -9, 4, 10, -3, 2, -7, -8, 6,
					-- layer=2 filter=160 channel=112
					-4, -26, -21, 7, 9, 10, 9, 5, -11,
					-- layer=2 filter=160 channel=113
					-11, -7, -38, 4, -31, -8, 3, 0, 22,
					-- layer=2 filter=160 channel=114
					11, 6, 5, 9, 6, 7, 1, 0, 2,
					-- layer=2 filter=160 channel=115
					5, 3, 4, 5, 1, 12, -2, -6, 1,
					-- layer=2 filter=160 channel=116
					20, -7, 0, -3, -13, 10, -15, -9, 0,
					-- layer=2 filter=160 channel=117
					18, -9, 10, 0, -18, -27, -12, -35, -8,
					-- layer=2 filter=160 channel=118
					-14, 14, 0, 14, -7, 1, 19, 21, 0,
					-- layer=2 filter=160 channel=119
					20, -49, -15, -12, -18, -28, -27, -1, -2,
					-- layer=2 filter=160 channel=120
					5, 4, 9, -4, -7, 0, -10, -4, -6,
					-- layer=2 filter=160 channel=121
					-7, -12, 4, -11, 2, 3, -8, 3, -4,
					-- layer=2 filter=160 channel=122
					21, 15, 0, -3, 7, -1, -6, 17, 3,
					-- layer=2 filter=160 channel=123
					-2, 24, 23, 2, -6, 11, 1, 9, -1,
					-- layer=2 filter=160 channel=124
					14, 29, -10, 31, 8, 19, 19, 12, 25,
					-- layer=2 filter=160 channel=125
					3, -5, -4, -2, 1, -1, -10, -10, -4,
					-- layer=2 filter=160 channel=126
					-6, -39, -7, -25, -99, -13, -11, -65, -83,
					-- layer=2 filter=160 channel=127
					4, 5, -12, -22, 4, -4, 19, 12, 13,
					-- layer=2 filter=161 channel=0
					-8, 19, 0, -1, 14, 13, -25, 15, 11,
					-- layer=2 filter=161 channel=1
					-36, 3, -17, -19, -31, -57, -17, -14, -6,
					-- layer=2 filter=161 channel=2
					-8, 2, 0, 0, 8, 6, 7, -1, 0,
					-- layer=2 filter=161 channel=3
					14, 7, 3, 26, -18, 5, -6, -14, 3,
					-- layer=2 filter=161 channel=4
					-14, -30, 0, -2, 5, 33, -14, 1, -11,
					-- layer=2 filter=161 channel=5
					-11, 31, 13, -9, 11, -7, -14, 11, -9,
					-- layer=2 filter=161 channel=6
					39, 58, 2, 76, 37, 44, 3, 22, 0,
					-- layer=2 filter=161 channel=7
					-16, -47, 16, -30, -106, -46, -10, -76, -28,
					-- layer=2 filter=161 channel=8
					4, -3, -3, 2, -4, 0, 8, -8, 3,
					-- layer=2 filter=161 channel=9
					-6, 0, 0, -1, -1, -12, 12, 21, 9,
					-- layer=2 filter=161 channel=10
					5, -2, 19, -2, 19, 29, -21, 9, -1,
					-- layer=2 filter=161 channel=11
					22, 15, 8, 11, -8, -1, -14, -7, 18,
					-- layer=2 filter=161 channel=12
					16, 2, 18, -11, -69, -71, 3, -7, -3,
					-- layer=2 filter=161 channel=13
					-2, 0, 7, -8, -4, -6, -7, 3, 0,
					-- layer=2 filter=161 channel=14
					0, -26, -24, -33, -68, -97, -5, -27, 8,
					-- layer=2 filter=161 channel=15
					45, -39, -23, 16, -19, -13, 16, -6, 10,
					-- layer=2 filter=161 channel=16
					-27, -14, -5, 21, -3, -21, 7, 19, -19,
					-- layer=2 filter=161 channel=17
					6, -4, -3, 5, 9, 0, -8, -10, -7,
					-- layer=2 filter=161 channel=18
					25, -21, -11, 14, 14, 3, -9, 0, 8,
					-- layer=2 filter=161 channel=19
					-60, -18, -17, -22, -32, 16, 11, -43, -54,
					-- layer=2 filter=161 channel=20
					-1, 0, 0, -5, -6, 10, -8, 3, 5,
					-- layer=2 filter=161 channel=21
					-3, -4, 14, 0, 0, 9, -3, 9, 1,
					-- layer=2 filter=161 channel=22
					3, 5, -3, -8, -5, -1, -1, -1, 1,
					-- layer=2 filter=161 channel=23
					4, 28, 11, -3, 29, 30, -14, -1, -23,
					-- layer=2 filter=161 channel=24
					-17, -5, -27, -2, 15, 7, -10, 35, 29,
					-- layer=2 filter=161 channel=25
					-34, -8, -21, -1, 14, 3, 6, 27, 17,
					-- layer=2 filter=161 channel=26
					9, 9, -12, 4, -9, 0, -3, -8, -7,
					-- layer=2 filter=161 channel=27
					-24, 22, 17, 8, 1, -11, -3, -9, -9,
					-- layer=2 filter=161 channel=28
					-19, -73, -51, -22, -67, -33, -72, -64, -60,
					-- layer=2 filter=161 channel=29
					4, -5, -7, 6, -4, 7, -5, 3, -3,
					-- layer=2 filter=161 channel=30
					-3, 0, 12, -12, -12, -5, 17, 23, -11,
					-- layer=2 filter=161 channel=31
					5, -19, -40, 7, 33, -34, 59, 72, -66,
					-- layer=2 filter=161 channel=32
					-8, -5, -2, -1, 10, 6, -8, -10, -10,
					-- layer=2 filter=161 channel=33
					35, -10, 2, 32, -94, -14, -2, -36, -7,
					-- layer=2 filter=161 channel=34
					3, 4, 85, 2, 62, 22, -19, -4, -41,
					-- layer=2 filter=161 channel=35
					22, -26, -13, -37, -40, -31, -107, -109, -95,
					-- layer=2 filter=161 channel=36
					3, 7, 7, -10, 15, -5, 0, 0, 7,
					-- layer=2 filter=161 channel=37
					3, 10, 8, 12, 18, -2, 7, 2, 13,
					-- layer=2 filter=161 channel=38
					0, 18, 15, 3, 5, -13, -23, -8, -16,
					-- layer=2 filter=161 channel=39
					34, 8, -7, 23, 8, -6, -8, -23, -23,
					-- layer=2 filter=161 channel=40
					29, 10, -6, 31, -28, -33, -33, -15, 35,
					-- layer=2 filter=161 channel=41
					4, -11, 5, 5, 4, 2, 0, 8, 0,
					-- layer=2 filter=161 channel=42
					29, 21, -3, 43, 4, -12, 14, -10, -7,
					-- layer=2 filter=161 channel=43
					15, 10, -7, -1, 21, 0, 16, -31, -7,
					-- layer=2 filter=161 channel=44
					4, 5, 0, -9, -5, -5, 4, 8, -5,
					-- layer=2 filter=161 channel=45
					-29, 0, -7, -36, -35, -21, 20, -30, 5,
					-- layer=2 filter=161 channel=46
					-2, 10, 0, -5, 19, 3, -2, 20, -11,
					-- layer=2 filter=161 channel=47
					-23, -76, -50, -6, -62, -39, -14, -12, 35,
					-- layer=2 filter=161 channel=48
					-4, -3, -9, 4, -3, 0, -4, -1, 4,
					-- layer=2 filter=161 channel=49
					7, -10, -17, 11, 2, 13, 24, 0, 18,
					-- layer=2 filter=161 channel=50
					0, 12, 0, -8, 11, 14, 11, 11, 3,
					-- layer=2 filter=161 channel=51
					1, 7, -7, 1, 12, 7, -4, -1, -5,
					-- layer=2 filter=161 channel=52
					7, 15, -9, -17, -16, -17, -2, -14, -4,
					-- layer=2 filter=161 channel=53
					30, 15, -18, 20, -33, 24, 26, 58, -56,
					-- layer=2 filter=161 channel=54
					7, 10, -12, -20, -19, 15, -25, -29, 1,
					-- layer=2 filter=161 channel=55
					-9, 0, 10, 4, -7, -6, -1, 6, -10,
					-- layer=2 filter=161 channel=56
					23, 12, 6, 20, -9, -3, -4, -9, 10,
					-- layer=2 filter=161 channel=57
					19, 10, -1, 4, 8, 0, 5, -9, 3,
					-- layer=2 filter=161 channel=58
					55, 26, 27, -17, -60, -57, 6, -29, -16,
					-- layer=2 filter=161 channel=59
					-23, -22, -23, -52, -63, -52, -60, -21, -18,
					-- layer=2 filter=161 channel=60
					-23, 13, 18, -64, -17, -19, -17, -26, -21,
					-- layer=2 filter=161 channel=61
					-36, 10, 22, -33, -8, 15, -21, -4, 24,
					-- layer=2 filter=161 channel=62
					-16, 35, 6, 22, 57, 44, 7, -9, -14,
					-- layer=2 filter=161 channel=63
					0, 0, -11, -8, -2, -13, -28, 4, -6,
					-- layer=2 filter=161 channel=64
					-4, -12, -3, 8, 18, -10, 5, 12, -8,
					-- layer=2 filter=161 channel=65
					-9, 26, 20, -9, 37, -5, -11, 2, 7,
					-- layer=2 filter=161 channel=66
					24, -1, 33, 1, -16, -8, -12, -13, 15,
					-- layer=2 filter=161 channel=67
					-1, 27, -9, -4, 27, 16, -23, 24, 23,
					-- layer=2 filter=161 channel=68
					2, 12, -8, 0, -5, -8, 8, 7, -6,
					-- layer=2 filter=161 channel=69
					-14, -1, -1, 24, 22, 7, 14, 7, 3,
					-- layer=2 filter=161 channel=70
					2, -29, 9, -10, -39, 2, -42, -42, -40,
					-- layer=2 filter=161 channel=71
					8, 22, -11, 16, -1, -35, 32, -24, -25,
					-- layer=2 filter=161 channel=72
					22, -4, -29, 6, -88, -47, -48, -45, -41,
					-- layer=2 filter=161 channel=73
					-26, 0, 24, -31, -33, 28, 12, 38, 44,
					-- layer=2 filter=161 channel=74
					16, 5, -9, -10, -23, -8, -23, 12, -1,
					-- layer=2 filter=161 channel=75
					59, 20, 24, 3, 28, -68, 77, 36, 108,
					-- layer=2 filter=161 channel=76
					26, 36, 23, -39, -21, 24, -13, 6, -16,
					-- layer=2 filter=161 channel=77
					-6, 6, 0, -5, 3, 1, 8, -7, 0,
					-- layer=2 filter=161 channel=78
					-5, 32, -4, 19, 11, 19, -1, -9, 5,
					-- layer=2 filter=161 channel=79
					-5, -6, -3, 10, 6, -7, 11, 4, -5,
					-- layer=2 filter=161 channel=80
					12, -14, -6, 16, 7, 3, 15, -14, 4,
					-- layer=2 filter=161 channel=81
					-3, 11, 7, 11, 14, -4, 16, 7, 2,
					-- layer=2 filter=161 channel=82
					-5, -6, 2, -7, -3, 6, 3, -5, -2,
					-- layer=2 filter=161 channel=83
					-15, 4, 0, 18, 7, 31, -4, 2, 4,
					-- layer=2 filter=161 channel=84
					6, -3, 7, 0, 8, -6, 0, -10, -4,
					-- layer=2 filter=161 channel=85
					-7, -1, -14, 5, -8, -4, -2, -1, 0,
					-- layer=2 filter=161 channel=86
					-10, -31, -13, -5, 1, -4, -12, -3, 3,
					-- layer=2 filter=161 channel=87
					20, 0, -10, -27, 22, 44, -58, -30, 12,
					-- layer=2 filter=161 channel=88
					-20, 11, 6, 2, -9, -21, -17, 14, 32,
					-- layer=2 filter=161 channel=89
					-6, -4, 12, -29, -47, -58, -18, -20, 0,
					-- layer=2 filter=161 channel=90
					0, 0, 1, 0, 2, 8, -2, -7, 4,
					-- layer=2 filter=161 channel=91
					55, 9, 17, 29, -4, -37, 3, -3, 9,
					-- layer=2 filter=161 channel=92
					-9, -2, -6, -23, -46, -67, -53, -26, -26,
					-- layer=2 filter=161 channel=93
					1, 50, -15, 34, 56, 39, 58, 24, -21,
					-- layer=2 filter=161 channel=94
					-44, 26, 31, -2, -22, 36, -35, 8, -26,
					-- layer=2 filter=161 channel=95
					9, -6, -4, 1, -10, -7, 6, 9, -14,
					-- layer=2 filter=161 channel=96
					24, 90, 20, -27, 53, 53, -23, 44, 25,
					-- layer=2 filter=161 channel=97
					4, -5, -12, 22, -15, -33, 47, -7, -1,
					-- layer=2 filter=161 channel=98
					-27, -70, -39, 4, -42, -15, -37, -66, -32,
					-- layer=2 filter=161 channel=99
					9, 38, 22, -4, -32, 5, 9, 7, 4,
					-- layer=2 filter=161 channel=100
					14, 27, 16, -1, -5, -3, -3, -20, -45,
					-- layer=2 filter=161 channel=101
					11, -13, -3, 2, -21, -10, 27, 9, -9,
					-- layer=2 filter=161 channel=102
					-20, 12, 11, -8, 4, 3, -17, 42, -2,
					-- layer=2 filter=161 channel=103
					4, 8, -1, 14, 2, -43, 42, 62, 79,
					-- layer=2 filter=161 channel=104
					-15, 9, -15, 7, 9, 43, -1, -22, -1,
					-- layer=2 filter=161 channel=105
					-11, 61, 74, -72, -12, -27, -45, -64, -39,
					-- layer=2 filter=161 channel=106
					-2, 0, 6, 7, -9, -34, 17, 20, 13,
					-- layer=2 filter=161 channel=107
					-27, -25, 0, -64, -44, 0, 5, -13, -12,
					-- layer=2 filter=161 channel=108
					-30, -18, -14, 4, -11, -19, 13, -7, 10,
					-- layer=2 filter=161 channel=109
					-9, 16, 2, 0, 8, -3, 0, 0, 6,
					-- layer=2 filter=161 channel=110
					-7, 16, 16, 0, 23, 1, -16, -8, -5,
					-- layer=2 filter=161 channel=111
					9, 4, -5, -12, -9, -12, 6, 8, 4,
					-- layer=2 filter=161 channel=112
					30, 4, -15, 10, 41, 1, 0, 13, 24,
					-- layer=2 filter=161 channel=113
					21, -10, -7, -22, -14, -35, -10, 8, -46,
					-- layer=2 filter=161 channel=114
					5, -5, 4, -6, 5, 7, -8, 15, 1,
					-- layer=2 filter=161 channel=115
					-2, -9, -3, 5, 4, -6, -6, 0, 7,
					-- layer=2 filter=161 channel=116
					12, 16, -17, -14, 20, 22, -42, 12, 24,
					-- layer=2 filter=161 channel=117
					-23, -14, 9, -42, -104, -49, 10, -59, 35,
					-- layer=2 filter=161 channel=118
					5, 1, -6, 9, 14, 15, 13, -6, 7,
					-- layer=2 filter=161 channel=119
					18, -36, 0, 14, 35, -4, 20, 36, 19,
					-- layer=2 filter=161 channel=120
					2, -9, -6, -3, -8, 7, 0, -9, 6,
					-- layer=2 filter=161 channel=121
					9, -1, 0, -11, -3, -5, 10, 6, 9,
					-- layer=2 filter=161 channel=122
					7, 5, 7, -2, -8, -7, 11, 1, 5,
					-- layer=2 filter=161 channel=123
					-33, -18, -12, -24, -72, -21, -26, -40, -51,
					-- layer=2 filter=161 channel=124
					-6, -27, -12, 13, -2, 26, 51, 7, -58,
					-- layer=2 filter=161 channel=125
					-6, 0, -5, -8, 5, 0, 6, -4, -5,
					-- layer=2 filter=161 channel=126
					-19, 44, 10, -31, 42, -28, 29, 55, -24,
					-- layer=2 filter=161 channel=127
					8, -18, 0, 4, -12, 3, -35, -12, -3,
					-- layer=2 filter=162 channel=0
					7, -4, 5, 2, -14, -18, 7, -33, -46,
					-- layer=2 filter=162 channel=1
					-22, 16, 10, -6, -5, 5, -14, 24, 26,
					-- layer=2 filter=162 channel=2
					0, 7, -10, 9, 7, -6, -7, 7, -8,
					-- layer=2 filter=162 channel=3
					-17, -37, -23, -20, -38, -60, 47, 8, -15,
					-- layer=2 filter=162 channel=4
					0, -8, -9, 11, 13, -31, -9, -21, 9,
					-- layer=2 filter=162 channel=5
					10, -15, -4, 35, 38, -9, 2, -4, 7,
					-- layer=2 filter=162 channel=6
					-17, 4, -48, -21, -11, -32, -37, 31, -25,
					-- layer=2 filter=162 channel=7
					-18, 3, 21, 33, 5, -18, -18, 38, -3,
					-- layer=2 filter=162 channel=8
					-9, 4, 4, 0, 0, -2, -4, 0, 7,
					-- layer=2 filter=162 channel=9
					-14, 0, 25, 12, -6, 2, 11, -26, -48,
					-- layer=2 filter=162 channel=10
					-17, -11, 8, -5, -44, -61, 6, -43, -40,
					-- layer=2 filter=162 channel=11
					23, 8, 13, 14, 6, 23, 0, -4, -18,
					-- layer=2 filter=162 channel=12
					19, 49, 26, -9, 1, 4, 7, 0, 35,
					-- layer=2 filter=162 channel=13
					-2, 7, -5, -6, -1, 1, 9, -9, 9,
					-- layer=2 filter=162 channel=14
					-13, 23, 27, -7, 1, 16, -18, -6, 5,
					-- layer=2 filter=162 channel=15
					32, -11, -13, 0, -11, -25, -15, -13, 0,
					-- layer=2 filter=162 channel=16
					-29, -56, -44, 0, 6, -10, 16, 9, 15,
					-- layer=2 filter=162 channel=17
					0, -6, -6, 12, 3, 10, 7, -7, 7,
					-- layer=2 filter=162 channel=18
					59, 28, 12, 7, 10, -6, -10, -11, 52,
					-- layer=2 filter=162 channel=19
					-19, -57, -21, 27, 6, -23, -3, 14, 16,
					-- layer=2 filter=162 channel=20
					9, 2, -2, 1, 11, -9, 5, 0, -3,
					-- layer=2 filter=162 channel=21
					-7, 9, 1, 10, 0, 5, 9, 3, 10,
					-- layer=2 filter=162 channel=22
					3, -2, -8, 6, 4, 8, -9, 4, 7,
					-- layer=2 filter=162 channel=23
					29, -25, -42, 25, -5, 12, 40, 28, 13,
					-- layer=2 filter=162 channel=24
					-20, -22, 24, 6, -27, -18, 35, -11, -7,
					-- layer=2 filter=162 channel=25
					6, 13, 20, -38, -37, -9, -6, -20, -38,
					-- layer=2 filter=162 channel=26
					3, -3, -6, 6, 4, 2, 2, 3, 9,
					-- layer=2 filter=162 channel=27
					-24, -7, 13, -2, 1, -1, 9, -13, -14,
					-- layer=2 filter=162 channel=28
					18, 24, -17, -9, -2, 3, 40, 15, 20,
					-- layer=2 filter=162 channel=29
					7, -1, 5, 6, 3, -6, -10, 4, -3,
					-- layer=2 filter=162 channel=30
					-14, 10, -27, 19, -20, 7, -1, -20, 21,
					-- layer=2 filter=162 channel=31
					-36, -23, -5, 72, 45, 30, 0, -30, -12,
					-- layer=2 filter=162 channel=32
					0, 2, 6, -3, -9, -2, -9, 8, -7,
					-- layer=2 filter=162 channel=33
					-6, -13, -21, 21, -49, -48, -12, 2, -17,
					-- layer=2 filter=162 channel=34
					8, -45, -102, -1, 2, -33, 6, 15, 43,
					-- layer=2 filter=162 channel=35
					17, 9, 10, -33, -19, 1, 16, -17, -10,
					-- layer=2 filter=162 channel=36
					1, 0, 10, 6, -10, 5, -10, 0, -9,
					-- layer=2 filter=162 channel=37
					25, 8, 5, 31, 0, 22, 12, -9, 0,
					-- layer=2 filter=162 channel=38
					26, 0, -7, 0, 8, 28, -3, -1, -18,
					-- layer=2 filter=162 channel=39
					5, -19, -23, 55, 17, -24, -17, 38, 0,
					-- layer=2 filter=162 channel=40
					59, -27, -63, -24, 4, 0, -13, 2, 65,
					-- layer=2 filter=162 channel=41
					0, -1, -5, 4, -1, -4, -1, -2, 9,
					-- layer=2 filter=162 channel=42
					12, -6, -32, 4, 36, 13, 35, 19, 16,
					-- layer=2 filter=162 channel=43
					0, -43, -19, -2, -25, -64, 42, -16, 20,
					-- layer=2 filter=162 channel=44
					-3, 6, -3, 0, 2, 7, 4, -7, -1,
					-- layer=2 filter=162 channel=45
					-10, 3, 21, -18, -24, -26, -12, -2, -49,
					-- layer=2 filter=162 channel=46
					-4, -33, -19, 2, -32, -38, 0, -32, -47,
					-- layer=2 filter=162 channel=47
					3, 23, -8, -5, -76, -40, 31, 46, 22,
					-- layer=2 filter=162 channel=48
					0, 6, -9, -7, 11, 6, -10, -11, -5,
					-- layer=2 filter=162 channel=49
					21, 40, -10, 23, 0, 14, 13, 24, 35,
					-- layer=2 filter=162 channel=50
					-11, -20, -5, -6, 29, 19, 16, 17, 31,
					-- layer=2 filter=162 channel=51
					24, 12, -3, 17, -4, 17, 9, 13, 0,
					-- layer=2 filter=162 channel=52
					25, -7, 5, 25, -33, -24, 41, 19, 35,
					-- layer=2 filter=162 channel=53
					-21, 7, -118, -20, -22, -40, -58, -17, -15,
					-- layer=2 filter=162 channel=54
					24, 15, 6, 8, -38, -12, 14, 32, 32,
					-- layer=2 filter=162 channel=55
					4, -7, -8, 3, -1, -2, 3, 0, -11,
					-- layer=2 filter=162 channel=56
					27, 4, -5, 24, 3, 12, -2, -28, -6,
					-- layer=2 filter=162 channel=57
					-3, -11, -6, -4, 7, -7, 3, -11, -5,
					-- layer=2 filter=162 channel=58
					35, 53, 21, 0, 21, 45, 20, -16, 20,
					-- layer=2 filter=162 channel=59
					-31, -51, -21, 4, 20, 14, -11, 19, -6,
					-- layer=2 filter=162 channel=60
					3, 11, 13, 8, 13, 25, -6, 43, 0,
					-- layer=2 filter=162 channel=61
					-1, 36, 54, -27, -20, 41, -23, 14, -4,
					-- layer=2 filter=162 channel=62
					-29, -30, -52, 0, 6, 21, -22, 20, 69,
					-- layer=2 filter=162 channel=63
					-9, -10, -7, 24, -21, -17, 26, 28, 0,
					-- layer=2 filter=162 channel=64
					-7, -25, -20, 13, 7, 11, 42, 38, 9,
					-- layer=2 filter=162 channel=65
					2, 11, 11, -20, 10, 36, -15, 40, 4,
					-- layer=2 filter=162 channel=66
					16, 17, 44, 37, 19, -1, 36, 14, 27,
					-- layer=2 filter=162 channel=67
					-19, -53, -22, 3, -3, -50, -16, -44, -3,
					-- layer=2 filter=162 channel=68
					5, -7, 0, 8, 2, -7, 1, 2, -1,
					-- layer=2 filter=162 channel=69
					-9, -4, -32, 3, 5, -5, 46, 34, 27,
					-- layer=2 filter=162 channel=70
					47, 27, 2, -22, 16, -4, 4, 8, -10,
					-- layer=2 filter=162 channel=71
					-16, -24, 0, 0, 16, 10, -26, -51, -12,
					-- layer=2 filter=162 channel=72
					17, 20, 23, 5, 12, 7, 19, 31, 11,
					-- layer=2 filter=162 channel=73
					35, 16, -17, 22, 12, -25, -23, 8, -11,
					-- layer=2 filter=162 channel=74
					5, 7, 7, 20, 28, -13, 7, -7, -32,
					-- layer=2 filter=162 channel=75
					-18, 0, -6, 2, 5, -4, -3, 12, 17,
					-- layer=2 filter=162 channel=76
					-31, -33, -65, -47, -10, -50, -22, -12, -1,
					-- layer=2 filter=162 channel=77
					7, 0, -7, 0, 3, -5, 5, 5, -9,
					-- layer=2 filter=162 channel=78
					31, -6, 5, 6, -30, 0, 8, -12, 0,
					-- layer=2 filter=162 channel=79
					7, 11, -1, -7, 8, -2, -5, 7, -6,
					-- layer=2 filter=162 channel=80
					-7, -36, -15, 0, 1, -70, -10, 3, -22,
					-- layer=2 filter=162 channel=81
					1, -1, 3, 6, 10, -1, -2, 3, -9,
					-- layer=2 filter=162 channel=82
					6, 1, 9, 0, 6, 5, -4, 3, 4,
					-- layer=2 filter=162 channel=83
					-21, -10, 0, -33, 17, 0, 9, 2, 3,
					-- layer=2 filter=162 channel=84
					1, 5, -6, 6, 8, 5, 2, 5, 8,
					-- layer=2 filter=162 channel=85
					4, 13, 1, 5, -7, 0, 3, 13, 0,
					-- layer=2 filter=162 channel=86
					2, 6, -17, 8, 12, 20, -6, 1, -11,
					-- layer=2 filter=162 channel=87
					-4, -25, -116, 1, -35, -39, -6, -27, 26,
					-- layer=2 filter=162 channel=88
					-22, -7, -2, -3, -2, 40, 15, 0, 0,
					-- layer=2 filter=162 channel=89
					-26, 2, -10, 4, 10, 30, -8, 0, 27,
					-- layer=2 filter=162 channel=90
					-6, 0, 7, 5, 2, -5, 10, -11, 4,
					-- layer=2 filter=162 channel=91
					-8, 17, 0, -10, 3, -20, -11, 9, -21,
					-- layer=2 filter=162 channel=92
					-12, 24, 24, -24, -4, 3, 6, 4, 19,
					-- layer=2 filter=162 channel=93
					-3, -45, -66, -9, 42, -7, -25, -50, -11,
					-- layer=2 filter=162 channel=94
					-51, 22, -12, -19, -14, -13, -13, 36, 15,
					-- layer=2 filter=162 channel=95
					14, 14, 4, 14, 11, 12, 14, 0, 16,
					-- layer=2 filter=162 channel=96
					30, -10, -66, 14, 0, -11, -28, -1, 8,
					-- layer=2 filter=162 channel=97
					34, -3, 22, 16, 1, -13, 10, 16, -1,
					-- layer=2 filter=162 channel=98
					18, 36, 3, -44, -38, -32, 34, 25, 10,
					-- layer=2 filter=162 channel=99
					10, -36, -37, 3, 5, 13, 17, 20, 2,
					-- layer=2 filter=162 channel=100
					15, -8, -41, 13, 15, 17, -8, 2, -5,
					-- layer=2 filter=162 channel=101
					-19, -14, 7, -28, -1, -13, -2, -23, -27,
					-- layer=2 filter=162 channel=102
					59, -15, 10, 8, -12, -25, 14, 10, 24,
					-- layer=2 filter=162 channel=103
					-52, 29, -3, -13, -7, -28, -13, -23, -33,
					-- layer=2 filter=162 channel=104
					-8, -3, -40, -5, -6, 14, -26, -13, 19,
					-- layer=2 filter=162 channel=105
					-54, -21, -37, -24, -16, 12, -14, 10, -6,
					-- layer=2 filter=162 channel=106
					-20, 19, -9, -1, 4, -37, -18, -23, -53,
					-- layer=2 filter=162 channel=107
					8, 5, 7, -46, 1, -13, -43, -25, -3,
					-- layer=2 filter=162 channel=108
					-26, -19, 25, -8, 0, 19, -14, -11, 18,
					-- layer=2 filter=162 channel=109
					5, 2, -3, -7, -4, 0, -7, -5, -6,
					-- layer=2 filter=162 channel=110
					4, -26, -1, 29, 32, 21, 35, 29, 23,
					-- layer=2 filter=162 channel=111
					0, 3, 7, 5, 8, -9, -2, 4, -1,
					-- layer=2 filter=162 channel=112
					-8, 28, 42, -3, -3, 13, -1, -14, -4,
					-- layer=2 filter=162 channel=113
					-11, 21, 11, -10, -13, 27, 17, 10, 15,
					-- layer=2 filter=162 channel=114
					7, -1, 0, -9, -1, -4, 9, 5, -7,
					-- layer=2 filter=162 channel=115
					-4, 0, 3, 2, 14, 5, -9, -5, 5,
					-- layer=2 filter=162 channel=116
					21, -18, -62, 14, -31, -35, 37, -8, 36,
					-- layer=2 filter=162 channel=117
					-31, -4, 28, -23, -8, -65, 19, -4, 27,
					-- layer=2 filter=162 channel=118
					0, -30, -44, 4, -38, -51, 8, 14, 3,
					-- layer=2 filter=162 channel=119
					0, -3, 0, -28, 3, -27, 17, -4, -3,
					-- layer=2 filter=162 channel=120
					-2, -2, 1, 2, 10, -5, 8, 0, 7,
					-- layer=2 filter=162 channel=121
					-6, 1, 7, 7, 8, -1, 11, -7, -3,
					-- layer=2 filter=162 channel=122
					10, 8, 7, 0, 9, 15, -10, 1, -7,
					-- layer=2 filter=162 channel=123
					-20, 5, -5, 26, -9, -12, 17, 52, 15,
					-- layer=2 filter=162 channel=124
					-5, -54, -26, 14, 0, 1, 12, 16, 20,
					-- layer=2 filter=162 channel=125
					-7, -7, -1, -2, 8, -4, 0, -1, -4,
					-- layer=2 filter=162 channel=126
					32, -33, -38, 34, -69, 13, -91, 17, 16,
					-- layer=2 filter=162 channel=127
					10, 40, -5, -18, 8, 2, 3, 34, 21,
					-- layer=2 filter=163 channel=0
					20, -18, 17, 4, 0, 12, 8, 9, 1,
					-- layer=2 filter=163 channel=1
					-8, 18, 16, 9, 22, 6, -15, 30, -5,
					-- layer=2 filter=163 channel=2
					-3, 4, -10, 4, -2, 6, 8, -6, -5,
					-- layer=2 filter=163 channel=3
					18, -17, -16, -11, -11, -24, 34, 28, 31,
					-- layer=2 filter=163 channel=4
					21, 17, -1, 35, -28, 28, 1, -4, -9,
					-- layer=2 filter=163 channel=5
					0, -14, 0, -8, -9, 16, -15, -38, -20,
					-- layer=2 filter=163 channel=6
					-10, 1, 3, -22, -14, -47, -42, -27, -35,
					-- layer=2 filter=163 channel=7
					52, -30, 13, 46, 33, 43, 49, 39, 50,
					-- layer=2 filter=163 channel=8
					0, 7, 3, 1, -4, 0, 3, 3, 1,
					-- layer=2 filter=163 channel=9
					28, 5, 15, -29, -36, -48, 12, 7, -32,
					-- layer=2 filter=163 channel=10
					5, -24, 4, 9, -10, -26, 17, 6, 17,
					-- layer=2 filter=163 channel=11
					9, 3, 6, 2, 1, 1, -6, 0, -2,
					-- layer=2 filter=163 channel=12
					-11, 8, 22, 34, 28, 26, 1, 56, 29,
					-- layer=2 filter=163 channel=13
					-2, 7, 3, -5, -1, -6, 7, 6, 0,
					-- layer=2 filter=163 channel=14
					-7, -13, 9, -1, 8, 0, -9, 21, 8,
					-- layer=2 filter=163 channel=15
					6, 15, 1, -7, -14, 48, 36, 11, 23,
					-- layer=2 filter=163 channel=16
					-24, 7, -25, -48, -30, -33, -30, -22, 3,
					-- layer=2 filter=163 channel=17
					-8, -5, -6, 2, 8, 3, 0, 4, 10,
					-- layer=2 filter=163 channel=18
					-35, 11, 13, -14, -24, 29, 7, -13, 4,
					-- layer=2 filter=163 channel=19
					17, 26, 8, -11, 33, 11, 14, 26, 11,
					-- layer=2 filter=163 channel=20
					7, 3, -7, 5, -2, 2, 6, 3, -10,
					-- layer=2 filter=163 channel=21
					2, -2, -15, -5, 11, -8, 8, -1, 9,
					-- layer=2 filter=163 channel=22
					7, -1, 5, 6, -8, -5, -7, -11, 2,
					-- layer=2 filter=163 channel=23
					3, -6, 1, 0, 2, 1, -2, 18, -21,
					-- layer=2 filter=163 channel=24
					7, -9, -24, 1, -5, -18, 30, 10, 34,
					-- layer=2 filter=163 channel=25
					-5, -25, -80, 16, -8, -37, 11, 11, -1,
					-- layer=2 filter=163 channel=26
					-8, 0, -5, -4, 0, 10, -4, -7, -11,
					-- layer=2 filter=163 channel=27
					22, 0, 5, 0, 2, 5, -2, -9, -2,
					-- layer=2 filter=163 channel=28
					-15, -24, -20, -3, 15, 31, -11, 19, 19,
					-- layer=2 filter=163 channel=29
					8, 8, -6, 0, -8, 1, 8, -7, 5,
					-- layer=2 filter=163 channel=30
					-22, -2, -2, -19, -22, -4, 3, -5, 0,
					-- layer=2 filter=163 channel=31
					6, -13, -4, -8, 9, -51, -8, 13, -28,
					-- layer=2 filter=163 channel=32
					8, 7, 5, 8, 4, -7, -9, -4, 1,
					-- layer=2 filter=163 channel=33
					39, -2, -18, 12, -3, 35, -21, 7, 13,
					-- layer=2 filter=163 channel=34
					-33, 8, 17, -69, -7, -8, -59, -47, 19,
					-- layer=2 filter=163 channel=35
					2, -13, 26, 0, -1, 16, -4, 16, 28,
					-- layer=2 filter=163 channel=36
					1, 6, -4, 16, 0, 6, 2, 11, 2,
					-- layer=2 filter=163 channel=37
					-4, 10, 19, 3, 4, -7, -10, -13, -1,
					-- layer=2 filter=163 channel=38
					-9, -4, 10, -9, 0, 30, 8, 0, -24,
					-- layer=2 filter=163 channel=39
					14, -6, 1, -12, -8, 3, -31, -29, 26,
					-- layer=2 filter=163 channel=40
					-5, -5, -27, -20, -58, -7, 43, -24, -10,
					-- layer=2 filter=163 channel=41
					-7, -8, -8, -11, 10, 0, -10, -10, 7,
					-- layer=2 filter=163 channel=42
					21, 17, 6, -12, -13, -3, -10, -2, -14,
					-- layer=2 filter=163 channel=43
					-41, -34, -27, -28, -41, -18, 13, 19, 29,
					-- layer=2 filter=163 channel=44
					0, 5, 7, -13, 6, -7, -3, -2, -8,
					-- layer=2 filter=163 channel=45
					30, 8, -16, 4, 3, 1, 31, 4, -14,
					-- layer=2 filter=163 channel=46
					-37, -5, 3, 4, -17, -8, 26, -5, -30,
					-- layer=2 filter=163 channel=47
					-4, 40, 20, 28, 44, 49, -2, 23, 25,
					-- layer=2 filter=163 channel=48
					1, 2, 0, -8, 3, -6, -10, 6, -6,
					-- layer=2 filter=163 channel=49
					11, 33, -7, 20, -48, -9, 57, 22, 29,
					-- layer=2 filter=163 channel=50
					-14, -8, 1, 6, 14, 7, -9, 15, 18,
					-- layer=2 filter=163 channel=51
					3, -16, 13, 0, -12, -12, -13, -7, -14,
					-- layer=2 filter=163 channel=52
					15, 20, 24, -18, -14, -1, -40, -4, 19,
					-- layer=2 filter=163 channel=53
					-52, -63, -9, 11, -18, -83, 3, -15, -33,
					-- layer=2 filter=163 channel=54
					8, 10, 27, 35, 17, 42, 13, 23, 6,
					-- layer=2 filter=163 channel=55
					10, -6, 0, 4, -8, -7, -4, -5, -2,
					-- layer=2 filter=163 channel=56
					17, -14, 10, 10, 0, 6, -15, -18, -1,
					-- layer=2 filter=163 channel=57
					12, -2, -3, 10, 1, 7, 1, -2, -8,
					-- layer=2 filter=163 channel=58
					-18, 9, 2, 23, 39, 48, 18, 52, 45,
					-- layer=2 filter=163 channel=59
					-8, -30, 6, -42, 8, -13, -1, 5, 49,
					-- layer=2 filter=163 channel=60
					-28, 10, 13, -13, 1, 47, -3, 23, -9,
					-- layer=2 filter=163 channel=61
					2, -16, -16, -4, -48, -6, 7, 18, -44,
					-- layer=2 filter=163 channel=62
					2, 34, 23, -10, 19, 19, 0, -12, 37,
					-- layer=2 filter=163 channel=63
					10, 18, 16, -9, 0, 2, -8, 0, -1,
					-- layer=2 filter=163 channel=64
					-5, 7, 23, -6, 14, -21, 17, 18, 8,
					-- layer=2 filter=163 channel=65
					-29, -13, 2, -6, -36, 13, -38, 12, -25,
					-- layer=2 filter=163 channel=66
					-14, 9, 8, 21, -20, 9, 62, 5, 6,
					-- layer=2 filter=163 channel=67
					11, -13, -18, -34, -48, -59, 22, 16, 2,
					-- layer=2 filter=163 channel=68
					1, 1, 7, -8, -6, -5, -3, 8, 4,
					-- layer=2 filter=163 channel=69
					0, 17, 21, -6, -2, -14, -19, -4, 0,
					-- layer=2 filter=163 channel=70
					-4, -28, 6, 16, 19, 17, 6, 16, 36,
					-- layer=2 filter=163 channel=71
					-5, 3, -21, 11, 2, 20, 20, 17, 26,
					-- layer=2 filter=163 channel=72
					8, -19, 2, 7, -4, 30, 19, 17, 30,
					-- layer=2 filter=163 channel=73
					8, -16, -11, 29, 16, -45, 15, -9, -8,
					-- layer=2 filter=163 channel=74
					17, -19, 2, -15, -19, -25, 22, -6, -5,
					-- layer=2 filter=163 channel=75
					-44, 5, 11, 14, 21, -21, -13, 14, 35,
					-- layer=2 filter=163 channel=76
					-29, -44, 26, -6, 9, -24, 6, 18, -37,
					-- layer=2 filter=163 channel=77
					-5, 13, 5, 3, -11, -9, 0, 0, -8,
					-- layer=2 filter=163 channel=78
					7, -17, -2, -8, -16, -2, 12, -3, 15,
					-- layer=2 filter=163 channel=79
					1, -8, 6, 6, 8, -8, -9, 0, -7,
					-- layer=2 filter=163 channel=80
					-13, 6, -10, 2, -2, -19, 5, -5, -6,
					-- layer=2 filter=163 channel=81
					8, 9, 23, 11, 11, 12, 15, 14, 11,
					-- layer=2 filter=163 channel=82
					3, -2, -3, 2, -5, -8, 11, -3, 5,
					-- layer=2 filter=163 channel=83
					-38, -13, -4, -7, 3, -3, -3, 16, -4,
					-- layer=2 filter=163 channel=84
					4, 3, 5, 0, -2, 1, 6, -4, 2,
					-- layer=2 filter=163 channel=85
					6, 2, 4, 4, 1, 6, 11, 0, 11,
					-- layer=2 filter=163 channel=86
					-12, 18, 7, 1, 3, 12, 7, -1, 4,
					-- layer=2 filter=163 channel=87
					-21, -23, 27, -45, -31, 37, -8, -33, -21,
					-- layer=2 filter=163 channel=88
					3, 30, 43, -10, -17, -9, -5, -7, -11,
					-- layer=2 filter=163 channel=89
					-18, -30, -1, -5, 0, -5, -10, 49, 31,
					-- layer=2 filter=163 channel=90
					-7, 1, 0, 9, 10, 10, 8, 2, 2,
					-- layer=2 filter=163 channel=91
					-14, 0, 8, 2, -9, 17, -7, 36, 29,
					-- layer=2 filter=163 channel=92
					4, 3, 11, 6, 13, 27, 11, 37, 14,
					-- layer=2 filter=163 channel=93
					-10, -1, -29, -17, 13, 25, -34, -16, 36,
					-- layer=2 filter=163 channel=94
					-18, -42, -32, -12, -47, -20, -35, 14, -58,
					-- layer=2 filter=163 channel=95
					1, 6, 3, 3, 0, -3, 10, -7, 5,
					-- layer=2 filter=163 channel=96
					18, -52, -22, -19, -9, -11, -60, -43, -30,
					-- layer=2 filter=163 channel=97
					16, 17, 7, -6, -44, -4, 20, 6, 4,
					-- layer=2 filter=163 channel=98
					2, 7, -1, 26, 35, 30, 0, 16, 13,
					-- layer=2 filter=163 channel=99
					2, -1, 40, -8, -11, -24, -12, 0, -35,
					-- layer=2 filter=163 channel=100
					-16, -12, -11, -22, -10, -2, 12, 5, 2,
					-- layer=2 filter=163 channel=101
					-12, -9, -28, 14, -8, -22, -11, 11, -2,
					-- layer=2 filter=163 channel=102
					-17, -19, 21, 2, -46, 36, -39, -29, -18,
					-- layer=2 filter=163 channel=103
					-3, -38, -10, -44, -48, -64, -21, 21, 2,
					-- layer=2 filter=163 channel=104
					-39, -8, -19, 11, -54, 8, -4, -33, -23,
					-- layer=2 filter=163 channel=105
					-9, -20, 35, -35, 8, -26, 24, 8, 26,
					-- layer=2 filter=163 channel=106
					-26, -26, -34, 1, -5, -36, -2, 7, -1,
					-- layer=2 filter=163 channel=107
					13, -12, -3, 9, -38, 1, 6, 10, -40,
					-- layer=2 filter=163 channel=108
					6, 16, 16, -19, -19, 10, -23, -22, -34,
					-- layer=2 filter=163 channel=109
					-3, -7, 9, -6, 0, 3, -5, -10, -4,
					-- layer=2 filter=163 channel=110
					-22, 13, 0, -17, 4, 13, 10, 14, -11,
					-- layer=2 filter=163 channel=111
					7, 3, 0, 8, -1, -4, -4, 5, -3,
					-- layer=2 filter=163 channel=112
					-16, 11, 3, -17, -45, -18, 2, 13, -28,
					-- layer=2 filter=163 channel=113
					-20, -4, -12, 5, 7, -6, -8, -1, 14,
					-- layer=2 filter=163 channel=114
					0, 12, 2, -10, -13, -17, -11, -12, -14,
					-- layer=2 filter=163 channel=115
					11, -8, 3, 4, -13, 8, -4, -8, 5,
					-- layer=2 filter=163 channel=116
					-18, -24, 22, -60, -33, 58, -27, -30, 2,
					-- layer=2 filter=163 channel=117
					14, -53, -21, 30, -14, 48, 42, 35, 9,
					-- layer=2 filter=163 channel=118
					13, 5, 8, 3, -16, 12, 13, 3, 21,
					-- layer=2 filter=163 channel=119
					-26, 50, 25, 11, -2, 18, -5, -7, -18,
					-- layer=2 filter=163 channel=120
					-3, 8, 3, 3, -7, -7, 0, 10, -3,
					-- layer=2 filter=163 channel=121
					-1, 6, 7, -6, 2, 8, 3, 1, 3,
					-- layer=2 filter=163 channel=122
					-1, -8, -10, 3, -16, -7, -14, -14, 3,
					-- layer=2 filter=163 channel=123
					18, -11, -6, 17, 21, 29, 23, 17, 34,
					-- layer=2 filter=163 channel=124
					-24, -27, -13, -48, -2, 16, 20, 19, -3,
					-- layer=2 filter=163 channel=125
					2, 0, 0, 3, 10, -2, 5, -2, -3,
					-- layer=2 filter=163 channel=126
					-6, 15, -12, -47, -3, -4, -51, 11, -12,
					-- layer=2 filter=163 channel=127
					-2, 20, 2, 7, -11, 11, -17, -4, 12,
					-- layer=2 filter=164 channel=0
					7, -20, -19, 1, 9, -1, -4, -6, -4,
					-- layer=2 filter=164 channel=1
					-22, -1, -20, 0, -11, -4, -17, -14, -10,
					-- layer=2 filter=164 channel=2
					2, 7, -6, 0, -8, 8, -3, 3, 6,
					-- layer=2 filter=164 channel=3
					-11, -12, -8, -3, 0, -19, -8, -5, 0,
					-- layer=2 filter=164 channel=4
					-5, 5, 20, 10, -5, 0, 10, 1, 17,
					-- layer=2 filter=164 channel=5
					-9, -9, -23, -4, 0, -5, -7, -1, -18,
					-- layer=2 filter=164 channel=6
					-11, -16, 17, -3, -10, 10, 7, -12, 8,
					-- layer=2 filter=164 channel=7
					-17, 0, -14, 9, -6, -14, -14, 0, -10,
					-- layer=2 filter=164 channel=8
					-9, -7, -7, -2, 4, 2, -9, -7, -11,
					-- layer=2 filter=164 channel=9
					-7, -13, -15, -6, -13, -8, -15, 7, 0,
					-- layer=2 filter=164 channel=10
					-12, 0, -15, -14, -1, 0, -14, 1, -1,
					-- layer=2 filter=164 channel=11
					0, 5, -9, -8, 0, -8, -3, -7, -3,
					-- layer=2 filter=164 channel=12
					-7, -12, -15, -26, -22, 2, -17, -8, -10,
					-- layer=2 filter=164 channel=13
					3, -6, -3, -8, 0, 4, -10, 4, 4,
					-- layer=2 filter=164 channel=14
					-14, -5, -6, -8, -12, -12, -11, -10, -19,
					-- layer=2 filter=164 channel=15
					-8, -26, 15, -13, -17, -7, -22, 0, -12,
					-- layer=2 filter=164 channel=16
					-4, -6, -17, 0, 0, -12, 10, 0, -14,
					-- layer=2 filter=164 channel=17
					8, -5, 7, -2, 8, 2, -3, -1, -5,
					-- layer=2 filter=164 channel=18
					-11, -10, 7, -13, -2, -14, -3, -6, -7,
					-- layer=2 filter=164 channel=19
					-11, 2, -27, -8, -21, 6, -27, -14, -19,
					-- layer=2 filter=164 channel=20
					-9, 1, 8, 2, 0, -11, -5, -7, 9,
					-- layer=2 filter=164 channel=21
					-7, -10, 3, -9, -2, -5, 4, -10, 3,
					-- layer=2 filter=164 channel=22
					-8, 9, 0, 0, 3, -3, 1, 7, -9,
					-- layer=2 filter=164 channel=23
					6, -3, 0, -3, -2, -5, 14, 0, -2,
					-- layer=2 filter=164 channel=24
					-22, -5, 3, -19, -19, -10, -12, 2, 1,
					-- layer=2 filter=164 channel=25
					-1, -22, -7, -12, -21, -12, -7, -3, -8,
					-- layer=2 filter=164 channel=26
					1, -1, -10, -5, -6, 2, -9, -3, -8,
					-- layer=2 filter=164 channel=27
					-3, -6, -13, -7, 1, -16, -18, -8, 0,
					-- layer=2 filter=164 channel=28
					11, -1, -6, 7, 7, -21, -8, 8, 6,
					-- layer=2 filter=164 channel=29
					4, -1, 6, -10, 4, 0, 5, 4, 2,
					-- layer=2 filter=164 channel=30
					3, -13, -6, 4, -5, -7, -3, 2, -3,
					-- layer=2 filter=164 channel=31
					-4, -3, 30, -28, -15, 22, -28, -12, 11,
					-- layer=2 filter=164 channel=32
					4, 5, 8, -10, -3, 2, -12, 6, 0,
					-- layer=2 filter=164 channel=33
					-8, 4, 2, -10, -18, -21, -9, 7, -18,
					-- layer=2 filter=164 channel=34
					-6, -16, 2, -12, -5, -17, -8, -11, -4,
					-- layer=2 filter=164 channel=35
					-6, -6, 2, -1, 0, -25, -6, -1, -1,
					-- layer=2 filter=164 channel=36
					1, -3, -4, 1, -8, 1, -1, 8, 7,
					-- layer=2 filter=164 channel=37
					-19, -11, -1, -15, -8, -12, -6, 0, -14,
					-- layer=2 filter=164 channel=38
					0, -12, -11, -8, -16, -13, 1, -22, -22,
					-- layer=2 filter=164 channel=39
					-22, -4, -21, -6, 6, -9, -7, -7, 1,
					-- layer=2 filter=164 channel=40
					14, 0, 40, -25, -17, 4, -21, -9, 1,
					-- layer=2 filter=164 channel=41
					-2, 7, -1, -9, -12, 8, 6, -6, -5,
					-- layer=2 filter=164 channel=42
					-13, 4, 22, -11, -13, -2, -3, -2, 2,
					-- layer=2 filter=164 channel=43
					-11, -31, 2, -4, -10, -14, -11, -18, -10,
					-- layer=2 filter=164 channel=44
					-1, -2, -7, 3, -1, 5, 6, -1, -5,
					-- layer=2 filter=164 channel=45
					-8, -21, -15, -31, -14, -4, -9, -19, -19,
					-- layer=2 filter=164 channel=46
					-2, -6, -16, 4, 2, -14, 10, 3, -17,
					-- layer=2 filter=164 channel=47
					8, -12, 0, -6, -5, -13, -24, -4, 7,
					-- layer=2 filter=164 channel=48
					3, 7, -8, 0, 7, -10, -5, 6, 8,
					-- layer=2 filter=164 channel=49
					-18, -15, 12, 3, -20, 7, 0, -14, 7,
					-- layer=2 filter=164 channel=50
					3, 6, -5, 1, 2, -7, -4, 8, -6,
					-- layer=2 filter=164 channel=51
					-10, -17, -13, -15, -10, -11, -16, -12, -13,
					-- layer=2 filter=164 channel=52
					-20, 10, -1, -8, -13, -21, -16, -9, -8,
					-- layer=2 filter=164 channel=53
					-4, -7, 15, 0, -16, 33, 1, 0, 21,
					-- layer=2 filter=164 channel=54
					-5, 7, 12, 0, -14, 4, -11, -5, -3,
					-- layer=2 filter=164 channel=55
					-9, -5, -6, -9, -8, -2, 5, 3, -6,
					-- layer=2 filter=164 channel=56
					-2, -1, 0, -3, 0, -15, -8, -2, -11,
					-- layer=2 filter=164 channel=57
					7, 8, -1, -8, -5, 8, -9, -3, 6,
					-- layer=2 filter=164 channel=58
					0, -11, -20, -28, 0, -1, -14, -8, -20,
					-- layer=2 filter=164 channel=59
					-1, 8, -33, -30, -16, -27, -13, -17, -13,
					-- layer=2 filter=164 channel=60
					4, -11, -14, 10, -11, 0, -12, 2, -10,
					-- layer=2 filter=164 channel=61
					0, -9, -16, 5, 11, -8, 9, 16, 12,
					-- layer=2 filter=164 channel=62
					-5, 4, 7, -10, -2, 5, 0, -3, 4,
					-- layer=2 filter=164 channel=63
					-1, -5, -11, 1, -5, -17, 2, 12, -7,
					-- layer=2 filter=164 channel=64
					3, 1, 12, 0, -6, 12, 10, 11, -7,
					-- layer=2 filter=164 channel=65
					14, 0, -1, -11, -16, 3, -2, -26, 15,
					-- layer=2 filter=164 channel=66
					25, -7, 0, 0, -27, -27, 15, -27, 21,
					-- layer=2 filter=164 channel=67
					-13, -4, -17, -10, -16, -17, -13, -17, 1,
					-- layer=2 filter=164 channel=68
					-5, -7, 4, 0, -10, 6, 5, -11, -4,
					-- layer=2 filter=164 channel=69
					3, -11, 8, -7, 2, 10, 3, 11, 6,
					-- layer=2 filter=164 channel=70
					-13, -5, -16, -17, -12, -14, 3, 5, -12,
					-- layer=2 filter=164 channel=71
					-15, -26, -15, -4, -8, -6, -10, -10, -10,
					-- layer=2 filter=164 channel=72
					-27, -5, 14, -9, -22, -22, -1, -4, -3,
					-- layer=2 filter=164 channel=73
					-7, -2, -14, -8, -6, -5, -6, 0, -8,
					-- layer=2 filter=164 channel=74
					3, -6, -14, -17, 4, 0, -7, -12, -6,
					-- layer=2 filter=164 channel=75
					-10, -3, -1, -13, -19, -19, -8, -7, -20,
					-- layer=2 filter=164 channel=76
					-11, 27, 20, 22, 2, 9, 0, 22, 12,
					-- layer=2 filter=164 channel=77
					-5, -8, -6, 8, 2, -11, 3, 10, 5,
					-- layer=2 filter=164 channel=78
					-21, -11, 0, -15, -5, -1, -3, -8, -6,
					-- layer=2 filter=164 channel=79
					-10, -7, -8, -7, -1, -9, -10, -9, 7,
					-- layer=2 filter=164 channel=80
					-6, -19, 12, -4, 0, 13, -12, -7, -2,
					-- layer=2 filter=164 channel=81
					-11, -4, -7, 9, 7, 8, -10, 0, -9,
					-- layer=2 filter=164 channel=82
					-6, 7, 7, 5, 3, 0, 6, 7, 8,
					-- layer=2 filter=164 channel=83
					8, -22, 5, -3, -1, 21, 15, 14, 1,
					-- layer=2 filter=164 channel=84
					-6, 9, -10, 6, 0, -1, 4, 7, 0,
					-- layer=2 filter=164 channel=85
					-5, -1, 2, -5, -10, 6, -5, 4, 6,
					-- layer=2 filter=164 channel=86
					-3, 4, 10, 0, -8, -2, 0, -3, -4,
					-- layer=2 filter=164 channel=87
					0, -16, 7, -4, -27, -6, -5, -11, -3,
					-- layer=2 filter=164 channel=88
					5, -4, -7, -6, -4, 5, -2, -3, 8,
					-- layer=2 filter=164 channel=89
					-10, 4, 0, -8, -19, -1, -14, -6, -6,
					-- layer=2 filter=164 channel=90
					3, 0, -1, -4, 10, 0, 9, 4, -7,
					-- layer=2 filter=164 channel=91
					-8, 0, -14, -34, -15, -11, -8, -10, -15,
					-- layer=2 filter=164 channel=92
					-22, 4, -8, -22, -3, 1, -16, -28, 3,
					-- layer=2 filter=164 channel=93
					7, -11, -1, 0, 0, 8, 4, -37, 5,
					-- layer=2 filter=164 channel=94
					7, 12, 9, 0, -7, -1, -6, 7, 18,
					-- layer=2 filter=164 channel=95
					2, -8, 2, -4, -3, 2, 0, 3, 7,
					-- layer=2 filter=164 channel=96
					6, -1, -22, 4, -4, -19, 7, 8, 6,
					-- layer=2 filter=164 channel=97
					-21, -5, 16, -13, -10, -3, 0, -13, -9,
					-- layer=2 filter=164 channel=98
					-6, 2, 3, -6, -17, -25, -7, -8, -3,
					-- layer=2 filter=164 channel=99
					1, 2, -5, -21, -5, -10, -4, 6, -10,
					-- layer=2 filter=164 channel=100
					-4, -3, -2, 5, 11, -12, -1, -1, -4,
					-- layer=2 filter=164 channel=101
					-2, -6, 0, -30, -6, 10, -9, -5, -2,
					-- layer=2 filter=164 channel=102
					-22, -1, -12, 13, -9, -5, 4, 14, 2,
					-- layer=2 filter=164 channel=103
					-7, 7, -4, -19, -9, -21, -1, 20, -30,
					-- layer=2 filter=164 channel=104
					-13, 0, 24, 19, -22, 21, 13, 3, 3,
					-- layer=2 filter=164 channel=105
					-8, 18, -27, 13, -7, -11, -9, 2, -17,
					-- layer=2 filter=164 channel=106
					-5, -9, -15, -26, -15, -7, -17, -3, -1,
					-- layer=2 filter=164 channel=107
					0, 1, 16, 4, 15, 20, 35, -8, 4,
					-- layer=2 filter=164 channel=108
					-25, -20, -18, -18, -22, 1, -22, -5, -14,
					-- layer=2 filter=164 channel=109
					-11, -2, -7, -7, 0, 0, -7, 3, -6,
					-- layer=2 filter=164 channel=110
					5, -4, -18, -19, -10, -27, -2, 5, -6,
					-- layer=2 filter=164 channel=111
					6, -8, -3, 0, 3, -6, 0, 1, 1,
					-- layer=2 filter=164 channel=112
					-2, -6, -6, 10, -16, 0, 6, -9, -2,
					-- layer=2 filter=164 channel=113
					5, -15, -16, 6, 2, 4, 18, 2, -2,
					-- layer=2 filter=164 channel=114
					7, -9, 3, 8, -3, 9, 2, 1, 6,
					-- layer=2 filter=164 channel=115
					10, 9, 3, 2, -4, 1, 2, -8, 3,
					-- layer=2 filter=164 channel=116
					-2, -13, -1, -1, -31, 0, 0, 5, -9,
					-- layer=2 filter=164 channel=117
					-3, 19, -4, 3, -13, -15, -12, 1, -14,
					-- layer=2 filter=164 channel=118
					-13, -21, 3, -7, -18, 7, -2, -13, -19,
					-- layer=2 filter=164 channel=119
					-19, 0, -5, -13, -1, 7, -11, -6, 12,
					-- layer=2 filter=164 channel=120
					9, -4, -8, -5, -2, 10, 4, 4, -5,
					-- layer=2 filter=164 channel=121
					4, -8, -1, 1, 2, -11, -10, 4, -6,
					-- layer=2 filter=164 channel=122
					5, -6, -9, 1, -8, -8, -6, 11, -1,
					-- layer=2 filter=164 channel=123
					2, -5, -15, -14, -5, -16, -12, -10, -11,
					-- layer=2 filter=164 channel=124
					-17, -19, 25, -20, -13, 1, 0, 3, -7,
					-- layer=2 filter=164 channel=125
					5, 2, -9, 0, 10, 6, 4, 4, 0,
					-- layer=2 filter=164 channel=126
					-8, 6, -19, 9, 4, -21, 5, 27, 14,
					-- layer=2 filter=164 channel=127
					0, -6, -8, 7, -3, -6, 16, -13, 17,
					-- layer=2 filter=165 channel=0
					-14, -11, -29, -25, 0, -28, -25, -5, 4,
					-- layer=2 filter=165 channel=1
					18, -8, 7, -2, -10, -2, 24, 40, -15,
					-- layer=2 filter=165 channel=2
					-2, 9, -4, 7, -9, -1, -10, 3, 0,
					-- layer=2 filter=165 channel=3
					-21, -9, 21, 3, 0, -19, 4, 5, 17,
					-- layer=2 filter=165 channel=4
					8, 42, -4, -21, -14, -19, -9, -51, -25,
					-- layer=2 filter=165 channel=5
					0, -5, -10, 7, -3, -10, -3, 1, -12,
					-- layer=2 filter=165 channel=6
					-11, 19, 17, 25, 20, 16, 22, 56, 51,
					-- layer=2 filter=165 channel=7
					18, 29, -14, -8, 19, 8, 4, 11, -4,
					-- layer=2 filter=165 channel=8
					7, 4, 5, 7, -12, 0, -7, 9, -3,
					-- layer=2 filter=165 channel=9
					14, 25, 15, 15, 53, 0, 13, -23, -5,
					-- layer=2 filter=165 channel=10
					-14, -24, -15, -31, -21, -19, -29, -15, 5,
					-- layer=2 filter=165 channel=11
					-2, 1, -13, -22, -5, -24, 18, 6, 12,
					-- layer=2 filter=165 channel=12
					10, -23, -4, -14, -10, -8, -4, 30, -34,
					-- layer=2 filter=165 channel=13
					-2, -1, 4, -7, 0, 8, -2, -2, 2,
					-- layer=2 filter=165 channel=14
					-2, -4, -7, -7, 8, -9, -6, 13, -30,
					-- layer=2 filter=165 channel=15
					-30, 30, 20, 39, -57, 4, 4, -19, -12,
					-- layer=2 filter=165 channel=16
					9, 14, 30, 46, 21, 17, -10, -17, -28,
					-- layer=2 filter=165 channel=17
					4, -7, -1, 2, 2, 7, 10, 11, 10,
					-- layer=2 filter=165 channel=18
					-21, 19, 13, -21, -41, -2, 0, -65, -23,
					-- layer=2 filter=165 channel=19
					5, 28, 17, 4, 17, 28, 21, 44, 25,
					-- layer=2 filter=165 channel=20
					1, -8, 0, 4, 11, -1, 5, 0, 0,
					-- layer=2 filter=165 channel=21
					-13, 8, -10, 3, -8, 4, -12, 1, 6,
					-- layer=2 filter=165 channel=22
					-2, 3, -11, -10, -5, -6, -6, -11, 1,
					-- layer=2 filter=165 channel=23
					17, 15, -2, 34, 12, -4, -15, -29, -25,
					-- layer=2 filter=165 channel=24
					4, -9, -5, -19, -4, -1, 0, 26, 32,
					-- layer=2 filter=165 channel=25
					0, 10, 3, -24, 6, 1, 27, 36, 22,
					-- layer=2 filter=165 channel=26
					-8, 9, -7, -9, -3, 7, 0, 0, -4,
					-- layer=2 filter=165 channel=27
					-2, 36, 13, 14, 8, 9, 0, 0, -4,
					-- layer=2 filter=165 channel=28
					4, -6, 10, -19, -27, -16, -23, -22, 9,
					-- layer=2 filter=165 channel=29
					2, -8, -7, 0, -3, 3, -4, 0, -10,
					-- layer=2 filter=165 channel=30
					-8, 29, -17, 18, 4, -12, -31, -36, -24,
					-- layer=2 filter=165 channel=31
					22, -19, 31, -18, -45, -50, 2, 8, 44,
					-- layer=2 filter=165 channel=32
					10, -5, 6, -8, 4, 0, 8, 4, -5,
					-- layer=2 filter=165 channel=33
					0, -23, 0, 47, -10, -1, 39, 3, -3,
					-- layer=2 filter=165 channel=34
					-6, 35, -24, -9, 8, -26, 16, 7, -6,
					-- layer=2 filter=165 channel=35
					14, 19, 4, -5, 43, -19, -4, -19, -11,
					-- layer=2 filter=165 channel=36
					-3, 2, 8, 0, -1, 9, -5, -9, -6,
					-- layer=2 filter=165 channel=37
					0, 0, 10, -2, 0, -6, 18, -3, -1,
					-- layer=2 filter=165 channel=38
					-10, 25, 31, 28, -19, 12, -9, -8, 0,
					-- layer=2 filter=165 channel=39
					17, 29, 12, 20, 21, 17, -20, -23, -31,
					-- layer=2 filter=165 channel=40
					-15, 14, 38, 22, 0, -4, -5, 35, -4,
					-- layer=2 filter=165 channel=41
					6, -6, 2, 0, 8, -6, 0, -7, 9,
					-- layer=2 filter=165 channel=42
					5, 14, 25, 49, 5, 14, -46, -13, -47,
					-- layer=2 filter=165 channel=43
					-15, -13, -17, -23, 26, -32, 4, 9, -25,
					-- layer=2 filter=165 channel=44
					4, 7, -5, 0, -7, -7, 4, 1, 4,
					-- layer=2 filter=165 channel=45
					-3, 26, 19, 4, -26, 11, -9, -19, -11,
					-- layer=2 filter=165 channel=46
					9, -5, -8, 18, -46, -44, -35, -40, -16,
					-- layer=2 filter=165 channel=47
					-2, -2, 3, -1, -29, -7, 5, -12, -6,
					-- layer=2 filter=165 channel=48
					2, 9, 9, 5, 9, 8, -3, 1, 1,
					-- layer=2 filter=165 channel=49
					6, -6, 14, -20, -57, 0, -19, -58, -8,
					-- layer=2 filter=165 channel=50
					-11, -8, -14, 0, 2, 1, 1, 0, -2,
					-- layer=2 filter=165 channel=51
					-9, -27, -22, -24, -23, -30, -7, -1, 3,
					-- layer=2 filter=165 channel=52
					-17, -5, 0, -25, 15, -3, 34, -2, 5,
					-- layer=2 filter=165 channel=53
					8, 38, 18, 37, -63, 33, 31, 29, 7,
					-- layer=2 filter=165 channel=54
					-18, -28, -14, -32, -6, -20, 5, 45, 9,
					-- layer=2 filter=165 channel=55
					-1, -6, -7, 0, -10, -3, -6, 0, -3,
					-- layer=2 filter=165 channel=56
					-2, 0, -14, -20, -12, -12, 5, 15, -12,
					-- layer=2 filter=165 channel=57
					-3, 4, 12, -7, 7, 0, 1, -2, -2,
					-- layer=2 filter=165 channel=58
					23, 8, 15, -14, -4, -3, -12, 6, -41,
					-- layer=2 filter=165 channel=59
					13, 28, -8, -37, 20, 27, 16, 16, -2,
					-- layer=2 filter=165 channel=60
					-20, -10, 38, -32, -18, -4, -6, -6, -35,
					-- layer=2 filter=165 channel=61
					1, 27, -19, -64, -15, -17, -25, -63, -36,
					-- layer=2 filter=165 channel=62
					-35, -13, -9, -13, 0, -15, 17, 25, 39,
					-- layer=2 filter=165 channel=63
					14, 7, -5, -8, -4, -7, -9, -20, -19,
					-- layer=2 filter=165 channel=64
					-4, -5, 1, -2, 38, -1, -15, 9, 8,
					-- layer=2 filter=165 channel=65
					17, 16, 31, -7, 6, 10, 8, -6, -5,
					-- layer=2 filter=165 channel=66
					4, -19, 13, -1, 15, -25, -25, -23, -33,
					-- layer=2 filter=165 channel=67
					6, 6, 15, 26, 29, 14, -50, -52, -21,
					-- layer=2 filter=165 channel=68
					5, -9, 4, -3, 5, -1, -4, -3, -1,
					-- layer=2 filter=165 channel=69
					10, 0, -2, 18, 38, -4, -2, 3, 4,
					-- layer=2 filter=165 channel=70
					19, 22, 14, -12, -7, -5, -28, -16, -10,
					-- layer=2 filter=165 channel=71
					-11, 25, -7, -4, 27, 6, 19, 23, 5,
					-- layer=2 filter=165 channel=72
					-23, -21, 13, -31, -9, -25, 0, -7, -21,
					-- layer=2 filter=165 channel=73
					52, 61, 15, -25, -7, 23, -11, -21, -20,
					-- layer=2 filter=165 channel=74
					7, 0, 10, 0, 24, 8, -62, -58, -56,
					-- layer=2 filter=165 channel=75
					-23, -26, 12, -15, 0, -17, -26, -45, -6,
					-- layer=2 filter=165 channel=76
					64, 61, 8, 6, -49, -15, 32, -13, -1,
					-- layer=2 filter=165 channel=77
					-4, -3, 6, -5, 4, -8, -2, -6, -3,
					-- layer=2 filter=165 channel=78
					-13, -19, -15, -32, -16, -17, -5, 6, 20,
					-- layer=2 filter=165 channel=79
					-5, -6, -4, 3, -1, 8, 4, 4, 10,
					-- layer=2 filter=165 channel=80
					-11, 8, 11, -7, -1, -15, -68, -65, -43,
					-- layer=2 filter=165 channel=81
					-10, -12, 1, -9, -7, -12, 0, -10, -8,
					-- layer=2 filter=165 channel=82
					8, 5, -4, -10, 8, -1, 7, -6, 2,
					-- layer=2 filter=165 channel=83
					-8, 17, 7, 3, 32, -20, -30, -62, -27,
					-- layer=2 filter=165 channel=84
					4, -11, -1, 10, -4, 6, -4, 1, -6,
					-- layer=2 filter=165 channel=85
					11, 15, 8, -12, 11, 6, -1, 7, -5,
					-- layer=2 filter=165 channel=86
					-5, 12, 16, -9, 13, -16, 1, -14, -3,
					-- layer=2 filter=165 channel=87
					4, 67, -21, 22, -31, -24, -5, -17, -6,
					-- layer=2 filter=165 channel=88
					16, 13, 1, 27, 35, 24, -16, -7, -31,
					-- layer=2 filter=165 channel=89
					9, -6, -18, -19, 20, -14, -7, 7, -13,
					-- layer=2 filter=165 channel=90
					-10, 2, -9, 10, -8, -4, -4, -1, -5,
					-- layer=2 filter=165 channel=91
					-5, -12, 13, -9, 8, 20, -6, 13, -27,
					-- layer=2 filter=165 channel=92
					11, -16, -5, -22, 0, 5, 0, 32, -25,
					-- layer=2 filter=165 channel=93
					-40, 44, 14, -56, -14, 9, -37, 67, 37,
					-- layer=2 filter=165 channel=94
					13, 10, 2, 28, 10, -9, 11, -18, -11,
					-- layer=2 filter=165 channel=95
					10, -7, 0, 0, -9, -2, -2, -8, -1,
					-- layer=2 filter=165 channel=96
					38, 17, -2, 20, 45, 44, 21, 74, 32,
					-- layer=2 filter=165 channel=97
					0, 11, 10, -3, -20, -15, -5, -14, 10,
					-- layer=2 filter=165 channel=98
					17, 9, -4, -38, -31, -13, 3, -10, -5,
					-- layer=2 filter=165 channel=99
					-2, 10, 12, -15, -3, 41, 27, -4, -12,
					-- layer=2 filter=165 channel=100
					47, 24, 27, 17, 3, -2, -80, -80, -68,
					-- layer=2 filter=165 channel=101
					-16, 0, -14, -16, -6, -4, 14, 23, 1,
					-- layer=2 filter=165 channel=102
					23, -8, -12, 5, 6, 12, 23, 20, 8,
					-- layer=2 filter=165 channel=103
					-15, -17, -54, -11, -14, 35, 11, -17, -23,
					-- layer=2 filter=165 channel=104
					20, 19, 4, 25, -20, 17, 10, -62, 28,
					-- layer=2 filter=165 channel=105
					9, 85, 32, 16, 16, -6, 21, 38, -3,
					-- layer=2 filter=165 channel=106
					-4, 3, 3, -8, -7, 5, 16, 9, 11,
					-- layer=2 filter=165 channel=107
					-37, 28, -50, -22, -20, -16, -12, 27, 4,
					-- layer=2 filter=165 channel=108
					-6, 11, 13, 1, 18, 7, -12, -6, 16,
					-- layer=2 filter=165 channel=109
					13, 4, -8, 2, -5, 0, -2, 8, -4,
					-- layer=2 filter=165 channel=110
					-22, 15, 2, 4, 53, 35, -30, 16, 21,
					-- layer=2 filter=165 channel=111
					4, 8, 1, 0, -5, 10, -3, 2, 5,
					-- layer=2 filter=165 channel=112
					20, 2, 10, -19, 1, 13, 29, -14, 1,
					-- layer=2 filter=165 channel=113
					10, 15, -5, -33, 3, -1, -39, -66, -37,
					-- layer=2 filter=165 channel=114
					0, 8, 0, 4, -1, -1, 23, 19, 8,
					-- layer=2 filter=165 channel=115
					-1, -6, -10, -4, -5, 12, 0, -6, -4,
					-- layer=2 filter=165 channel=116
					4, 45, -2, 17, -39, -2, 19, -25, -6,
					-- layer=2 filter=165 channel=117
					-19, -2, -62, -37, 23, 24, 2, 16, 12,
					-- layer=2 filter=165 channel=118
					-21, 7, 7, -16, -18, 2, -7, -29, 0,
					-- layer=2 filter=165 channel=119
					6, 24, -12, 6, -17, -13, 0, -66, -21,
					-- layer=2 filter=165 channel=120
					-5, 1, 0, -6, -8, 0, 5, -1, -9,
					-- layer=2 filter=165 channel=121
					2, 0, -1, -3, 6, 8, 3, 11, -3,
					-- layer=2 filter=165 channel=122
					6, 5, 14, 11, -6, -8, 3, -3, 14,
					-- layer=2 filter=165 channel=123
					4, -8, -5, -32, -8, -9, 28, 0, 26,
					-- layer=2 filter=165 channel=124
					-25, 17, -5, 8, -41, -15, -19, -4, -25,
					-- layer=2 filter=165 channel=125
					-11, -5, 11, 5, 4, -1, 0, -7, 4,
					-- layer=2 filter=165 channel=126
					46, 34, -21, 9, -27, 18, 24, 24, -36,
					-- layer=2 filter=165 channel=127
					-8, -1, -3, 12, 23, 8, -1, -11, -10,
					-- layer=2 filter=166 channel=0
					-12, -11, -7, 0, -3, -8, -15, -14, -11,
					-- layer=2 filter=166 channel=1
					1, -6, -3, -11, -1, 5, -13, -13, 0,
					-- layer=2 filter=166 channel=2
					-5, -11, 7, 8, -8, 3, -8, -9, 4,
					-- layer=2 filter=166 channel=3
					-7, -3, -3, -7, -8, 4, 3, -11, -8,
					-- layer=2 filter=166 channel=4
					-4, 7, 4, -3, 0, 8, -3, -1, 6,
					-- layer=2 filter=166 channel=5
					0, -5, 0, 0, 4, 0, 4, -11, -2,
					-- layer=2 filter=166 channel=6
					-14, -12, 2, -15, 0, -2, -7, -6, 1,
					-- layer=2 filter=166 channel=7
					-11, -6, -8, 1, -2, -14, 1, -7, 2,
					-- layer=2 filter=166 channel=8
					1, -7, -9, 4, -7, -2, -4, -10, 6,
					-- layer=2 filter=166 channel=9
					-2, -1, -7, -8, -13, -8, -13, -8, 4,
					-- layer=2 filter=166 channel=10
					-9, -1, 4, -13, 4, -8, -3, -14, 3,
					-- layer=2 filter=166 channel=11
					0, -9, 5, -12, 0, 1, -12, -9, -6,
					-- layer=2 filter=166 channel=12
					12, -8, 9, 4, -5, -3, -17, -10, -10,
					-- layer=2 filter=166 channel=13
					0, 4, -3, 3, -11, 0, 1, 3, -3,
					-- layer=2 filter=166 channel=14
					-2, 6, -11, -8, -1, -4, -8, 4, -5,
					-- layer=2 filter=166 channel=15
					1, 2, -1, -13, 1, 4, -2, -6, -5,
					-- layer=2 filter=166 channel=16
					4, -9, -9, -4, -5, 9, -6, -13, -6,
					-- layer=2 filter=166 channel=17
					-3, 3, -8, 10, -6, 7, 0, -3, 3,
					-- layer=2 filter=166 channel=18
					-6, -3, 12, -10, 6, -3, -4, 11, 8,
					-- layer=2 filter=166 channel=19
					3, -7, -6, -3, -4, 1, 1, 0, -2,
					-- layer=2 filter=166 channel=20
					1, -1, -1, 5, 2, -7, 3, -6, 4,
					-- layer=2 filter=166 channel=21
					8, -4, -6, 5, -1, -9, -4, -8, -6,
					-- layer=2 filter=166 channel=22
					-5, -1, -6, -2, -4, 10, -10, 0, -7,
					-- layer=2 filter=166 channel=23
					9, -7, 7, -4, -5, 0, -2, 4, 0,
					-- layer=2 filter=166 channel=24
					-2, -13, -14, -16, -8, -16, -4, 0, -12,
					-- layer=2 filter=166 channel=25
					5, 1, -15, 0, 3, -1, -1, -2, -9,
					-- layer=2 filter=166 channel=26
					-5, 8, -4, -6, 0, 9, 2, -3, 0,
					-- layer=2 filter=166 channel=27
					-10, -2, -14, -14, 0, 3, -8, -5, 6,
					-- layer=2 filter=166 channel=28
					-7, -8, 4, -10, -14, 3, -7, -2, -8,
					-- layer=2 filter=166 channel=29
					6, -10, 2, -10, -7, -1, 3, -8, 10,
					-- layer=2 filter=166 channel=30
					-2, 3, 6, 2, 2, 1, -5, 1, 3,
					-- layer=2 filter=166 channel=31
					0, 4, 5, -13, 1, -8, -4, -6, -9,
					-- layer=2 filter=166 channel=32
					9, -10, -10, 10, -5, 7, 0, -11, 3,
					-- layer=2 filter=166 channel=33
					-2, 4, 10, -2, 0, -11, -5, -10, 2,
					-- layer=2 filter=166 channel=34
					-12, 0, -9, -1, 0, 0, -2, -4, -5,
					-- layer=2 filter=166 channel=35
					-1, -14, 3, 1, -11, 1, 0, 8, -2,
					-- layer=2 filter=166 channel=36
					8, -2, -2, 0, 6, 10, -5, -7, 10,
					-- layer=2 filter=166 channel=37
					-9, -14, -6, -1, -7, 0, -5, -11, 2,
					-- layer=2 filter=166 channel=38
					0, 1, 7, -1, -9, -3, 4, 4, 4,
					-- layer=2 filter=166 channel=39
					8, -4, 4, 0, -1, 13, 2, -11, -3,
					-- layer=2 filter=166 channel=40
					11, -2, -1, -7, 8, -7, -1, 1, -9,
					-- layer=2 filter=166 channel=41
					-3, 10, -5, 8, 0, 0, 7, 8, -7,
					-- layer=2 filter=166 channel=42
					2, -11, -8, -9, 8, 0, 1, 7, 4,
					-- layer=2 filter=166 channel=43
					3, -13, -4, 2, -6, -12, 0, -12, -7,
					-- layer=2 filter=166 channel=44
					-10, -10, 0, 2, 0, 10, -1, 3, 5,
					-- layer=2 filter=166 channel=45
					-4, -8, -2, -16, 1, -6, -10, -3, -6,
					-- layer=2 filter=166 channel=46
					1, 0, 2, -6, -15, 8, -8, -11, -1,
					-- layer=2 filter=166 channel=47
					3, -17, 0, -2, 1, 4, 6, 0, 13,
					-- layer=2 filter=166 channel=48
					9, -7, -3, -7, 7, 0, 3, 8, -8,
					-- layer=2 filter=166 channel=49
					-11, -9, 4, -13, -3, -2, -7, 0, -13,
					-- layer=2 filter=166 channel=50
					-1, 6, -2, -4, 8, -8, -1, 0, -9,
					-- layer=2 filter=166 channel=51
					-14, -14, -6, -9, 1, 4, -7, -2, 7,
					-- layer=2 filter=166 channel=52
					-9, -10, -6, -5, 7, 3, -11, -3, -12,
					-- layer=2 filter=166 channel=53
					0, -20, 6, 0, -5, -8, -1, -3, -5,
					-- layer=2 filter=166 channel=54
					-3, -10, -8, -14, -8, -4, -7, 1, 1,
					-- layer=2 filter=166 channel=55
					1, 5, -7, -5, -1, -4, 0, -9, 2,
					-- layer=2 filter=166 channel=56
					-6, -16, -8, -1, -7, 5, 0, 0, 0,
					-- layer=2 filter=166 channel=57
					6, 3, -8, -5, -2, 3, -6, 1, -3,
					-- layer=2 filter=166 channel=58
					3, -1, 4, -1, -4, 0, -13, 1, -15,
					-- layer=2 filter=166 channel=59
					0, -2, 2, -12, -3, 2, -11, -7, 1,
					-- layer=2 filter=166 channel=60
					-1, -8, -15, -9, 4, 1, -3, -2, -6,
					-- layer=2 filter=166 channel=61
					-2, -3, 3, 0, 2, -13, -12, -8, -1,
					-- layer=2 filter=166 channel=62
					-1, 0, -5, -8, -6, 4, 0, 6, -2,
					-- layer=2 filter=166 channel=63
					-3, -12, 6, -6, 0, 4, -8, 0, 0,
					-- layer=2 filter=166 channel=64
					2, -4, -11, 5, -5, 3, 2, 2, 10,
					-- layer=2 filter=166 channel=65
					-2, -10, 1, 4, -13, 0, 10, 3, -14,
					-- layer=2 filter=166 channel=66
					-1, 0, 4, -3, -5, 6, -7, 10, 0,
					-- layer=2 filter=166 channel=67
					-9, 3, 3, -13, -16, 8, -2, 0, 5,
					-- layer=2 filter=166 channel=68
					-8, 6, 4, 2, -1, 8, 9, -1, -5,
					-- layer=2 filter=166 channel=69
					1, 5, 10, -5, -8, -9, -3, 8, 2,
					-- layer=2 filter=166 channel=70
					0, -4, 7, -2, -3, 3, -2, 0, -3,
					-- layer=2 filter=166 channel=71
					-11, 0, -7, -5, 0, 5, -6, -2, 7,
					-- layer=2 filter=166 channel=72
					-1, 0, -8, -15, -4, -14, -3, -12, -9,
					-- layer=2 filter=166 channel=73
					-16, 0, 1, -20, -17, -5, -11, -9, -4,
					-- layer=2 filter=166 channel=74
					-4, -5, -6, 1, 1, 2, -1, -5, -5,
					-- layer=2 filter=166 channel=75
					9, 6, -11, 6, 4, -4, 7, -4, 2,
					-- layer=2 filter=166 channel=76
					0, -7, -1, -4, 9, -5, 0, -3, -6,
					-- layer=2 filter=166 channel=77
					0, -10, -3, -10, 2, -3, -8, 0, -1,
					-- layer=2 filter=166 channel=78
					-15, -1, 0, 4, 5, 4, -12, -11, 8,
					-- layer=2 filter=166 channel=79
					4, -3, -3, -5, 6, 2, -7, 6, 0,
					-- layer=2 filter=166 channel=80
					5, 7, -1, 5, -1, -5, 5, -9, 13,
					-- layer=2 filter=166 channel=81
					1, 6, -2, -8, 6, 0, 0, 2, 4,
					-- layer=2 filter=166 channel=82
					-9, 3, 9, -8, 8, 9, 0, 0, 3,
					-- layer=2 filter=166 channel=83
					3, 1, -2, -8, 5, 4, -9, 3, -5,
					-- layer=2 filter=166 channel=84
					2, 5, 8, 5, 2, 0, -9, -1, 7,
					-- layer=2 filter=166 channel=85
					-7, 2, -8, 7, -1, 6, 9, 3, 7,
					-- layer=2 filter=166 channel=86
					8, 4, 7, 2, -1, -6, 0, 7, 0,
					-- layer=2 filter=166 channel=87
					0, -6, -9, 3, -7, -8, -1, 8, -5,
					-- layer=2 filter=166 channel=88
					-1, -2, -9, 1, -6, -7, -5, -4, 10,
					-- layer=2 filter=166 channel=89
					0, 1, 8, -4, 0, 0, -18, -10, 8,
					-- layer=2 filter=166 channel=90
					1, 2, 10, 8, 0, 3, -6, 0, 4,
					-- layer=2 filter=166 channel=91
					7, -10, -7, 2, -1, 5, -12, -8, -1,
					-- layer=2 filter=166 channel=92
					-7, 0, 3, -11, 0, -3, 3, 7, 0,
					-- layer=2 filter=166 channel=93
					-3, 3, 3, -11, 4, -3, -3, -17, -9,
					-- layer=2 filter=166 channel=94
					1, 3, -10, -2, -5, -3, -4, -13, 3,
					-- layer=2 filter=166 channel=95
					-12, -9, -6, 3, -7, 2, 8, 5, 8,
					-- layer=2 filter=166 channel=96
					4, -6, -21, -2, -11, -6, -15, -16, -9,
					-- layer=2 filter=166 channel=97
					-5, -14, 5, -9, 3, -5, -6, -10, -12,
					-- layer=2 filter=166 channel=98
					-14, -8, 3, -12, -11, -6, -9, -4, 13,
					-- layer=2 filter=166 channel=99
					2, -14, -10, 3, -13, -14, -11, -6, -5,
					-- layer=2 filter=166 channel=100
					-4, -11, 1, -3, -18, -1, 4, -10, -2,
					-- layer=2 filter=166 channel=101
					-2, -8, -11, -12, -8, 6, -1, -1, -14,
					-- layer=2 filter=166 channel=102
					-1, 2, -6, -8, -9, 0, -6, 0, 0,
					-- layer=2 filter=166 channel=103
					4, 9, 4, -10, -2, -3, -9, 4, -2,
					-- layer=2 filter=166 channel=104
					9, -5, -2, -5, -8, 4, -9, 2, 5,
					-- layer=2 filter=166 channel=105
					-2, -9, -4, 7, -10, 5, -10, 3, 9,
					-- layer=2 filter=166 channel=106
					-15, -6, 2, 0, 0, -3, 4, 3, -10,
					-- layer=2 filter=166 channel=107
					5, 6, -4, -1, -4, 1, 2, -10, -1,
					-- layer=2 filter=166 channel=108
					5, -4, -3, 1, -10, -7, -11, -11, -4,
					-- layer=2 filter=166 channel=109
					7, -11, 5, -9, 7, 6, -4, -4, 1,
					-- layer=2 filter=166 channel=110
					-7, 3, -6, -4, -14, 0, 7, -7, 6,
					-- layer=2 filter=166 channel=111
					8, 6, 0, -9, 9, 0, 9, 0, -7,
					-- layer=2 filter=166 channel=112
					-15, 0, -13, -14, -9, -3, 1, 1, -8,
					-- layer=2 filter=166 channel=113
					-3, -12, 0, 8, -3, -1, -4, 0, 3,
					-- layer=2 filter=166 channel=114
					3, 2, 1, 6, -6, -6, -5, 1, -2,
					-- layer=2 filter=166 channel=115
					5, 0, -1, 4, 7, 4, 8, 5, 0,
					-- layer=2 filter=166 channel=116
					2, 0, 7, -6, -9, 7, 4, 2, -7,
					-- layer=2 filter=166 channel=117
					-4, -14, -7, -8, -9, 3, -18, -3, 0,
					-- layer=2 filter=166 channel=118
					0, 5, -2, -14, -3, -11, -12, -6, 1,
					-- layer=2 filter=166 channel=119
					-7, 6, 11, 3, 2, 10, 3, 7, -1,
					-- layer=2 filter=166 channel=120
					-8, -1, -6, 7, 2, 3, -3, -8, -7,
					-- layer=2 filter=166 channel=121
					-9, 2, -7, -8, 0, -5, -6, 6, 2,
					-- layer=2 filter=166 channel=122
					-3, -9, 4, 1, 6, 1, -1, -10, -3,
					-- layer=2 filter=166 channel=123
					-13, -11, 6, -10, -15, -16, -14, -6, -8,
					-- layer=2 filter=166 channel=124
					-10, -8, 1, -3, -11, -7, 0, -13, -11,
					-- layer=2 filter=166 channel=125
					-7, 0, -3, 0, -10, 7, -1, 2, -5,
					-- layer=2 filter=166 channel=126
					6, -5, -5, -6, -7, -9, -2, 9, 4,
					-- layer=2 filter=166 channel=127
					-4, -5, -3, -8, -16, -6, -10, -1, -7,
					-- layer=2 filter=167 channel=0
					0, -7, -13, -6, -14, -6, -11, -11, -3,
					-- layer=2 filter=167 channel=1
					-7, -13, -1, -9, -7, -16, 7, -11, 0,
					-- layer=2 filter=167 channel=2
					-7, 0, -2, 8, 0, 3, -9, -5, 2,
					-- layer=2 filter=167 channel=3
					5, -14, -3, -14, 1, 4, -15, 1, -11,
					-- layer=2 filter=167 channel=4
					3, -4, 2, -2, -7, -1, -1, 4, 2,
					-- layer=2 filter=167 channel=5
					2, 5, -5, -14, -3, 0, -8, -3, -11,
					-- layer=2 filter=167 channel=6
					3, -17, -9, -11, 4, -3, -18, 7, -12,
					-- layer=2 filter=167 channel=7
					-11, -12, -4, -11, -1, -6, 2, -9, -9,
					-- layer=2 filter=167 channel=8
					9, -9, 0, 2, -7, -4, 7, 0, 0,
					-- layer=2 filter=167 channel=9
					-9, 1, -3, -11, -7, 2, -15, 2, 12,
					-- layer=2 filter=167 channel=10
					0, -12, -4, 1, 0, -7, -17, 0, 6,
					-- layer=2 filter=167 channel=11
					-2, -7, -12, 4, -7, -9, -13, 0, -15,
					-- layer=2 filter=167 channel=12
					4, -4, -13, 0, -12, -19, 3, -15, -8,
					-- layer=2 filter=167 channel=13
					-7, 5, 8, -6, -7, 0, -4, -9, -2,
					-- layer=2 filter=167 channel=14
					-10, -6, -2, 7, -16, 1, 6, 6, -12,
					-- layer=2 filter=167 channel=15
					-6, -5, 0, 10, -6, -5, -11, 10, -13,
					-- layer=2 filter=167 channel=16
					-7, 2, -8, -3, 0, 0, 13, -2, 12,
					-- layer=2 filter=167 channel=17
					8, 4, -8, -2, 9, 6, 8, -3, 3,
					-- layer=2 filter=167 channel=18
					3, -13, 7, 10, -6, -2, 7, 5, -3,
					-- layer=2 filter=167 channel=19
					-7, 6, -2, -3, -5, -4, 8, -9, -6,
					-- layer=2 filter=167 channel=20
					-7, -5, 3, 9, 0, -6, 6, 5, -7,
					-- layer=2 filter=167 channel=21
					-3, -9, 9, 1, 1, -6, -9, 3, -5,
					-- layer=2 filter=167 channel=22
					7, 8, -1, -3, -8, 7, 7, 0, -6,
					-- layer=2 filter=167 channel=23
					-13, -2, -4, -10, 0, 6, -3, -3, 9,
					-- layer=2 filter=167 channel=24
					-12, -18, -15, -5, -4, -7, -12, 0, -14,
					-- layer=2 filter=167 channel=25
					4, 3, -7, 7, 3, -4, 1, -2, 0,
					-- layer=2 filter=167 channel=26
					0, -1, -3, -4, -6, 4, 5, 4, 0,
					-- layer=2 filter=167 channel=27
					12, 1, -10, -7, -2, -13, -2, -8, 3,
					-- layer=2 filter=167 channel=28
					-2, -7, 2, -4, 12, -1, -9, -14, -13,
					-- layer=2 filter=167 channel=29
					-10, -11, 5, -6, -6, 4, -8, -5, -5,
					-- layer=2 filter=167 channel=30
					2, -5, 3, -12, -4, 3, -3, 1, 6,
					-- layer=2 filter=167 channel=31
					-9, -3, 1, -2, -4, -16, 2, -13, -1,
					-- layer=2 filter=167 channel=32
					-9, -9, 0, -5, 2, 5, 7, 7, -1,
					-- layer=2 filter=167 channel=33
					-15, -17, 0, 2, -8, 0, 0, -4, -7,
					-- layer=2 filter=167 channel=34
					-11, 1, 3, -17, -7, -4, 6, 1, -14,
					-- layer=2 filter=167 channel=35
					2, 4, 0, 1, -1, -4, 2, -8, -8,
					-- layer=2 filter=167 channel=36
					-13, -10, -15, 3, -15, 0, -11, -14, -9,
					-- layer=2 filter=167 channel=37
					5, -12, -3, -14, -5, -3, 3, -6, -2,
					-- layer=2 filter=167 channel=38
					8, -11, 5, -2, 3, 2, -6, 2, 1,
					-- layer=2 filter=167 channel=39
					-8, -4, -6, 5, 1, 0, 3, 11, -9,
					-- layer=2 filter=167 channel=40
					-11, -8, 2, -10, -5, -5, -4, 4, 9,
					-- layer=2 filter=167 channel=41
					-5, 0, 1, -7, 7, 6, -5, -6, -3,
					-- layer=2 filter=167 channel=42
					0, -12, -2, 4, 3, -11, 6, 11, -3,
					-- layer=2 filter=167 channel=43
					-14, -9, 0, -10, 7, -6, -7, -17, 2,
					-- layer=2 filter=167 channel=44
					4, -9, 6, 4, 3, -2, 9, -4, 1,
					-- layer=2 filter=167 channel=45
					-8, -4, 2, -9, -2, -15, 6, -1, 6,
					-- layer=2 filter=167 channel=46
					-7, -1, 0, -7, -13, 2, 4, 2, 4,
					-- layer=2 filter=167 channel=47
					-4, 4, 1, 3, 3, -3, -13, 2, -14,
					-- layer=2 filter=167 channel=48
					-1, -8, -8, 0, 1, 6, 0, 4, 10,
					-- layer=2 filter=167 channel=49
					-10, 6, -1, 10, -1, -2, 0, -6, -9,
					-- layer=2 filter=167 channel=50
					-4, 0, 9, -6, -10, -9, -10, -10, 10,
					-- layer=2 filter=167 channel=51
					2, -14, -10, 1, 2, -6, -3, -11, -1,
					-- layer=2 filter=167 channel=52
					-9, 0, -10, -10, -8, -13, -7, -10, -6,
					-- layer=2 filter=167 channel=53
					0, -10, 0, 7, -14, -3, 0, -9, -16,
					-- layer=2 filter=167 channel=54
					-4, -4, -3, -8, 4, -2, -9, -10, 0,
					-- layer=2 filter=167 channel=55
					-1, -7, 8, -9, 6, -9, -6, 3, 1,
					-- layer=2 filter=167 channel=56
					-6, -11, -13, 0, 0, -13, -1, -15, -14,
					-- layer=2 filter=167 channel=57
					-2, 7, 9, -4, -7, -10, -1, 0, -4,
					-- layer=2 filter=167 channel=58
					2, -5, -7, 4, -2, -18, 4, 1, -10,
					-- layer=2 filter=167 channel=59
					6, 2, -3, 5, -10, 3, 0, -10, -14,
					-- layer=2 filter=167 channel=60
					-16, 7, 0, 5, -5, -8, 4, 0, -18,
					-- layer=2 filter=167 channel=61
					-5, 3, 2, -11, 8, 3, -13, -2, 0,
					-- layer=2 filter=167 channel=62
					-2, 2, -6, 2, 0, 3, -3, 8, 2,
					-- layer=2 filter=167 channel=63
					-7, -2, -15, -3, -7, 3, 6, 4, -1,
					-- layer=2 filter=167 channel=64
					3, 6, -10, -11, -3, -10, 0, 3, 6,
					-- layer=2 filter=167 channel=65
					0, -15, -14, -5, -2, 1, -14, -15, -12,
					-- layer=2 filter=167 channel=66
					1, -4, -3, 3, -9, 6, -3, 4, -1,
					-- layer=2 filter=167 channel=67
					-7, -1, -2, 0, -6, -4, -6, 5, 4,
					-- layer=2 filter=167 channel=68
					4, 1, -3, 0, -7, 6, 0, 3, -11,
					-- layer=2 filter=167 channel=69
					-11, 6, -5, -14, -10, -14, -5, 10, -8,
					-- layer=2 filter=167 channel=70
					2, -13, 3, 6, 6, 8, -12, -2, -14,
					-- layer=2 filter=167 channel=71
					7, -5, 0, 0, 9, -6, 0, 1, -5,
					-- layer=2 filter=167 channel=72
					3, -11, 1, -11, 0, -3, -9, -10, 0,
					-- layer=2 filter=167 channel=73
					-8, -14, -6, 3, -3, -10, 1, -6, 1,
					-- layer=2 filter=167 channel=74
					5, -4, -7, 7, 7, 8, 8, -2, -4,
					-- layer=2 filter=167 channel=75
					3, -3, -13, -11, -11, 0, -14, -12, -14,
					-- layer=2 filter=167 channel=76
					10, -3, 16, -4, -5, 9, 2, 0, -1,
					-- layer=2 filter=167 channel=77
					1, -10, 1, -5, 6, -6, -7, 0, -9,
					-- layer=2 filter=167 channel=78
					-9, -1, -16, -5, -1, -9, -8, -11, -14,
					-- layer=2 filter=167 channel=79
					-4, -3, 0, 1, 7, 6, -5, -2, 8,
					-- layer=2 filter=167 channel=80
					0, -6, -9, 5, 2, 3, 10, -6, 11,
					-- layer=2 filter=167 channel=81
					1, 0, -9, -7, 4, -5, 6, -10, -2,
					-- layer=2 filter=167 channel=82
					2, 10, -2, 6, 7, 0, -6, -1, -1,
					-- layer=2 filter=167 channel=83
					-1, -7, 2, -1, 2, -10, 2, -1, 3,
					-- layer=2 filter=167 channel=84
					4, 9, -2, -6, -2, 6, -2, 3, 1,
					-- layer=2 filter=167 channel=85
					-8, 5, -4, -2, -2, -6, -6, 8, 1,
					-- layer=2 filter=167 channel=86
					-2, -1, 10, 5, -3, 8, 1, -2, 7,
					-- layer=2 filter=167 channel=87
					11, 8, -1, 5, -6, 9, -12, 7, 2,
					-- layer=2 filter=167 channel=88
					-9, -2, 0, 2, 3, -11, -2, 8, -9,
					-- layer=2 filter=167 channel=89
					3, -3, -7, 4, -9, -7, -3, 2, -9,
					-- layer=2 filter=167 channel=90
					5, -3, 9, 8, -4, 4, 0, -7, 10,
					-- layer=2 filter=167 channel=91
					6, 7, -12, -9, 5, -1, 0, -11, -1,
					-- layer=2 filter=167 channel=92
					-2, -12, -16, -10, -10, -6, -6, -2, -3,
					-- layer=2 filter=167 channel=93
					-2, -18, -13, -10, -4, -10, 0, -10, -15,
					-- layer=2 filter=167 channel=94
					-4, -2, -4, -12, -9, -9, 5, -9, -15,
					-- layer=2 filter=167 channel=95
					-8, 7, 5, 2, 4, -9, 7, 7, 5,
					-- layer=2 filter=167 channel=96
					-8, -3, -13, -7, -5, 1, -1, 5, -9,
					-- layer=2 filter=167 channel=97
					-16, -3, -13, 0, -2, -12, -3, 1, -5,
					-- layer=2 filter=167 channel=98
					0, 4, -1, -7, -7, 3, -6, -5, -6,
					-- layer=2 filter=167 channel=99
					-5, -11, 8, -7, 3, -9, -6, -1, -4,
					-- layer=2 filter=167 channel=100
					-5, 0, -4, -7, -10, -8, 7, -1, -11,
					-- layer=2 filter=167 channel=101
					9, 1, -5, 3, -2, -4, 8, 8, -4,
					-- layer=2 filter=167 channel=102
					4, -10, 7, 0, 1, 1, 7, 2, -2,
					-- layer=2 filter=167 channel=103
					-5, -4, -9, -8, -5, -3, 5, 0, 9,
					-- layer=2 filter=167 channel=104
					-13, -8, -6, 0, 2, 0, -5, -4, -4,
					-- layer=2 filter=167 channel=105
					7, -2, 0, -6, 3, 0, -3, -5, -12,
					-- layer=2 filter=167 channel=106
					-5, 6, -5, -10, -5, -8, -10, -7, 5,
					-- layer=2 filter=167 channel=107
					-1, 2, -7, -7, 3, -13, -7, -1, 3,
					-- layer=2 filter=167 channel=108
					-7, -6, -1, -5, -1, 1, -2, 6, -3,
					-- layer=2 filter=167 channel=109
					4, 1, 0, -9, 6, -4, -5, -7, 0,
					-- layer=2 filter=167 channel=110
					-3, 1, 2, 0, 1, -15, 7, 0, 4,
					-- layer=2 filter=167 channel=111
					-8, -6, -4, -10, -10, -3, -5, 7, 6,
					-- layer=2 filter=167 channel=112
					3, -14, -10, -7, -5, -3, -5, -9, -6,
					-- layer=2 filter=167 channel=113
					-7, -12, -14, -8, -12, -5, 2, -9, -2,
					-- layer=2 filter=167 channel=114
					1, 0, -5, -3, -4, 5, 6, 9, 3,
					-- layer=2 filter=167 channel=115
					9, -5, 7, 3, -3, 1, 7, -1, 4,
					-- layer=2 filter=167 channel=116
					3, 2, 4, 5, 3, 11, 3, -7, 0,
					-- layer=2 filter=167 channel=117
					-11, 0, -4, -6, 4, 8, -8, 1, 3,
					-- layer=2 filter=167 channel=118
					0, -10, 2, -5, -5, -7, -17, 0, -2,
					-- layer=2 filter=167 channel=119
					3, -1, 3, 2, -2, 3, 9, 6, 5,
					-- layer=2 filter=167 channel=120
					7, -7, 3, 1, -7, 3, 4, 9, -2,
					-- layer=2 filter=167 channel=121
					9, 0, 9, -4, -10, 5, -4, 6, 9,
					-- layer=2 filter=167 channel=122
					5, 6, -7, 1, 1, 5, 4, -8, 5,
					-- layer=2 filter=167 channel=123
					-11, -11, -2, -7, 0, -5, -1, -8, -7,
					-- layer=2 filter=167 channel=124
					-5, 4, -5, 1, 0, -11, -7, 0, 3,
					-- layer=2 filter=167 channel=125
					6, -4, -8, 6, -8, 1, 10, -6, -6,
					-- layer=2 filter=167 channel=126
					-10, 3, 4, -4, -4, -3, -1, 0, -3,
					-- layer=2 filter=167 channel=127
					-14, 2, -2, -14, -9, 4, 2, 8, -1,
					-- layer=2 filter=168 channel=0
					-21, 4, -5, -7, -7, -5, -24, -17, -9,
					-- layer=2 filter=168 channel=1
					-21, 4, -16, -21, -7, -18, -14, -11, -6,
					-- layer=2 filter=168 channel=2
					-3, -6, 4, 5, 5, -4, -10, 7, -4,
					-- layer=2 filter=168 channel=3
					-1, -16, -18, -17, -10, -4, -11, -2, -20,
					-- layer=2 filter=168 channel=4
					5, -5, -17, -15, -2, 13, -4, -15, -26,
					-- layer=2 filter=168 channel=5
					-19, 16, -1, -17, 0, -6, 0, -14, -9,
					-- layer=2 filter=168 channel=6
					21, 9, -31, 16, 12, 0, 11, 12, 0,
					-- layer=2 filter=168 channel=7
					-10, -11, -27, -22, -9, 1, -12, -1, -8,
					-- layer=2 filter=168 channel=8
					-11, -1, -1, 2, -8, -2, -3, 8, -1,
					-- layer=2 filter=168 channel=9
					-4, -8, 1, -9, -11, -13, 2, -7, -16,
					-- layer=2 filter=168 channel=10
					-8, -4, -9, -8, -15, -2, -4, -19, -12,
					-- layer=2 filter=168 channel=11
					-19, -1, -27, -20, -7, -22, -25, -11, 0,
					-- layer=2 filter=168 channel=12
					3, -13, -26, -13, -5, -10, 1, -23, -20,
					-- layer=2 filter=168 channel=13
					4, -2, -10, -4, 0, 8, 7, 5, -2,
					-- layer=2 filter=168 channel=14
					-27, -23, -8, -18, -4, -15, 2, -6, -8,
					-- layer=2 filter=168 channel=15
					0, -13, 2, -2, -22, -10, 0, -7, 0,
					-- layer=2 filter=168 channel=16
					-6, -5, -4, -1, -9, 7, -9, -9, -6,
					-- layer=2 filter=168 channel=17
					0, 5, -3, 3, 5, -1, 4, -9, -8,
					-- layer=2 filter=168 channel=18
					-22, 8, -19, 2, 1, -15, 3, -11, -14,
					-- layer=2 filter=168 channel=19
					-17, -14, -18, -31, -26, -17, -15, -24, -21,
					-- layer=2 filter=168 channel=20
					-9, 0, 7, 6, -3, 0, 7, -1, 2,
					-- layer=2 filter=168 channel=21
					-7, -5, 7, 1, 8, 8, -1, -5, 10,
					-- layer=2 filter=168 channel=22
					-1, -1, 5, 7, -7, -3, -10, 11, -3,
					-- layer=2 filter=168 channel=23
					1, -4, -21, 10, -12, -18, 0, 2, -20,
					-- layer=2 filter=168 channel=24
					-17, -6, -3, -21, -10, 0, 0, -18, -19,
					-- layer=2 filter=168 channel=25
					-31, -16, -3, -8, -11, -18, -24, -20, -24,
					-- layer=2 filter=168 channel=26
					-7, 8, -9, 8, -2, -1, -1, 6, -3,
					-- layer=2 filter=168 channel=27
					-22, -3, -9, -18, 1, 0, -13, -9, -15,
					-- layer=2 filter=168 channel=28
					-17, -8, 7, 4, -12, -26, -7, -21, -16,
					-- layer=2 filter=168 channel=29
					-10, 5, -4, 0, -1, -11, -9, -1, 0,
					-- layer=2 filter=168 channel=30
					-12, -3, 5, 0, 9, 3, -14, -8, 0,
					-- layer=2 filter=168 channel=31
					-13, -5, 7, -10, -15, -12, -2, -7, -13,
					-- layer=2 filter=168 channel=32
					-3, -5, 5, 0, 8, -2, 11, -5, -8,
					-- layer=2 filter=168 channel=33
					1, -12, -21, -16, -7, 10, -13, -22, -10,
					-- layer=2 filter=168 channel=34
					-14, 20, -10, -13, -6, -1, -17, -16, -7,
					-- layer=2 filter=168 channel=35
					-32, 0, 1, -11, -15, -23, -17, -15, -17,
					-- layer=2 filter=168 channel=36
					0, -8, -1, 1, 4, -2, -6, -4, 4,
					-- layer=2 filter=168 channel=37
					-2, -14, -23, -15, -5, 1, -20, -23, 1,
					-- layer=2 filter=168 channel=38
					-8, -5, -5, -12, 14, 1, 0, -17, 2,
					-- layer=2 filter=168 channel=39
					19, 3, -11, 7, -7, -14, -4, -18, -3,
					-- layer=2 filter=168 channel=40
					-8, 3, -17, -11, -13, -1, -12, -14, -2,
					-- layer=2 filter=168 channel=41
					-7, 5, 5, -7, -12, 3, -11, -8, -8,
					-- layer=2 filter=168 channel=42
					2, -13, 2, -1, -22, -19, -8, -23, -2,
					-- layer=2 filter=168 channel=43
					-3, 24, 1, 3, 0, -22, 0, -14, -3,
					-- layer=2 filter=168 channel=44
					7, 3, -3, 5, 1, -5, -7, -5, 5,
					-- layer=2 filter=168 channel=45
					-1, -4, 1, -10, -5, -12, 0, -14, -11,
					-- layer=2 filter=168 channel=46
					-13, -12, -16, -21, -1, -5, -17, -8, -15,
					-- layer=2 filter=168 channel=47
					-25, -1, -23, -7, -7, -4, -1, -10, -13,
					-- layer=2 filter=168 channel=48
					9, 8, 7, -5, 9, -10, 6, -2, 9,
					-- layer=2 filter=168 channel=49
					-14, 10, 12, -23, 3, -6, 11, 7, -16,
					-- layer=2 filter=168 channel=50
					8, -7, -6, -4, -3, -4, -2, -8, 10,
					-- layer=2 filter=168 channel=51
					-8, -5, 2, -19, -21, -16, -6, -15, 0,
					-- layer=2 filter=168 channel=52
					-8, 1, -8, -15, -18, -10, -8, -26, -13,
					-- layer=2 filter=168 channel=53
					-3, -18, 13, -19, -4, -1, -16, -4, -6,
					-- layer=2 filter=168 channel=54
					-11, -5, -21, -20, -11, -9, -5, -15, -15,
					-- layer=2 filter=168 channel=55
					-5, -4, 6, 0, -5, -5, -5, -2, 5,
					-- layer=2 filter=168 channel=56
					-16, 14, -10, -3, -16, 2, -2, -22, -7,
					-- layer=2 filter=168 channel=57
					-10, -4, 4, 11, -1, -10, 8, 7, -9,
					-- layer=2 filter=168 channel=58
					-21, -18, 3, -16, -6, -14, -9, -10, -1,
					-- layer=2 filter=168 channel=59
					21, -8, -16, -20, 5, -13, -22, 11, -31,
					-- layer=2 filter=168 channel=60
					-8, -12, -19, -17, -5, -10, -20, -6, -17,
					-- layer=2 filter=168 channel=61
					13, -6, -2, 8, -7, -5, -18, -5, -5,
					-- layer=2 filter=168 channel=62
					-3, 3, -30, -2, -10, -18, 7, 7, -25,
					-- layer=2 filter=168 channel=63
					-2, -16, -24, 0, 5, -21, -4, -7, -19,
					-- layer=2 filter=168 channel=64
					0, -10, -2, 16, -4, -10, 11, -8, -4,
					-- layer=2 filter=168 channel=65
					19, -14, 0, 2, 5, 6, 0, 18, 23,
					-- layer=2 filter=168 channel=66
					8, 7, -10, -11, -10, -6, -7, 8, 0,
					-- layer=2 filter=168 channel=67
					-7, -7, -2, 0, -10, 2, 0, 0, 3,
					-- layer=2 filter=168 channel=68
					3, 8, 7, 8, -3, -2, -3, 3, 6,
					-- layer=2 filter=168 channel=69
					0, -12, -10, 14, -5, -13, 2, -11, -6,
					-- layer=2 filter=168 channel=70
					-17, 2, -14, -6, -23, -31, -30, -26, -4,
					-- layer=2 filter=168 channel=71
					-9, -12, -5, -14, 8, -7, -14, -8, -5,
					-- layer=2 filter=168 channel=72
					-24, -13, -18, -23, -14, 7, 8, -16, -27,
					-- layer=2 filter=168 channel=73
					-11, -3, -7, -24, -12, -1, -8, -15, -11,
					-- layer=2 filter=168 channel=74
					-4, -16, 9, -16, 3, -10, 0, -12, -4,
					-- layer=2 filter=168 channel=75
					-16, -15, 6, 15, -20, 0, -2, 15, 5,
					-- layer=2 filter=168 channel=76
					0, -7, -7, -12, -19, -4, -4, -13, -12,
					-- layer=2 filter=168 channel=77
					-1, -6, -11, 5, -9, -7, 5, 2, -8,
					-- layer=2 filter=168 channel=78
					-2, -6, -3, -6, 0, 0, 1, 6, -14,
					-- layer=2 filter=168 channel=79
					-1, -8, -8, 6, 0, 0, 5, -2, -10,
					-- layer=2 filter=168 channel=80
					1, 4, -8, 10, 10, -7, 19, 4, -21,
					-- layer=2 filter=168 channel=81
					-5, -3, 1, 7, -4, -6, -11, -1, 6,
					-- layer=2 filter=168 channel=82
					9, -1, 6, 5, 7, 1, 0, 7, 6,
					-- layer=2 filter=168 channel=83
					7, -12, 3, 9, -12, -15, -10, -9, -10,
					-- layer=2 filter=168 channel=84
					0, 5, 0, 6, 8, 0, -11, 7, 2,
					-- layer=2 filter=168 channel=85
					0, -5, -1, 0, 0, 9, 6, 0, -1,
					-- layer=2 filter=168 channel=86
					-10, -7, 9, -11, 7, 11, -2, 9, 10,
					-- layer=2 filter=168 channel=87
					-16, -17, -11, -7, -13, 4, -10, -3, -15,
					-- layer=2 filter=168 channel=88
					-6, -14, -7, 5, 12, 3, 6, 5, 9,
					-- layer=2 filter=168 channel=89
					-18, -34, -15, -8, -10, -10, -27, -6, -16,
					-- layer=2 filter=168 channel=90
					-6, 3, 0, 7, -2, -7, -6, -8, -3,
					-- layer=2 filter=168 channel=91
					-13, -21, -20, -16, -4, -17, -19, -6, -7,
					-- layer=2 filter=168 channel=92
					-19, -20, -13, -25, -8, -18, -1, -25, -19,
					-- layer=2 filter=168 channel=93
					1, -1, -24, 2, 11, -17, -6, 7, -8,
					-- layer=2 filter=168 channel=94
					12, -2, -15, -8, -22, 15, -32, -13, -6,
					-- layer=2 filter=168 channel=95
					-4, 10, 3, 0, -8, -2, 3, -7, -11,
					-- layer=2 filter=168 channel=96
					-30, -3, -5, -1, -1, 2, -5, 0, -5,
					-- layer=2 filter=168 channel=97
					-16, -9, -2, -10, 0, -11, -3, -13, -21,
					-- layer=2 filter=168 channel=98
					-15, -5, -19, -22, -28, -20, -13, -24, -24,
					-- layer=2 filter=168 channel=99
					-9, -2, -6, -39, -6, -22, -21, -9, -5,
					-- layer=2 filter=168 channel=100
					-10, -10, -3, -4, 3, -8, -21, -16, 6,
					-- layer=2 filter=168 channel=101
					-13, -26, -1, 1, 8, 1, 0, -7, -9,
					-- layer=2 filter=168 channel=102
					-5, -11, -14, 8, 0, 2, 1, 8, -6,
					-- layer=2 filter=168 channel=103
					-15, -7, -9, -2, -2, 2, 1, 0, -13,
					-- layer=2 filter=168 channel=104
					-22, -5, -12, -20, 4, 12, -2, 7, -22,
					-- layer=2 filter=168 channel=105
					1, -8, 2, -20, -4, 12, -4, 4, 0,
					-- layer=2 filter=168 channel=106
					-11, -7, 7, -5, -5, -15, 2, -4, -6,
					-- layer=2 filter=168 channel=107
					-17, -12, -6, 3, -17, -11, -7, -13, -9,
					-- layer=2 filter=168 channel=108
					-15, -16, -6, 0, -13, 0, 0, -19, -6,
					-- layer=2 filter=168 channel=109
					-10, -8, 5, -2, -1, 6, -8, -9, -3,
					-- layer=2 filter=168 channel=110
					4, -17, -26, 5, -25, -27, 12, -3, -27,
					-- layer=2 filter=168 channel=111
					-7, 3, 5, -6, 4, -11, 3, 0, 3,
					-- layer=2 filter=168 channel=112
					-13, -8, -4, 0, -9, 0, -18, -12, 14,
					-- layer=2 filter=168 channel=113
					-2, 1, 20, 15, -17, -2, -6, -18, 18,
					-- layer=2 filter=168 channel=114
					2, 1, -8, -8, 0, -10, 5, -8, -3,
					-- layer=2 filter=168 channel=115
					-3, 5, 0, -2, -11, -6, -6, 0, 7,
					-- layer=2 filter=168 channel=116
					-7, -4, -15, -23, -18, 15, -14, -4, -15,
					-- layer=2 filter=168 channel=117
					-14, -19, -13, -37, 0, -16, 8, -5, -21,
					-- layer=2 filter=168 channel=118
					8, 10, -11, 2, 16, 2, 16, -5, -17,
					-- layer=2 filter=168 channel=119
					-20, 9, 0, 8, -15, -22, 1, -7, -8,
					-- layer=2 filter=168 channel=120
					2, 0, 6, 6, 0, -8, 6, -3, -6,
					-- layer=2 filter=168 channel=121
					0, 8, -1, 2, -3, 2, 7, -7, -5,
					-- layer=2 filter=168 channel=122
					0, 0, -1, 7, -1, -9, -5, -6, -3,
					-- layer=2 filter=168 channel=123
					8, -36, -34, -5, -8, 12, -4, -15, 0,
					-- layer=2 filter=168 channel=124
					-5, -23, -9, -13, -30, -3, 3, -7, -14,
					-- layer=2 filter=168 channel=125
					-2, 9, -10, -7, -7, 5, 4, -5, 1,
					-- layer=2 filter=168 channel=126
					-9, 4, 4, -7, -3, -2, -13, -7, -4,
					-- layer=2 filter=168 channel=127
					-9, -20, -10, 2, -12, -22, 0, -7, -18,
					-- layer=2 filter=169 channel=0
					-7, -7, -10, -11, -20, -6, 3, 5, 16,
					-- layer=2 filter=169 channel=1
					-51, -23, -4, -22, -34, 28, -20, -20, -14,
					-- layer=2 filter=169 channel=2
					0, 7, 3, 7, -9, -1, -8, 2, -8,
					-- layer=2 filter=169 channel=3
					24, -26, -60, 24, 18, -52, 0, -4, -7,
					-- layer=2 filter=169 channel=4
					32, 26, -19, -28, -10, -4, -9, -39, -1,
					-- layer=2 filter=169 channel=5
					-7, -16, 21, -21, -6, 7, 8, -2, 22,
					-- layer=2 filter=169 channel=6
					-33, -1, 16, -29, 23, 36, 6, 30, 54,
					-- layer=2 filter=169 channel=7
					36, 21, 20, -8, 35, 34, -1, -44, -13,
					-- layer=2 filter=169 channel=8
					4, 2, -9, 1, 11, -8, 6, 0, 1,
					-- layer=2 filter=169 channel=9
					22, 12, -56, 33, -6, -46, 10, -36, -20,
					-- layer=2 filter=169 channel=10
					18, 20, -48, 48, 19, -53, -2, -9, 13,
					-- layer=2 filter=169 channel=11
					-18, -4, -3, 3, 0, 32, -3, 9, 22,
					-- layer=2 filter=169 channel=12
					-26, -4, -3, -14, -5, 21, -15, -5, -43,
					-- layer=2 filter=169 channel=13
					-1, 2, 9, 1, -6, 7, 2, -7, 2,
					-- layer=2 filter=169 channel=14
					-44, -26, 9, -2, -29, 7, -16, -24, -39,
					-- layer=2 filter=169 channel=15
					-33, 21, -27, -4, 8, -8, 9, -20, -9,
					-- layer=2 filter=169 channel=16
					12, 0, -8, -2, 8, -24, 9, -4, -4,
					-- layer=2 filter=169 channel=17
					3, 9, -8, 6, 9, 9, 7, 0, -2,
					-- layer=2 filter=169 channel=18
					-6, 10, 23, -33, -6, 51, 31, 12, -4,
					-- layer=2 filter=169 channel=19
					-37, -20, 2, 16, -18, 16, 1, 13, 21,
					-- layer=2 filter=169 channel=20
					-5, -7, 4, 7, 8, -8, 3, -2, 2,
					-- layer=2 filter=169 channel=21
					-5, 13, 6, 2, -4, -4, -2, 15, 0,
					-- layer=2 filter=169 channel=22
					9, 1, -4, -8, 4, 7, -8, -14, 4,
					-- layer=2 filter=169 channel=23
					19, -6, -2, -1, -20, -3, -14, -22, 34,
					-- layer=2 filter=169 channel=24
					51, 24, -71, 24, -21, -52, 11, -41, -31,
					-- layer=2 filter=169 channel=25
					19, 28, -34, 25, 11, -51, 3, -21, -34,
					-- layer=2 filter=169 channel=26
					-4, -7, -6, -3, 7, 0, -5, 6, 2,
					-- layer=2 filter=169 channel=27
					-14, -38, 16, 10, -4, 26, -19, -1, 13,
					-- layer=2 filter=169 channel=28
					9, 16, 42, 1, -10, 10, 40, 12, 7,
					-- layer=2 filter=169 channel=29
					-9, -1, -2, -4, 4, -8, -8, -8, -2,
					-- layer=2 filter=169 channel=30
					-1, -19, -15, 16, 0, -14, 4, 7, -34,
					-- layer=2 filter=169 channel=31
					43, 41, -22, -42, 0, 20, 7, 56, -15,
					-- layer=2 filter=169 channel=32
					2, 0, -5, -7, 4, -5, 4, -3, -9,
					-- layer=2 filter=169 channel=33
					-1, -5, 23, 0, -35, -10, 27, 13, -5,
					-- layer=2 filter=169 channel=34
					-32, 23, 0, 20, 43, -17, 63, 86, 9,
					-- layer=2 filter=169 channel=35
					-2, 28, 14, 1, -5, -21, 24, 17, -23,
					-- layer=2 filter=169 channel=36
					-6, -9, -2, -4, 0, 2, -3, 5, 0,
					-- layer=2 filter=169 channel=37
					-9, -10, 10, -8, 0, 22, 1, -6, 29,
					-- layer=2 filter=169 channel=38
					-22, -15, -5, 12, -22, 27, 6, 30, 34,
					-- layer=2 filter=169 channel=39
					50, 20, 19, -7, -1, -20, 31, -1, -16,
					-- layer=2 filter=169 channel=40
					0, 34, 6, -4, -16, -33, 18, 19, -38,
					-- layer=2 filter=169 channel=41
					0, 5, 7, 8, -2, 2, 9, 2, 8,
					-- layer=2 filter=169 channel=42
					-9, 1, 20, 14, 35, 25, -5, 6, -6,
					-- layer=2 filter=169 channel=43
					0, 1, -64, -17, -15, 3, -11, 7, -30,
					-- layer=2 filter=169 channel=44
					2, 4, -9, -3, 0, 2, -1, -9, 0,
					-- layer=2 filter=169 channel=45
					4, -9, 5, -10, -28, -9, -6, -5, -29,
					-- layer=2 filter=169 channel=46
					-10, 24, -19, 39, 13, -44, -11, -18, -34,
					-- layer=2 filter=169 channel=47
					32, 32, 7, 24, -3, -11, 43, 18, -12,
					-- layer=2 filter=169 channel=48
					-7, 5, 3, 6, -2, -7, 3, 8, -1,
					-- layer=2 filter=169 channel=49
					-37, -14, -4, -67, -9, 13, -36, -40, -7,
					-- layer=2 filter=169 channel=50
					-6, -2, -9, 3, -4, 0, 13, -9, 19,
					-- layer=2 filter=169 channel=51
					-9, 3, 15, -11, -12, -10, -10, 19, 5,
					-- layer=2 filter=169 channel=52
					-36, -4, -1, -31, 6, 10, -8, 24, 9,
					-- layer=2 filter=169 channel=53
					12, 3, 10, 25, 18, 10, 14, 3, -37,
					-- layer=2 filter=169 channel=54
					4, 31, 25, -3, -7, 5, 20, 3, 19,
					-- layer=2 filter=169 channel=55
					0, 0, 0, 0, 13, -1, -2, 13, 1,
					-- layer=2 filter=169 channel=56
					-4, -3, -3, -2, 2, 23, -12, 10, 9,
					-- layer=2 filter=169 channel=57
					7, 4, 4, -6, -14, -8, -8, -3, 3,
					-- layer=2 filter=169 channel=58
					0, 2, 5, 23, 8, 26, -18, 8, -18,
					-- layer=2 filter=169 channel=59
					-11, 8, -45, 29, 8, 32, -14, 3, 1,
					-- layer=2 filter=169 channel=60
					-9, 12, 0, 25, 11, -36, -17, -10, -1,
					-- layer=2 filter=169 channel=61
					-33, -2, 19, 4, 31, 12, -33, -25, -2,
					-- layer=2 filter=169 channel=62
					-22, -21, 12, 2, -13, 31, 16, 29, 50,
					-- layer=2 filter=169 channel=63
					5, 0, 6, -4, -7, -23, -45, -23, -14,
					-- layer=2 filter=169 channel=64
					22, 10, -14, 26, 14, -9, 6, -13, -41,
					-- layer=2 filter=169 channel=65
					-63, -29, 22, 13, 13, 31, 4, 1, 21,
					-- layer=2 filter=169 channel=66
					6, -29, 32, 21, -2, -12, -32, 19, -39,
					-- layer=2 filter=169 channel=67
					-6, -13, -67, 60, 35, -14, 23, 52, 7,
					-- layer=2 filter=169 channel=68
					1, 4, 6, 0, 6, 8, 6, -4, -3,
					-- layer=2 filter=169 channel=69
					6, 4, -7, -7, -22, -32, 2, -17, -20,
					-- layer=2 filter=169 channel=70
					10, -3, 58, 0, -9, -21, 8, 8, -8,
					-- layer=2 filter=169 channel=71
					-2, -37, 16, 20, 41, 39, 14, 18, 21,
					-- layer=2 filter=169 channel=72
					-1, -6, 41, -54, -16, 26, -10, -24, -57,
					-- layer=2 filter=169 channel=73
					-16, 18, -13, -38, -14, 5, -7, 28, -12,
					-- layer=2 filter=169 channel=74
					7, -10, -46, 49, 8, -28, -6, 47, -55,
					-- layer=2 filter=169 channel=75
					-76, -19, 66, 41, 28, 21, 32, -36, -54,
					-- layer=2 filter=169 channel=76
					-1, -38, -13, -1, 18, -17, -10, -19, -7,
					-- layer=2 filter=169 channel=77
					-1, 8, 8, -6, -6, -8, 9, 0, 6,
					-- layer=2 filter=169 channel=78
					8, -12, -14, -23, -2, 14, -4, 0, -3,
					-- layer=2 filter=169 channel=79
					9, 11, -5, 5, -3, 8, -7, -1, 3,
					-- layer=2 filter=169 channel=80
					22, -9, -31, 2, 3, -37, -9, -9, 9,
					-- layer=2 filter=169 channel=81
					-6, 2, -2, -2, -3, 5, 0, 6, -4,
					-- layer=2 filter=169 channel=82
					10, -10, 10, 10, 3, 7, 11, 3, -3,
					-- layer=2 filter=169 channel=83
					-5, -33, 32, -17, 3, 9, -13, -40, 17,
					-- layer=2 filter=169 channel=84
					9, 7, 3, 4, 6, 4, 4, 0, -8,
					-- layer=2 filter=169 channel=85
					1, -4, 4, 9, 13, -2, 9, 1, 7,
					-- layer=2 filter=169 channel=86
					7, -12, -14, 1, -12, 0, -3, -16, -21,
					-- layer=2 filter=169 channel=87
					21, 30, -29, 42, 50, 13, 27, 67, 12,
					-- layer=2 filter=169 channel=88
					-6, 3, -13, 22, -41, 22, 21, 46, -61,
					-- layer=2 filter=169 channel=89
					-39, -2, -23, 0, 2, 22, -42, -18, -30,
					-- layer=2 filter=169 channel=90
					1, -6, 0, -5, -10, 4, 11, 6, -3,
					-- layer=2 filter=169 channel=91
					-30, -5, -11, 20, 11, 0, -14, -7, -45,
					-- layer=2 filter=169 channel=92
					-22, -16, 10, -35, -5, 45, -29, -34, -21,
					-- layer=2 filter=169 channel=93
					-22, 3, -24, 6, -5, 7, 50, 23, 2,
					-- layer=2 filter=169 channel=94
					-51, 9, 18, -63, 0, 47, 4, 1, 36,
					-- layer=2 filter=169 channel=95
					1, 9, 13, 1, -8, -3, -6, 5, 6,
					-- layer=2 filter=169 channel=96
					-3, -39, -23, -18, 13, 25, -53, 42, 26,
					-- layer=2 filter=169 channel=97
					19, 12, -6, 28, -11, -5, 23, -3, -33,
					-- layer=2 filter=169 channel=98
					-2, 2, 0, -17, -20, 5, -8, -13, -22,
					-- layer=2 filter=169 channel=99
					-25, -19, 26, 13, 51, 23, 38, 9, 30,
					-- layer=2 filter=169 channel=100
					-29, 8, 18, 24, 19, 14, -9, 20, 42,
					-- layer=2 filter=169 channel=101
					-4, -6, 15, 23, 9, -39, 27, -19, -11,
					-- layer=2 filter=169 channel=102
					-9, -31, -13, -27, 21, 26, 10, 45, 2,
					-- layer=2 filter=169 channel=103
					-23, -25, 14, -17, -30, -69, -17, -57, 37,
					-- layer=2 filter=169 channel=104
					39, -1, 24, -62, 11, 36, -52, -4, 9,
					-- layer=2 filter=169 channel=105
					10, -28, -21, 38, -6, 6, -10, -24, 30,
					-- layer=2 filter=169 channel=106
					20, 19, -55, 46, -36, -36, 42, -19, -51,
					-- layer=2 filter=169 channel=107
					-27, 48, 10, -13, -21, 16, -31, 28, -15,
					-- layer=2 filter=169 channel=108
					-39, -37, -13, -27, 59, 38, -17, 10, 16,
					-- layer=2 filter=169 channel=109
					0, 3, -7, -5, 6, -2, 4, 0, 3,
					-- layer=2 filter=169 channel=110
					28, 22, -3, 32, 39, 17, 25, -7, -76,
					-- layer=2 filter=169 channel=111
					-3, 7, -4, 7, 1, -1, -6, -2, 0,
					-- layer=2 filter=169 channel=112
					4, 22, -25, 39, -21, -6, -2, -41, 28,
					-- layer=2 filter=169 channel=113
					-9, -27, 22, -1, -13, 0, -40, -43, -34,
					-- layer=2 filter=169 channel=114
					0, -5, 7, -3, -5, -4, 4, -8, 0,
					-- layer=2 filter=169 channel=115
					-1, 2, -8, 7, 4, 8, -3, -4, -12,
					-- layer=2 filter=169 channel=116
					-7, 2, -33, -11, 15, 9, 18, 54, 14,
					-- layer=2 filter=169 channel=117
					-24, -23, 40, -15, -8, -12, 10, -28, -9,
					-- layer=2 filter=169 channel=118
					0, -40, -34, 3, -6, 12, -51, 28, 13,
					-- layer=2 filter=169 channel=119
					-3, 20, 2, 2, 32, -1, 19, 27, -7,
					-- layer=2 filter=169 channel=120
					-1, 8, -8, -6, 5, -7, 10, 8, -7,
					-- layer=2 filter=169 channel=121
					-2, -3, 6, -1, -7, -6, -6, -3, 6,
					-- layer=2 filter=169 channel=122
					6, 0, -10, 4, 1, 13, -5, -7, 4,
					-- layer=2 filter=169 channel=123
					26, -4, 25, 10, 28, 19, 16, 0, -33,
					-- layer=2 filter=169 channel=124
					-3, 7, 33, 14, -6, 11, 7, 21, 30,
					-- layer=2 filter=169 channel=125
					-1, -2, -9, 12, -5, 10, -11, 4, 4,
					-- layer=2 filter=169 channel=126
					17, -8, -44, 48, -23, -3, 5, -8, 7,
					-- layer=2 filter=169 channel=127
					-11, -13, 8, 1, -25, 16, -53, -18, -2,
					-- layer=2 filter=170 channel=0
					-17, -45, -20, 5, -12, -17, 2, -25, -12,
					-- layer=2 filter=170 channel=1
					-25, -53, -3, -45, -28, 26, 35, -32, 1,
					-- layer=2 filter=170 channel=2
					8, 0, 1, 3, -7, 9, -8, 3, 6,
					-- layer=2 filter=170 channel=3
					20, 4, 11, -22, -1, -18, -35, -8, -29,
					-- layer=2 filter=170 channel=4
					30, 31, -20, 26, -23, 8, -27, -53, 5,
					-- layer=2 filter=170 channel=5
					-16, 0, -18, -17, -5, 6, -47, -13, 7,
					-- layer=2 filter=170 channel=6
					-7, -6, -17, 13, 0, -47, -5, -5, -41,
					-- layer=2 filter=170 channel=7
					54, -30, -24, -16, 11, 48, -34, -17, -10,
					-- layer=2 filter=170 channel=8
					-2, 9, -7, -7, 4, -4, 5, 4, -7,
					-- layer=2 filter=170 channel=9
					-34, -10, 1, -5, -65, 43, 24, -12, 78,
					-- layer=2 filter=170 channel=10
					-11, -11, 10, 10, -34, 11, 3, -32, -30,
					-- layer=2 filter=170 channel=11
					-19, -10, -4, -57, -1, 1, -52, -29, 1,
					-- layer=2 filter=170 channel=12
					-11, -5, 0, -21, 17, 29, 15, -7, 27,
					-- layer=2 filter=170 channel=13
					3, 0, 6, 7, -8, -1, 4, 2, -9,
					-- layer=2 filter=170 channel=14
					-7, -37, 11, -12, -11, -3, 23, 2, -27,
					-- layer=2 filter=170 channel=15
					-9, -35, -14, 7, 19, 16, 4, 9, -35,
					-- layer=2 filter=170 channel=16
					38, 15, 18, -35, -35, 36, -58, -28, 34,
					-- layer=2 filter=170 channel=17
					-4, 0, 7, -4, 0, 4, -6, 9, 6,
					-- layer=2 filter=170 channel=18
					18, 5, -5, -49, -8, 8, -48, 18, 1,
					-- layer=2 filter=170 channel=19
					-7, 16, -14, -3, -7, 33, -26, -46, -3,
					-- layer=2 filter=170 channel=20
					5, 12, 0, 8, -9, 1, 11, 0, 0,
					-- layer=2 filter=170 channel=21
					-8, 2, -4, -1, 7, 0, 12, 3, -12,
					-- layer=2 filter=170 channel=22
					-6, -2, -5, -10, -6, -9, -8, -10, -8,
					-- layer=2 filter=170 channel=23
					37, -6, 17, 31, -13, -2, 0, 2, -4,
					-- layer=2 filter=170 channel=24
					-29, -48, -61, -90, -26, -32, -41, 25, -11,
					-- layer=2 filter=170 channel=25
					-50, -48, -64, -62, 16, -47, -89, -26, -79,
					-- layer=2 filter=170 channel=26
					1, 0, 7, 0, -8, -3, -1, 6, 6,
					-- layer=2 filter=170 channel=27
					-35, 0, 8, -79, -24, 0, -38, -6, 14,
					-- layer=2 filter=170 channel=28
					37, 36, 39, 33, 23, -27, -34, -42, -21,
					-- layer=2 filter=170 channel=29
					-10, 6, -7, 8, 5, -4, -3, 5, 8,
					-- layer=2 filter=170 channel=30
					-49, -9, -13, 15, -10, 18, 20, -54, 9,
					-- layer=2 filter=170 channel=31
					88, 76, 35, 40, 66, 55, 46, 4, 40,
					-- layer=2 filter=170 channel=32
					-10, -11, -5, 7, -8, -9, 3, 3, -9,
					-- layer=2 filter=170 channel=33
					43, -3, -53, 32, 20, -14, 0, -3, -30,
					-- layer=2 filter=170 channel=34
					36, 45, 22, -29, 1, 18, -20, -3, -39,
					-- layer=2 filter=170 channel=35
					48, 37, 13, 29, -1, 13, -33, -52, -12,
					-- layer=2 filter=170 channel=36
					-1, -10, -3, 6, 2, -6, 5, -6, 6,
					-- layer=2 filter=170 channel=37
					-21, -10, 7, -25, -16, 22, -36, -17, 10,
					-- layer=2 filter=170 channel=38
					-80, -34, 12, -39, 25, -4, 30, -42, -9,
					-- layer=2 filter=170 channel=39
					31, -56, 11, -31, -31, 66, 26, 39, 38,
					-- layer=2 filter=170 channel=40
					69, -67, -40, 42, 67, 34, 19, 46, 15,
					-- layer=2 filter=170 channel=41
					-10, 4, 4, -6, 0, -1, 8, -3, -9,
					-- layer=2 filter=170 channel=42
					17, -7, 18, 3, -4, 41, -20, 9, 27,
					-- layer=2 filter=170 channel=43
					4, 22, -32, 12, -47, 28, -1, -30, -22,
					-- layer=2 filter=170 channel=44
					-6, -6, 4, 10, -9, -7, -3, 1, 12,
					-- layer=2 filter=170 channel=45
					22, 37, -28, -1, -23, 14, -20, 0, 17,
					-- layer=2 filter=170 channel=46
					-42, -11, 0, -17, -32, 6, 16, -17, -13,
					-- layer=2 filter=170 channel=47
					61, 9, 8, 45, 9, -12, 0, -32, -16,
					-- layer=2 filter=170 channel=48
					-1, 3, 9, -1, -7, 0, 4, 1, 2,
					-- layer=2 filter=170 channel=49
					0, 17, -24, -52, 6, 13, -45, 15, 33,
					-- layer=2 filter=170 channel=50
					14, -1, -11, 9, 8, 33, 13, -8, -9,
					-- layer=2 filter=170 channel=51
					-21, 2, 13, -21, -19, 1, -42, -35, -8,
					-- layer=2 filter=170 channel=52
					27, -42, -27, -52, -36, -12, -50, 16, 38,
					-- layer=2 filter=170 channel=53
					-11, 59, -14, 42, -21, 14, -43, -48, -2,
					-- layer=2 filter=170 channel=54
					32, 40, -8, -9, 13, 23, -52, -59, 0,
					-- layer=2 filter=170 channel=55
					2, -9, -8, -7, -9, 6, -7, 3, -3,
					-- layer=2 filter=170 channel=56
					-31, -10, -6, -53, -26, 17, -37, -34, -12,
					-- layer=2 filter=170 channel=57
					1, -4, -10, -3, 0, 9, -2, -1, 7,
					-- layer=2 filter=170 channel=58
					-17, 18, 22, 32, 34, 17, 16, -7, 21,
					-- layer=2 filter=170 channel=59
					-19, -20, -27, -2, 15, -8, 48, 23, -42,
					-- layer=2 filter=170 channel=60
					-22, 4, -13, 25, 62, 7, 61, -38, -33,
					-- layer=2 filter=170 channel=61
					14, -27, -55, -2, 30, -34, 17, 1, -40,
					-- layer=2 filter=170 channel=62
					-7, 9, -10, -31, -4, 0, -32, -25, -14,
					-- layer=2 filter=170 channel=63
					6, -30, -13, 31, 15, -10, 32, 18, 8,
					-- layer=2 filter=170 channel=64
					10, -9, -17, 7, -24, 5, 24, -1, 23,
					-- layer=2 filter=170 channel=65
					-49, -3, -47, -9, 28, -31, 24, 5, -36,
					-- layer=2 filter=170 channel=66
					6, 25, 17, 43, -10, 4, -7, -30, 7,
					-- layer=2 filter=170 channel=67
					-62, -35, 0, -18, 3, -1, -25, 1, 34,
					-- layer=2 filter=170 channel=68
					-3, -9, -4, 0, 4, -5, 2, -8, -7,
					-- layer=2 filter=170 channel=69
					3, -37, -5, 10, -19, 21, 7, -5, 43,
					-- layer=2 filter=170 channel=70
					44, 24, 9, 55, 6, 0, -49, -44, 6,
					-- layer=2 filter=170 channel=71
					-30, 60, 27, -31, -40, 30, -95, -20, -2,
					-- layer=2 filter=170 channel=72
					20, -10, 23, -39, -6, 1, 23, 3, -62,
					-- layer=2 filter=170 channel=73
					17, 40, 6, 6, 18, -38, -19, -43, -15,
					-- layer=2 filter=170 channel=74
					-17, -50, -23, 3, -11, -45, 28, -2, 18,
					-- layer=2 filter=170 channel=75
					-26, 0, -4, 5, -4, -25, -23, 0, 17,
					-- layer=2 filter=170 channel=76
					26, 27, -19, 41, 0, 30, 43, -44, 22,
					-- layer=2 filter=170 channel=77
					0, 4, -1, 8, 5, -11, 3, 0, -11,
					-- layer=2 filter=170 channel=78
					-1, 1, -48, -62, -14, 9, -53, -16, 4,
					-- layer=2 filter=170 channel=79
					0, 11, 2, 5, 8, 5, 0, 5, 3,
					-- layer=2 filter=170 channel=80
					35, -18, 10, 17, -7, 10, -17, -10, 37,
					-- layer=2 filter=170 channel=81
					-11, -8, 7, 6, -2, -5, -4, 2, -11,
					-- layer=2 filter=170 channel=82
					8, -2, 7, 6, -3, 0, 8, 4, 0,
					-- layer=2 filter=170 channel=83
					11, -3, 31, 39, -11, 16, -19, -39, 1,
					-- layer=2 filter=170 channel=84
					11, 0, -11, -8, 5, 3, 3, 0, -11,
					-- layer=2 filter=170 channel=85
					1, 4, 9, 2, 5, -6, -5, 7, 8,
					-- layer=2 filter=170 channel=86
					-9, 0, -11, -5, -11, -12, 5, 6, -15,
					-- layer=2 filter=170 channel=87
					16, -14, -8, 12, 12, 30, -64, 31, -6,
					-- layer=2 filter=170 channel=88
					-22, -23, -52, 6, -19, -16, 58, -12, 0,
					-- layer=2 filter=170 channel=89
					-37, -29, 9, -14, 11, 25, 41, -2, -21,
					-- layer=2 filter=170 channel=90
					4, -8, 2, 0, 1, -7, -7, 3, 2,
					-- layer=2 filter=170 channel=91
					-51, 11, 34, 7, 26, 16, 21, -19, 1,
					-- layer=2 filter=170 channel=92
					2, -51, 14, -39, 0, 28, 52, -5, 1,
					-- layer=2 filter=170 channel=93
					38, 25, -3, 5, 31, -35, -18, -26, -35,
					-- layer=2 filter=170 channel=94
					-11, -5, 0, -18, 26, 37, 2, -1, -41,
					-- layer=2 filter=170 channel=95
					-6, -12, 1, 5, 4, -2, -1, -3, 7,
					-- layer=2 filter=170 channel=96
					33, 21, -1, -28, 33, -29, -36, 17, -19,
					-- layer=2 filter=170 channel=97
					-15, -11, -42, -23, -47, -12, -53, -30, 22,
					-- layer=2 filter=170 channel=98
					37, 8, 1, 59, 3, 3, -13, -11, -27,
					-- layer=2 filter=170 channel=99
					-6, -47, 21, 2, -10, 33, -15, -33, 30,
					-- layer=2 filter=170 channel=100
					-20, -2, 2, 0, 42, -1, 13, -33, -8,
					-- layer=2 filter=170 channel=101
					-63, -25, -27, -75, -30, -24, -131, -130, -43,
					-- layer=2 filter=170 channel=102
					-21, 18, 6, -47, -23, 14, -82, 0, 45,
					-- layer=2 filter=170 channel=103
					45, 17, 50, -43, -1, 32, 22, 6, 59,
					-- layer=2 filter=170 channel=104
					-23, 40, 15, -65, 44, 4, -71, -2, -12,
					-- layer=2 filter=170 channel=105
					-39, 5, 37, 48, -60, 24, -33, -36, -6,
					-- layer=2 filter=170 channel=106
					-70, -28, -43, -47, -4, -50, -72, -47, -22,
					-- layer=2 filter=170 channel=107
					26, 16, 23, 7, 20, 33, 20, 7, 15,
					-- layer=2 filter=170 channel=108
					5, 8, 8, -42, -42, 6, -7, -24, 17,
					-- layer=2 filter=170 channel=109
					9, 7, -1, 7, 12, 1, -12, 5, -6,
					-- layer=2 filter=170 channel=110
					30, -25, 11, 10, 20, -22, -23, 28, -8,
					-- layer=2 filter=170 channel=111
					2, 4, -6, -10, 3, -10, -8, 1, -11,
					-- layer=2 filter=170 channel=112
					-20, -25, -74, -26, 6, 4, -38, -34, -18,
					-- layer=2 filter=170 channel=113
					-24, 2, 5, 36, 8, 2, 26, -20, 34,
					-- layer=2 filter=170 channel=114
					7, 3, -1, -4, 18, -5, 1, 8, 2,
					-- layer=2 filter=170 channel=115
					-2, 9, -6, -7, 4, -10, 0, 7, 0,
					-- layer=2 filter=170 channel=116
					21, -32, -3, -2, 36, 29, -26, 26, 0,
					-- layer=2 filter=170 channel=117
					40, -7, 2, -58, -23, 32, -39, -66, -22,
					-- layer=2 filter=170 channel=118
					-10, 10, -18, 30, 2, -19, -37, -33, -16,
					-- layer=2 filter=170 channel=119
					28, 16, -3, -42, -23, -4, -78, -16, -6,
					-- layer=2 filter=170 channel=120
					5, 2, -9, 3, -2, 2, 6, 0, 4,
					-- layer=2 filter=170 channel=121
					-11, -5, 1, -8, -2, 4, 7, 1, -6,
					-- layer=2 filter=170 channel=122
					-7, 1, -4, 10, 3, -7, 1, 3, -6,
					-- layer=2 filter=170 channel=123
					25, -29, -18, 18, -1, -1, -10, 17, -34,
					-- layer=2 filter=170 channel=124
					2, -15, -36, -10, 11, 11, -39, -12, -15,
					-- layer=2 filter=170 channel=125
					-2, 4, -10, -2, -11, 2, -11, 0, -9,
					-- layer=2 filter=170 channel=126
					21, 17, 14, 26, 39, -71, 48, 0, -107,
					-- layer=2 filter=170 channel=127
					-50, -4, 6, 32, 11, -20, 47, 1, -14,
					-- layer=2 filter=171 channel=0
					-2, -7, 0, -2, -14, -14, -10, -13, -7,
					-- layer=2 filter=171 channel=1
					0, -8, 1, -21, -16, -23, -5, -19, -9,
					-- layer=2 filter=171 channel=2
					-4, 1, 7, 0, 7, 0, 7, 5, -1,
					-- layer=2 filter=171 channel=3
					-4, -13, -17, 10, -13, -17, -24, -6, 0,
					-- layer=2 filter=171 channel=4
					-11, -28, 4, -2, 1, -9, 5, 1, 17,
					-- layer=2 filter=171 channel=5
					-6, 5, 8, 4, -27, 8, 0, -3, -18,
					-- layer=2 filter=171 channel=6
					-4, -20, -3, -6, -30, -22, -14, 9, 9,
					-- layer=2 filter=171 channel=7
					0, -20, 21, 0, 0, -10, -10, -29, 4,
					-- layer=2 filter=171 channel=8
					-3, 0, -11, 9, 0, 1, 4, -3, -3,
					-- layer=2 filter=171 channel=9
					-16, -4, -11, 11, -22, -18, 3, 8, -15,
					-- layer=2 filter=171 channel=10
					-17, 9, -17, 4, -15, -2, 12, -11, -15,
					-- layer=2 filter=171 channel=11
					-13, -5, 24, -9, -6, -22, -20, -14, -1,
					-- layer=2 filter=171 channel=12
					-5, -16, 7, 6, -2, 6, -5, 8, -7,
					-- layer=2 filter=171 channel=13
					-7, 8, -5, 0, -7, -8, 8, 7, 7,
					-- layer=2 filter=171 channel=14
					-9, -4, -1, -6, -10, -3, -12, -7, 2,
					-- layer=2 filter=171 channel=15
					-5, -10, -11, -11, -8, 10, -9, -10, 16,
					-- layer=2 filter=171 channel=16
					-7, 14, -9, -8, 3, 7, -7, 7, -2,
					-- layer=2 filter=171 channel=17
					-10, 1, 1, 1, 9, -5, -1, 0, -1,
					-- layer=2 filter=171 channel=18
					4, -13, 0, -12, -21, -26, -13, -7, -2,
					-- layer=2 filter=171 channel=19
					-17, -12, -2, -10, -2, -7, -3, -17, -14,
					-- layer=2 filter=171 channel=20
					-5, -4, 8, 8, 3, -2, 1, -1, 11,
					-- layer=2 filter=171 channel=21
					9, 8, -8, -4, 7, 4, 5, 6, -1,
					-- layer=2 filter=171 channel=22
					-3, -8, 2, -6, 9, -10, 9, -6, 1,
					-- layer=2 filter=171 channel=23
					-17, -10, 2, -12, -28, -10, -18, -18, -15,
					-- layer=2 filter=171 channel=24
					0, -1, -10, -11, -15, -7, 4, -4, -5,
					-- layer=2 filter=171 channel=25
					12, -9, -9, 1, -9, -4, -13, 4, 4,
					-- layer=2 filter=171 channel=26
					-7, -8, 7, 4, 9, 9, -9, 3, 1,
					-- layer=2 filter=171 channel=27
					-12, -24, -8, 8, 10, -13, 1, -3, -32,
					-- layer=2 filter=171 channel=28
					26, 8, -1, -3, -18, 7, -17, -30, 0,
					-- layer=2 filter=171 channel=29
					-5, 9, 0, -2, 3, 2, 4, -3, 8,
					-- layer=2 filter=171 channel=30
					-9, -6, -4, -21, 4, 16, -3, -17, 0,
					-- layer=2 filter=171 channel=31
					0, 1, -12, 0, 4, 5, 8, -10, -10,
					-- layer=2 filter=171 channel=32
					0, -8, 7, 3, -6, -11, -4, 10, -3,
					-- layer=2 filter=171 channel=33
					-2, -4, 15, -14, 3, 2, -20, -22, 18,
					-- layer=2 filter=171 channel=34
					6, -5, -18, -7, -25, 7, -3, -6, -6,
					-- layer=2 filter=171 channel=35
					15, 11, 9, -7, -23, 4, -7, -16, -7,
					-- layer=2 filter=171 channel=36
					0, 2, -3, -9, 8, -7, -5, -3, 8,
					-- layer=2 filter=171 channel=37
					12, -17, -15, 4, -18, 12, -14, -8, -9,
					-- layer=2 filter=171 channel=38
					1, -4, -12, 9, -20, -5, 0, -27, -13,
					-- layer=2 filter=171 channel=39
					-12, -18, -12, 17, 6, -7, -3, 4, 8,
					-- layer=2 filter=171 channel=40
					-3, -14, -7, -7, -1, -9, -4, -8, -3,
					-- layer=2 filter=171 channel=41
					5, 8, -6, -6, 2, -11, 7, -4, 3,
					-- layer=2 filter=171 channel=42
					7, -6, -4, -14, -9, 0, -10, 0, -1,
					-- layer=2 filter=171 channel=43
					-9, -16, -18, -1, -8, 5, 0, -10, -7,
					-- layer=2 filter=171 channel=44
					-10, -1, -7, 0, 2, 4, -4, 8, 6,
					-- layer=2 filter=171 channel=45
					-2, -4, 0, -12, -10, -9, -8, 2, -8,
					-- layer=2 filter=171 channel=46
					-22, -24, -20, -7, -7, 3, 6, 12, -5,
					-- layer=2 filter=171 channel=47
					2, 1, -14, -10, -21, 1, -21, 0, 4,
					-- layer=2 filter=171 channel=48
					-10, -4, 4, -4, -1, 4, -9, -5, -4,
					-- layer=2 filter=171 channel=49
					-16, -13, -8, -1, -9, -9, -19, -2, -2,
					-- layer=2 filter=171 channel=50
					-3, -3, 4, -2, -9, 3, -2, -3, 7,
					-- layer=2 filter=171 channel=51
					-6, 4, -4, -8, -16, 10, -23, -11, 9,
					-- layer=2 filter=171 channel=52
					-22, -23, -6, -8, -18, 5, -1, -4, 4,
					-- layer=2 filter=171 channel=53
					-2, -4, 1, 1, -11, -8, 0, -4, -12,
					-- layer=2 filter=171 channel=54
					-29, -19, 3, -11, -21, -25, -9, 0, -22,
					-- layer=2 filter=171 channel=55
					-7, 0, -6, 0, 6, -9, 2, 9, -1,
					-- layer=2 filter=171 channel=56
					-3, 2, 1, -12, -18, 1, -13, -18, 14,
					-- layer=2 filter=171 channel=57
					4, -4, -2, 2, 0, -1, -3, -9, 2,
					-- layer=2 filter=171 channel=58
					-8, -15, -6, 6, -12, 1, -9, 11, -16,
					-- layer=2 filter=171 channel=59
					-6, -18, 8, 13, -6, -19, -13, 2, 4,
					-- layer=2 filter=171 channel=60
					-2, 7, -32, 11, -7, 10, -2, 4, -9,
					-- layer=2 filter=171 channel=61
					-10, -9, -16, -8, -16, -10, 7, -18, -11,
					-- layer=2 filter=171 channel=62
					-14, -9, -3, -3, -7, -44, -10, -19, 6,
					-- layer=2 filter=171 channel=63
					-14, -10, -12, -10, -19, -27, 0, 7, -5,
					-- layer=2 filter=171 channel=64
					-15, -11, -9, -1, -14, -17, -2, 0, -17,
					-- layer=2 filter=171 channel=65
					-7, 11, 2, 0, -21, -9, -17, -6, -5,
					-- layer=2 filter=171 channel=66
					2, -3, 3, 2, 2, -3, 7, -8, 6,
					-- layer=2 filter=171 channel=67
					-12, -23, -17, 10, -9, -22, 12, -6, -9,
					-- layer=2 filter=171 channel=68
					-4, -2, -1, 4, -6, 6, 0, -1, 0,
					-- layer=2 filter=171 channel=69
					-17, -4, 5, -13, -16, 11, -10, 5, 0,
					-- layer=2 filter=171 channel=70
					6, 0, -5, -25, -7, 8, -14, -16, -25,
					-- layer=2 filter=171 channel=71
					-12, -21, -13, -11, -14, -12, -5, 11, 7,
					-- layer=2 filter=171 channel=72
					25, -26, 10, -10, 9, -11, -28, -17, 3,
					-- layer=2 filter=171 channel=73
					-16, -7, -4, -19, 7, 0, 7, 0, -1,
					-- layer=2 filter=171 channel=74
					-18, -16, -10, 23, -17, -9, 2, 0, -4,
					-- layer=2 filter=171 channel=75
					12, -17, -2, -6, -4, 3, -11, 5, 0,
					-- layer=2 filter=171 channel=76
					1, -3, 7, -4, 0, -2, 0, -8, -19,
					-- layer=2 filter=171 channel=77
					-4, 3, 1, -4, -9, -8, 0, 5, 4,
					-- layer=2 filter=171 channel=78
					-4, -23, 10, -1, -9, -13, -12, -11, 1,
					-- layer=2 filter=171 channel=79
					5, 6, 1, -7, 2, 9, -2, -7, 0,
					-- layer=2 filter=171 channel=80
					-24, -6, -2, 8, 18, -6, -3, 8, 1,
					-- layer=2 filter=171 channel=81
					2, 2, 6, -5, 3, -3, -11, 2, 3,
					-- layer=2 filter=171 channel=82
					-10, -10, 3, 5, 0, 0, -1, -11, 1,
					-- layer=2 filter=171 channel=83
					-27, -18, -11, -12, -14, 16, -4, -16, 5,
					-- layer=2 filter=171 channel=84
					1, -1, -10, 4, -4, 4, -3, -2, -10,
					-- layer=2 filter=171 channel=85
					5, -10, -3, 4, 2, 8, 5, -6, 8,
					-- layer=2 filter=171 channel=86
					-4, 7, 1, -2, -7, 6, -5, -10, -6,
					-- layer=2 filter=171 channel=87
					4, -21, 12, -6, 13, 0, -13, -1, -1,
					-- layer=2 filter=171 channel=88
					-1, -4, -5, -16, -16, -6, -7, 3, -8,
					-- layer=2 filter=171 channel=89
					-21, -11, 16, -14, 1, -3, -8, 10, 6,
					-- layer=2 filter=171 channel=90
					-4, -3, 5, 4, -9, -5, -5, 8, 2,
					-- layer=2 filter=171 channel=91
					9, -9, -24, 1, -7, -6, -16, 9, -17,
					-- layer=2 filter=171 channel=92
					8, -6, 8, 21, 0, -12, -6, 10, -6,
					-- layer=2 filter=171 channel=93
					-1, 6, -9, -12, -6, -7, -2, 0, -17,
					-- layer=2 filter=171 channel=94
					-4, -21, 17, -9, -21, -15, -1, -8, 7,
					-- layer=2 filter=171 channel=95
					-9, -8, 7, 6, 1, -4, -7, -11, -11,
					-- layer=2 filter=171 channel=96
					4, 8, 13, -10, 3, -8, -16, -1, -17,
					-- layer=2 filter=171 channel=97
					-9, -4, -17, -1, -20, -5, -17, 5, 10,
					-- layer=2 filter=171 channel=98
					10, 6, -11, -13, -4, -12, -12, -1, 7,
					-- layer=2 filter=171 channel=99
					-6, -4, -6, -13, -2, -17, 8, -5, -13,
					-- layer=2 filter=171 channel=100
					-16, 0, -18, 4, -19, 15, -3, 4, -18,
					-- layer=2 filter=171 channel=101
					-17, -17, 0, 2, 0, 0, 10, 11, -5,
					-- layer=2 filter=171 channel=102
					12, -6, 8, -28, 3, -1, -1, 8, -7,
					-- layer=2 filter=171 channel=103
					-8, 7, -7, -1, 8, -2, -8, -13, 7,
					-- layer=2 filter=171 channel=104
					-2, -21, 22, -18, 0, -1, -6, -1, 13,
					-- layer=2 filter=171 channel=105
					0, -12, -5, -18, -6, -1, 0, 4, 21,
					-- layer=2 filter=171 channel=106
					2, 10, -13, -6, -10, -18, -28, -16, -25,
					-- layer=2 filter=171 channel=107
					11, -14, -8, -4, -8, -9, -9, 2, 3,
					-- layer=2 filter=171 channel=108
					-16, 0, -32, -15, -22, -12, -7, -1, -16,
					-- layer=2 filter=171 channel=109
					8, 0, -6, 2, 2, -2, -4, -5, -2,
					-- layer=2 filter=171 channel=110
					-25, -20, -21, -6, -5, -10, -7, -1, -9,
					-- layer=2 filter=171 channel=111
					4, 7, 9, 7, -5, -6, -8, 4, 7,
					-- layer=2 filter=171 channel=112
					-10, 3, -12, -1, -16, -15, 0, -12, -20,
					-- layer=2 filter=171 channel=113
					-11, 4, -31, -21, -22, 9, -9, -18, 0,
					-- layer=2 filter=171 channel=114
					10, -1, 5, 11, 1, 7, 5, -9, 3,
					-- layer=2 filter=171 channel=115
					-8, -6, -8, 8, 4, -7, 5, -6, 3,
					-- layer=2 filter=171 channel=116
					20, -26, 18, -5, -4, -14, -12, -10, -8,
					-- layer=2 filter=171 channel=117
					-8, -16, -14, -16, -24, -3, -9, 2, 1,
					-- layer=2 filter=171 channel=118
					-5, -19, -24, 2, 2, -6, -6, 0, -6,
					-- layer=2 filter=171 channel=119
					-15, -22, -5, -18, -10, -9, -25, -8, -20,
					-- layer=2 filter=171 channel=120
					7, -2, 7, 9, 7, -4, 6, -4, -1,
					-- layer=2 filter=171 channel=121
					-5, 7, 3, 2, 2, -1, 7, -2, -10,
					-- layer=2 filter=171 channel=122
					7, 5, 10, 7, 4, -8, 1, 1, 8,
					-- layer=2 filter=171 channel=123
					-10, -20, -10, -24, -18, -29, -14, 3, -1,
					-- layer=2 filter=171 channel=124
					-13, -11, -4, -6, -11, 6, -4, -10, 18,
					-- layer=2 filter=171 channel=125
					1, 5, -9, 8, -9, 8, 0, 0, -1,
					-- layer=2 filter=171 channel=126
					-12, -7, -6, -11, -6, 1, -10, -1, -5,
					-- layer=2 filter=171 channel=127
					2, -21, -7, -10, -21, 6, -16, -4, -10,
					-- layer=2 filter=172 channel=0
					-15, 1, 6, -12, 2, 4, 12, 10, 29,
					-- layer=2 filter=172 channel=1
					15, -30, -32, 26, -6, -47, 24, -14, -21,
					-- layer=2 filter=172 channel=2
					6, 1, 1, -9, 0, 9, 5, 5, -7,
					-- layer=2 filter=172 channel=3
					-15, 16, 40, -23, 13, 17, -50, -2, 26,
					-- layer=2 filter=172 channel=4
					-8, -30, -8, 3, -12, -23, 9, 4, 28,
					-- layer=2 filter=172 channel=5
					-13, -29, 23, -46, 1, -10, 0, 0, 8,
					-- layer=2 filter=172 channel=6
					-24, -32, -10, -14, -51, -36, 17, -37, -42,
					-- layer=2 filter=172 channel=7
					-6, -5, 7, 47, -1, 4, 1, 40, 20,
					-- layer=2 filter=172 channel=8
					-6, -9, 8, 10, 5, 4, -1, 5, 3,
					-- layer=2 filter=172 channel=9
					0, 10, -13, -9, 5, 0, -12, 12, 0,
					-- layer=2 filter=172 channel=10
					9, 12, 23, -19, 22, 27, -15, 13, 39,
					-- layer=2 filter=172 channel=11
					-16, 1, 19, -11, 7, 12, -8, 20, 13,
					-- layer=2 filter=172 channel=12
					-26, -22, 5, 32, -27, -29, 19, -24, -19,
					-- layer=2 filter=172 channel=13
					-1, -1, 6, -6, 7, -5, 0, -6, 3,
					-- layer=2 filter=172 channel=14
					0, -13, -7, 11, 28, -2, 31, 25, 21,
					-- layer=2 filter=172 channel=15
					-26, -2, 18, 6, -21, -20, -5, -38, -36,
					-- layer=2 filter=172 channel=16
					-4, -10, -19, 25, -11, -4, 26, 10, 1,
					-- layer=2 filter=172 channel=17
					-4, 0, 2, -4, 7, -11, 9, -3, -2,
					-- layer=2 filter=172 channel=18
					19, -13, -11, 26, 6, -18, 10, 8, -31,
					-- layer=2 filter=172 channel=19
					6, -29, -14, 39, 4, -34, 42, 12, -41,
					-- layer=2 filter=172 channel=20
					1, 9, -11, 9, 8, -4, -1, -6, -4,
					-- layer=2 filter=172 channel=21
					13, -20, -18, -6, -6, -15, -2, 6, -19,
					-- layer=2 filter=172 channel=22
					-9, -7, 0, -1, -6, -7, -2, 6, -6,
					-- layer=2 filter=172 channel=23
					15, -15, -12, 11, -20, -18, 28, -14, 19,
					-- layer=2 filter=172 channel=24
					0, 14, 11, -13, 23, 22, -11, 13, 4,
					-- layer=2 filter=172 channel=25
					-34, 14, 15, -25, -7, 5, -32, -6, 2,
					-- layer=2 filter=172 channel=26
					4, 3, 5, 5, 3, -6, 1, 2, 7,
					-- layer=2 filter=172 channel=27
					16, 23, 34, -13, 13, 15, -19, 10, 3,
					-- layer=2 filter=172 channel=28
					15, 6, 27, 29, -5, 21, 22, 17, 14,
					-- layer=2 filter=172 channel=29
					6, -4, 11, 11, 3, 6, -5, -9, 9,
					-- layer=2 filter=172 channel=30
					14, 14, -55, 34, 41, -5, 22, 22, -21,
					-- layer=2 filter=172 channel=31
					30, 19, 14, 31, -40, -40, 20, -37, -31,
					-- layer=2 filter=172 channel=32
					-4, -8, 0, -2, -3, -6, -4, -9, 6,
					-- layer=2 filter=172 channel=33
					0, -20, 31, 9, -52, -37, -22, -42, -9,
					-- layer=2 filter=172 channel=34
					36, -77, -88, 46, -63, -32, 34, -51, -95,
					-- layer=2 filter=172 channel=35
					15, -11, 0, -2, 2, 17, -14, -21, -17,
					-- layer=2 filter=172 channel=36
					2, 4, 0, 8, -12, 1, -7, 0, 0,
					-- layer=2 filter=172 channel=37
					-19, 0, 21, 0, 3, 14, -13, -10, 24,
					-- layer=2 filter=172 channel=38
					-1, -22, -40, -33, 6, -10, -28, -3, -1,
					-- layer=2 filter=172 channel=39
					-12, -1, -25, 0, -11, 3, -3, 19, 25,
					-- layer=2 filter=172 channel=40
					36, 38, -28, 10, -33, -51, -5, -74, -38,
					-- layer=2 filter=172 channel=41
					-5, 10, 6, 8, -9, 0, -12, 10, -10,
					-- layer=2 filter=172 channel=42
					-4, -4, 2, 18, -5, 3, 10, -8, 4,
					-- layer=2 filter=172 channel=43
					-7, 18, 56, -40, 22, 36, -60, -33, -9,
					-- layer=2 filter=172 channel=44
					-10, 8, 0, -3, -5, 5, 6, 4, 3,
					-- layer=2 filter=172 channel=45
					-6, -9, 43, -49, -1, 45, -12, 21, 15,
					-- layer=2 filter=172 channel=46
					-3, -16, -25, -6, 2, -8, -14, 21, 4,
					-- layer=2 filter=172 channel=47
					-2, 18, 10, 22, -12, -6, 36, 36, 26,
					-- layer=2 filter=172 channel=48
					-9, 0, 7, 2, -4, 5, -1, 8, -10,
					-- layer=2 filter=172 channel=49
					18, -9, 5, 55, 37, -20, 48, 43, -21,
					-- layer=2 filter=172 channel=50
					0, 3, -20, 1, 11, 7, 16, 18, 13,
					-- layer=2 filter=172 channel=51
					-9, -3, 15, -1, 15, 22, 10, -10, 9,
					-- layer=2 filter=172 channel=52
					-17, -9, -21, 4, 1, 50, 28, -11, -9,
					-- layer=2 filter=172 channel=53
					-26, 20, -21, -4, -31, -26, -16, 11, -5,
					-- layer=2 filter=172 channel=54
					-15, -14, 19, 17, -22, -39, 62, 8, 12,
					-- layer=2 filter=172 channel=55
					0, -10, 7, 12, -11, -4, 9, 8, 2,
					-- layer=2 filter=172 channel=56
					-17, -1, 24, -35, -6, 19, -21, 8, 11,
					-- layer=2 filter=172 channel=57
					-6, -3, 14, -5, 3, 10, 4, -5, 6,
					-- layer=2 filter=172 channel=58
					0, -68, -19, 1, -51, -67, -30, -45, -4,
					-- layer=2 filter=172 channel=59
					-6, -61, -23, -38, -102, -88, -50, -44, -22,
					-- layer=2 filter=172 channel=60
					-30, -28, -37, -27, -19, -64, 8, -20, -17,
					-- layer=2 filter=172 channel=61
					33, 35, 20, 24, 53, 44, 50, 13, -22,
					-- layer=2 filter=172 channel=62
					-1, -51, -53, 14, -27, -48, 36, -1, -45,
					-- layer=2 filter=172 channel=63
					1, -7, -7, -21, -2, -26, 22, 19, 27,
					-- layer=2 filter=172 channel=64
					17, -20, -32, 50, 2, -18, 42, 2, -2,
					-- layer=2 filter=172 channel=65
					36, 37, -37, 31, 28, 20, 67, -30, -43,
					-- layer=2 filter=172 channel=66
					-44, 36, 20, 20, 4, -4, 37, -6, 0,
					-- layer=2 filter=172 channel=67
					3, -14, -15, -41, -18, 3, -47, -10, 0,
					-- layer=2 filter=172 channel=68
					-2, 2, 7, 3, -9, 0, -6, -4, 0,
					-- layer=2 filter=172 channel=69
					-7, -2, -22, 30, 12, -9, 25, 6, -9,
					-- layer=2 filter=172 channel=70
					19, 23, 17, 15, -1, 28, 2, 12, 20,
					-- layer=2 filter=172 channel=71
					22, 22, 52, -46, -23, 9, -49, -8, -5,
					-- layer=2 filter=172 channel=72
					2, 0, 26, 43, 1, -18, 19, 19, 26,
					-- layer=2 filter=172 channel=73
					-2, 9, 26, 27, -5, 50, 27, 51, 33,
					-- layer=2 filter=172 channel=74
					-34, -9, -26, -21, -23, -4, -51, -14, 0,
					-- layer=2 filter=172 channel=75
					48, -39, -20, 12, -19, 39, -19, 9, -35,
					-- layer=2 filter=172 channel=76
					-2, -26, 4, 7, -48, -1, -26, -36, 2,
					-- layer=2 filter=172 channel=77
					2, -4, -5, 0, 3, 0, -4, 3, -9,
					-- layer=2 filter=172 channel=78
					-17, -17, 0, 5, 30, 25, 5, -7, -12,
					-- layer=2 filter=172 channel=79
					-5, 7, 9, 8, 9, 7, 0, 5, 8,
					-- layer=2 filter=172 channel=80
					20, -7, -22, 28, 7, -18, 25, 8, -5,
					-- layer=2 filter=172 channel=81
					14, 12, 9, 8, 13, 7, 6, 1, 10,
					-- layer=2 filter=172 channel=82
					0, 7, 2, 6, -5, -5, -4, -1, 3,
					-- layer=2 filter=172 channel=83
					20, -8, 3, 27, 5, -6, 39, 18, 13,
					-- layer=2 filter=172 channel=84
					8, 10, 0, 6, 11, 7, -2, -6, 2,
					-- layer=2 filter=172 channel=85
					3, 3, -12, 14, -10, 0, 2, 0, 1,
					-- layer=2 filter=172 channel=86
					-6, 2, -8, -5, -5, 11, 9, 1, 16,
					-- layer=2 filter=172 channel=87
					-44, -81, -114, -43, -111, -89, -98, -141, -67,
					-- layer=2 filter=172 channel=88
					-13, 8, -18, 22, -9, -16, 25, -52, 2,
					-- layer=2 filter=172 channel=89
					-16, -57, -59, 26, -9, -29, 3, -23, -23,
					-- layer=2 filter=172 channel=90
					3, 0, -2, 0, -10, 0, 8, 7, 2,
					-- layer=2 filter=172 channel=91
					-24, -16, -17, -17, -43, -27, -80, -54, -34,
					-- layer=2 filter=172 channel=92
					-6, -20, -17, 2, -26, -53, -3, -31, -22,
					-- layer=2 filter=172 channel=93
					17, -3, -20, -16, 2, -23, 40, -23, -52,
					-- layer=2 filter=172 channel=94
					48, 16, 38, 61, 13, -35, 57, 71, -8,
					-- layer=2 filter=172 channel=95
					-14, -12, -9, 1, 3, -8, -15, 8, 0,
					-- layer=2 filter=172 channel=96
					22, -23, -45, 7, -28, -59, 48, -43, -25,
					-- layer=2 filter=172 channel=97
					11, 5, -6, 0, -16, 12, -20, -7, -8,
					-- layer=2 filter=172 channel=98
					17, 44, 12, 48, 35, 17, 45, 21, 29,
					-- layer=2 filter=172 channel=99
					59, 8, 11, 33, 18, 35, 21, 42, -7,
					-- layer=2 filter=172 channel=100
					-18, -26, -35, 6, -34, -1, -33, -5, -10,
					-- layer=2 filter=172 channel=101
					30, 38, 41, -17, -6, 8, -29, -8, 5,
					-- layer=2 filter=172 channel=102
					29, -32, -40, 21, -10, -75, 70, 7, -3,
					-- layer=2 filter=172 channel=103
					-10, -3, -17, -52, -21, 42, -6, -19, 45,
					-- layer=2 filter=172 channel=104
					13, -14, 26, 45, 11, -24, 39, 23, -15,
					-- layer=2 filter=172 channel=105
					-12, 14, -20, 37, 17, 26, -43, 18, 2,
					-- layer=2 filter=172 channel=106
					-32, 2, -2, -34, -6, -20, -48, -9, -14,
					-- layer=2 filter=172 channel=107
					-17, 36, 4, -11, -17, 18, -13, -1, -14,
					-- layer=2 filter=172 channel=108
					-4, -28, 11, 0, 9, -13, 52, 45, 32,
					-- layer=2 filter=172 channel=109
					8, -3, 15, -18, 4, 32, -1, -17, 14,
					-- layer=2 filter=172 channel=110
					20, -8, -19, 74, 5, 0, 50, -25, -28,
					-- layer=2 filter=172 channel=111
					10, 5, 9, -3, -2, -10, -2, 4, 8,
					-- layer=2 filter=172 channel=112
					-2, 23, 1, -11, 30, 10, -6, -7, -3,
					-- layer=2 filter=172 channel=113
					48, 25, -46, 15, 64, -7, 17, 22, -17,
					-- layer=2 filter=172 channel=114
					0, 32, -9, -2, 3, 6, -6, -5, 2,
					-- layer=2 filter=172 channel=115
					-9, -6, -2, 8, -7, 7, -10, 9, -4,
					-- layer=2 filter=172 channel=116
					-24, -19, -93, -22, -70, -118, -15, -82, -77,
					-- layer=2 filter=172 channel=117
					-12, 0, 10, 54, 35, 10, 26, 40, -7,
					-- layer=2 filter=172 channel=118
					-10, 23, 31, 4, 22, 19, -8, 6, 30,
					-- layer=2 filter=172 channel=119
					-11, -23, -4, -8, -15, -22, 16, 22, -19,
					-- layer=2 filter=172 channel=120
					6, 7, 3, -6, -1, 2, 2, 9, -5,
					-- layer=2 filter=172 channel=121
					-2, -7, -7, -9, 8, -4, -1, -10, -7,
					-- layer=2 filter=172 channel=122
					15, 0, 1, 5, 5, 10, -4, 9, 0,
					-- layer=2 filter=172 channel=123
					-13, -24, -15, 14, -12, -36, -6, 13, 12,
					-- layer=2 filter=172 channel=124
					-26, -48, -43, 42, -41, -63, 10, -58, -39,
					-- layer=2 filter=172 channel=125
					-3, -8, 1, 0, 4, 1, -8, 4, 9,
					-- layer=2 filter=172 channel=126
					24, -39, -42, -40, 7, -34, -13, 19, -25,
					-- layer=2 filter=172 channel=127
					14, 0, -27, -11, -4, -19, 35, -2, -10,
					-- layer=2 filter=173 channel=0
					6, -6, -5, -6, -4, 0, 1, 9, 0,
					-- layer=2 filter=173 channel=1
					0, -3, -4, -4, 6, 6, 7, 6, -8,
					-- layer=2 filter=173 channel=2
					-2, 5, -2, 5, 2, 8, -5, -1, -3,
					-- layer=2 filter=173 channel=3
					0, -4, -13, -2, -7, 3, 5, -7, -4,
					-- layer=2 filter=173 channel=4
					-6, -8, 9, -5, -8, -3, 8, -8, -7,
					-- layer=2 filter=173 channel=5
					-2, -10, 3, 0, -9, -6, -10, -2, -12,
					-- layer=2 filter=173 channel=6
					-4, -3, 7, 0, -9, -9, -5, 4, -9,
					-- layer=2 filter=173 channel=7
					-4, -4, -9, 8, -11, -6, -11, -6, 0,
					-- layer=2 filter=173 channel=8
					0, -2, 9, -6, 1, -7, -6, -7, 0,
					-- layer=2 filter=173 channel=9
					-1, 1, -5, -7, -7, -3, 1, -7, -1,
					-- layer=2 filter=173 channel=10
					6, 8, -14, -8, 3, -11, -6, -3, 7,
					-- layer=2 filter=173 channel=11
					-6, 4, -1, -11, 5, -12, -11, -7, -13,
					-- layer=2 filter=173 channel=12
					0, -12, 7, -5, 7, 0, -6, 0, -11,
					-- layer=2 filter=173 channel=13
					-3, -1, 8, -4, -11, 4, 6, -1, 0,
					-- layer=2 filter=173 channel=14
					6, 6, -6, -2, 0, -1, 9, -9, -9,
					-- layer=2 filter=173 channel=15
					2, 0, -2, -2, 5, 1, -1, 1, 6,
					-- layer=2 filter=173 channel=16
					2, 5, 3, 2, 6, -8, 0, -7, -3,
					-- layer=2 filter=173 channel=17
					4, 3, 2, 7, -10, 5, 6, 2, 7,
					-- layer=2 filter=173 channel=18
					-10, 0, 4, -7, 5, 8, 8, 2, -11,
					-- layer=2 filter=173 channel=19
					10, -11, 10, -8, 6, 1, 1, 6, 3,
					-- layer=2 filter=173 channel=20
					-2, 2, -5, 8, 5, 1, -7, 9, -1,
					-- layer=2 filter=173 channel=21
					-5, -4, 5, -8, -7, 9, -2, -6, -9,
					-- layer=2 filter=173 channel=22
					-2, -2, 7, -5, 2, 8, -5, -12, -1,
					-- layer=2 filter=173 channel=23
					-6, -2, 7, 9, 8, 4, 7, 5, -3,
					-- layer=2 filter=173 channel=24
					-12, -11, -6, -8, 2, -8, 0, -5, -7,
					-- layer=2 filter=173 channel=25
					4, -2, 1, 0, -10, -2, -3, 6, -4,
					-- layer=2 filter=173 channel=26
					8, -7, 4, 4, -8, 6, 2, 9, -10,
					-- layer=2 filter=173 channel=27
					-1, -9, 9, 6, 4, -10, -6, -6, 3,
					-- layer=2 filter=173 channel=28
					12, -1, -5, 2, 5, 3, -6, 1, -1,
					-- layer=2 filter=173 channel=29
					-4, -8, 8, 4, -11, -9, -10, -11, -9,
					-- layer=2 filter=173 channel=30
					-9, 5, -12, -3, -9, -2, -6, -5, -10,
					-- layer=2 filter=173 channel=31
					6, -11, 8, 3, 7, 3, -8, 4, -6,
					-- layer=2 filter=173 channel=32
					3, 7, -8, 1, -3, 0, 2, -4, 4,
					-- layer=2 filter=173 channel=33
					5, 7, 3, -6, -11, -8, 6, 4, 3,
					-- layer=2 filter=173 channel=34
					-10, 4, -11, -3, -8, -9, -1, -7, 4,
					-- layer=2 filter=173 channel=35
					-6, -1, 6, -3, -7, -13, -11, -10, 0,
					-- layer=2 filter=173 channel=36
					-8, 2, 2, -3, -2, 1, -5, -4, 9,
					-- layer=2 filter=173 channel=37
					1, -4, 0, -2, -1, 2, 5, -3, -1,
					-- layer=2 filter=173 channel=38
					-11, -5, -11, 6, -11, -6, 5, -4, -3,
					-- layer=2 filter=173 channel=39
					-1, 4, -9, -3, -9, -10, 1, -10, -9,
					-- layer=2 filter=173 channel=40
					-3, -10, -1, -7, -8, 4, -2, -6, 5,
					-- layer=2 filter=173 channel=41
					-6, -9, 2, -8, -9, -5, -2, -9, -1,
					-- layer=2 filter=173 channel=42
					0, -10, -2, -2, 8, -7, 1, -11, 7,
					-- layer=2 filter=173 channel=43
					-2, -8, 5, 8, -4, -2, 5, -5, 3,
					-- layer=2 filter=173 channel=44
					4, -2, -2, -4, 9, -7, 4, -5, 0,
					-- layer=2 filter=173 channel=45
					-1, 7, -1, -6, -4, -2, -8, 5, 5,
					-- layer=2 filter=173 channel=46
					-7, -10, 7, 1, 0, 4, 1, -3, 8,
					-- layer=2 filter=173 channel=47
					-7, 2, 4, 9, 8, -8, -9, -3, -3,
					-- layer=2 filter=173 channel=48
					8, -8, 9, -2, 5, -5, 4, -4, -8,
					-- layer=2 filter=173 channel=49
					-7, -9, -2, -9, 1, -2, 3, -9, 0,
					-- layer=2 filter=173 channel=50
					-4, 0, -4, 4, -2, -2, -3, -4, 2,
					-- layer=2 filter=173 channel=51
					3, -1, -6, 4, -3, -9, -6, -1, -5,
					-- layer=2 filter=173 channel=52
					8, 1, -13, 0, -6, -4, -8, 5, -4,
					-- layer=2 filter=173 channel=53
					-5, -7, -9, -2, -1, 7, 1, 6, -3,
					-- layer=2 filter=173 channel=54
					5, 0, 0, -6, -7, -5, -11, -12, 0,
					-- layer=2 filter=173 channel=55
					-2, 8, 8, -2, -10, 7, -4, -2, 2,
					-- layer=2 filter=173 channel=56
					-8, -7, 5, 0, -3, -10, -9, 8, 4,
					-- layer=2 filter=173 channel=57
					-7, 0, -6, -2, 7, -10, -6, -11, 0,
					-- layer=2 filter=173 channel=58
					1, 2, 6, 8, -9, -7, 8, -10, -12,
					-- layer=2 filter=173 channel=59
					-3, 2, 1, -10, 2, 7, -3, -9, -1,
					-- layer=2 filter=173 channel=60
					0, 0, -2, -9, 4, -3, -7, -4, -5,
					-- layer=2 filter=173 channel=61
					-7, 3, -6, -7, 5, -8, 7, -2, -6,
					-- layer=2 filter=173 channel=62
					-15, -2, 5, -9, -2, 5, 4, -12, 4,
					-- layer=2 filter=173 channel=63
					-3, 4, -9, 9, 3, -4, 2, -5, -4,
					-- layer=2 filter=173 channel=64
					0, -7, -5, -11, -5, -10, 3, -4, -4,
					-- layer=2 filter=173 channel=65
					3, -3, -6, -12, -10, -1, -11, -9, -2,
					-- layer=2 filter=173 channel=66
					-12, -1, 7, 7, -4, 8, 0, 0, -10,
					-- layer=2 filter=173 channel=67
					-10, 7, 1, 7, 7, 0, 4, -6, 0,
					-- layer=2 filter=173 channel=68
					6, 0, -9, 1, 5, 4, 2, 7, 7,
					-- layer=2 filter=173 channel=69
					-6, -3, 7, 0, -10, 1, -9, 3, 3,
					-- layer=2 filter=173 channel=70
					7, 4, 1, -10, 0, -5, 6, 0, 4,
					-- layer=2 filter=173 channel=71
					-6, 0, 8, -4, 7, -10, 0, -9, -9,
					-- layer=2 filter=173 channel=72
					9, 8, -4, 6, -3, 3, -1, -5, -3,
					-- layer=2 filter=173 channel=73
					0, -2, 5, 1, -9, -2, 4, 4, -4,
					-- layer=2 filter=173 channel=74
					-4, -2, 6, 6, -5, 8, -9, -3, -1,
					-- layer=2 filter=173 channel=75
					-9, -11, -5, -12, 8, 5, 7, -10, -4,
					-- layer=2 filter=173 channel=76
					6, -8, -1, -5, 0, 3, 5, -6, -6,
					-- layer=2 filter=173 channel=77
					4, 1, 1, -11, 8, 6, -7, 3, -11,
					-- layer=2 filter=173 channel=78
					8, 0, -11, 6, 0, 3, -5, 6, -5,
					-- layer=2 filter=173 channel=79
					-6, 4, -4, 0, 4, -9, -8, -2, 1,
					-- layer=2 filter=173 channel=80
					2, -6, 5, -6, -2, -2, 6, 1, -3,
					-- layer=2 filter=173 channel=81
					7, 6, 5, -6, 0, 6, 4, -1, -3,
					-- layer=2 filter=173 channel=82
					10, 0, 3, 3, -6, -6, -5, 5, 6,
					-- layer=2 filter=173 channel=83
					-9, -9, -4, -11, -6, -5, -5, 3, 5,
					-- layer=2 filter=173 channel=84
					-10, 5, 2, 3, -8, -1, -6, 8, -1,
					-- layer=2 filter=173 channel=85
					5, 0, -8, 7, -7, 6, 3, 5, -12,
					-- layer=2 filter=173 channel=86
					-10, 7, -7, -5, -7, 5, -2, 8, -8,
					-- layer=2 filter=173 channel=87
					-1, 2, -7, -6, 7, 1, -3, -1, 7,
					-- layer=2 filter=173 channel=88
					-7, 7, -10, -2, 2, -6, -6, 6, 2,
					-- layer=2 filter=173 channel=89
					0, -7, 8, -4, -9, 0, -9, 4, 4,
					-- layer=2 filter=173 channel=90
					6, -9, 1, -10, 0, -10, -6, -9, -1,
					-- layer=2 filter=173 channel=91
					0, -1, 1, 0, -4, 4, -5, 2, 4,
					-- layer=2 filter=173 channel=92
					-4, -4, 2, -9, -2, 8, 10, -3, -2,
					-- layer=2 filter=173 channel=93
					8, -9, 4, -9, -10, 2, -7, -1, 5,
					-- layer=2 filter=173 channel=94
					11, -7, -1, 0, -4, 7, -3, -1, -2,
					-- layer=2 filter=173 channel=95
					-12, -5, 8, -8, -2, 2, -5, -11, -7,
					-- layer=2 filter=173 channel=96
					5, 4, -10, -8, -1, -6, 6, -7, -10,
					-- layer=2 filter=173 channel=97
					5, 2, 6, 7, 7, -2, 2, 5, -12,
					-- layer=2 filter=173 channel=98
					10, -8, 10, 5, -13, -13, -12, 5, 3,
					-- layer=2 filter=173 channel=99
					3, 0, -4, 0, 3, 10, 0, -2, 2,
					-- layer=2 filter=173 channel=100
					-6, 1, -12, -9, 3, 2, -5, -1, 7,
					-- layer=2 filter=173 channel=101
					0, 5, 6, -11, -10, 5, 0, -2, -10,
					-- layer=2 filter=173 channel=102
					-1, 2, 8, 2, 0, -7, -7, 7, -9,
					-- layer=2 filter=173 channel=103
					2, 8, -9, -10, -6, 3, -10, -4, -11,
					-- layer=2 filter=173 channel=104
					-5, 3, -9, -10, -4, -1, 9, -7, 0,
					-- layer=2 filter=173 channel=105
					-5, -9, -12, 8, 6, 2, -2, 6, -2,
					-- layer=2 filter=173 channel=106
					3, -4, 5, -3, -8, 2, 5, -4, -3,
					-- layer=2 filter=173 channel=107
					8, 0, 1, 9, 0, 6, 2, -1, -9,
					-- layer=2 filter=173 channel=108
					-11, -8, 5, 6, 4, 1, -7, 2, -1,
					-- layer=2 filter=173 channel=109
					-7, -3, 0, -4, -8, 4, 4, 7, 2,
					-- layer=2 filter=173 channel=110
					-11, -1, -9, -2, 0, 5, 3, 6, 0,
					-- layer=2 filter=173 channel=111
					-8, -9, 3, -7, 1, 1, 0, -2, -6,
					-- layer=2 filter=173 channel=112
					0, -6, -5, -1, -9, 0, 0, 8, -10,
					-- layer=2 filter=173 channel=113
					-11, -12, 6, 6, 7, -2, -8, -1, 2,
					-- layer=2 filter=173 channel=114
					11, -6, 10, 3, 4, 0, -7, -6, 8,
					-- layer=2 filter=173 channel=115
					0, -5, -10, -1, -6, -10, 0, 9, 2,
					-- layer=2 filter=173 channel=116
					-12, -6, 7, 4, -1, -7, -6, -1, -3,
					-- layer=2 filter=173 channel=117
					-11, -7, 2, -1, -15, -3, -14, -13, 0,
					-- layer=2 filter=173 channel=118
					2, 6, -2, -1, 6, 3, -7, -2, 2,
					-- layer=2 filter=173 channel=119
					-11, -6, 0, -3, 5, 8, -6, -2, 6,
					-- layer=2 filter=173 channel=120
					-8, 5, -5, -7, 4, 6, 3, 7, -10,
					-- layer=2 filter=173 channel=121
					-5, 4, -2, -3, 0, 5, 7, 7, -5,
					-- layer=2 filter=173 channel=122
					-4, 0, -10, 6, 7, 8, -9, -9, 4,
					-- layer=2 filter=173 channel=123
					4, -2, -6, -2, -5, -2, 1, -9, 5,
					-- layer=2 filter=173 channel=124
					6, 5, -1, 1, 7, 5, 2, -9, -4,
					-- layer=2 filter=173 channel=125
					-3, 7, 0, -6, -11, -5, 3, -1, -5,
					-- layer=2 filter=173 channel=126
					-3, 0, -2, -7, 0, 3, -3, -11, 0,
					-- layer=2 filter=173 channel=127
					-10, -9, 5, 1, 0, -10, 9, -1, -6,
					-- layer=2 filter=174 channel=0
					1, 27, -33, -17, 7, -14, 4, -7, -6,
					-- layer=2 filter=174 channel=1
					5, 21, 21, 2, -16, 2, -1, -30, -45,
					-- layer=2 filter=174 channel=2
					3, -1, -8, -1, 0, 2, 0, 5, 6,
					-- layer=2 filter=174 channel=3
					4, -1, 6, 39, 23, 1, 11, -42, -39,
					-- layer=2 filter=174 channel=4
					-48, -31, -20, -44, -12, -13, -10, -15, -27,
					-- layer=2 filter=174 channel=5
					19, 25, 13, -8, 29, -15, -12, -6, -11,
					-- layer=2 filter=174 channel=6
					-95, 16, -26, -62, 14, 6, 5, 23, 31,
					-- layer=2 filter=174 channel=7
					3, 11, -64, 13, 50, 32, 22, 34, 26,
					-- layer=2 filter=174 channel=8
					0, -10, -6, -10, 5, -3, 2, -5, 0,
					-- layer=2 filter=174 channel=9
					53, 34, 36, 19, 34, 17, 14, -43, 15,
					-- layer=2 filter=174 channel=10
					-14, -9, -20, -6, 17, 3, -5, -17, 0,
					-- layer=2 filter=174 channel=11
					-5, 15, -7, 12, 5, -6, 16, 0, -8,
					-- layer=2 filter=174 channel=12
					8, 21, 18, 7, -24, -10, 21, 6, 0,
					-- layer=2 filter=174 channel=13
					-4, -7, 9, 4, 9, 1, -3, 2, 0,
					-- layer=2 filter=174 channel=14
					8, 11, 9, -32, -13, -36, -20, -34, -60,
					-- layer=2 filter=174 channel=15
					-4, 32, 14, 50, -1, 28, 0, -3, 5,
					-- layer=2 filter=174 channel=16
					4, -19, 2, 11, 0, -15, -19, 23, 18,
					-- layer=2 filter=174 channel=17
					0, -8, 1, 0, 2, 1, -2, -4, 0,
					-- layer=2 filter=174 channel=18
					-16, -15, 35, -4, 0, 3, 8, -17, -11,
					-- layer=2 filter=174 channel=19
					-40, -15, -53, 8, 18, 6, 2, 27, 0,
					-- layer=2 filter=174 channel=20
					-10, -10, 5, 5, -8, 2, -13, -11, -4,
					-- layer=2 filter=174 channel=21
					8, -7, 4, 12, 13, 11, 0, -10, -12,
					-- layer=2 filter=174 channel=22
					0, -8, 0, -2, 5, -5, -2, 7, 6,
					-- layer=2 filter=174 channel=23
					-4, 19, -24, 0, 0, -35, 12, 19, 0,
					-- layer=2 filter=174 channel=24
					27, 12, 7, 16, 20, 23, 0, -43, -28,
					-- layer=2 filter=174 channel=25
					-21, -26, -33, 9, -2, -1, -3, -19, -16,
					-- layer=2 filter=174 channel=26
					5, -2, -5, 0, 2, -10, -5, -8, 0,
					-- layer=2 filter=174 channel=27
					3, 16, 4, 31, 29, 0, -4, -14, -10,
					-- layer=2 filter=174 channel=28
					-58, -92, -22, 6, 22, -12, 49, 15, 18,
					-- layer=2 filter=174 channel=29
					-9, 3, 0, -2, -9, -3, -2, 0, -2,
					-- layer=2 filter=174 channel=30
					-3, -21, -14, -19, -89, -8, -49, 3, 4,
					-- layer=2 filter=174 channel=31
					-16, -1, -11, -22, -1, -11, 5, 9, -4,
					-- layer=2 filter=174 channel=32
					-3, -4, 4, 4, 10, 10, -6, -8, 9,
					-- layer=2 filter=174 channel=33
					13, 30, -6, 38, 42, 23, 28, 0, -30,
					-- layer=2 filter=174 channel=34
					-53, -116, 3, -4, 20, 13, 23, 15, 19,
					-- layer=2 filter=174 channel=35
					-43, -60, -51, 5, 16, 16, 51, 29, 16,
					-- layer=2 filter=174 channel=36
					5, 4, -8, 10, -9, -9, 0, -1, 13,
					-- layer=2 filter=174 channel=37
					8, 9, -3, 5, 7, 11, 17, -19, -8,
					-- layer=2 filter=174 channel=38
					-4, 17, -12, 15, -11, -26, -8, -13, -18,
					-- layer=2 filter=174 channel=39
					35, 4, 14, 63, 31, 14, 31, -10, 3,
					-- layer=2 filter=174 channel=40
					-43, -63, -12, 35, -32, 33, 14, -47, 10,
					-- layer=2 filter=174 channel=41
					8, -8, -10, -2, 0, 2, 3, -6, 9,
					-- layer=2 filter=174 channel=42
					42, 19, 7, -13, -44, -4, 21, 12, -1,
					-- layer=2 filter=174 channel=43
					8, -12, 9, 18, 13, 18, 0, -6, -13,
					-- layer=2 filter=174 channel=44
					-9, -1, -5, -6, 1, 0, -8, 3, 1,
					-- layer=2 filter=174 channel=45
					-68, 0, -39, -3, 28, 8, -1, 32, 15,
					-- layer=2 filter=174 channel=46
					-28, -47, -27, 34, -30, 45, -9, -5, -4,
					-- layer=2 filter=174 channel=47
					-29, -34, -45, 15, 20, 10, 45, 9, -2,
					-- layer=2 filter=174 channel=48
					-2, -1, -1, -1, 2, -2, 4, 9, 7,
					-- layer=2 filter=174 channel=49
					-46, -14, 21, 15, 27, 26, -4, -6, 28,
					-- layer=2 filter=174 channel=50
					11, -10, -16, -10, 16, 0, -5, 0, 13,
					-- layer=2 filter=174 channel=51
					3, 3, -14, 5, 18, -24, 16, -5, -6,
					-- layer=2 filter=174 channel=52
					5, 2, 7, -5, -2, 0, 32, -2, -17,
					-- layer=2 filter=174 channel=53
					-9, 38, 49, -62, 18, 16, -9, -7, 27,
					-- layer=2 filter=174 channel=54
					-57, -74, -67, -31, -4, -33, 35, 27, -8,
					-- layer=2 filter=174 channel=55
					5, -2, 5, -8, 0, 10, -2, -3, 0,
					-- layer=2 filter=174 channel=56
					30, 17, 16, 9, 9, 2, 5, -18, -18,
					-- layer=2 filter=174 channel=57
					6, 0, -9, -4, -7, -14, -5, 3, -7,
					-- layer=2 filter=174 channel=58
					-9, -3, -2, -5, -26, -32, 30, 24, 21,
					-- layer=2 filter=174 channel=59
					-25, 42, -42, 25, 24, 0, 32, -36, -66,
					-- layer=2 filter=174 channel=60
					2, 21, -20, -24, 0, 3, -24, 5, -30,
					-- layer=2 filter=174 channel=61
					-29, 11, -42, 3, 34, 23, -57, 27, 2,
					-- layer=2 filter=174 channel=62
					-80, -20, 5, -59, -4, -6, 16, 41, -1,
					-- layer=2 filter=174 channel=63
					16, 10, -17, -4, -37, -27, -12, -47, -47,
					-- layer=2 filter=174 channel=64
					25, -10, -22, 7, -29, -10, 12, -14, -13,
					-- layer=2 filter=174 channel=65
					-24, 26, -12, 13, 0, 29, -55, 14, -1,
					-- layer=2 filter=174 channel=66
					1, 10, -12, -14, 18, 26, -5, -7, -3,
					-- layer=2 filter=174 channel=67
					0, 9, -28, -16, -5, -4, -6, -12, -34,
					-- layer=2 filter=174 channel=68
					-6, 0, -6, -7, -7, -11, -8, 0, -8,
					-- layer=2 filter=174 channel=69
					15, 2, 8, -22, -43, -20, 0, -44, 9,
					-- layer=2 filter=174 channel=70
					-65, -75, -26, -10, 7, -5, 36, 40, 16,
					-- layer=2 filter=174 channel=71
					8, 18, -11, 15, 0, -63, -8, -42, -22,
					-- layer=2 filter=174 channel=72
					49, 49, 3, 19, 0, 24, -39, -26, -45,
					-- layer=2 filter=174 channel=73
					5, -5, -15, 36, 35, 37, 28, 43, 65,
					-- layer=2 filter=174 channel=74
					0, -3, -40, -17, -48, -27, -34, 17, -15,
					-- layer=2 filter=174 channel=75
					-24, -21, -23, -66, -114, -74, -14, 3, -41,
					-- layer=2 filter=174 channel=76
					-34, -2, 2, 24, 57, 9, 36, 42, 73,
					-- layer=2 filter=174 channel=77
					4, 10, 10, 0, 9, 6, -9, -4, 5,
					-- layer=2 filter=174 channel=78
					-43, -9, -7, 10, 20, -9, -1, 8, -16,
					-- layer=2 filter=174 channel=79
					-2, -9, -4, -5, -10, 9, 6, -2, 7,
					-- layer=2 filter=174 channel=80
					-17, -34, -50, 16, 13, -12, 14, -9, -13,
					-- layer=2 filter=174 channel=81
					5, 11, 2, 4, -2, 14, 11, -7, -9,
					-- layer=2 filter=174 channel=82
					4, 13, 5, -6, -10, -1, -6, 7, -5,
					-- layer=2 filter=174 channel=83
					-29, -9, -50, -45, -34, -48, -21, 0, 29,
					-- layer=2 filter=174 channel=84
					6, 0, 7, -5, 0, -10, -9, -4, 5,
					-- layer=2 filter=174 channel=85
					-10, 13, 6, -5, 1, -1, -10, -5, 0,
					-- layer=2 filter=174 channel=86
					0, 17, 3, -5, 15, 12, 4, 6, 3,
					-- layer=2 filter=174 channel=87
					-99, 47, 38, 30, 23, 15, 0, 21, 7,
					-- layer=2 filter=174 channel=88
					12, 3, -19, -8, -41, -49, -31, 2, -5,
					-- layer=2 filter=174 channel=89
					-1, 26, -8, -5, 4, 4, -13, -47, -42,
					-- layer=2 filter=174 channel=90
					6, -7, -5, 0, -5, -4, 5, -9, -6,
					-- layer=2 filter=174 channel=91
					29, 26, 16, -31, -31, -6, 11, 26, -25,
					-- layer=2 filter=174 channel=92
					0, 19, 17, 18, -6, 15, 10, -31, -28,
					-- layer=2 filter=174 channel=93
					-43, -50, -47, 36, 46, -4, 34, 47, -16,
					-- layer=2 filter=174 channel=94
					-45, 35, 46, 2, 27, 29, -15, 8, 17,
					-- layer=2 filter=174 channel=95
					-26, -27, -23, -19, -30, -10, 1, -25, -10,
					-- layer=2 filter=174 channel=96
					-57, 34, -34, -79, 13, -22, 5, 27, 42,
					-- layer=2 filter=174 channel=97
					17, -10, -11, 36, -14, 9, -4, -35, 4,
					-- layer=2 filter=174 channel=98
					-48, -76, -49, 21, 7, 28, 43, 35, 20,
					-- layer=2 filter=174 channel=99
					-33, -8, -42, -14, -13, 34, -11, 25, 0,
					-- layer=2 filter=174 channel=100
					-1, 34, -6, -13, -24, -23, -39, -6, -6,
					-- layer=2 filter=174 channel=101
					-6, -19, -30, 31, 1, -28, -2, -35, -39,
					-- layer=2 filter=174 channel=102
					3, 11, -1, -68, 10, 35, -16, 24, 3,
					-- layer=2 filter=174 channel=103
					-18, 17, 3, 15, 68, -27, 1, 11, 12,
					-- layer=2 filter=174 channel=104
					-49, 43, 34, -1, 19, 1, 9, 29, 20,
					-- layer=2 filter=174 channel=105
					-54, 49, -15, 41, 90, -53, 39, 81, 14,
					-- layer=2 filter=174 channel=106
					1, -15, -27, 13, -6, -30, 9, -31, -56,
					-- layer=2 filter=174 channel=107
					-21, -23, 35, -34, 39, 31, 10, 3, -1,
					-- layer=2 filter=174 channel=108
					20, 52, 12, -17, 14, 3, -52, -29, -3,
					-- layer=2 filter=174 channel=109
					-21, 19, 16, 1, 7, 27, 0, 6, 5,
					-- layer=2 filter=174 channel=110
					25, 6, -13, 0, -35, 9, -34, 2, 1,
					-- layer=2 filter=174 channel=111
					0, -9, 5, -2, 3, 5, 3, -5, 6,
					-- layer=2 filter=174 channel=112
					24, 6, -32, 17, 46, 28, -14, -3, -23,
					-- layer=2 filter=174 channel=113
					17, -5, 21, 14, -66, -14, -31, -7, -7,
					-- layer=2 filter=174 channel=114
					-3, -6, -17, 3, -21, -16, -11, 3, -7,
					-- layer=2 filter=174 channel=115
					2, -6, -7, 5, -13, 1, 0, -2, -3,
					-- layer=2 filter=174 channel=116
					-44, 26, 51, -17, 45, 13, -2, 11, 13,
					-- layer=2 filter=174 channel=117
					-6, -1, -23, -19, 50, 11, 17, 9, 7,
					-- layer=2 filter=174 channel=118
					-23, -20, 11, 23, 34, 33, -11, -8, 8,
					-- layer=2 filter=174 channel=119
					-22, -41, -17, -37, -18, 2, -26, -9, -20,
					-- layer=2 filter=174 channel=120
					0, 0, -3, -4, 3, -5, -1, 3, 1,
					-- layer=2 filter=174 channel=121
					10, 1, -8, 2, -1, 0, 8, 9, 0,
					-- layer=2 filter=174 channel=122
					-12, -7, -12, -6, 1, -2, -6, 3, 5,
					-- layer=2 filter=174 channel=123
					-3, 11, -28, 27, 9, 20, 36, 18, 17,
					-- layer=2 filter=174 channel=124
					-49, 30, -1, 15, 11, -4, -1, 0, -30,
					-- layer=2 filter=174 channel=125
					-5, 10, -10, 2, 0, -3, -15, 3, -5,
					-- layer=2 filter=174 channel=126
					21, 18, -35, 62, 23, 28, -35, -19, 15,
					-- layer=2 filter=174 channel=127
					-3, 8, -2, 4, -6, -46, -24, -16, -57,
					-- layer=2 filter=175 channel=0
					7, 0, -5, 2, -4, -8, -11, 7, -6,
					-- layer=2 filter=175 channel=1
					9, -9, 7, 1, -5, 4, 8, -5, -4,
					-- layer=2 filter=175 channel=2
					4, -1, -9, 7, 7, -8, -5, 12, -9,
					-- layer=2 filter=175 channel=3
					7, 3, -6, -7, 1, -3, 0, -1, -5,
					-- layer=2 filter=175 channel=4
					-1, 4, -10, 3, 4, 2, 4, -12, -12,
					-- layer=2 filter=175 channel=5
					-8, 1, -17, -10, -14, 0, 2, 2, -9,
					-- layer=2 filter=175 channel=6
					-4, -6, 0, -1, 9, -6, -3, -2, -6,
					-- layer=2 filter=175 channel=7
					0, 2, 8, 3, -10, -3, -4, -5, -4,
					-- layer=2 filter=175 channel=8
					-3, 11, -2, 8, 8, 2, 3, 0, -8,
					-- layer=2 filter=175 channel=9
					-3, -4, -11, 4, -9, 2, -11, -1, -12,
					-- layer=2 filter=175 channel=10
					3, -6, -2, 0, 5, -12, 8, 4, 4,
					-- layer=2 filter=175 channel=11
					-8, 3, -3, 1, 3, 1, 0, -2, 0,
					-- layer=2 filter=175 channel=12
					0, 5, -11, 0, 3, 0, 3, 1, 3,
					-- layer=2 filter=175 channel=13
					-1, 12, 1, 10, -2, 5, -6, 8, 10,
					-- layer=2 filter=175 channel=14
					-3, -9, -8, -6, 0, -8, 2, -1, -8,
					-- layer=2 filter=175 channel=15
					-4, 0, 2, 5, -6, -11, 1, -7, 5,
					-- layer=2 filter=175 channel=16
					-1, 3, 6, -10, -3, 7, -8, -10, 0,
					-- layer=2 filter=175 channel=17
					-3, 10, -4, 4, 0, -3, 10, 7, -5,
					-- layer=2 filter=175 channel=18
					2, 3, -3, -4, 1, -2, 4, -5, -6,
					-- layer=2 filter=175 channel=19
					-7, -12, -12, -7, 3, 0, -4, 4, -9,
					-- layer=2 filter=175 channel=20
					1, 8, -8, -5, 2, 0, -3, -4, 10,
					-- layer=2 filter=175 channel=21
					0, 0, -8, 2, 7, 3, 2, 9, -10,
					-- layer=2 filter=175 channel=22
					6, 6, -8, -3, 5, 6, 6, 3, -4,
					-- layer=2 filter=175 channel=23
					-12, 2, 0, 2, -9, 1, -2, -6, 1,
					-- layer=2 filter=175 channel=24
					-7, 6, -9, 1, 3, 0, -3, 4, 7,
					-- layer=2 filter=175 channel=25
					-11, -3, -12, -11, -3, -10, -18, -3, -6,
					-- layer=2 filter=175 channel=26
					-2, 1, 0, 5, -10, -7, -4, 3, -5,
					-- layer=2 filter=175 channel=27
					7, -5, 4, 0, -4, 2, -6, -1, -3,
					-- layer=2 filter=175 channel=28
					-1, -3, 7, 7, -7, -14, -3, -11, 3,
					-- layer=2 filter=175 channel=29
					-7, -6, -7, 0, 7, -2, 0, 2, -3,
					-- layer=2 filter=175 channel=30
					-8, -6, 0, -5, 0, -5, 1, -3, 4,
					-- layer=2 filter=175 channel=31
					1, -9, 0, -2, -7, 6, -2, 8, 5,
					-- layer=2 filter=175 channel=32
					7, -5, -4, -2, -5, 0, 0, 3, 2,
					-- layer=2 filter=175 channel=33
					-4, -1, -14, 2, -11, -3, 5, -3, -4,
					-- layer=2 filter=175 channel=34
					-14, 1, -11, -8, -3, 0, -7, -2, 3,
					-- layer=2 filter=175 channel=35
					3, -3, -12, -6, 9, -5, -6, 0, -11,
					-- layer=2 filter=175 channel=36
					-1, 4, 5, 5, 2, 2, 0, 0, -4,
					-- layer=2 filter=175 channel=37
					-1, -9, -4, -3, -12, -13, 3, -12, -11,
					-- layer=2 filter=175 channel=38
					11, -11, -5, -6, -2, -4, -14, 8, -10,
					-- layer=2 filter=175 channel=39
					-2, 0, 6, 0, 5, -2, -1, 0, -3,
					-- layer=2 filter=175 channel=40
					2, 6, 6, -14, 11, -2, 1, -5, -3,
					-- layer=2 filter=175 channel=41
					11, 2, 2, 0, 0, -7, -3, 9, -9,
					-- layer=2 filter=175 channel=42
					-5, -7, -3, -12, 2, -5, -5, -1, 0,
					-- layer=2 filter=175 channel=43
					-12, -9, -9, -8, 3, -12, -7, 2, -2,
					-- layer=2 filter=175 channel=44
					9, 2, -5, 5, -5, -2, 5, 8, -9,
					-- layer=2 filter=175 channel=45
					7, -7, 0, 0, -4, 0, 1, 10, -2,
					-- layer=2 filter=175 channel=46
					-9, -8, 4, -3, -5, -10, -7, 2, 8,
					-- layer=2 filter=175 channel=47
					-5, 3, -4, -11, -9, -3, -7, 3, -4,
					-- layer=2 filter=175 channel=48
					-8, 4, 4, 0, -11, -5, -3, 9, 1,
					-- layer=2 filter=175 channel=49
					-6, -11, 8, 2, -15, -16, -2, -4, -11,
					-- layer=2 filter=175 channel=50
					10, 0, -3, 8, -3, 7, -6, 6, 5,
					-- layer=2 filter=175 channel=51
					-7, -8, -1, 2, 0, -16, -10, -11, -17,
					-- layer=2 filter=175 channel=52
					2, 0, -3, -10, 2, -7, -4, 6, -3,
					-- layer=2 filter=175 channel=53
					8, 4, 1, 5, 8, 3, -4, 4, -16,
					-- layer=2 filter=175 channel=54
					-5, -2, -10, 0, 4, -5, -8, 5, -19,
					-- layer=2 filter=175 channel=55
					-6, 9, 6, 4, -7, -5, 5, -4, 2,
					-- layer=2 filter=175 channel=56
					-13, -6, -5, 6, -8, -8, -9, 4, 6,
					-- layer=2 filter=175 channel=57
					3, 3, 10, -10, 0, 3, 6, 4, 9,
					-- layer=2 filter=175 channel=58
					7, -11, 6, 6, 0, -12, 3, -1, 6,
					-- layer=2 filter=175 channel=59
					-11, -11, 0, 5, 1, -2, -8, -9, 6,
					-- layer=2 filter=175 channel=60
					-6, -14, 7, -9, -14, 6, -13, -4, -10,
					-- layer=2 filter=175 channel=61
					-14, -5, -7, -2, -3, -3, 3, -2, -15,
					-- layer=2 filter=175 channel=62
					-12, -6, 1, -2, -4, -7, -12, -4, -2,
					-- layer=2 filter=175 channel=63
					-4, -2, -9, -2, 5, 3, -3, 7, 0,
					-- layer=2 filter=175 channel=64
					-1, -9, -10, 6, -9, -7, 6, -5, 6,
					-- layer=2 filter=175 channel=65
					6, -11, 8, 1, -4, 7, -11, 0, -6,
					-- layer=2 filter=175 channel=66
					1, -5, -1, 6, -10, 7, 8, -1, 5,
					-- layer=2 filter=175 channel=67
					1, 4, -7, -8, 1, -5, -2, -6, 6,
					-- layer=2 filter=175 channel=68
					-2, -8, 9, 5, -8, -11, -10, 5, -1,
					-- layer=2 filter=175 channel=69
					5, 8, -4, -11, -3, 4, 2, -9, -11,
					-- layer=2 filter=175 channel=70
					-8, -11, 8, -7, -2, 1, -7, 2, 5,
					-- layer=2 filter=175 channel=71
					-15, 0, -11, -17, 3, -5, 0, -8, -7,
					-- layer=2 filter=175 channel=72
					1, -11, -7, -4, -7, -12, -1, -5, -12,
					-- layer=2 filter=175 channel=73
					-6, 0, 0, 0, -7, -11, 9, -13, 5,
					-- layer=2 filter=175 channel=74
					-7, 2, -2, 0, -1, 6, -5, -8, -9,
					-- layer=2 filter=175 channel=75
					-11, -1, 4, -10, -9, -3, -7, 7, 0,
					-- layer=2 filter=175 channel=76
					-4, 8, -8, -7, -8, -1, -4, 3, 7,
					-- layer=2 filter=175 channel=77
					10, 10, 2, 6, -4, -9, -7, 4, -5,
					-- layer=2 filter=175 channel=78
					-2, -2, -14, 0, -13, -13, 1, 6, -12,
					-- layer=2 filter=175 channel=79
					3, 9, 0, -7, 10, 3, 1, 3, 8,
					-- layer=2 filter=175 channel=80
					-6, 1, 5, 1, -4, -8, -6, -9, 0,
					-- layer=2 filter=175 channel=81
					-6, 2, -10, 1, -9, -7, 7, 2, -2,
					-- layer=2 filter=175 channel=82
					0, -9, -4, 9, 0, -6, -10, 0, -3,
					-- layer=2 filter=175 channel=83
					-11, -6, -3, 6, -9, 0, 8, 1, 0,
					-- layer=2 filter=175 channel=84
					1, 12, -5, 0, -9, 1, 10, 5, -4,
					-- layer=2 filter=175 channel=85
					5, -2, -1, 1, 7, 0, 6, -7, 4,
					-- layer=2 filter=175 channel=86
					-6, 8, -5, -2, -4, -7, -6, -6, 0,
					-- layer=2 filter=175 channel=87
					-3, 0, -1, -4, 1, -7, -8, -2, -10,
					-- layer=2 filter=175 channel=88
					6, 7, 8, -2, -11, -9, -5, 8, 8,
					-- layer=2 filter=175 channel=89
					-11, 3, -13, -4, -5, 7, -7, 0, 0,
					-- layer=2 filter=175 channel=90
					-5, -2, -1, -2, 7, 5, -1, 6, -9,
					-- layer=2 filter=175 channel=91
					3, 4, 1, 0, -3, -7, 5, 4, 4,
					-- layer=2 filter=175 channel=92
					0, -1, -2, -8, -4, -9, -7, -11, -8,
					-- layer=2 filter=175 channel=93
					-14, -5, -5, -2, -8, 9, 5, 3, -7,
					-- layer=2 filter=175 channel=94
					0, 0, -16, 3, 0, -9, -14, -1, -16,
					-- layer=2 filter=175 channel=95
					-2, 7, -4, -4, -8, 1, -10, -11, 0,
					-- layer=2 filter=175 channel=96
					-7, 4, -11, 0, 5, -2, -8, -20, 0,
					-- layer=2 filter=175 channel=97
					5, 8, 8, 3, 4, 3, 0, -6, -11,
					-- layer=2 filter=175 channel=98
					-1, -12, 1, -13, -1, -13, 1, -6, 5,
					-- layer=2 filter=175 channel=99
					-16, -5, 0, 1, -2, -3, -10, 4, 1,
					-- layer=2 filter=175 channel=100
					-11, 4, -5, 0, 0, 4, 3, -11, -6,
					-- layer=2 filter=175 channel=101
					-13, -10, 1, -15, 0, -2, -17, 0, -20,
					-- layer=2 filter=175 channel=102
					10, 3, -1, -5, -7, -10, 5, -3, -11,
					-- layer=2 filter=175 channel=103
					-4, 2, 3, 2, 8, -6, -5, 4, -10,
					-- layer=2 filter=175 channel=104
					-7, -7, -10, 3, 8, 0, -5, 2, -1,
					-- layer=2 filter=175 channel=105
					-12, -8, 2, 8, 4, 0, 3, -6, 3,
					-- layer=2 filter=175 channel=106
					7, -5, -14, -8, 0, -9, -2, -7, -12,
					-- layer=2 filter=175 channel=107
					-1, 3, 11, 6, -8, 0, 0, -9, -10,
					-- layer=2 filter=175 channel=108
					-11, 0, -9, 1, -2, -4, 3, 7, -2,
					-- layer=2 filter=175 channel=109
					-7, 2, -2, -3, -5, 8, 9, 6, 6,
					-- layer=2 filter=175 channel=110
					-1, 6, 2, -13, -9, -3, 1, -1, -3,
					-- layer=2 filter=175 channel=111
					-6, -10, 8, -7, 3, 0, 7, 2, -4,
					-- layer=2 filter=175 channel=112
					2, -8, -6, 0, -8, 8, -10, -10, 0,
					-- layer=2 filter=175 channel=113
					-12, -10, -8, -8, 8, 3, 0, 1, -8,
					-- layer=2 filter=175 channel=114
					-9, 3, 1, 2, 5, 0, 3, -2, -6,
					-- layer=2 filter=175 channel=115
					7, -4, 7, -3, 8, 1, 6, 4, 8,
					-- layer=2 filter=175 channel=116
					0, -6, 0, -9, -12, -1, -13, -12, -12,
					-- layer=2 filter=175 channel=117
					-2, -13, 5, 3, -8, -8, 1, -2, -15,
					-- layer=2 filter=175 channel=118
					0, 5, 3, 4, -4, -9, 2, 2, -11,
					-- layer=2 filter=175 channel=119
					-2, -4, 1, 1, 2, -13, -5, 2, -7,
					-- layer=2 filter=175 channel=120
					-5, 7, -5, 0, -7, 6, -1, 1, -2,
					-- layer=2 filter=175 channel=121
					-7, -8, -8, -2, 8, -1, -4, 10, 10,
					-- layer=2 filter=175 channel=122
					-2, 8, -6, -2, -9, 4, -7, -5, 8,
					-- layer=2 filter=175 channel=123
					2, -5, -9, -5, -5, -9, 0, -10, -8,
					-- layer=2 filter=175 channel=124
					10, -7, 3, -10, 2, -5, 1, 0, 6,
					-- layer=2 filter=175 channel=125
					-6, -6, -8, 1, 8, -4, 2, 7, -10,
					-- layer=2 filter=175 channel=126
					-6, -1, 6, 0, -9, -3, 7, -5, 8,
					-- layer=2 filter=175 channel=127
					6, -7, -3, -11, 0, 0, -10, -11, -3,
					-- layer=2 filter=176 channel=0
					11, 5, -32, -35, 5, 20, -28, -22, -9,
					-- layer=2 filter=176 channel=1
					-5, -7, 13, -21, -20, 3, 13, 16, 16,
					-- layer=2 filter=176 channel=2
					-3, -8, 0, 7, -6, -3, 6, -2, -9,
					-- layer=2 filter=176 channel=3
					-26, 5, -10, -2, -7, -10, -41, -11, -4,
					-- layer=2 filter=176 channel=4
					-9, -8, 31, -21, -11, 26, 11, 20, -37,
					-- layer=2 filter=176 channel=5
					-12, -11, -21, -44, 3, 24, -26, -17, -4,
					-- layer=2 filter=176 channel=6
					16, -12, -23, 14, -15, -10, -14, 27, 29,
					-- layer=2 filter=176 channel=7
					11, 40, 0, 2, -2, 6, 2, 5, -6,
					-- layer=2 filter=176 channel=8
					-8, -2, 0, -9, 3, 2, 1, 4, -10,
					-- layer=2 filter=176 channel=9
					-12, -10, 6, -20, -11, -8, 7, 4, -16,
					-- layer=2 filter=176 channel=10
					15, -18, -10, -4, 19, 14, -2, -10, -2,
					-- layer=2 filter=176 channel=11
					-7, -12, -2, -11, -39, -11, -27, -25, 4,
					-- layer=2 filter=176 channel=12
					11, 1, 8, 8, -29, -3, 0, 20, 11,
					-- layer=2 filter=176 channel=13
					3, 5, 9, 0, -9, 0, 5, 4, 3,
					-- layer=2 filter=176 channel=14
					-12, -17, -9, -27, -19, -14, -3, 4, 8,
					-- layer=2 filter=176 channel=15
					-20, 3, 6, -3, -4, -17, -39, -23, -18,
					-- layer=2 filter=176 channel=16
					-1, 15, 10, 17, 9, 7, 12, -16, -28,
					-- layer=2 filter=176 channel=17
					10, 3, -7, 4, -8, 5, -2, -4, 10,
					-- layer=2 filter=176 channel=18
					-22, -3, 26, -32, 13, -6, -4, -24, -15,
					-- layer=2 filter=176 channel=19
					2, -13, -14, -18, -36, 15, -34, -15, 16,
					-- layer=2 filter=176 channel=20
					-5, 1, -5, -1, -9, 6, -7, 0, 4,
					-- layer=2 filter=176 channel=21
					-3, -11, -6, 8, -11, -4, 1, -6, -1,
					-- layer=2 filter=176 channel=22
					-2, 8, 11, -11, 1, 1, 7, -3, -5,
					-- layer=2 filter=176 channel=23
					10, 2, 8, -1, 25, 6, 14, -9, -29,
					-- layer=2 filter=176 channel=24
					-13, -4, -36, -23, -35, -35, -25, -40, -41,
					-- layer=2 filter=176 channel=25
					-16, -4, -37, -44, -46, -22, -37, -30, -10,
					-- layer=2 filter=176 channel=26
					-5, 5, 1, 4, 6, 6, 8, -2, 1,
					-- layer=2 filter=176 channel=27
					-15, 8, -9, -31, -25, -3, -16, -25, -3,
					-- layer=2 filter=176 channel=28
					-11, 0, -15, -3, 12, 19, -1, -31, -5,
					-- layer=2 filter=176 channel=29
					0, 1, 1, -12, 0, 7, 3, -5, -8,
					-- layer=2 filter=176 channel=30
					-2, -28, -12, 15, 21, -9, 22, 18, -19,
					-- layer=2 filter=176 channel=31
					-14, 49, 40, -9, 11, -3, 2, 0, 20,
					-- layer=2 filter=176 channel=32
					4, -7, 5, -4, -3, -7, -11, -5, 5,
					-- layer=2 filter=176 channel=33
					-27, 4, -8, -1, 2, -23, -4, 9, 6,
					-- layer=2 filter=176 channel=34
					-31, -10, 9, -16, 18, 15, -3, -30, 23,
					-- layer=2 filter=176 channel=35
					11, 1, -16, 1, 34, 6, 5, -15, -16,
					-- layer=2 filter=176 channel=36
					4, -8, -7, -7, -11, -9, 7, -2, -2,
					-- layer=2 filter=176 channel=37
					-29, -28, 5, -16, -38, 2, -23, -8, 2,
					-- layer=2 filter=176 channel=38
					9, -24, -22, -30, -25, -16, -7, 18, -8,
					-- layer=2 filter=176 channel=39
					5, 14, -14, 17, 0, -28, 5, 3, -16,
					-- layer=2 filter=176 channel=40
					-23, -26, 6, -3, -11, -17, -27, -15, 6,
					-- layer=2 filter=176 channel=41
					-2, -1, 1, 2, -7, 7, -6, 0, 1,
					-- layer=2 filter=176 channel=42
					4, 13, 6, 27, 5, 10, 14, 1, 15,
					-- layer=2 filter=176 channel=43
					-30, -9, -18, -26, 22, -26, 3, -37, -24,
					-- layer=2 filter=176 channel=44
					7, 6, -4, -6, -10, -6, -3, 2, -8,
					-- layer=2 filter=176 channel=45
					-17, 4, -35, -4, -8, -25, 10, 5, 0,
					-- layer=2 filter=176 channel=46
					-12, -18, -14, 11, 16, -6, 13, 10, 24,
					-- layer=2 filter=176 channel=47
					-5, -3, 0, -25, -20, 1, 17, 9, 22,
					-- layer=2 filter=176 channel=48
					8, -9, -2, 0, -5, 3, 7, 4, -2,
					-- layer=2 filter=176 channel=49
					-16, -11, 34, -20, -4, -1, 3, 0, -9,
					-- layer=2 filter=176 channel=50
					-8, 7, -5, 0, 0, 7, -7, -8, -1,
					-- layer=2 filter=176 channel=51
					0, -6, 2, -11, -18, -9, -10, -24, 2,
					-- layer=2 filter=176 channel=52
					-44, -3, 9, -3, -35, -10, -9, -31, 12,
					-- layer=2 filter=176 channel=53
					2, 8, 34, -31, -30, 7, -21, -7, 3,
					-- layer=2 filter=176 channel=54
					10, 0, -1, -11, 10, 14, 0, 10, 3,
					-- layer=2 filter=176 channel=55
					1, 1, -6, 2, -11, -5, -2, 8, -6,
					-- layer=2 filter=176 channel=56
					-22, -16, -19, -13, 1, 12, -14, -29, 0,
					-- layer=2 filter=176 channel=57
					1, -7, 4, -11, 0, -2, 2, 6, -5,
					-- layer=2 filter=176 channel=58
					28, 2, -23, 4, -20, -10, -12, 18, -3,
					-- layer=2 filter=176 channel=59
					27, 7, -17, 3, -10, -27, -3, 21, -9,
					-- layer=2 filter=176 channel=60
					27, 2, -30, -20, -18, 4, 0, 13, -5,
					-- layer=2 filter=176 channel=61
					48, 22, -34, -20, 24, 15, -21, -13, 20,
					-- layer=2 filter=176 channel=62
					7, -6, -12, 43, -11, -2, -18, 6, 39,
					-- layer=2 filter=176 channel=63
					33, 14, -19, 5, 2, 10, 13, -7, 11,
					-- layer=2 filter=176 channel=64
					0, -8, -1, 10, -4, -20, 13, 6, -6,
					-- layer=2 filter=176 channel=65
					31, -15, -21, 18, -3, -18, -20, 12, 13,
					-- layer=2 filter=176 channel=66
					-6, 37, -4, 30, -3, 0, 6, 0, 28,
					-- layer=2 filter=176 channel=67
					-17, -20, -21, -21, -16, -16, -18, 7, -27,
					-- layer=2 filter=176 channel=68
					-4, -5, -9, 4, 5, 8, 0, -3, 5,
					-- layer=2 filter=176 channel=69
					0, -1, 17, -5, -1, -4, 0, 13, 8,
					-- layer=2 filter=176 channel=70
					-9, -16, -10, -10, 34, -5, -8, 0, -25,
					-- layer=2 filter=176 channel=71
					-11, -11, -19, -28, -10, -2, -37, -15, -5,
					-- layer=2 filter=176 channel=72
					-24, -24, -15, -10, -25, -12, -29, -13, -24,
					-- layer=2 filter=176 channel=73
					-20, 33, 1, -7, -2, -23, -10, 17, -1,
					-- layer=2 filter=176 channel=74
					-3, -33, -6, 0, -14, -7, 0, 15, -3,
					-- layer=2 filter=176 channel=75
					-14, -23, -19, -16, -12, -1, -11, -28, 24,
					-- layer=2 filter=176 channel=76
					21, 51, 37, -27, -20, -15, -10, 12, -9,
					-- layer=2 filter=176 channel=77
					-3, -3, 7, 0, 0, 5, 0, -5, 2,
					-- layer=2 filter=176 channel=78
					-43, -13, 0, -24, -53, -26, -7, -13, 0,
					-- layer=2 filter=176 channel=79
					-1, -7, -4, 4, -7, -1, 4, 6, 3,
					-- layer=2 filter=176 channel=80
					-17, -18, -8, 6, -7, -3, 10, -2, -23,
					-- layer=2 filter=176 channel=81
					-8, -7, 0, 8, -2, -9, -9, 8, -7,
					-- layer=2 filter=176 channel=82
					-6, 2, 5, 3, 8, -3, 3, 7, 0,
					-- layer=2 filter=176 channel=83
					13, -17, 1, 8, 15, 19, -6, 0, -16,
					-- layer=2 filter=176 channel=84
					2, -11, 0, -6, -7, -6, -7, -3, -2,
					-- layer=2 filter=176 channel=85
					10, -3, -10, -12, 9, -6, -7, 5, 8,
					-- layer=2 filter=176 channel=86
					-5, 0, -7, 5, 4, -8, -7, -8, 7,
					-- layer=2 filter=176 channel=87
					-22, 0, 12, 16, -18, -12, -6, -56, -9,
					-- layer=2 filter=176 channel=88
					4, -17, 0, -7, -9, -21, 14, 14, 6,
					-- layer=2 filter=176 channel=89
					-6, -33, -17, -37, -18, -3, -21, -3, 10,
					-- layer=2 filter=176 channel=90
					-5, 9, -1, -4, 10, -3, -8, 0, 8,
					-- layer=2 filter=176 channel=91
					0, -5, -13, 1, -19, 0, -12, -9, -1,
					-- layer=2 filter=176 channel=92
					16, -10, -14, 0, -37, 3, -13, 7, -8,
					-- layer=2 filter=176 channel=93
					-2, -22, 0, 37, 0, -18, 7, 16, 42,
					-- layer=2 filter=176 channel=94
					44, 32, -15, -5, -19, 25, -2, -9, 24,
					-- layer=2 filter=176 channel=95
					3, 7, 8, 0, 6, 6, -1, 0, -5,
					-- layer=2 filter=176 channel=96
					6, -5, 11, -26, -12, -1, 6, -2, -36,
					-- layer=2 filter=176 channel=97
					-28, 0, -5, -8, -20, -17, -5, 12, 7,
					-- layer=2 filter=176 channel=98
					17, 19, -38, -32, -1, -4, -19, -27, -7,
					-- layer=2 filter=176 channel=99
					-15, -6, -3, -39, -40, -15, -27, -21, -13,
					-- layer=2 filter=176 channel=100
					-9, -19, -23, -14, -10, -11, -10, -11, -16,
					-- layer=2 filter=176 channel=101
					-23, -13, -21, -29, -29, -26, -11, -22, -33,
					-- layer=2 filter=176 channel=102
					-24, -12, 37, -43, 3, -11, -11, -23, -47,
					-- layer=2 filter=176 channel=103
					6, 8, -11, 14, -18, 30, 26, 23, 7,
					-- layer=2 filter=176 channel=104
					5, 5, 23, -16, -20, 32, 0, -4, -1,
					-- layer=2 filter=176 channel=105
					17, 35, 17, -34, 10, -29, 11, -26, -12,
					-- layer=2 filter=176 channel=106
					-19, 6, -22, -47, -40, -40, -16, -3, -42,
					-- layer=2 filter=176 channel=107
					-11, 1, 0, 1, 3, 38, 6, 73, 0,
					-- layer=2 filter=176 channel=108
					-40, -37, -3, -25, -35, -16, -21, -22, -13,
					-- layer=2 filter=176 channel=109
					8, 1, 1, -6, -4, -6, 0, -4, 2,
					-- layer=2 filter=176 channel=110
					14, 8, -29, 24, 15, -15, -3, -9, -9,
					-- layer=2 filter=176 channel=111
					-1, -5, 2, -5, -11, -11, 7, -8, -2,
					-- layer=2 filter=176 channel=112
					39, 3, -35, -33, 0, 0, -25, -10, 20,
					-- layer=2 filter=176 channel=113
					35, -5, -3, 12, 41, 18, 7, 3, 14,
					-- layer=2 filter=176 channel=114
					-5, -7, 0, 8, 2, -6, -8, 2, -6,
					-- layer=2 filter=176 channel=115
					-7, 9, 5, 6, -4, 7, 9, -7, 3,
					-- layer=2 filter=176 channel=116
					-10, -4, 18, -12, -8, -2, -21, -41, -7,
					-- layer=2 filter=176 channel=117
					-14, 15, 10, -19, -23, 8, -9, 11, -12,
					-- layer=2 filter=176 channel=118
					-38, -6, 10, 2, -13, -8, -2, -17, -34,
					-- layer=2 filter=176 channel=119
					-20, -1, 14, -32, -4, -5, -14, 1, -10,
					-- layer=2 filter=176 channel=120
					-5, 2, 6, -4, 6, 0, 8, 0, -8,
					-- layer=2 filter=176 channel=121
					-8, -10, -8, -8, -2, 9, 3, -6, 3,
					-- layer=2 filter=176 channel=122
					-6, 8, 0, 8, 2, 6, 3, -2, 5,
					-- layer=2 filter=176 channel=123
					21, 11, -11, -4, -1, -17, 4, -13, 7,
					-- layer=2 filter=176 channel=124
					-2, 13, 20, 2, -10, -12, -14, 15, 7,
					-- layer=2 filter=176 channel=125
					0, 8, 3, 7, 0, 9, -8, -1, 8,
					-- layer=2 filter=176 channel=126
					18, 15, -16, -22, -4, 2, 20, -6, -8,
					-- layer=2 filter=176 channel=127
					-6, -15, 0, 10, 15, -14, 1, 21, -8,
					-- layer=2 filter=177 channel=0
					-4, -13, 2, -4, 0, 3, 2, -7, 2,
					-- layer=2 filter=177 channel=1
					2, -4, 5, -16, -19, -7, -9, -6, -11,
					-- layer=2 filter=177 channel=2
					-8, 4, -9, -10, 0, -7, -7, 3, 8,
					-- layer=2 filter=177 channel=3
					-12, -8, -10, -1, 2, -6, -16, -1, -13,
					-- layer=2 filter=177 channel=4
					-3, -3, -14, -1, 0, 3, 1, 2, -7,
					-- layer=2 filter=177 channel=5
					-10, -22, -1, -16, 0, 0, -19, -13, -12,
					-- layer=2 filter=177 channel=6
					3, -4, -10, 3, -4, 10, -6, -4, -2,
					-- layer=2 filter=177 channel=7
					-7, -10, -9, -5, -21, -10, -19, -9, -7,
					-- layer=2 filter=177 channel=8
					2, 0, -5, -8, 8, 0, 8, 6, 3,
					-- layer=2 filter=177 channel=9
					-6, -7, 0, -6, -4, -9, 3, 7, -11,
					-- layer=2 filter=177 channel=10
					-4, -10, -12, -13, -10, -15, -3, -11, -2,
					-- layer=2 filter=177 channel=11
					-13, 0, -7, -16, -1, -12, -14, -8, -5,
					-- layer=2 filter=177 channel=12
					-10, -13, -8, -3, -13, 7, -7, -16, 4,
					-- layer=2 filter=177 channel=13
					3, 4, -10, 0, -9, 0, -10, -7, -8,
					-- layer=2 filter=177 channel=14
					5, -6, -11, -6, 3, -1, -6, 3, -3,
					-- layer=2 filter=177 channel=15
					-11, 6, -7, 7, -13, -5, 3, -1, 6,
					-- layer=2 filter=177 channel=16
					9, 8, -8, 6, 1, 0, -5, -2, -12,
					-- layer=2 filter=177 channel=17
					2, -8, 1, 8, 5, -7, 0, 8, 1,
					-- layer=2 filter=177 channel=18
					-18, -14, 0, -13, -6, -6, -1, 1, 2,
					-- layer=2 filter=177 channel=19
					-15, -2, 3, 0, -19, -11, -15, 2, 0,
					-- layer=2 filter=177 channel=20
					-2, -12, 6, -4, -11, -9, 0, 6, 5,
					-- layer=2 filter=177 channel=21
					0, 9, -7, 0, -6, 0, 9, 5, 0,
					-- layer=2 filter=177 channel=22
					5, -8, -2, 8, 0, -6, 5, -6, 1,
					-- layer=2 filter=177 channel=23
					-4, -11, -13, 0, -13, -2, -8, -17, 1,
					-- layer=2 filter=177 channel=24
					-3, 7, 1, -10, -9, 3, -3, -10, -9,
					-- layer=2 filter=177 channel=25
					-11, 1, -3, -16, -3, -5, -9, -9, 9,
					-- layer=2 filter=177 channel=26
					-9, -8, 0, -4, -9, -7, -5, 9, -9,
					-- layer=2 filter=177 channel=27
					-11, -13, -3, -3, -14, -3, -16, -8, -9,
					-- layer=2 filter=177 channel=28
					-6, -10, -12, 1, -18, -15, -7, -4, -2,
					-- layer=2 filter=177 channel=29
					0, -6, -3, -4, 3, 6, -10, 0, 6,
					-- layer=2 filter=177 channel=30
					8, 4, -1, 4, 4, -13, -13, 2, 3,
					-- layer=2 filter=177 channel=31
					-9, -4, -16, 1, -8, -1, 2, -6, 5,
					-- layer=2 filter=177 channel=32
					-8, -6, -5, 4, -4, 3, 7, 6, 0,
					-- layer=2 filter=177 channel=33
					5, -1, 5, 5, -13, -3, -8, 4, 5,
					-- layer=2 filter=177 channel=34
					-1, 1, -11, -6, 0, -13, -14, -13, -10,
					-- layer=2 filter=177 channel=35
					-2, -17, -4, -12, 3, -2, -10, -12, -18,
					-- layer=2 filter=177 channel=36
					7, -3, -4, 8, -9, 5, 8, -9, 8,
					-- layer=2 filter=177 channel=37
					-15, -14, -6, -6, -13, 1, -20, -7, -13,
					-- layer=2 filter=177 channel=38
					-9, -17, -5, -15, -10, -8, -8, 2, -5,
					-- layer=2 filter=177 channel=39
					-8, 0, 7, -6, 0, 0, 2, -12, 4,
					-- layer=2 filter=177 channel=40
					6, -8, 0, -10, 3, -2, 10, -12, 6,
					-- layer=2 filter=177 channel=41
					-2, -3, 0, -12, -1, 11, -10, 4, 5,
					-- layer=2 filter=177 channel=42
					-6, 4, 2, -4, -12, -9, 4, -1, 6,
					-- layer=2 filter=177 channel=43
					-15, -12, -8, -12, -9, -10, -8, -5, -7,
					-- layer=2 filter=177 channel=44
					-2, -6, 8, 1, 7, -2, 4, 3, 0,
					-- layer=2 filter=177 channel=45
					-2, -7, 0, 4, -12, -8, -4, 8, -11,
					-- layer=2 filter=177 channel=46
					-9, -10, -1, 2, -2, 0, -8, -6, -6,
					-- layer=2 filter=177 channel=47
					-15, -8, 0, -9, -5, -7, -10, -15, -4,
					-- layer=2 filter=177 channel=48
					9, -3, -4, 4, 6, 4, -9, 2, 0,
					-- layer=2 filter=177 channel=49
					3, 4, -9, 5, 0, 5, 7, 5, 3,
					-- layer=2 filter=177 channel=50
					-4, -11, 0, -3, -1, -4, -2, 4, 0,
					-- layer=2 filter=177 channel=51
					-12, -3, -2, -11, -14, -2, -5, -8, -11,
					-- layer=2 filter=177 channel=52
					-11, -12, -8, -16, -16, -17, -19, -17, -10,
					-- layer=2 filter=177 channel=53
					4, -12, -8, -11, -6, -2, -6, -14, -7,
					-- layer=2 filter=177 channel=54
					-3, -5, 1, -1, -8, -3, -3, -14, -3,
					-- layer=2 filter=177 channel=55
					1, -4, 9, 8, -5, -5, 5, 6, 0,
					-- layer=2 filter=177 channel=56
					-18, -7, -17, 5, -4, -5, -5, -1, -17,
					-- layer=2 filter=177 channel=57
					-2, 8, -9, 0, -5, -5, -6, -3, -5,
					-- layer=2 filter=177 channel=58
					-15, -3, -17, -16, -7, -11, -15, -16, -13,
					-- layer=2 filter=177 channel=59
					-7, -12, -15, -19, -5, -12, -5, -8, 0,
					-- layer=2 filter=177 channel=60
					-17, -4, -19, -8, -18, -7, 3, -10, -14,
					-- layer=2 filter=177 channel=61
					-15, 4, -1, -16, -5, -1, -14, -8, 2,
					-- layer=2 filter=177 channel=62
					-10, -7, 0, -2, -7, 3, -6, -10, 1,
					-- layer=2 filter=177 channel=63
					-14, 3, -12, -5, -3, -11, -9, 0, -17,
					-- layer=2 filter=177 channel=64
					-4, 0, -11, -12, 4, -8, 0, 5, 5,
					-- layer=2 filter=177 channel=65
					-11, -11, 4, 5, -8, -4, -9, 0, 9,
					-- layer=2 filter=177 channel=66
					8, -1, 7, 2, 1, 8, -10, -9, 11,
					-- layer=2 filter=177 channel=67
					-3, 7, 0, -5, 2, 3, 4, 5, 4,
					-- layer=2 filter=177 channel=68
					1, 6, -11, 4, 4, -1, -1, -11, -3,
					-- layer=2 filter=177 channel=69
					3, 14, -2, -10, 7, 0, -7, 2, -10,
					-- layer=2 filter=177 channel=70
					-10, -13, -7, -11, -2, -7, -1, -13, -7,
					-- layer=2 filter=177 channel=71
					0, -12, -12, -15, -5, 7, -9, -4, -2,
					-- layer=2 filter=177 channel=72
					-5, -6, -8, -14, -6, -7, -10, -22, -14,
					-- layer=2 filter=177 channel=73
					5, -2, -3, 7, 1, -5, -3, 4, 6,
					-- layer=2 filter=177 channel=74
					-8, -3, 4, -13, -10, -2, 0, 2, -8,
					-- layer=2 filter=177 channel=75
					-10, -6, -2, -11, 3, -2, -4, -10, 4,
					-- layer=2 filter=177 channel=76
					-13, -1, -7, -4, 1, 2, 2, -9, -4,
					-- layer=2 filter=177 channel=77
					6, 8, 5, 7, -7, -1, 7, 0, 0,
					-- layer=2 filter=177 channel=78
					-10, -15, -8, -8, -11, 5, -3, -8, -4,
					-- layer=2 filter=177 channel=79
					-9, 4, 2, 0, 5, -1, 6, 6, -1,
					-- layer=2 filter=177 channel=80
					-9, -5, -10, -13, -11, 5, -7, -3, 7,
					-- layer=2 filter=177 channel=81
					7, -8, 8, -9, -3, 0, 0, 0, -5,
					-- layer=2 filter=177 channel=82
					0, 4, 7, -10, 1, 1, 0, -1, -1,
					-- layer=2 filter=177 channel=83
					-1, -6, 0, -1, 2, -7, 2, -6, -3,
					-- layer=2 filter=177 channel=84
					0, 2, -8, 3, -6, 7, -5, -6, -4,
					-- layer=2 filter=177 channel=85
					-10, 4, 5, -8, -5, -6, 7, 6, 8,
					-- layer=2 filter=177 channel=86
					3, 0, 4, -6, -7, 11, -10, -2, -1,
					-- layer=2 filter=177 channel=87
					-7, -12, -18, -6, -11, 1, 2, -12, -2,
					-- layer=2 filter=177 channel=88
					2, -3, -6, -15, 0, 1, 0, -9, 0,
					-- layer=2 filter=177 channel=89
					-9, 1, -2, -18, -20, -16, -4, 7, -8,
					-- layer=2 filter=177 channel=90
					7, 7, -5, 3, 10, 6, -6, 10, -2,
					-- layer=2 filter=177 channel=91
					0, 2, -3, -7, -13, 2, -4, -9, 7,
					-- layer=2 filter=177 channel=92
					7, 5, -8, -15, -6, -2, 4, 5, 0,
					-- layer=2 filter=177 channel=93
					5, -12, 0, 11, -10, 6, 3, -10, 2,
					-- layer=2 filter=177 channel=94
					-4, 10, 1, 2, -13, -6, 1, -11, -4,
					-- layer=2 filter=177 channel=95
					5, 2, -8, 3, -7, -11, 5, 0, -3,
					-- layer=2 filter=177 channel=96
					-13, -2, 13, -11, 3, 5, -6, -18, 10,
					-- layer=2 filter=177 channel=97
					-9, 2, -11, 4, 4, -10, -2, 0, -8,
					-- layer=2 filter=177 channel=98
					-5, -17, 3, -2, -18, -12, -13, -6, 0,
					-- layer=2 filter=177 channel=99
					-5, -6, -5, 0, -5, -6, -19, -24, 3,
					-- layer=2 filter=177 channel=100
					-6, -14, 0, -13, -10, 2, -2, -7, -1,
					-- layer=2 filter=177 channel=101
					-14, 1, -16, -19, 0, -5, -14, -10, -10,
					-- layer=2 filter=177 channel=102
					-5, -10, 15, -13, -2, -3, -1, -2, -18,
					-- layer=2 filter=177 channel=103
					8, 11, 7, 1, 4, -9, 7, -8, -8,
					-- layer=2 filter=177 channel=104
					-3, 4, -1, 2, -3, 4, 9, -14, 5,
					-- layer=2 filter=177 channel=105
					7, -12, 2, -7, -8, 2, -3, -6, 9,
					-- layer=2 filter=177 channel=106
					-9, -2, -12, 1, -5, -5, 0, -2, -11,
					-- layer=2 filter=177 channel=107
					-6, 10, -9, -5, 0, 8, 9, -7, 0,
					-- layer=2 filter=177 channel=108
					-4, -7, -10, -10, 11, -3, -11, -9, 5,
					-- layer=2 filter=177 channel=109
					1, -7, 2, 10, 1, -3, 9, -7, 0,
					-- layer=2 filter=177 channel=110
					15, 4, 1, 11, -2, -8, -6, 9, -15,
					-- layer=2 filter=177 channel=111
					1, -4, 3, -1, 8, -7, -6, 1, 0,
					-- layer=2 filter=177 channel=112
					-9, -14, 4, -10, -9, -8, 0, -10, 2,
					-- layer=2 filter=177 channel=113
					0, -8, -9, 0, -11, 5, 2, -9, -12,
					-- layer=2 filter=177 channel=114
					0, 9, -7, 5, 2, -7, 0, 11, 7,
					-- layer=2 filter=177 channel=115
					-8, 7, 10, 1, 2, -9, 4, 2, 0,
					-- layer=2 filter=177 channel=116
					-8, -4, -16, 4, 11, -5, 6, -11, 2,
					-- layer=2 filter=177 channel=117
					-6, -4, -6, -15, -17, -22, -2, -14, 0,
					-- layer=2 filter=177 channel=118
					2, -4, 1, -1, 3, 1, -3, 0, -6,
					-- layer=2 filter=177 channel=119
					-10, -12, -15, -12, -9, 2, -2, 0, 1,
					-- layer=2 filter=177 channel=120
					-5, -7, -7, -2, 8, 5, 2, -3, 3,
					-- layer=2 filter=177 channel=121
					-6, -7, 10, -5, 6, 3, 2, -1, -6,
					-- layer=2 filter=177 channel=122
					-4, -5, 8, 0, 8, -5, 4, -10, -5,
					-- layer=2 filter=177 channel=123
					-18, -6, -1, -14, -10, -15, -18, -8, -12,
					-- layer=2 filter=177 channel=124
					-1, 11, -6, 12, -10, -4, 1, 1, -1,
					-- layer=2 filter=177 channel=125
					-5, 2, 4, 9, -4, 5, 8, -8, -4,
					-- layer=2 filter=177 channel=126
					-2, -5, -6, -5, -9, 3, -1, -12, -6,
					-- layer=2 filter=177 channel=127
					-14, -3, -7, -3, -20, -14, -16, -16, -17,
					-- layer=2 filter=178 channel=0
					2, -8, -5, 2, -9, -17, 18, -2, 1,
					-- layer=2 filter=178 channel=1
					5, -8, 36, 31, -21, -9, -24, 20, -14,
					-- layer=2 filter=178 channel=2
					6, -10, 2, 0, 7, -7, 8, 0, -6,
					-- layer=2 filter=178 channel=3
					49, -54, -35, -28, -17, 0, 10, -5, 23,
					-- layer=2 filter=178 channel=4
					7, 19, 19, -7, -4, 0, -5, 2, 26,
					-- layer=2 filter=178 channel=5
					-14, -19, 22, -6, -10, -3, 14, 7, 41,
					-- layer=2 filter=178 channel=6
					-21, 25, 33, 8, -12, -6, 31, -73, -36,
					-- layer=2 filter=178 channel=7
					3, -13, 15, 13, 28, 1, 5, -8, -4,
					-- layer=2 filter=178 channel=8
					0, 0, 0, 9, 5, 2, 8, -7, -4,
					-- layer=2 filter=178 channel=9
					72, -21, -5, 16, -73, -20, 0, 44, 8,
					-- layer=2 filter=178 channel=10
					23, -25, -17, 4, 14, 2, 14, 6, 35,
					-- layer=2 filter=178 channel=11
					7, 5, -8, -15, -17, -6, -7, -1, 22,
					-- layer=2 filter=178 channel=12
					-18, -2, 18, -7, -15, -1, -2, 4, -22,
					-- layer=2 filter=178 channel=13
					3, 7, 0, 8, 4, -3, 5, 1, 0,
					-- layer=2 filter=178 channel=14
					-15, -4, 19, 22, -36, -31, -27, 10, -32,
					-- layer=2 filter=178 channel=15
					-3, 40, -44, 3, -33, 8, -12, -30, -11,
					-- layer=2 filter=178 channel=16
					10, -9, -32, -8, 21, -23, 19, 9, -22,
					-- layer=2 filter=178 channel=17
					8, -4, -3, 0, -3, 1, -4, -6, -4,
					-- layer=2 filter=178 channel=18
					51, 2, 44, 18, 16, -23, -20, -39, 6,
					-- layer=2 filter=178 channel=19
					16, 35, 37, 22, 13, 4, -17, -14, -32,
					-- layer=2 filter=178 channel=20
					0, 0, -2, 6, -10, -10, 5, 7, -10,
					-- layer=2 filter=178 channel=21
					8, 11, -8, 3, -4, -1, 29, 9, 0,
					-- layer=2 filter=178 channel=22
					9, -7, -8, -2, -7, -10, -6, 3, 3,
					-- layer=2 filter=178 channel=23
					-5, 23, 6, -15, -20, 1, 36, 15, 6,
					-- layer=2 filter=178 channel=24
					44, 0, -55, -30, -58, -45, -2, 5, 1,
					-- layer=2 filter=178 channel=25
					19, 19, -44, -18, -5, -5, -25, 0, 13,
					-- layer=2 filter=178 channel=26
					4, -5, -2, -8, -4, -4, 3, 10, -1,
					-- layer=2 filter=178 channel=27
					-2, -10, -3, -32, -63, -37, -35, -18, -6,
					-- layer=2 filter=178 channel=28
					13, 6, 2, 27, 36, 18, 22, 4, 38,
					-- layer=2 filter=178 channel=29
					4, 7, 2, 10, -1, 2, -5, 5, 3,
					-- layer=2 filter=178 channel=30
					20, -16, 1, -53, -32, -20, -13, 25, -22,
					-- layer=2 filter=178 channel=31
					-9, -71, -45, 6, -35, 74, -9, 47, -8,
					-- layer=2 filter=178 channel=32
					-6, -9, -1, -6, 4, -8, -4, 5, 5,
					-- layer=2 filter=178 channel=33
					-51, -25, -4, 6, -28, -11, -41, -3, 26,
					-- layer=2 filter=178 channel=34
					17, 15, 35, 21, 66, 22, 2, 14, -19,
					-- layer=2 filter=178 channel=35
					44, 20, 18, 30, 38, -9, 43, -6, 13,
					-- layer=2 filter=178 channel=36
					-11, 7, 0, -3, -14, 3, 10, -7, 1,
					-- layer=2 filter=178 channel=37
					11, 3, 12, -18, -13, 13, -3, 6, 18,
					-- layer=2 filter=178 channel=38
					-15, -9, -12, -20, -78, 11, 18, 12, 26,
					-- layer=2 filter=178 channel=39
					19, 8, -22, 3, 32, -19, -62, -12, 0,
					-- layer=2 filter=178 channel=40
					51, 37, -57, 18, 19, 30, -5, 39, 2,
					-- layer=2 filter=178 channel=41
					-6, 6, 4, 1, -8, 8, 9, 5, 0,
					-- layer=2 filter=178 channel=42
					13, 32, -23, -10, 14, -23, 33, 6, -42,
					-- layer=2 filter=178 channel=43
					56, -18, -3, 12, -9, -29, 21, -3, 25,
					-- layer=2 filter=178 channel=44
					1, -3, 8, -4, -3, 6, -12, -8, -5,
					-- layer=2 filter=178 channel=45
					56, -22, -32, 27, -46, -37, -5, -4, -29,
					-- layer=2 filter=178 channel=46
					1, -6, -25, -1, -16, -16, -8, 19, 1,
					-- layer=2 filter=178 channel=47
					0, -1, -25, 2, 18, -2, -3, 14, 16,
					-- layer=2 filter=178 channel=48
					-1, -7, 8, -7, 0, 2, -6, -9, -9,
					-- layer=2 filter=178 channel=49
					-4, -2, -14, 1, -29, -62, -30, -90, -62,
					-- layer=2 filter=178 channel=50
					4, 1, -13, -13, -13, -15, 0, 2, -3,
					-- layer=2 filter=178 channel=51
					-13, 0, -24, -12, -26, -22, -5, 7, 2,
					-- layer=2 filter=178 channel=52
					16, 37, -25, -22, -31, -26, -27, 41, 25,
					-- layer=2 filter=178 channel=53
					-11, 22, 0, -19, -16, 22, 20, -40, -8,
					-- layer=2 filter=178 channel=54
					9, 5, 9, 12, 32, 17, 12, 0, 18,
					-- layer=2 filter=178 channel=55
					-3, 5, -3, -11, -3, 5, 0, -4, 0,
					-- layer=2 filter=178 channel=56
					-3, 5, 5, -1, 5, -5, 8, 0, 24,
					-- layer=2 filter=178 channel=57
					-8, 13, 1, 11, 3, 1, 15, -3, -2,
					-- layer=2 filter=178 channel=58
					-8, 28, 3, 13, -18, 12, -15, -1, 7,
					-- layer=2 filter=178 channel=59
					-43, 9, 19, 21, 31, -12, 8, -40, 53,
					-- layer=2 filter=178 channel=60
					17, 28, -4, 8, 0, -10, 20, -8, -41,
					-- layer=2 filter=178 channel=61
					-7, -37, -38, 23, -18, -41, 34, -41, -35,
					-- layer=2 filter=178 channel=62
					-24, 4, 7, 29, 18, 26, 14, -50, -29,
					-- layer=2 filter=178 channel=63
					-13, -7, 0, 1, 0, 3, 26, 6, -1,
					-- layer=2 filter=178 channel=64
					-3, 1, -20, -25, -24, -21, -29, -3, -43,
					-- layer=2 filter=178 channel=65
					-34, 4, 1, 13, -22, -25, 33, -50, -41,
					-- layer=2 filter=178 channel=66
					-38, -13, 38, -21, 54, -6, 25, -12, -12,
					-- layer=2 filter=178 channel=67
					7, 21, 3, 0, -21, 9, 7, 30, 41,
					-- layer=2 filter=178 channel=68
					-3, 8, 8, -2, -4, 0, -1, -9, -6,
					-- layer=2 filter=178 channel=69
					6, 17, -18, 2, -10, -18, -24, -7, -33,
					-- layer=2 filter=178 channel=70
					18, 0, 16, 16, 29, 15, 11, -3, 11,
					-- layer=2 filter=178 channel=71
					25, 4, -30, 20, 12, -34, 6, -11, 24,
					-- layer=2 filter=178 channel=72
					-23, -6, 23, 5, -3, 10, 12, -14, -22,
					-- layer=2 filter=178 channel=73
					-23, -65, -85, -29, -13, -26, 3, 13, 30,
					-- layer=2 filter=178 channel=74
					-5, -38, -26, -11, -26, 3, -2, 2, -5,
					-- layer=2 filter=178 channel=75
					-48, -27, 3, -2, 5, -8, -3, -20, -50,
					-- layer=2 filter=178 channel=76
					-19, -31, -29, -27, -27, 37, 5, -7, 48,
					-- layer=2 filter=178 channel=77
					0, 10, 2, -8, -8, -7, -4, 2, 3,
					-- layer=2 filter=178 channel=78
					9, -10, -2, -32, -23, 5, -24, -21, 30,
					-- layer=2 filter=178 channel=79
					-3, -6, -3, -9, 1, -3, -5, -4, 5,
					-- layer=2 filter=178 channel=80
					25, 16, -14, -1, -9, -24, -20, 16, -21,
					-- layer=2 filter=178 channel=81
					6, 12, 4, 1, 12, 10, 8, -7, -6,
					-- layer=2 filter=178 channel=82
					0, 10, -2, -9, -10, -1, 4, 0, 5,
					-- layer=2 filter=178 channel=83
					24, 30, 18, -24, -8, 5, 42, -20, 6,
					-- layer=2 filter=178 channel=84
					-4, -1, 2, -4, 3, -6, 0, 8, 9,
					-- layer=2 filter=178 channel=85
					1, 2, 3, 2, 3, 3, 10, 0, 9,
					-- layer=2 filter=178 channel=86
					-9, -5, 1, 0, 1, -10, -7, -19, -9,
					-- layer=2 filter=178 channel=87
					38, 30, 5, 8, 42, 21, -5, 12, 25,
					-- layer=2 filter=178 channel=88
					9, -8, -2, 8, -1, 9, 8, 9, -7,
					-- layer=2 filter=178 channel=89
					-9, 4, 39, 18, -16, -16, -3, 5, -34,
					-- layer=2 filter=178 channel=90
					1, -4, -10, 6, 1, 7, -1, -9, 7,
					-- layer=2 filter=178 channel=91
					3, 28, 19, 35, 3, -16, 2, -6, -46,
					-- layer=2 filter=178 channel=92
					3, 17, 32, 16, -17, -2, -17, -19, -23,
					-- layer=2 filter=178 channel=93
					0, 47, 16, -3, -41, -3, 21, -13, -39,
					-- layer=2 filter=178 channel=94
					-6, 28, 23, 3, 0, 3, 20, -33, 5,
					-- layer=2 filter=178 channel=95
					7, 2, 11, 5, 5, 0, -4, -5, 3,
					-- layer=2 filter=178 channel=96
					-37, 24, -3, 2, 17, -23, 4, -36, -23,
					-- layer=2 filter=178 channel=97
					31, 4, -5, -13, -68, -13, -64, -24, -11,
					-- layer=2 filter=178 channel=98
					25, -27, -32, 24, 28, -1, 29, -3, 0,
					-- layer=2 filter=178 channel=99
					3, 32, -5, -3, 6, -13, 10, -49, 26,
					-- layer=2 filter=178 channel=100
					-10, -3, -1, -50, 5, 25, 39, 44, 31,
					-- layer=2 filter=178 channel=101
					36, -30, -14, 31, -41, -22, -13, -2, -14,
					-- layer=2 filter=178 channel=102
					-23, 7, -9, 4, 21, -86, -20, -21, -34,
					-- layer=2 filter=178 channel=103
					7, 7, 34, 27, 10, 26, 24, -11, -15,
					-- layer=2 filter=178 channel=104
					-25, 0, 15, -19, -2, -29, -52, -88, -10,
					-- layer=2 filter=178 channel=105
					65, -19, 71, 0, 30, 39, 14, -8, 19,
					-- layer=2 filter=178 channel=106
					4, 40, -16, 20, -25, -40, 6, 12, 26,
					-- layer=2 filter=178 channel=107
					-5, -1, -17, 31, -6, 7, 13, 5, -13,
					-- layer=2 filter=178 channel=108
					9, -4, 0, 0, -38, -43, -12, -9, -50,
					-- layer=2 filter=178 channel=109
					-4, 1, -4, -9, 15, 0, -8, 17, -2,
					-- layer=2 filter=178 channel=110
					-2, -7, -13, -13, 6, 0, 24, 0, -37,
					-- layer=2 filter=178 channel=111
					7, -6, -9, 7, 4, 9, -1, 3, 2,
					-- layer=2 filter=178 channel=112
					12, -1, -38, 26, -33, -1, 9, -17, 18,
					-- layer=2 filter=178 channel=113
					1, 8, -11, -28, -10, -14, 9, -7, 10,
					-- layer=2 filter=178 channel=114
					17, 9, -5, -9, 2, 11, 3, 15, 5,
					-- layer=2 filter=178 channel=115
					1, -10, -5, 12, -2, -6, -6, -3, 8,
					-- layer=2 filter=178 channel=116
					5, 61, 2, -7, 28, 2, -43, -4, 33,
					-- layer=2 filter=178 channel=117
					-7, -61, -8, 28, -16, 4, 0, 11, -18,
					-- layer=2 filter=178 channel=118
					0, -18, -17, -28, -11, 6, -13, -20, 15,
					-- layer=2 filter=178 channel=119
					32, 18, 7, 50, 28, -11, 11, -12, 43,
					-- layer=2 filter=178 channel=120
					-7, -3, 0, -3, 6, 5, -4, 0, 1,
					-- layer=2 filter=178 channel=121
					5, -6, -7, -5, 0, -1, -7, -3, 8,
					-- layer=2 filter=178 channel=122
					-3, -3, -2, -2, 5, -18, 0, 3, 4,
					-- layer=2 filter=178 channel=123
					-5, -21, -10, -11, 12, 19, 0, 6, -3,
					-- layer=2 filter=178 channel=124
					-9, 0, 20, -18, -15, 22, 6, -13, 62,
					-- layer=2 filter=178 channel=125
					-11, 0, 2, -2, -9, 9, -9, -7, 9,
					-- layer=2 filter=178 channel=126
					-26, -2, -32, 2, -14, -47, -3, -44, 1,
					-- layer=2 filter=178 channel=127
					-17, 13, 30, 9, -35, 8, 7, 26, 22,
					-- layer=2 filter=179 channel=0
					-13, -17, 3, -7, -6, 2, -11, 5, -10,
					-- layer=2 filter=179 channel=1
					-7, 3, -14, -8, -9, -4, -5, -9, -4,
					-- layer=2 filter=179 channel=2
					0, -8, 6, 7, 4, 6, 6, -4, 7,
					-- layer=2 filter=179 channel=3
					10, -10, -3, 0, 12, -8, -12, -3, -6,
					-- layer=2 filter=179 channel=4
					-6, -4, 9, 0, -6, 1, -3, 2, 1,
					-- layer=2 filter=179 channel=5
					-4, -10, 1, 3, -14, -6, 5, 6, -8,
					-- layer=2 filter=179 channel=6
					3, -8, 3, 6, -16, -11, -2, -8, 0,
					-- layer=2 filter=179 channel=7
					-2, 11, 4, 0, -8, -6, -12, 5, -13,
					-- layer=2 filter=179 channel=8
					0, 6, -1, 0, -2, -6, 0, 3, 5,
					-- layer=2 filter=179 channel=9
					-14, -3, -12, -14, 1, -13, -13, -4, 4,
					-- layer=2 filter=179 channel=10
					4, -9, 4, -2, -6, 0, -6, -2, 3,
					-- layer=2 filter=179 channel=11
					-7, 0, 6, 2, 7, 1, 0, -12, -2,
					-- layer=2 filter=179 channel=12
					-6, -8, -9, 0, 0, -10, 5, 5, 3,
					-- layer=2 filter=179 channel=13
					-3, -11, -6, 9, -3, 1, -6, -10, 9,
					-- layer=2 filter=179 channel=14
					-8, -13, -15, -7, 2, 6, -10, 5, -12,
					-- layer=2 filter=179 channel=15
					-2, 6, -8, 4, -2, -1, 0, -3, -2,
					-- layer=2 filter=179 channel=16
					-4, -10, -1, -7, -5, -10, 6, -8, 4,
					-- layer=2 filter=179 channel=17
					11, 4, -5, 0, -2, -2, 10, 6, 8,
					-- layer=2 filter=179 channel=18
					6, 4, -3, 3, -9, -1, -4, 7, 6,
					-- layer=2 filter=179 channel=19
					8, -9, -1, -10, -5, -10, -11, -2, -13,
					-- layer=2 filter=179 channel=20
					3, -7, -1, 11, -5, -7, 1, -4, 0,
					-- layer=2 filter=179 channel=21
					-1, -10, -8, -7, 7, 6, -5, 2, -4,
					-- layer=2 filter=179 channel=22
					-4, 6, 9, 7, 7, 0, -10, 9, -4,
					-- layer=2 filter=179 channel=23
					-15, -9, -11, -9, 8, 0, -11, 3, 5,
					-- layer=2 filter=179 channel=24
					0, -16, -8, 2, -10, -9, 7, -6, 2,
					-- layer=2 filter=179 channel=25
					-5, -4, -3, 4, -4, 0, -7, -5, -5,
					-- layer=2 filter=179 channel=26
					8, -5, 0, -3, 10, 2, -1, 9, 4,
					-- layer=2 filter=179 channel=27
					-3, -11, -14, -3, -4, 6, -3, 4, 4,
					-- layer=2 filter=179 channel=28
					-3, -8, 4, -4, 10, -4, 7, -4, -3,
					-- layer=2 filter=179 channel=29
					0, 0, -1, 8, 6, -6, 0, -7, 3,
					-- layer=2 filter=179 channel=30
					-16, 0, 5, -15, 0, -8, -5, -9, -1,
					-- layer=2 filter=179 channel=31
					1, -5, 0, 4, 0, -4, -6, 0, -3,
					-- layer=2 filter=179 channel=32
					4, 0, -6, -2, -2, 11, 11, 8, 6,
					-- layer=2 filter=179 channel=33
					-5, -4, 0, 2, 8, -7, 7, 5, -11,
					-- layer=2 filter=179 channel=34
					-17, -9, -9, -14, -13, 4, 4, -4, -6,
					-- layer=2 filter=179 channel=35
					-1, -10, -9, -6, 1, 7, -4, -4, 9,
					-- layer=2 filter=179 channel=36
					0, -2, 0, 8, 11, -8, 5, -12, 5,
					-- layer=2 filter=179 channel=37
					-1, -3, -4, 7, -5, -6, -5, 7, 0,
					-- layer=2 filter=179 channel=38
					-4, -14, -7, 3, 0, -5, -6, -3, -1,
					-- layer=2 filter=179 channel=39
					-7, -3, 4, -12, -4, -9, 2, -9, -2,
					-- layer=2 filter=179 channel=40
					-3, -7, -14, -13, -13, -7, 3, -7, -12,
					-- layer=2 filter=179 channel=41
					6, 0, -1, -6, -8, 2, 8, -12, -10,
					-- layer=2 filter=179 channel=42
					2, -12, 8, -13, -9, -11, -6, -4, 7,
					-- layer=2 filter=179 channel=43
					-1, 0, 0, -12, -7, -14, -5, 2, -7,
					-- layer=2 filter=179 channel=44
					-6, 2, 3, 10, -3, 0, -1, -3, -10,
					-- layer=2 filter=179 channel=45
					-4, -5, -4, -9, -2, -9, -12, -12, -14,
					-- layer=2 filter=179 channel=46
					-14, -6, 3, -12, -5, 6, -4, -10, 0,
					-- layer=2 filter=179 channel=47
					8, 3, 0, -14, 1, -7, -9, -3, 1,
					-- layer=2 filter=179 channel=48
					5, -6, 0, 7, -3, -6, -5, 4, 5,
					-- layer=2 filter=179 channel=49
					-7, 4, 5, 5, -9, -6, 1, 1, 3,
					-- layer=2 filter=179 channel=50
					5, 9, 1, 3, 1, 1, 0, 10, 0,
					-- layer=2 filter=179 channel=51
					-14, -12, -10, -8, -4, 0, -17, 7, -11,
					-- layer=2 filter=179 channel=52
					3, -8, -4, 1, 0, -6, -5, -3, -5,
					-- layer=2 filter=179 channel=53
					7, -12, 1, 0, -13, 6, -7, -18, -7,
					-- layer=2 filter=179 channel=54
					8, -14, -6, -13, -1, 4, -10, 2, -10,
					-- layer=2 filter=179 channel=55
					4, -7, -7, 8, -4, -8, 9, 0, -1,
					-- layer=2 filter=179 channel=56
					0, -3, -8, -1, 2, -10, 1, -6, -12,
					-- layer=2 filter=179 channel=57
					-1, -4, 2, 4, 9, 7, 3, 7, 1,
					-- layer=2 filter=179 channel=58
					-2, -1, -15, -5, 0, -8, 0, 0, -11,
					-- layer=2 filter=179 channel=59
					-9, 0, -6, -6, -14, -6, -7, 0, -8,
					-- layer=2 filter=179 channel=60
					-10, -4, -6, -18, -4, -5, -7, -4, -2,
					-- layer=2 filter=179 channel=61
					-16, 0, 6, -4, -3, 1, -5, -6, -8,
					-- layer=2 filter=179 channel=62
					-15, 3, -4, -14, -7, 0, -3, 6, -14,
					-- layer=2 filter=179 channel=63
					-4, -6, 0, 1, -19, -13, -2, -15, 8,
					-- layer=2 filter=179 channel=64
					-9, -6, 3, -1, -13, 1, -8, -14, 4,
					-- layer=2 filter=179 channel=65
					-5, -13, -9, -19, -9, -1, -7, 2, 0,
					-- layer=2 filter=179 channel=66
					0, -8, 9, 6, -8, -1, 0, -3, -9,
					-- layer=2 filter=179 channel=67
					-3, 7, 0, -5, -12, 1, -5, -2, -16,
					-- layer=2 filter=179 channel=68
					5, 0, 8, -10, -9, -1, -10, 8, 3,
					-- layer=2 filter=179 channel=69
					-13, -6, 3, 0, 1, -4, -9, 8, -6,
					-- layer=2 filter=179 channel=70
					-13, -6, -10, 1, -6, -2, -2, -10, 0,
					-- layer=2 filter=179 channel=71
					-9, -3, -13, -3, 0, 1, 5, -1, 3,
					-- layer=2 filter=179 channel=72
					-2, -6, -1, -5, 2, 11, -15, -11, -5,
					-- layer=2 filter=179 channel=73
					-3, 0, -1, 4, -6, -10, 1, -5, -17,
					-- layer=2 filter=179 channel=74
					-11, -6, -4, -11, -8, -10, -4, 4, 0,
					-- layer=2 filter=179 channel=75
					-10, 5, -12, -3, -2, -5, -8, 11, 0,
					-- layer=2 filter=179 channel=76
					-7, -2, 1, -16, -6, -9, -14, -9, -11,
					-- layer=2 filter=179 channel=77
					-10, 4, 0, 5, 0, -1, 3, -9, -4,
					-- layer=2 filter=179 channel=78
					-5, -3, 0, -9, 5, -11, 4, 5, -10,
					-- layer=2 filter=179 channel=79
					1, -1, -1, -3, 7, -8, 10, 6, 5,
					-- layer=2 filter=179 channel=80
					-8, -8, 4, -12, -4, 0, -9, -4, 1,
					-- layer=2 filter=179 channel=81
					3, -3, -2, -2, -6, 6, 8, -8, 3,
					-- layer=2 filter=179 channel=82
					4, -7, -2, 5, 9, -2, -2, 5, 5,
					-- layer=2 filter=179 channel=83
					2, -7, -5, 4, 4, -3, 3, -8, 6,
					-- layer=2 filter=179 channel=84
					1, 3, -1, 4, 2, -11, 6, -3, 5,
					-- layer=2 filter=179 channel=85
					-8, -6, 6, 6, 5, 8, 7, -9, 6,
					-- layer=2 filter=179 channel=86
					-3, 3, 2, -1, -9, -5, 0, 6, 0,
					-- layer=2 filter=179 channel=87
					2, 4, 0, -11, -1, 3, -2, -15, 9,
					-- layer=2 filter=179 channel=88
					-7, 4, 6, 1, 0, 4, 1, -16, 8,
					-- layer=2 filter=179 channel=89
					-5, 1, -10, -9, -9, -3, -7, -2, -3,
					-- layer=2 filter=179 channel=90
					-7, 1, 0, -8, -3, -2, 3, -3, -1,
					-- layer=2 filter=179 channel=91
					1, -1, -4, -3, -14, 1, -9, -12, -11,
					-- layer=2 filter=179 channel=92
					0, -8, 5, -8, 0, 0, 2, 9, -8,
					-- layer=2 filter=179 channel=93
					5, 6, 9, 3, 0, -11, -16, -13, -5,
					-- layer=2 filter=179 channel=94
					4, -5, 1, -11, -9, -5, 0, -6, 2,
					-- layer=2 filter=179 channel=95
					0, -3, -6, 2, 8, 3, 2, 7, 0,
					-- layer=2 filter=179 channel=96
					-1, 0, -14, -11, -2, -2, 4, -7, -1,
					-- layer=2 filter=179 channel=97
					-6, -4, -6, -2, -4, -7, 0, -8, -5,
					-- layer=2 filter=179 channel=98
					5, -14, -8, -5, 0, -3, -10, -1, 6,
					-- layer=2 filter=179 channel=99
					-8, -11, -18, -5, -14, -19, -11, -6, -7,
					-- layer=2 filter=179 channel=100
					-5, 0, 0, -15, 1, -5, 1, -12, -6,
					-- layer=2 filter=179 channel=101
					8, 2, -2, 0, -5, 0, 0, -2, 0,
					-- layer=2 filter=179 channel=102
					-4, -15, -7, 6, 5, 0, -11, -2, -8,
					-- layer=2 filter=179 channel=103
					-8, -11, 0, 2, -11, 0, 9, 3, 0,
					-- layer=2 filter=179 channel=104
					4, -12, 8, 4, -14, -6, 2, -10, 5,
					-- layer=2 filter=179 channel=105
					-7, -15, 3, -9, 4, -2, -5, -5, -2,
					-- layer=2 filter=179 channel=106
					-4, -3, 7, -11, -15, -8, -3, 5, 0,
					-- layer=2 filter=179 channel=107
					-6, -6, -7, -2, 2, -8, 5, 2, -6,
					-- layer=2 filter=179 channel=108
					-1, -12, -7, 2, -4, -1, 3, -11, -11,
					-- layer=2 filter=179 channel=109
					5, -1, 2, -9, 0, 8, -3, -9, -6,
					-- layer=2 filter=179 channel=110
					-17, -4, -4, -10, -3, 1, -3, -8, -11,
					-- layer=2 filter=179 channel=111
					-6, -2, -4, 3, 4, 0, 5, 7, -2,
					-- layer=2 filter=179 channel=112
					-10, -16, -3, -6, -4, -6, -2, 8, -8,
					-- layer=2 filter=179 channel=113
					-21, -1, 9, -4, -3, -4, -11, -4, 0,
					-- layer=2 filter=179 channel=114
					-2, 4, -5, 5, 4, -1, 1, -8, 0,
					-- layer=2 filter=179 channel=115
					-1, 6, 6, 0, 4, -10, -9, 3, 9,
					-- layer=2 filter=179 channel=116
					-4, 3, 2, 1, 5, -7, -13, -6, -6,
					-- layer=2 filter=179 channel=117
					-15, -2, -7, -19, 1, 0, -13, -16, -16,
					-- layer=2 filter=179 channel=118
					4, 5, -11, 0, -6, -10, 5, -12, -12,
					-- layer=2 filter=179 channel=119
					0, -4, 6, -11, -1, 5, -11, -9, -10,
					-- layer=2 filter=179 channel=120
					8, 6, -4, 8, -2, 6, 7, -4, 5,
					-- layer=2 filter=179 channel=121
					0, 8, 10, -7, 10, 1, -1, -3, 7,
					-- layer=2 filter=179 channel=122
					9, 10, 0, -3, -4, 0, 3, -5, 5,
					-- layer=2 filter=179 channel=123
					2, 7, -4, 0, 7, 7, -7, -2, 2,
					-- layer=2 filter=179 channel=124
					-4, 7, -3, -4, -2, 0, 0, -7, 0,
					-- layer=2 filter=179 channel=125
					2, 4, -5, -3, -10, -9, -1, -1, 8,
					-- layer=2 filter=179 channel=126
					-5, -5, 6, 11, 1, 7, 4, -11, 10,
					-- layer=2 filter=179 channel=127
					2, 1, -16, -1, 4, -1, -15, 4, -4,
					-- layer=2 filter=180 channel=0
					-2, -13, -7, -12, -10, 0, -11, 2, 0,
					-- layer=2 filter=180 channel=1
					6, -2, -11, 0, 1, 5, -2, -2, -17,
					-- layer=2 filter=180 channel=2
					-3, 7, 1, 7, 8, -7, -11, -6, 5,
					-- layer=2 filter=180 channel=3
					-12, 1, 3, 6, 1, 4, -5, 7, -12,
					-- layer=2 filter=180 channel=4
					-8, -11, -4, -4, -1, 8, -3, -5, 0,
					-- layer=2 filter=180 channel=5
					-10, -12, 6, -1, -1, 5, 6, -9, -5,
					-- layer=2 filter=180 channel=6
					-3, -3, -8, 6, -9, -6, 3, 1, -6,
					-- layer=2 filter=180 channel=7
					2, -11, 3, -8, -4, -14, -10, -14, -11,
					-- layer=2 filter=180 channel=8
					6, 10, 2, -9, 2, -9, -8, 1, -2,
					-- layer=2 filter=180 channel=9
					1, 0, -6, -5, -1, -6, 2, -5, -7,
					-- layer=2 filter=180 channel=10
					3, -8, -5, 1, 5, -5, 0, -5, 8,
					-- layer=2 filter=180 channel=11
					-11, -5, -1, 0, -3, -11, -17, -11, -2,
					-- layer=2 filter=180 channel=12
					4, -11, -4, 3, 5, -2, 4, 6, 2,
					-- layer=2 filter=180 channel=13
					5, 10, -1, -8, -5, -2, 10, -1, -6,
					-- layer=2 filter=180 channel=14
					-3, -9, 0, 4, 0, 1, -3, -9, -16,
					-- layer=2 filter=180 channel=15
					8, 4, 5, 7, -4, -10, 3, -1, 1,
					-- layer=2 filter=180 channel=16
					2, 2, 6, 5, -10, 8, 4, -1, -5,
					-- layer=2 filter=180 channel=17
					10, 5, -7, 7, 6, 5, 9, -7, 4,
					-- layer=2 filter=180 channel=18
					-11, -9, -1, 5, -8, 2, 4, 1, 1,
					-- layer=2 filter=180 channel=19
					2, 9, -9, -5, 2, -8, -3, -10, 4,
					-- layer=2 filter=180 channel=20
					-4, -9, 4, 7, 7, -5, -11, 1, -1,
					-- layer=2 filter=180 channel=21
					-2, -1, 2, 6, 6, -3, 2, -3, -2,
					-- layer=2 filter=180 channel=22
					8, 11, 7, 0, -2, 0, -6, 0, 0,
					-- layer=2 filter=180 channel=23
					4, 0, -4, 0, -9, -10, 2, 1, -2,
					-- layer=2 filter=180 channel=24
					-4, 2, 0, 6, 0, -8, -4, 7, -1,
					-- layer=2 filter=180 channel=25
					5, 1, 6, -5, -3, -8, 0, -12, 6,
					-- layer=2 filter=180 channel=26
					8, -9, -1, -8, -9, 5, 1, 5, -4,
					-- layer=2 filter=180 channel=27
					-8, 5, -10, -5, 0, 6, 1, -8, 8,
					-- layer=2 filter=180 channel=28
					-7, -3, -8, -1, 6, -16, 3, 0, -5,
					-- layer=2 filter=180 channel=29
					-7, -1, -6, 0, 4, -3, 5, -8, 0,
					-- layer=2 filter=180 channel=30
					-16, -3, -4, -1, 5, 3, -3, 3, -13,
					-- layer=2 filter=180 channel=31
					-3, -8, -9, 1, 3, -5, -4, 1, -11,
					-- layer=2 filter=180 channel=32
					-2, 2, 0, 6, 4, 6, 1, 2, 0,
					-- layer=2 filter=180 channel=33
					3, 8, 4, -7, 1, -12, -1, 7, 0,
					-- layer=2 filter=180 channel=34
					-5, -8, -8, -2, -11, 6, -1, -7, 6,
					-- layer=2 filter=180 channel=35
					5, -8, -3, 7, -14, -8, -9, 2, 0,
					-- layer=2 filter=180 channel=36
					-7, -5, 7, -3, 4, -3, 5, -6, -7,
					-- layer=2 filter=180 channel=37
					-11, -15, -5, 3, -13, -1, 2, -9, -5,
					-- layer=2 filter=180 channel=38
					2, -11, 6, 3, -10, -7, 1, -13, -2,
					-- layer=2 filter=180 channel=39
					7, 2, 1, 1, 0, -12, 6, -11, -5,
					-- layer=2 filter=180 channel=40
					4, 3, -9, -7, -8, 3, -5, 3, 10,
					-- layer=2 filter=180 channel=41
					10, -3, -7, -4, 10, -1, 5, -7, -7,
					-- layer=2 filter=180 channel=42
					-10, 3, -9, 4, -4, 4, 2, 2, -3,
					-- layer=2 filter=180 channel=43
					-8, -11, 0, -8, 3, -1, 3, -3, 3,
					-- layer=2 filter=180 channel=44
					0, 9, 2, 8, -3, -8, -5, 4, 1,
					-- layer=2 filter=180 channel=45
					5, -7, -11, -1, -9, 6, 1, 1, -7,
					-- layer=2 filter=180 channel=46
					-5, -10, -6, -11, -6, -14, -11, -1, 6,
					-- layer=2 filter=180 channel=47
					4, 3, 9, -2, -5, -9, -6, -10, -4,
					-- layer=2 filter=180 channel=48
					-5, 5, -8, 8, 3, 3, 9, -6, 2,
					-- layer=2 filter=180 channel=49
					-2, -7, -8, -2, -11, 8, -9, -2, -3,
					-- layer=2 filter=180 channel=50
					4, -9, -1, -2, 0, 0, 6, 2, 4,
					-- layer=2 filter=180 channel=51
					0, -7, -10, -15, -9, 0, -12, -6, -12,
					-- layer=2 filter=180 channel=52
					4, -11, 3, 0, -14, -7, -6, 8, -2,
					-- layer=2 filter=180 channel=53
					-11, -4, 4, 4, -3, -8, -10, 4, -11,
					-- layer=2 filter=180 channel=54
					-5, 1, -1, -10, -17, -8, 3, -1, 6,
					-- layer=2 filter=180 channel=55
					9, -1, 4, -6, 11, 4, 2, 7, -7,
					-- layer=2 filter=180 channel=56
					4, 4, -7, -6, 2, 6, -5, -11, 1,
					-- layer=2 filter=180 channel=57
					-7, -1, 5, -1, 4, 5, -6, -6, 4,
					-- layer=2 filter=180 channel=58
					6, -12, 4, 2, -9, 2, 0, 1, -1,
					-- layer=2 filter=180 channel=59
					-16, 2, -9, -9, -4, -8, -7, 0, 10,
					-- layer=2 filter=180 channel=60
					0, 3, 3, -5, -6, 8, 5, -6, 0,
					-- layer=2 filter=180 channel=61
					-6, -1, -11, -5, 3, -6, 6, 5, 2,
					-- layer=2 filter=180 channel=62
					-8, -15, -10, -9, -6, -9, -1, 3, -4,
					-- layer=2 filter=180 channel=63
					-12, -5, -15, 0, -5, -7, -4, -10, -9,
					-- layer=2 filter=180 channel=64
					-11, -8, 3, -4, -4, 0, 3, -11, -7,
					-- layer=2 filter=180 channel=65
					0, 5, -1, 3, -12, -2, -11, 0, -8,
					-- layer=2 filter=180 channel=66
					0, 1, -4, -7, 6, 3, -2, 2, 0,
					-- layer=2 filter=180 channel=67
					7, 6, -4, 6, -8, -5, 1, 1, -1,
					-- layer=2 filter=180 channel=68
					2, -7, -10, -1, -8, 0, -12, -8, 6,
					-- layer=2 filter=180 channel=69
					4, 2, 4, -2, -12, 4, -8, 1, -10,
					-- layer=2 filter=180 channel=70
					-14, -11, -11, -12, -15, 0, 4, -18, -14,
					-- layer=2 filter=180 channel=71
					-5, 6, -6, -8, 0, 4, -9, 2, 2,
					-- layer=2 filter=180 channel=72
					-8, -6, 3, -16, -13, 1, -11, -7, -9,
					-- layer=2 filter=180 channel=73
					-3, 0, 4, -8, -6, -1, -4, 2, 2,
					-- layer=2 filter=180 channel=74
					-10, -2, 2, 2, -6, 2, 1, -6, -9,
					-- layer=2 filter=180 channel=75
					-8, 5, 8, 11, 4, -4, 6, 3, 3,
					-- layer=2 filter=180 channel=76
					8, -17, 5, -3, 0, -4, 0, 9, -1,
					-- layer=2 filter=180 channel=77
					0, 0, 7, 0, -6, -3, 1, 5, 10,
					-- layer=2 filter=180 channel=78
					-2, -8, -9, -7, 5, 0, 0, -1, 2,
					-- layer=2 filter=180 channel=79
					6, -4, -1, -3, 1, -9, 7, -11, 1,
					-- layer=2 filter=180 channel=80
					7, 8, 0, -5, 8, -12, -5, 6, -3,
					-- layer=2 filter=180 channel=81
					0, -3, 4, -9, -8, -1, -5, -2, 4,
					-- layer=2 filter=180 channel=82
					-8, -4, -8, 3, -5, -1, 2, 8, -1,
					-- layer=2 filter=180 channel=83
					3, -13, -11, -1, 0, 7, -3, -15, -13,
					-- layer=2 filter=180 channel=84
					-10, 9, 3, -8, 2, 3, -4, -9, 3,
					-- layer=2 filter=180 channel=85
					0, 0, -8, -5, 1, 0, -6, -4, 5,
					-- layer=2 filter=180 channel=86
					7, 0, 8, -5, 1, 9, -2, 0, -10,
					-- layer=2 filter=180 channel=87
					-5, -3, 7, 1, -16, -7, 0, -5, -5,
					-- layer=2 filter=180 channel=88
					-9, -1, 4, -6, 3, -6, 8, -11, -11,
					-- layer=2 filter=180 channel=89
					-5, -8, 3, 3, -8, -9, -5, -4, -1,
					-- layer=2 filter=180 channel=90
					2, -4, -6, -9, 5, 0, 7, -2, 4,
					-- layer=2 filter=180 channel=91
					-6, -5, 6, -16, 8, -7, -2, 1, -11,
					-- layer=2 filter=180 channel=92
					-6, -11, 1, -11, -2, -4, -1, 4, -5,
					-- layer=2 filter=180 channel=93
					6, -2, 4, 3, 0, 2, -4, 3, -3,
					-- layer=2 filter=180 channel=94
					0, -6, -4, -12, -9, -11, -4, -10, 1,
					-- layer=2 filter=180 channel=95
					5, 4, 2, 0, 2, -10, -9, -7, 9,
					-- layer=2 filter=180 channel=96
					5, -4, -2, -7, 0, -8, -3, 7, 5,
					-- layer=2 filter=180 channel=97
					-8, -1, 8, -8, -6, -6, -12, -9, -10,
					-- layer=2 filter=180 channel=98
					4, -20, -10, -16, -14, 0, -8, -10, -3,
					-- layer=2 filter=180 channel=99
					-3, 2, -10, 1, -9, -3, -2, 2, 3,
					-- layer=2 filter=180 channel=100
					7, -9, -1, -9, -11, -5, -3, 2, 2,
					-- layer=2 filter=180 channel=101
					-10, 6, -9, -6, 2, 0, 2, 4, 6,
					-- layer=2 filter=180 channel=102
					-5, -10, -2, 9, -5, -8, -13, -9, -3,
					-- layer=2 filter=180 channel=103
					3, -1, -12, -10, -7, 5, -5, 6, -1,
					-- layer=2 filter=180 channel=104
					0, -8, 8, -3, -7, 4, -5, 3, -5,
					-- layer=2 filter=180 channel=105
					-9, 3, -10, 6, 0, -9, 0, -8, 7,
					-- layer=2 filter=180 channel=106
					0, 2, 1, -5, 0, -1, -4, -3, -11,
					-- layer=2 filter=180 channel=107
					0, -8, -5, 4, 3, 2, -2, 5, -4,
					-- layer=2 filter=180 channel=108
					4, -1, 2, 1, -1, -2, -5, 9, -11,
					-- layer=2 filter=180 channel=109
					5, -6, 7, 5, -3, 5, 5, 6, -8,
					-- layer=2 filter=180 channel=110
					5, -6, -2, 2, -1, 0, 4, -6, 2,
					-- layer=2 filter=180 channel=111
					-4, -4, -8, -2, 3, 2, 1, -2, -3,
					-- layer=2 filter=180 channel=112
					-2, 0, -3, 1, 3, -9, -7, 3, 1,
					-- layer=2 filter=180 channel=113
					2, 3, -7, -8, -2, 1, -12, -5, -6,
					-- layer=2 filter=180 channel=114
					4, -1, 10, 7, -9, -10, -6, 10, 2,
					-- layer=2 filter=180 channel=115
					-1, -7, 5, -2, 1, 5, 9, 1, -6,
					-- layer=2 filter=180 channel=116
					0, -5, 3, -7, 1, -10, 2, -1, 0,
					-- layer=2 filter=180 channel=117
					-12, 2, -12, 2, -13, -8, -1, -11, 0,
					-- layer=2 filter=180 channel=118
					2, -9, -12, -5, -5, 4, 5, 6, 0,
					-- layer=2 filter=180 channel=119
					-1, -8, -7, -5, 2, -13, -3, 0, 9,
					-- layer=2 filter=180 channel=120
					1, -3, 5, -4, -8, 3, -5, -9, 10,
					-- layer=2 filter=180 channel=121
					7, 0, -11, -4, 5, 3, 2, 0, 1,
					-- layer=2 filter=180 channel=122
					0, -7, 5, 4, 6, 8, -3, -1, -9,
					-- layer=2 filter=180 channel=123
					6, -4, -10, -12, -16, 10, -2, 2, 6,
					-- layer=2 filter=180 channel=124
					4, 5, 6, -10, -6, -5, -13, 4, 7,
					-- layer=2 filter=180 channel=125
					-5, 2, 11, -1, 11, -1, 0, -4, -8,
					-- layer=2 filter=180 channel=126
					-3, 6, -5, -1, 6, -4, -9, -5, 4,
					-- layer=2 filter=180 channel=127
					3, 1, -3, -2, 1, -4, -1, 0, 4,
					-- layer=2 filter=181 channel=0
					2, -9, -4, -21, 19, 5, 0, 10, -19,
					-- layer=2 filter=181 channel=1
					0, 20, -11, 2, 0, 13, -36, -25, -37,
					-- layer=2 filter=181 channel=2
					1, -4, -6, 0, -10, 4, 0, -3, -1,
					-- layer=2 filter=181 channel=3
					-59, -6, -16, 15, 18, -8, -22, -17, 12,
					-- layer=2 filter=181 channel=4
					45, -30, 20, 43, -26, -39, 1, -32, 48,
					-- layer=2 filter=181 channel=5
					-12, -31, 5, 17, 20, -11, -13, -8, -45,
					-- layer=2 filter=181 channel=6
					-8, -11, -13, -12, -40, 15, 2, 21, -7,
					-- layer=2 filter=181 channel=7
					31, 4, -42, -22, -38, -3, -16, 24, 44,
					-- layer=2 filter=181 channel=8
					8, -6, -6, 0, -5, -9, -5, -3, 0,
					-- layer=2 filter=181 channel=9
					-37, -69, -57, -19, -86, -23, -6, 1, -9,
					-- layer=2 filter=181 channel=10
					-39, -20, 0, 8, 13, -15, 30, 13, -17,
					-- layer=2 filter=181 channel=11
					-6, -14, 11, 6, -2, -21, -39, -24, -13,
					-- layer=2 filter=181 channel=12
					-20, 20, 4, -28, -23, 23, -31, -34, -10,
					-- layer=2 filter=181 channel=13
					1, -9, -2, 1, 7, -11, -3, 8, -1,
					-- layer=2 filter=181 channel=14
					-21, -31, -11, -13, -13, 3, -30, -58, -57,
					-- layer=2 filter=181 channel=15
					25, -26, -23, 5, 24, 7, -22, -101, -6,
					-- layer=2 filter=181 channel=16
					-3, 4, -39, -14, -40, -12, 0, -23, 6,
					-- layer=2 filter=181 channel=17
					10, 5, -4, 6, 0, 9, -8, -1, 3,
					-- layer=2 filter=181 channel=18
					-9, -39, -17, 7, -33, -4, -23, -2, -3,
					-- layer=2 filter=181 channel=19
					33, 20, 21, 30, 19, 4, 3, 14, -35,
					-- layer=2 filter=181 channel=20
					7, 9, 8, 0, 1, -2, -5, -2, 10,
					-- layer=2 filter=181 channel=21
					7, -7, 8, 6, 0, -4, 6, -10, -4,
					-- layer=2 filter=181 channel=22
					2, 1, -3, -5, -4, 9, 2, 6, -2,
					-- layer=2 filter=181 channel=23
					-12, -33, -42, -3, -30, -39, 18, -3, 40,
					-- layer=2 filter=181 channel=24
					-68, -39, -59, -24, -50, -58, 6, 41, 18,
					-- layer=2 filter=181 channel=25
					0, -44, -66, -34, -28, -68, -42, 16, 25,
					-- layer=2 filter=181 channel=26
					-10, -6, 5, 8, -10, -1, 7, 4, 8,
					-- layer=2 filter=181 channel=27
					51, 29, 27, 25, 37, 11, -29, -42, -38,
					-- layer=2 filter=181 channel=28
					-40, -2, 8, 19, 3, 10, 56, -19, -25,
					-- layer=2 filter=181 channel=29
					0, -7, 0, 6, -5, -5, -4, -10, 8,
					-- layer=2 filter=181 channel=30
					7, 17, -15, 28, -14, -31, 20, 17, -22,
					-- layer=2 filter=181 channel=31
					17, 8, -6, 34, 33, -19, 16, -35, -12,
					-- layer=2 filter=181 channel=32
					0, -7, 5, -1, 8, -7, 6, 3, -4,
					-- layer=2 filter=181 channel=33
					31, -6, -32, 4, -38, -6, -88, 0, 1,
					-- layer=2 filter=181 channel=34
					-13, -16, -51, -11, -2, -28, 2, -21, -34,
					-- layer=2 filter=181 channel=35
					19, 5, 27, 30, 32, 28, 54, 22, 18,
					-- layer=2 filter=181 channel=36
					-2, -8, 6, -12, -3, 8, -8, 7, 5,
					-- layer=2 filter=181 channel=37
					-5, 1, 7, 8, 21, -9, -37, -22, -30,
					-- layer=2 filter=181 channel=38
					30, 12, 21, 22, 24, -4, -31, -39, -48,
					-- layer=2 filter=181 channel=39
					-49, -16, -63, -23, -33, -51, 3, 1, 9,
					-- layer=2 filter=181 channel=40
					-58, 62, -19, 41, 31, -59, 26, -23, 8,
					-- layer=2 filter=181 channel=41
					6, -8, 5, -2, -7, 5, 8, 4, -5,
					-- layer=2 filter=181 channel=42
					-29, -17, -9, -30, -13, 1, 19, -9, 35,
					-- layer=2 filter=181 channel=43
					-11, -34, 42, 20, -2, 30, -18, -78, -18,
					-- layer=2 filter=181 channel=44
					-7, -1, 6, -8, 7, 1, -7, -10, 4,
					-- layer=2 filter=181 channel=45
					68, 58, 73, 30, 42, 32, -3, -21, 25,
					-- layer=2 filter=181 channel=46
					13, 0, -29, 40, 0, -7, -2, 14, -12,
					-- layer=2 filter=181 channel=47
					13, 21, 26, -5, -37, 6, 11, -11, -6,
					-- layer=2 filter=181 channel=48
					-10, 4, -1, 1, 4, 1, -7, 0, 0,
					-- layer=2 filter=181 channel=49
					-21, -64, -16, 3, -35, 20, -1, -48, -15,
					-- layer=2 filter=181 channel=50
					-4, 9, 10, 19, 1, 2, -13, -18, 16,
					-- layer=2 filter=181 channel=51
					-11, -17, -14, -9, -8, -22, -21, -3, -10,
					-- layer=2 filter=181 channel=52
					-21, 20, 4, -14, -5, -21, -25, 8, -34,
					-- layer=2 filter=181 channel=53
					-26, -29, -11, -7, -55, -26, 21, -18, -39,
					-- layer=2 filter=181 channel=54
					-10, -19, 3, 15, -17, -38, -15, 8, 12,
					-- layer=2 filter=181 channel=55
					-6, 9, -2, -2, 0, -5, -1, -8, -6,
					-- layer=2 filter=181 channel=56
					0, -21, 12, -6, -12, -20, -17, -29, -14,
					-- layer=2 filter=181 channel=57
					1, 9, -3, -9, -2, -2, 3, -9, -2,
					-- layer=2 filter=181 channel=58
					-6, 3, 4, 9, 6, -8, -12, -2, -4,
					-- layer=2 filter=181 channel=59
					27, 14, 2, 14, 18, 1, -58, -3, -45,
					-- layer=2 filter=181 channel=60
					-13, -33, -35, 16, 33, -29, -8, 42, -22,
					-- layer=2 filter=181 channel=61
					-1, -13, -22, 15, 32, 10, -7, 46, 46,
					-- layer=2 filter=181 channel=62
					-12, -37, -8, 17, -25, 12, -31, -11, -4,
					-- layer=2 filter=181 channel=63
					-15, -10, -37, -12, -25, -28, -1, 27, 7,
					-- layer=2 filter=181 channel=64
					-26, -60, -25, 5, -4, -2, 69, 34, 30,
					-- layer=2 filter=181 channel=65
					-4, 27, -27, 6, 29, 22, 2, 28, 22,
					-- layer=2 filter=181 channel=66
					1, -15, 16, -32, -37, -11, -2, -4, 14,
					-- layer=2 filter=181 channel=67
					-35, -39, -14, -9, -39, -55, 11, 19, -33,
					-- layer=2 filter=181 channel=68
					-9, -10, -10, 8, 6, -5, -10, 7, -7,
					-- layer=2 filter=181 channel=69
					-22, -17, -16, 0, -47, 0, 36, 38, 25,
					-- layer=2 filter=181 channel=70
					21, 19, 41, 13, 33, 11, 56, 16, -5,
					-- layer=2 filter=181 channel=71
					4, 25, 22, 9, 9, -4, -23, -48, -35,
					-- layer=2 filter=181 channel=72
					-1, -38, -58, -20, -31, -1, -8, -28, -14,
					-- layer=2 filter=181 channel=73
					40, 27, 15, -6, -35, -31, -38, -3, -41,
					-- layer=2 filter=181 channel=74
					-39, -14, -55, 26, -5, -75, 25, 36, -24,
					-- layer=2 filter=181 channel=75
					-21, -13, 44, 5, 1, 17, 35, -5, -30,
					-- layer=2 filter=181 channel=76
					26, -6, -31, 46, -57, -42, 1, 27, 32,
					-- layer=2 filter=181 channel=77
					0, -4, -1, 4, 8, 0, 4, -3, -7,
					-- layer=2 filter=181 channel=78
					9, -19, -16, 12, -23, -43, -33, -24, 0,
					-- layer=2 filter=181 channel=79
					8, 2, -8, 2, 4, 9, -6, -8, -7,
					-- layer=2 filter=181 channel=80
					6, -48, -35, 15, 2, -15, 31, -5, -21,
					-- layer=2 filter=181 channel=81
					-5, 2, -2, 1, 8, -3, 6, -2, -5,
					-- layer=2 filter=181 channel=82
					2, -8, -2, 4, 2, 10, 2, 1, 0,
					-- layer=2 filter=181 channel=83
					48, 40, 41, 11, 30, 22, 53, -3, 13,
					-- layer=2 filter=181 channel=84
					7, 1, 1, -11, -2, 3, 0, 5, 0,
					-- layer=2 filter=181 channel=85
					10, 0, -14, 2, 11, 11, -5, 4, -11,
					-- layer=2 filter=181 channel=86
					-6, 5, -1, 9, 14, 0, 7, 11, -1,
					-- layer=2 filter=181 channel=87
					3, -34, -36, 39, -19, -24, -15, -17, -2,
					-- layer=2 filter=181 channel=88
					-24, 20, -26, 10, -2, -23, 21, 43, 29,
					-- layer=2 filter=181 channel=89
					-29, -27, -25, 18, -13, 19, -3, -27, -27,
					-- layer=2 filter=181 channel=90
					-8, 1, -5, -7, -5, -8, 8, -9, -1,
					-- layer=2 filter=181 channel=91
					-15, -1, -4, 6, -7, 32, -42, -13, -2,
					-- layer=2 filter=181 channel=92
					-8, 25, -16, -20, 16, 35, -58, -32, -32,
					-- layer=2 filter=181 channel=93
					9, 42, 11, 46, -2, 33, -9, 1, -2,
					-- layer=2 filter=181 channel=94
					63, -42, -11, 15, -21, 43, 3, 53, 42,
					-- layer=2 filter=181 channel=95
					5, -2, 2, 15, 4, 10, 12, 13, 10,
					-- layer=2 filter=181 channel=96
					0, -56, -23, 25, 17, -67, 19, 47, -14,
					-- layer=2 filter=181 channel=97
					-3, -48, -18, 6, -7, 3, 18, 2, 4,
					-- layer=2 filter=181 channel=98
					3, -1, 6, 0, -11, -8, 26, 32, 3,
					-- layer=2 filter=181 channel=99
					29, 1, 5, -17, -6, -52, 8, 28, -36,
					-- layer=2 filter=181 channel=100
					30, 17, 14, 33, 53, 27, 14, 9, -55,
					-- layer=2 filter=181 channel=101
					-4, -17, -20, -48, -54, -57, -26, -92, -38,
					-- layer=2 filter=181 channel=102
					-23, -18, 17, 45, -27, -15, 10, 30, -13,
					-- layer=2 filter=181 channel=103
					50, 12, -21, -50, -1, 33, -5, -41, 29,
					-- layer=2 filter=181 channel=104
					-20, -40, 5, 10, -23, 8, 26, -39, 7,
					-- layer=2 filter=181 channel=105
					13, -51, -24, 1, -66, -12, 33, 9, -46,
					-- layer=2 filter=181 channel=106
					-26, -83, -40, -47, -57, -61, -14, -28, -4,
					-- layer=2 filter=181 channel=107
					-44, -43, -80, -21, -22, 20, -18, -9, 12,
					-- layer=2 filter=181 channel=108
					7, -4, 24, 13, 13, -7, -6, -37, -35,
					-- layer=2 filter=181 channel=109
					16, 3, 0, 7, -16, -3, 20, 5, 7,
					-- layer=2 filter=181 channel=110
					0, -19, -47, -75, 13, 3, 24, 49, 48,
					-- layer=2 filter=181 channel=111
					-6, 1, -7, 5, -3, -1, 3, -6, 0,
					-- layer=2 filter=181 channel=112
					-9, 12, -54, 27, 4, 1, 11, 23, 14,
					-- layer=2 filter=181 channel=113
					5, 20, -50, -1, 15, -2, 56, 26, 23,
					-- layer=2 filter=181 channel=114
					-11, 13, 7, -6, 10, -8, 3, 0, 0,
					-- layer=2 filter=181 channel=115
					0, -5, -7, -8, -5, 9, -7, -8, 9,
					-- layer=2 filter=181 channel=116
					-27, 0, -41, 35, -11, -35, -28, 14, -22,
					-- layer=2 filter=181 channel=117
					15, 27, -11, 3, -47, -54, -46, -12, 28,
					-- layer=2 filter=181 channel=118
					-22, 1, 22, -6, -10, -15, -19, -72, 4,
					-- layer=2 filter=181 channel=119
					45, 1, 60, 20, -15, 6, 2, 33, -11,
					-- layer=2 filter=181 channel=120
					4, -6, -7, -10, -4, 5, 7, -8, -8,
					-- layer=2 filter=181 channel=121
					9, -4, -7, 1, -6, -6, 10, 3, 0,
					-- layer=2 filter=181 channel=122
					7, -4, 7, 13, 10, 4, -6, -9, -5,
					-- layer=2 filter=181 channel=123
					14, 13, -33, -8, -51, -9, -11, 21, 16,
					-- layer=2 filter=181 channel=124
					11, -48, -45, 63, -52, -19, -6, -45, -12,
					-- layer=2 filter=181 channel=125
					-2, 1, -3, -4, 6, -5, 0, -4, 5,
					-- layer=2 filter=181 channel=126
					19, -22, -18, -9, 60, -85, -36, 82, -20,
					-- layer=2 filter=181 channel=127
					53, 65, 13, -7, 7, -9, 46, -2, -7,
					-- layer=2 filter=182 channel=0
					6, -36, -17, 1, -38, -28, -15, -26, -23,
					-- layer=2 filter=182 channel=1
					-16, 3, -36, -6, 4, -35, -29, -18, -29,
					-- layer=2 filter=182 channel=2
					-1, 0, -9, -4, 5, 7, -8, 10, -8,
					-- layer=2 filter=182 channel=3
					-43, -37, -7, -5, -21, 20, 13, 20, -7,
					-- layer=2 filter=182 channel=4
					-3, 26, -40, 1, -30, -22, -18, -46, -28,
					-- layer=2 filter=182 channel=5
					7, -5, -10, -33, -5, -21, -26, -14, 37,
					-- layer=2 filter=182 channel=6
					38, 30, 4, -3, 26, -31, 8, 15, -50,
					-- layer=2 filter=182 channel=7
					-24, -34, -43, 29, -24, 31, 2, -39, -67,
					-- layer=2 filter=182 channel=8
					7, 1, -4, -5, 3, -5, -10, 2, 5,
					-- layer=2 filter=182 channel=9
					-79, -41, -54, -48, -39, -40, -17, -6, -19,
					-- layer=2 filter=182 channel=10
					-60, -66, -28, -15, -46, -1, 8, -25, -22,
					-- layer=2 filter=182 channel=11
					9, 6, -11, -8, -20, 3, -29, -16, 22,
					-- layer=2 filter=182 channel=12
					-19, -22, 0, 3, -4, -20, -25, -24, 7,
					-- layer=2 filter=182 channel=13
					-7, -5, -1, 0, -8, -2, 9, -10, 8,
					-- layer=2 filter=182 channel=14
					-1, 2, -6, -2, 2, -35, -3, 7, -5,
					-- layer=2 filter=182 channel=15
					-3, 11, 68, 13, 21, 35, -24, 19, 33,
					-- layer=2 filter=182 channel=16
					3, -3, -4, 0, 10, 22, 0, 4, 22,
					-- layer=2 filter=182 channel=17
					0, -7, -7, -6, -5, 8, -8, 1, -5,
					-- layer=2 filter=182 channel=18
					18, -7, 24, 3, -32, -6, -29, 8, -33,
					-- layer=2 filter=182 channel=19
					7, 35, -26, -2, 30, -21, -26, -51, -39,
					-- layer=2 filter=182 channel=20
					-1, -2, 5, 10, -2, -2, 5, 6, -9,
					-- layer=2 filter=182 channel=21
					5, 9, 6, 0, 8, 5, -4, -1, -6,
					-- layer=2 filter=182 channel=22
					0, 7, 7, -7, 9, -4, -8, -3, 0,
					-- layer=2 filter=182 channel=23
					-58, -16, -15, -33, -39, -24, -7, -26, -27,
					-- layer=2 filter=182 channel=24
					-11, -34, 8, -2, -12, 25, 24, -10, -7,
					-- layer=2 filter=182 channel=25
					4, -17, 6, 6, -3, 15, 6, 13, 27,
					-- layer=2 filter=182 channel=26
					-1, 8, 9, 9, 3, -5, -6, 5, 2,
					-- layer=2 filter=182 channel=27
					-54, -29, -86, -32, -43, -16, -61, -39, -22,
					-- layer=2 filter=182 channel=28
					-18, 14, 11, 18, 9, -7, 2, 24, 14,
					-- layer=2 filter=182 channel=29
					0, -2, -10, -9, -9, 0, -2, 0, 7,
					-- layer=2 filter=182 channel=30
					-25, -8, -13, -20, -17, -13, 26, -12, -29,
					-- layer=2 filter=182 channel=31
					97, 39, 18, 60, 35, 37, 13, -22, 26,
					-- layer=2 filter=182 channel=32
					-6, 3, -7, 6, 2, 0, 0, -8, 6,
					-- layer=2 filter=182 channel=33
					-32, -28, 2, 9, -2, 57, -18, -30, -24,
					-- layer=2 filter=182 channel=34
					-11, 56, -30, 13, -7, 11, 18, 8, -19,
					-- layer=2 filter=182 channel=35
					-39, 0, -9, -4, -58, -20, 17, -18, 2,
					-- layer=2 filter=182 channel=36
					3, 2, 4, 0, -1, -4, -1, 0, -6,
					-- layer=2 filter=182 channel=37
					3, 15, -16, -32, 0, 2, -26, 8, 21,
					-- layer=2 filter=182 channel=38
					-11, -13, -35, -33, -15, 2, -9, -11, -25,
					-- layer=2 filter=182 channel=39
					-76, -38, 2, 11, 2, 13, 17, -27, -46,
					-- layer=2 filter=182 channel=40
					18, 18, 37, 46, 4, 34, 16, 71, 14,
					-- layer=2 filter=182 channel=41
					-10, -2, -7, 5, -5, -9, -8, -1, 2,
					-- layer=2 filter=182 channel=42
					-20, -34, 28, -9, 5, -19, 15, 10, 10,
					-- layer=2 filter=182 channel=43
					-30, -22, 7, -15, -51, 30, -49, -13, 9,
					-- layer=2 filter=182 channel=44
					1, 3, 10, -4, -8, 0, -6, 0, -6,
					-- layer=2 filter=182 channel=45
					27, -13, -20, 18, 0, 25, -31, -63, -22,
					-- layer=2 filter=182 channel=46
					1, -49, -28, 9, -10, -18, -2, -47, -4,
					-- layer=2 filter=182 channel=47
					-45, -31, -21, 15, -20, 24, -11, 2, -9,
					-- layer=2 filter=182 channel=48
					-2, 5, 4, -6, 10, -9, -9, -5, -3,
					-- layer=2 filter=182 channel=49
					50, -25, 33, 18, 2, -8, 0, -4, 0,
					-- layer=2 filter=182 channel=50
					-8, -7, -14, -8, -13, -9, -4, -2, -12,
					-- layer=2 filter=182 channel=51
					14, -11, -42, -24, 0, -28, -6, -18, -6,
					-- layer=2 filter=182 channel=52
					7, 20, -36, 1, -4, -10, -33, -2, -8,
					-- layer=2 filter=182 channel=53
					37, -44, 19, 32, 29, 2, 24, 8, -37,
					-- layer=2 filter=182 channel=54
					10, 0, 0, 27, 2, 5, -11, -18, 10,
					-- layer=2 filter=182 channel=55
					-1, -3, 8, 0, -5, 8, 6, -9, 10,
					-- layer=2 filter=182 channel=56
					21, -4, -10, -18, -36, -6, -49, -3, 16,
					-- layer=2 filter=182 channel=57
					3, 10, -2, 7, -4, 9, 0, 5, -9,
					-- layer=2 filter=182 channel=58
					-18, -31, -9, -18, 10, -24, -3, -32, 6,
					-- layer=2 filter=182 channel=59
					4, -35, 1, -21, 10, 1, -25, -34, -25,
					-- layer=2 filter=182 channel=60
					-11, 57, -9, 3, 26, -77, -7, 9, -14,
					-- layer=2 filter=182 channel=61
					-14, -26, 9, 13, -11, -44, -1, -3, -72,
					-- layer=2 filter=182 channel=62
					46, 54, -13, -9, 21, 1, 0, -1, -21,
					-- layer=2 filter=182 channel=63
					-51, -36, 5, -24, -20, -19, -4, -28, -32,
					-- layer=2 filter=182 channel=64
					-58, -17, -1, -37, -59, 1, 5, 0, -8,
					-- layer=2 filter=182 channel=65
					18, 28, -14, -12, 9, -64, -20, -5, -77,
					-- layer=2 filter=182 channel=66
					1, -15, 43, -3, 49, -2, 19, 27, 2,
					-- layer=2 filter=182 channel=67
					-46, -49, -71, -24, -21, -18, -12, -25, -10,
					-- layer=2 filter=182 channel=68
					2, -3, 0, 3, 7, 7, 6, 3, -11,
					-- layer=2 filter=182 channel=69
					-59, -10, -18, -33, -29, -54, -1, -14, -12,
					-- layer=2 filter=182 channel=70
					-21, 0, 20, -10, -29, -29, 1, -8, -3,
					-- layer=2 filter=182 channel=71
					-25, -26, -37, 1, -31, -6, -22, -17, -29,
					-- layer=2 filter=182 channel=72
					-45, -20, 12, 9, 16, -2, -10, 24, -28,
					-- layer=2 filter=182 channel=73
					21, 6, 0, 25, 28, 53, -7, -28, -32,
					-- layer=2 filter=182 channel=74
					-54, -36, -7, -18, -35, -6, 38, -1, 7,
					-- layer=2 filter=182 channel=75
					36, 7, 10, 17, 43, -28, 11, 31, 7,
					-- layer=2 filter=182 channel=76
					17, -19, -11, 18, 31, -4, 22, -16, 12,
					-- layer=2 filter=182 channel=77
					1, 7, -7, -10, 4, -10, -3, -12, 5,
					-- layer=2 filter=182 channel=78
					17, 3, -3, -21, -3, 10, -22, 9, 8,
					-- layer=2 filter=182 channel=79
					1, -4, 1, 10, -9, -8, 9, -8, -9,
					-- layer=2 filter=182 channel=80
					1, -33, -25, -8, -11, -5, -9, -4, 14,
					-- layer=2 filter=182 channel=81
					-1, 7, 8, -5, 0, 5, -2, -5, 0,
					-- layer=2 filter=182 channel=82
					-1, -4, 9, 7, -8, 11, -10, 5, -9,
					-- layer=2 filter=182 channel=83
					-23, -58, -34, -24, -14, -63, 0, -27, -36,
					-- layer=2 filter=182 channel=84
					2, 0, 4, -5, 10, 9, -2, -7, 0,
					-- layer=2 filter=182 channel=85
					0, -1, 2, 0, 2, 5, -10, -5, -4,
					-- layer=2 filter=182 channel=86
					-1, -6, 7, 4, 0, 6, -4, 0, -2,
					-- layer=2 filter=182 channel=87
					-5, 22, 15, 35, -27, 11, -4, 33, -16,
					-- layer=2 filter=182 channel=88
					-50, -52, -16, -35, -44, -27, -10, -35, -20,
					-- layer=2 filter=182 channel=89
					-12, -17, -9, -16, 16, -47, -16, -11, -22,
					-- layer=2 filter=182 channel=90
					-6, 9, 10, 1, -4, 1, 4, 3, -8,
					-- layer=2 filter=182 channel=91
					-39, 8, 10, -2, 15, 1, -3, 29, 31,
					-- layer=2 filter=182 channel=92
					-32, -13, -18, -3, -11, -42, -12, -7, -37,
					-- layer=2 filter=182 channel=93
					47, 86, -38, -1, 53, -35, -6, 14, -12,
					-- layer=2 filter=182 channel=94
					6, -24, 5, 2, -30, -25, 16, 15, -71,
					-- layer=2 filter=182 channel=95
					6, 0, -4, -4, 3, 3, -2, -6, 2,
					-- layer=2 filter=182 channel=96
					10, -5, -17, -1, 4, -31, -34, -8, -18,
					-- layer=2 filter=182 channel=97
					-26, -7, 5, 0, -20, 36, -14, -10, -9,
					-- layer=2 filter=182 channel=98
					-26, -6, -22, 4, -18, 21, -9, 20, -9,
					-- layer=2 filter=182 channel=99
					12, 29, -18, -18, 27, -2, -24, 10, -14,
					-- layer=2 filter=182 channel=100
					5, 0, -3, -17, 19, 18, 2, -21, 5,
					-- layer=2 filter=182 channel=101
					-5, -40, -50, 7, -56, 2, 16, 1, 7,
					-- layer=2 filter=182 channel=102
					5, 28, -15, -26, -37, -40, -23, -4, -36,
					-- layer=2 filter=182 channel=103
					-35, 13, 1, 0, -16, 12, -69, -13, 10,
					-- layer=2 filter=182 channel=104
					27, -31, 14, 7, 11, -12, 1, -5, -23,
					-- layer=2 filter=182 channel=105
					11, -3, -73, 9, -37, -37, 21, 47, 35,
					-- layer=2 filter=182 channel=106
					5, -18, -6, -5, -10, 1, 35, -4, 5,
					-- layer=2 filter=182 channel=107
					20, 46, -2, -29, 37, -8, -12, 3, -35,
					-- layer=2 filter=182 channel=108
					-12, 2, -55, -12, -18, -61, -20, -4, -74,
					-- layer=2 filter=182 channel=109
					3, -5, 6, -3, -1, 7, 9, 3, -2,
					-- layer=2 filter=182 channel=110
					-41, 3, 24, -19, -12, 19, -9, -11, -22,
					-- layer=2 filter=182 channel=111
					-3, -1, 7, -11, -11, -10, 3, -2, 0,
					-- layer=2 filter=182 channel=112
					-24, -27, -6, 10, -25, -36, 0, -22, -76,
					-- layer=2 filter=182 channel=113
					-40, -22, -25, -16, 2, -30, -7, -12, -70,
					-- layer=2 filter=182 channel=114
					2, 0, -6, 8, 9, -8, 13, 5, 7,
					-- layer=2 filter=182 channel=115
					-6, -8, -3, 2, -8, -3, 9, 2, 0,
					-- layer=2 filter=182 channel=116
					-21, 26, 29, 16, -20, 10, -11, 51, -32,
					-- layer=2 filter=182 channel=117
					10, -24, -20, 43, 32, 12, -40, -22, -32,
					-- layer=2 filter=182 channel=118
					-32, -49, -14, -14, -36, -3, -53, -14, -7,
					-- layer=2 filter=182 channel=119
					-17, 0, 23, -8, 4, 0, -27, -22, -19,
					-- layer=2 filter=182 channel=120
					5, -1, 1, 1, -6, 0, 8, 6, 9,
					-- layer=2 filter=182 channel=121
					7, -6, -9, -9, 4, 5, 8, 2, -9,
					-- layer=2 filter=182 channel=122
					-1, 8, -9, 7, -2, 1, -6, 1, -5,
					-- layer=2 filter=182 channel=123
					-33, -35, -13, 4, 17, 30, 0, -17, -9,
					-- layer=2 filter=182 channel=124
					38, 0, 43, 0, 12, 34, 5, -11, 14,
					-- layer=2 filter=182 channel=125
					-6, -6, -6, -7, -5, 4, -8, 0, -1,
					-- layer=2 filter=182 channel=126
					11, 2, 42, 25, 19, -11, -19, 38, -39,
					-- layer=2 filter=182 channel=127
					-21, 17, -33, -20, 10, -48, -7, -10, -60,
					-- layer=2 filter=183 channel=0
					-9, -4, 6, -15, -5, -1, -25, -16, 4,
					-- layer=2 filter=183 channel=1
					-25, -28, -20, -17, -20, -8, 1, -24, -13,
					-- layer=2 filter=183 channel=2
					-10, 10, 0, 7, -8, -4, 8, 9, -5,
					-- layer=2 filter=183 channel=3
					10, -7, -1, -34, -30, -14, -24, -38, 0,
					-- layer=2 filter=183 channel=4
					-31, 10, -7, 7, 17, -39, -8, -6, -31,
					-- layer=2 filter=183 channel=5
					9, 18, 10, 2, 22, 32, 21, 24, 26,
					-- layer=2 filter=183 channel=6
					0, -21, 3, 0, 25, -1, 18, -26, 10,
					-- layer=2 filter=183 channel=7
					-13, -7, -1, -27, -26, -16, -18, -12, 21,
					-- layer=2 filter=183 channel=8
					-8, 4, 1, -3, 0, 2, 2, -5, -6,
					-- layer=2 filter=183 channel=9
					5, -25, -20, -25, -9, -37, -26, -23, -32,
					-- layer=2 filter=183 channel=10
					-1, 3, -13, -24, 0, -16, -27, 2, 5,
					-- layer=2 filter=183 channel=11
					-12, -1, -2, 0, 17, 3, 14, -12, -18,
					-- layer=2 filter=183 channel=12
					-33, -13, 1, -31, -23, 5, 1, -15, -12,
					-- layer=2 filter=183 channel=13
					-1, 1, 10, -3, 3, -6, -1, 7, 3,
					-- layer=2 filter=183 channel=14
					-49, -28, -19, -20, -27, -10, -2, -35, -11,
					-- layer=2 filter=183 channel=15
					-3, 13, -2, -10, -36, -14, 2, -40, -6,
					-- layer=2 filter=183 channel=16
					-20, -7, -4, 5, -24, -15, -8, 4, 1,
					-- layer=2 filter=183 channel=17
					6, -6, 1, 9, -9, 4, 3, -2, 8,
					-- layer=2 filter=183 channel=18
					-24, 6, -41, 32, 17, -24, 12, 12, -35,
					-- layer=2 filter=183 channel=19
					2, -10, -25, -13, 0, -13, -19, -17, -13,
					-- layer=2 filter=183 channel=20
					-7, -6, -1, -9, 0, -7, 1, 3, -8,
					-- layer=2 filter=183 channel=21
					7, -6, 2, 4, 9, -4, 5, 5, -7,
					-- layer=2 filter=183 channel=22
					-6, 0, 4, 2, -7, 0, 2, 3, -9,
					-- layer=2 filter=183 channel=23
					-38, -8, -6, -1, 11, 1, -13, 9, 16,
					-- layer=2 filter=183 channel=24
					9, -17, -31, -1, -31, -6, -23, -13, -8,
					-- layer=2 filter=183 channel=25
					16, -21, -22, -6, -33, -4, -25, -9, -7,
					-- layer=2 filter=183 channel=26
					4, -2, -2, 1, -5, -9, 1, 3, 2,
					-- layer=2 filter=183 channel=27
					3, 4, 2, 8, 15, 7, 22, 5, -4,
					-- layer=2 filter=183 channel=28
					-23, 5, -19, -26, -6, 6, -18, -4, 1,
					-- layer=2 filter=183 channel=29
					6, 0, 5, -5, 2, 0, 6, 5, 0,
					-- layer=2 filter=183 channel=30
					0, -10, 23, -15, 0, -2, 12, 11, -33,
					-- layer=2 filter=183 channel=31
					15, -27, -2, 15, -3, -12, 1, -7, -18,
					-- layer=2 filter=183 channel=32
					4, -6, 6, -6, 8, 9, 0, 1, 0,
					-- layer=2 filter=183 channel=33
					-21, -5, 9, 3, -18, 5, 10, -4, -18,
					-- layer=2 filter=183 channel=34
					-29, 25, -66, 11, -10, -22, 36, 18, -31,
					-- layer=2 filter=183 channel=35
					-6, 12, -17, -2, -15, 5, 4, -27, -5,
					-- layer=2 filter=183 channel=36
					3, -4, -8, 6, 6, 0, -2, -10, 7,
					-- layer=2 filter=183 channel=37
					11, -9, -2, -1, 19, 7, 18, 17, -7,
					-- layer=2 filter=183 channel=38
					-16, -15, 31, -32, 19, 2, 13, -2, -16,
					-- layer=2 filter=183 channel=39
					-45, -18, 1, 1, -29, -23, 0, 13, 29,
					-- layer=2 filter=183 channel=40
					14, 33, -35, 8, 13, -45, 28, -11, -5,
					-- layer=2 filter=183 channel=41
					5, 7, 3, 6, -5, 3, -8, -3, 0,
					-- layer=2 filter=183 channel=42
					-17, -21, -7, -23, 14, -12, 3, 6, 5,
					-- layer=2 filter=183 channel=43
					-1, 7, -21, 15, -16, -18, 11, -38, -10,
					-- layer=2 filter=183 channel=44
					-9, -8, 0, 1, 3, 6, 9, 5, -9,
					-- layer=2 filter=183 channel=45
					15, -1, 19, 0, -29, 15, 5, -36, -6,
					-- layer=2 filter=183 channel=46
					0, -21, -27, -6, -26, -28, -41, -18, -16,
					-- layer=2 filter=183 channel=47
					-1, 8, -24, -19, -18, -9, -3, -5, 2,
					-- layer=2 filter=183 channel=48
					3, 1, 3, 2, -8, 6, 0, -7, -9,
					-- layer=2 filter=183 channel=49
					-11, -5, -48, 12, -15, -35, 3, -18, -14,
					-- layer=2 filter=183 channel=50
					6, 3, 0, 1, 2, 3, 8, 1, 7,
					-- layer=2 filter=183 channel=51
					4, -19, 9, -10, 0, 9, -7, -18, -5,
					-- layer=2 filter=183 channel=52
					1, 3, 10, -4, 2, -5, 0, -7, 0,
					-- layer=2 filter=183 channel=53
					9, 7, -24, -34, -29, -32, 8, -21, -32,
					-- layer=2 filter=183 channel=54
					-22, 8, -15, -9, -8, -20, 7, -18, -6,
					-- layer=2 filter=183 channel=55
					0, -2, -10, 2, 1, 5, 2, 1, 4,
					-- layer=2 filter=183 channel=56
					1, 11, 7, 21, 11, 1, 14, -2, 9,
					-- layer=2 filter=183 channel=57
					0, 4, 0, -7, -5, -5, -3, 8, 3,
					-- layer=2 filter=183 channel=58
					-19, -22, 24, 3, -7, 3, 9, -20, -20,
					-- layer=2 filter=183 channel=59
					-5, -31, 32, 1, -41, -2, 1, 15, -2,
					-- layer=2 filter=183 channel=60
					-10, -19, 8, -18, 15, -2, 1, -28, -2,
					-- layer=2 filter=183 channel=61
					-24, -16, 12, -17, 4, 10, -33, -19, 3,
					-- layer=2 filter=183 channel=62
					0, -14, -11, 6, 13, -13, 30, -19, 7,
					-- layer=2 filter=183 channel=63
					-28, -5, 4, -16, 1, -3, -31, 0, 31,
					-- layer=2 filter=183 channel=64
					18, -3, -21, 5, -11, -13, -15, -1, -19,
					-- layer=2 filter=183 channel=65
					-11, -29, 20, -24, 18, 8, 2, -11, -2,
					-- layer=2 filter=183 channel=66
					14, 8, 7, -5, -9, -14, -18, 14, 22,
					-- layer=2 filter=183 channel=67
					0, 0, -5, -8, -7, 6, -23, -6, -25,
					-- layer=2 filter=183 channel=68
					4, 0, -4, 6, 5, 9, 11, 6, -8,
					-- layer=2 filter=183 channel=69
					-12, -1, -13, -8, 5, -11, 26, 3, 8,
					-- layer=2 filter=183 channel=70
					-18, 12, 10, -11, 0, 1, 9, -22, 5,
					-- layer=2 filter=183 channel=71
					1, 1, -24, 1, -25, -5, -13, -20, -17,
					-- layer=2 filter=183 channel=72
					-11, 3, -17, -31, -18, -7, -20, 4, 14,
					-- layer=2 filter=183 channel=73
					18, -4, -26, -11, -37, -16, -2, -50, -28,
					-- layer=2 filter=183 channel=74
					-7, 7, 18, -9, 0, 1, -23, 10, -11,
					-- layer=2 filter=183 channel=75
					-42, -13, -17, -17, -20, 14, 1, -14, 16,
					-- layer=2 filter=183 channel=76
					0, 27, 0, -16, -18, -20, 6, -31, -10,
					-- layer=2 filter=183 channel=77
					2, 0, -4, 9, -8, -7, -4, -4, 5,
					-- layer=2 filter=183 channel=78
					-2, -22, -27, -18, 7, -15, -26, -21, -8,
					-- layer=2 filter=183 channel=79
					-8, 0, -11, -3, -2, -8, -10, 5, -10,
					-- layer=2 filter=183 channel=80
					-24, -7, -26, 6, 9, -24, 10, -19, -18,
					-- layer=2 filter=183 channel=81
					3, 0, 0, -8, -7, 3, -5, -9, -13,
					-- layer=2 filter=183 channel=82
					8, -5, -8, 1, -2, -2, 3, 7, -3,
					-- layer=2 filter=183 channel=83
					-48, -19, 1, -15, 34, 32, -18, 15, 17,
					-- layer=2 filter=183 channel=84
					8, 1, 0, 5, -3, 3, -8, -10, 9,
					-- layer=2 filter=183 channel=85
					4, -5, -6, 0, 5, 4, -2, 7, 1,
					-- layer=2 filter=183 channel=86
					-3, 6, 7, 6, 0, -11, 8, -4, 5,
					-- layer=2 filter=183 channel=87
					-46, 20, 1, 25, -14, -17, -25, -12, -13,
					-- layer=2 filter=183 channel=88
					-15, 0, 25, -25, 6, 10, -25, -10, -1,
					-- layer=2 filter=183 channel=89
					-34, -18, 18, -13, -30, -19, 4, -12, -6,
					-- layer=2 filter=183 channel=90
					2, -7, -9, 0, 10, 0, 3, 1, -4,
					-- layer=2 filter=183 channel=91
					-30, -29, -16, -23, -32, 16, 4, -25, -13,
					-- layer=2 filter=183 channel=92
					-39, -43, 6, -6, -36, 2, 0, -5, -7,
					-- layer=2 filter=183 channel=93
					-3, -14, -9, -18, 7, -16, 29, -19, -5,
					-- layer=2 filter=183 channel=94
					-32, -3, 0, -24, 0, 5, -21, -11, 14,
					-- layer=2 filter=183 channel=95
					11, -5, 6, 1, -3, 5, 0, -1, -2,
					-- layer=2 filter=183 channel=96
					-38, 53, -4, -14, 2, -28, -42, 3, 11,
					-- layer=2 filter=183 channel=97
					9, -48, -11, -3, -15, -27, -9, -40, -33,
					-- layer=2 filter=183 channel=98
					0, -7, -34, -8, -3, -10, -18, -11, -10,
					-- layer=2 filter=183 channel=99
					17, -13, -22, -43, -24, 6, -23, -11, -19,
					-- layer=2 filter=183 channel=100
					-14, 17, 5, -15, 34, 30, 51, -16, -25,
					-- layer=2 filter=183 channel=101
					-7, -31, -26, -20, -40, -9, -36, -45, -4,
					-- layer=2 filter=183 channel=102
					-8, 33, -34, 17, 32, -39, -3, 3, -3,
					-- layer=2 filter=183 channel=103
					-2, -11, 6, 18, 7, -13, 9, 7, 0,
					-- layer=2 filter=183 channel=104
					-22, -17, -17, -1, -6, -31, -10, -10, 1,
					-- layer=2 filter=183 channel=105
					0, -10, 22, 4, -17, -8, -18, -34, 16,
					-- layer=2 filter=183 channel=106
					-1, -21, -11, -16, -32, 15, -7, -23, -7,
					-- layer=2 filter=183 channel=107
					-3, -22, 0, 12, -35, -21, -13, 6, 7,
					-- layer=2 filter=183 channel=108
					-32, 5, -34, -15, -3, -27, 1, 17, 8,
					-- layer=2 filter=183 channel=109
					4, -9, 0, -7, 5, 0, -5, 6, 0,
					-- layer=2 filter=183 channel=110
					-11, -30, -53, -25, -34, -30, -27, -12, -16,
					-- layer=2 filter=183 channel=111
					9, -9, 8, 3, 5, 5, -1, 2, 7,
					-- layer=2 filter=183 channel=112
					-5, -36, -4, -11, -17, 5, -9, -2, 0,
					-- layer=2 filter=183 channel=113
					3, -33, 17, -21, 2, -3, -22, 19, -11,
					-- layer=2 filter=183 channel=114
					-10, -1, -11, 10, -5, -7, 3, 7, 0,
					-- layer=2 filter=183 channel=115
					1, -6, -9, 3, 4, 7, -6, 2, -4,
					-- layer=2 filter=183 channel=116
					-16, 39, -23, 22, 1, -18, -25, -36, -4,
					-- layer=2 filter=183 channel=117
					4, 14, -26, -42, -36, -39, -41, -34, -37,
					-- layer=2 filter=183 channel=118
					-1, -14, -35, -5, -29, -16, -7, -23, -41,
					-- layer=2 filter=183 channel=119
					-31, 19, -17, 30, -13, 21, 32, 0, -16,
					-- layer=2 filter=183 channel=120
					0, 8, 7, 4, 3, -7, -3, 0, -4,
					-- layer=2 filter=183 channel=121
					5, -5, 0, 5, 9, 6, -5, -2, 4,
					-- layer=2 filter=183 channel=122
					-2, -1, 2, 7, -5, -1, 3, -2, -1,
					-- layer=2 filter=183 channel=123
					-5, -3, 4, -7, -18, -13, -16, -13, 15,
					-- layer=2 filter=183 channel=124
					-2, -15, 8, 8, -30, -2, -11, -51, -35,
					-- layer=2 filter=183 channel=125
					-7, 3, 2, -8, 4, 0, 4, -7, -5,
					-- layer=2 filter=183 channel=126
					-21, 5, 3, -18, -12, -20, -19, -12, -9,
					-- layer=2 filter=183 channel=127
					-29, -24, 24, -41, 7, 13, 21, 6, -15,
					-- layer=2 filter=184 channel=0
					37, 9, 8, -2, -3, 1, 2, 18, 12,
					-- layer=2 filter=184 channel=1
					-37, -13, 16, -16, -36, -31, -30, -35, -55,
					-- layer=2 filter=184 channel=2
					8, -7, 5, -2, -12, -7, -9, -1, 10,
					-- layer=2 filter=184 channel=3
					22, -21, 1, -1, -8, -36, -10, -7, 19,
					-- layer=2 filter=184 channel=4
					-16, -4, -17, -3, -13, -18, -17, -10, -12,
					-- layer=2 filter=184 channel=5
					30, 14, -37, -11, -26, 39, 16, -16, -11,
					-- layer=2 filter=184 channel=6
					23, 52, -15, 31, 70, 27, 56, 7, 58,
					-- layer=2 filter=184 channel=7
					-22, 0, 54, 6, -25, -4, 10, 7, 20,
					-- layer=2 filter=184 channel=8
					5, 9, -3, 2, -8, -10, -3, 7, -3,
					-- layer=2 filter=184 channel=9
					7, -13, -14, 2, -21, -27, -17, -20, -28,
					-- layer=2 filter=184 channel=10
					23, -22, 1, -17, -14, 3, 19, 9, -5,
					-- layer=2 filter=184 channel=11
					2, 0, 11, 6, -1, 2, 18, 8, 11,
					-- layer=2 filter=184 channel=12
					-16, 6, 21, 1, -11, -23, -26, -52, -40,
					-- layer=2 filter=184 channel=13
					2, -1, 7, 4, 7, 3, -1, 8, 9,
					-- layer=2 filter=184 channel=14
					3, -15, 35, -20, -31, -27, -1, -18, -30,
					-- layer=2 filter=184 channel=15
					-40, -37, -43, 80, -8, -8, -1, -49, -33,
					-- layer=2 filter=184 channel=16
					-18, 1, 4, -15, 15, 0, -28, -1, -14,
					-- layer=2 filter=184 channel=17
					-5, 5, 10, -5, -9, -6, 5, -11, -4,
					-- layer=2 filter=184 channel=18
					-10, 55, 9, -17, 8, -4, -26, 3, -17,
					-- layer=2 filter=184 channel=19
					1, 8, -7, -10, -40, -16, 22, -8, -65,
					-- layer=2 filter=184 channel=20
					2, 4, 0, -1, 7, 1, -8, -3, 2,
					-- layer=2 filter=184 channel=21
					-15, 11, -7, -5, -16, -9, -20, -5, -13,
					-- layer=2 filter=184 channel=22
					1, 0, -8, -4, 2, 1, 9, 0, -11,
					-- layer=2 filter=184 channel=23
					-27, 8, -15, 16, 0, 20, -11, -16, 11,
					-- layer=2 filter=184 channel=24
					48, 8, 24, 21, 1, 5, 20, -5, -22,
					-- layer=2 filter=184 channel=25
					34, 5, 26, 21, 12, -11, 22, 1, -13,
					-- layer=2 filter=184 channel=26
					0, 5, 1, -2, 4, 6, -2, 5, -5,
					-- layer=2 filter=184 channel=27
					79, 16, -2, 17, -7, 7, 23, -10, -38,
					-- layer=2 filter=184 channel=28
					30, -20, 0, 20, 12, -12, -15, -11, 15,
					-- layer=2 filter=184 channel=29
					8, 2, -4, 0, 0, -5, -8, -3, -4,
					-- layer=2 filter=184 channel=30
					-11, -5, -20, -11, -10, 18, -34, -13, -15,
					-- layer=2 filter=184 channel=31
					33, 22, -40, 102, -8, 20, 20, 12, 58,
					-- layer=2 filter=184 channel=32
					9, 4, -1, -11, -9, 2, -3, -1, -2,
					-- layer=2 filter=184 channel=33
					6, -13, 31, 16, -23, -28, 79, 2, -14,
					-- layer=2 filter=184 channel=34
					-32, 44, 19, -35, 31, 2, -6, -11, -36,
					-- layer=2 filter=184 channel=35
					31, 21, -27, 26, 7, -17, -12, -33, -15,
					-- layer=2 filter=184 channel=36
					-19, -3, -12, -3, -11, 7, -17, -3, -8,
					-- layer=2 filter=184 channel=37
					2, 0, 11, -6, -3, 9, 11, 12, -7,
					-- layer=2 filter=184 channel=38
					35, 11, -32, 19, -32, -4, 40, -21, -35,
					-- layer=2 filter=184 channel=39
					-17, -10, -20, 16, 14, -5, 2, -14, -8,
					-- layer=2 filter=184 channel=40
					-23, 25, -21, 11, -5, 61, -2, 24, -14,
					-- layer=2 filter=184 channel=41
					7, 0, -3, -7, -7, -5, 3, -3, -1,
					-- layer=2 filter=184 channel=42
					2, 16, 1, 28, 14, 28, 0, 5, -4,
					-- layer=2 filter=184 channel=43
					37, 0, -22, -6, -13, -40, -26, -40, -34,
					-- layer=2 filter=184 channel=44
					-8, 2, -4, 7, 0, -8, 3, -3, -11,
					-- layer=2 filter=184 channel=45
					25, 0, 3, 27, -16, -16, -5, -19, -20,
					-- layer=2 filter=184 channel=46
					-6, -3, 4, -19, -29, 2, -18, 12, -12,
					-- layer=2 filter=184 channel=47
					0, -52, 47, 2, 12, 13, 45, 4, 4,
					-- layer=2 filter=184 channel=48
					9, 2, 3, -9, 4, -6, -8, 3, -9,
					-- layer=2 filter=184 channel=49
					0, 33, 26, -35, 51, 21, -15, 35, 22,
					-- layer=2 filter=184 channel=50
					-19, -8, 1, -8, 0, -14, 15, -11, -15,
					-- layer=2 filter=184 channel=51
					-1, -11, 0, 11, 15, 0, 14, 0, -3,
					-- layer=2 filter=184 channel=52
					-53, 12, 28, -3, -6, -1, 29, 5, -23,
					-- layer=2 filter=184 channel=53
					44, 22, 3, 20, -17, -7, 24, -5, -3,
					-- layer=2 filter=184 channel=54
					-8, -11, -17, -11, -1, 11, 35, 1, 16,
					-- layer=2 filter=184 channel=55
					9, 10, 5, 7, 0, 4, -3, 1, -1,
					-- layer=2 filter=184 channel=56
					22, 7, 12, 1, 11, 15, 0, 10, 5,
					-- layer=2 filter=184 channel=57
					5, 6, 2, -3, -10, -6, -1, -16, 1,
					-- layer=2 filter=184 channel=58
					-1, 5, 20, 17, -11, -23, -16, -64, -5,
					-- layer=2 filter=184 channel=59
					20, 44, -29, 5, -6, -54, 0, -89, -50,
					-- layer=2 filter=184 channel=60
					17, 23, -17, -28, -32, -4, -32, -69, -10,
					-- layer=2 filter=184 channel=61
					9, 26, -12, -36, 9, -12, 0, 1, -21,
					-- layer=2 filter=184 channel=62
					-23, 57, 2, 12, 35, 0, 21, -11, 37,
					-- layer=2 filter=184 channel=63
					-16, 0, 10, -13, -1, 11, 9, -8, -8,
					-- layer=2 filter=184 channel=64
					-5, -19, 0, 22, 15, 29, -5, 5, 16,
					-- layer=2 filter=184 channel=65
					8, 12, -33, -33, 15, 17, 13, -4, 16,
					-- layer=2 filter=184 channel=66
					40, -12, 16, 4, -24, -4, -14, 30, -25,
					-- layer=2 filter=184 channel=67
					-36, 8, 14, -13, -38, -34, -45, -45, -60,
					-- layer=2 filter=184 channel=68
					-9, 1, -4, -11, -5, -2, -6, 2, 10,
					-- layer=2 filter=184 channel=69
					-23, -13, 16, 0, 16, -5, -14, 31, 30,
					-- layer=2 filter=184 channel=70
					24, -6, -41, 16, 3, 13, -11, -23, 0,
					-- layer=2 filter=184 channel=71
					10, -15, -14, -2, -26, -34, -5, -13, -31,
					-- layer=2 filter=184 channel=72
					1, -18, 20, -2, -30, -24, 21, -22, -18,
					-- layer=2 filter=184 channel=73
					15, 0, 23, -1, -31, -14, 10, -15, 6,
					-- layer=2 filter=184 channel=74
					-13, 20, 7, 41, -38, -33, 10, 9, -23,
					-- layer=2 filter=184 channel=75
					-13, -8, 31, 11, 18, 16, -2, -13, 26,
					-- layer=2 filter=184 channel=76
					6, -40, -4, 35, -5, 1, 57, 13, -5,
					-- layer=2 filter=184 channel=77
					-5, 0, -11, 7, 7, 9, 4, 1, 2,
					-- layer=2 filter=184 channel=78
					6, 10, 4, 1, 5, 0, 25, -3, 18,
					-- layer=2 filter=184 channel=79
					3, -7, 7, 2, 4, 11, -11, 11, 7,
					-- layer=2 filter=184 channel=80
					-24, -20, 0, -18, 1, -6, -7, 9, 5,
					-- layer=2 filter=184 channel=81
					-12, 0, -13, -4, 12, -18, -6, 0, 0,
					-- layer=2 filter=184 channel=82
					3, 5, 3, -8, -1, -6, -3, 1, 0,
					-- layer=2 filter=184 channel=83
					11, -2, -21, 23, 43, 49, -25, 0, 1,
					-- layer=2 filter=184 channel=84
					8, 0, 6, -2, -5, 5, -1, -4, -1,
					-- layer=2 filter=184 channel=85
					-1, -9, -18, -1, -2, -3, 0, 7, 4,
					-- layer=2 filter=184 channel=86
					-2, 4, 5, 21, 8, 1, 7, 15, -3,
					-- layer=2 filter=184 channel=87
					-12, 47, -10, 5, -5, 17, -17, 7, -12,
					-- layer=2 filter=184 channel=88
					-21, -9, 13, -4, -37, 8, -30, -8, 0,
					-- layer=2 filter=184 channel=89
					-4, 4, 29, -14, -35, -18, -23, -78, -62,
					-- layer=2 filter=184 channel=90
					0, 4, -8, -2, 9, 9, -9, -7, 9,
					-- layer=2 filter=184 channel=91
					8, 23, -2, 27, -6, 2, -12, -53, -19,
					-- layer=2 filter=184 channel=92
					-3, -18, 20, 8, -3, -9, -19, -53, -25,
					-- layer=2 filter=184 channel=93
					-21, 8, -24, -37, -23, 0, 14, 11, 22,
					-- layer=2 filter=184 channel=94
					-11, 51, -32, -38, 2, 27, 32, 15, -18,
					-- layer=2 filter=184 channel=95
					1, -7, -9, -2, 0, -7, -4, 1, -18,
					-- layer=2 filter=184 channel=96
					5, 60, 18, 19, 42, 40, 16, 24, 33,
					-- layer=2 filter=184 channel=97
					-1, -3, 51, -2, 10, -13, 3, 0, 17,
					-- layer=2 filter=184 channel=98
					-10, -38, 6, 8, -3, 29, -4, 27, 5,
					-- layer=2 filter=184 channel=99
					-13, 12, -21, 11, 1, 12, 32, 18, -32,
					-- layer=2 filter=184 channel=100
					17, 15, -28, 28, 11, 39, -26, -47, -34,
					-- layer=2 filter=184 channel=101
					22, -35, 25, -3, -31, -26, 0, -39, -39,
					-- layer=2 filter=184 channel=102
					-2, 40, -6, -3, 11, -28, -1, -10, 14,
					-- layer=2 filter=184 channel=103
					-36, -3, -15, 9, -9, -6, 12, 42, 5,
					-- layer=2 filter=184 channel=104
					21, 55, 13, 27, 14, 12, 1, 27, 24,
					-- layer=2 filter=184 channel=105
					-28, -8, 32, -4, -34, -1, -11, -9, 51,
					-- layer=2 filter=184 channel=106
					7, 0, 30, 39, -31, -26, 29, -31, -46,
					-- layer=2 filter=184 channel=107
					-28, 19, 29, 6, -36, 1, 13, -28, -39,
					-- layer=2 filter=184 channel=108
					12, 29, 2, 0, 0, -20, -4, -10, -34,
					-- layer=2 filter=184 channel=109
					-7, -4, -12, 0, 15, 14, 0, -4, 7,
					-- layer=2 filter=184 channel=110
					8, 9, 29, 24, 6, 50, -17, -13, 15,
					-- layer=2 filter=184 channel=111
					5, 1, 0, 3, -8, 3, 7, 4, 5,
					-- layer=2 filter=184 channel=112
					28, 8, -14, -14, -6, 16, -15, 0, -1,
					-- layer=2 filter=184 channel=113
					14, -31, -2, -31, 5, 20, -31, 2, 7,
					-- layer=2 filter=184 channel=114
					-8, -6, 0, 10, 8, -5, 2, 7, 17,
					-- layer=2 filter=184 channel=115
					3, 6, 8, 6, 4, 4, -2, -8, 3,
					-- layer=2 filter=184 channel=116
					-6, 24, -18, 0, -29, -20, -44, -8, -9,
					-- layer=2 filter=184 channel=117
					-67, -9, 49, -13, -10, -24, 26, -5, -26,
					-- layer=2 filter=184 channel=118
					17, -17, 16, -1, 7, 7, 3, 25, 45,
					-- layer=2 filter=184 channel=119
					-14, 37, 7, 21, 13, -15, -13, 26, -15,
					-- layer=2 filter=184 channel=120
					8, -3, 5, 0, -1, 1, 8, 8, -9,
					-- layer=2 filter=184 channel=121
					2, -3, 10, -2, -2, 1, 2, 6, -8,
					-- layer=2 filter=184 channel=122
					11, 15, 13, -10, 11, 5, 0, -5, 0,
					-- layer=2 filter=184 channel=123
					-28, -3, 27, -21, -15, -9, 25, -13, 16,
					-- layer=2 filter=184 channel=124
					-24, -14, -25, 39, -33, -9, -4, -29, -20,
					-- layer=2 filter=184 channel=125
					7, -1, 1, 5, -10, -6, -1, -5, -1,
					-- layer=2 filter=184 channel=126
					43, 8, -25, 36, 29, -28, 74, -8, -7,
					-- layer=2 filter=184 channel=127
					-15, 13, -22, -1, 7, -15, 6, -12, -11,
					-- layer=2 filter=185 channel=0
					-26, -11, -12, -33, -26, -20, -14, -11, 2,
					-- layer=2 filter=185 channel=1
					-17, 17, 1, -11, 6, 17, -57, -53, -31,
					-- layer=2 filter=185 channel=2
					9, 5, 8, 0, 10, -5, 2, -5, 10,
					-- layer=2 filter=185 channel=3
					0, -4, -5, 0, 0, -39, -26, -5, 3,
					-- layer=2 filter=185 channel=4
					-8, -5, 41, -14, -22, -20, -11, -27, 0,
					-- layer=2 filter=185 channel=5
					0, -11, 36, -28, 9, 5, 44, 0, 9,
					-- layer=2 filter=185 channel=6
					-21, -29, -1, -8, -52, -22, -50, -28, 7,
					-- layer=2 filter=185 channel=7
					-12, -7, -4, 19, -11, -24, 10, -15, -28,
					-- layer=2 filter=185 channel=8
					-1, 3, -10, 5, -2, -2, 4, -1, 5,
					-- layer=2 filter=185 channel=9
					-16, 7, 9, -18, -19, -15, -28, -24, -45,
					-- layer=2 filter=185 channel=10
					7, 0, -8, -32, -19, -13, -28, -12, -6,
					-- layer=2 filter=185 channel=11
					-23, -24, 13, -14, -38, -4, -1, -25, -3,
					-- layer=2 filter=185 channel=12
					-33, -11, -14, 6, 18, 28, -61, -57, -36,
					-- layer=2 filter=185 channel=13
					-3, -11, 3, -2, -7, 8, -5, -4, 4,
					-- layer=2 filter=185 channel=14
					-32, 7, -2, -4, 3, 25, -10, -20, -8,
					-- layer=2 filter=185 channel=15
					24, 18, 5, 30, 5, 18, 22, 12, 49,
					-- layer=2 filter=185 channel=16
					-16, -7, 17, -13, -12, -38, 15, 23, 24,
					-- layer=2 filter=185 channel=17
					-6, 4, 0, -9, 6, 10, 7, 2, -2,
					-- layer=2 filter=185 channel=18
					36, -34, -19, 4, -25, 22, 38, -27, 1,
					-- layer=2 filter=185 channel=19
					0, 0, 19, -1, 2, -10, -27, -39, -11,
					-- layer=2 filter=185 channel=20
					8, 0, 0, 0, -5, 7, -1, 0, -7,
					-- layer=2 filter=185 channel=21
					-7, 3, 5, -6, -8, -2, -3, -4, -12,
					-- layer=2 filter=185 channel=22
					4, 3, -5, -2, 5, 2, 5, 2, 8,
					-- layer=2 filter=185 channel=23
					20, -37, 8, -19, -37, -6, -31, -1, 39,
					-- layer=2 filter=185 channel=24
					-8, -9, 13, -2, -18, -15, -28, 1, -16,
					-- layer=2 filter=185 channel=25
					-25, -9, -17, 0, 10, -13, -3, 0, -2,
					-- layer=2 filter=185 channel=26
					-8, 0, -7, -8, 0, 2, -9, -4, -5,
					-- layer=2 filter=185 channel=27
					0, 29, 43, -22, 13, 15, -14, 2, 2,
					-- layer=2 filter=185 channel=28
					-21, -34, -39, -59, -4, 0, -4, 10, 24,
					-- layer=2 filter=185 channel=29
					-10, 1, -7, -9, 5, 5, -1, -9, 8,
					-- layer=2 filter=185 channel=30
					-9, 22, -14, -26, -31, -15, 8, -24, -41,
					-- layer=2 filter=185 channel=31
					18, 27, 56, -26, 14, 61, 2, 6, 34,
					-- layer=2 filter=185 channel=32
					11, 7, 5, 8, 9, -3, -8, 0, -3,
					-- layer=2 filter=185 channel=33
					-29, -12, -25, 22, -32, -29, 51, 27, 9,
					-- layer=2 filter=185 channel=34
					52, -13, -28, 2, -32, -31, 38, -50, -6,
					-- layer=2 filter=185 channel=35
					-29, -48, -30, 11, 45, 8, -8, -19, 15,
					-- layer=2 filter=185 channel=36
					4, 1, -3, 3, 2, 3, -2, 2, 0,
					-- layer=2 filter=185 channel=37
					11, 6, 31, -10, -16, -11, -2, -20, 0,
					-- layer=2 filter=185 channel=38
					-9, 1, 34, -38, -13, 16, -1, 7, -7,
					-- layer=2 filter=185 channel=39
					14, -7, -5, 23, -4, -19, 15, 3, 5,
					-- layer=2 filter=185 channel=40
					31, 36, 8, -28, -51, -37, 59, 17, 23,
					-- layer=2 filter=185 channel=41
					-10, 0, -6, 3, 8, -10, 0, 8, 5,
					-- layer=2 filter=185 channel=42
					-10, -38, 0, 15, -1, -7, -36, -9, 36,
					-- layer=2 filter=185 channel=43
					33, 17, 17, 1, 0, -8, 36, 33, 20,
					-- layer=2 filter=185 channel=44
					4, 0, -3, 9, 6, -3, 0, 1, 1,
					-- layer=2 filter=185 channel=45
					2, 14, 37, -32, -7, -14, 30, 25, 33,
					-- layer=2 filter=185 channel=46
					0, -13, 28, -9, 18, -16, 10, 26, 26,
					-- layer=2 filter=185 channel=47
					-5, -31, -26, -25, -27, -30, 35, 22, 31,
					-- layer=2 filter=185 channel=48
					6, 0, 10, 4, -2, -10, 3, -6, -8,
					-- layer=2 filter=185 channel=49
					28, 13, 5, 14, -26, -3, -23, -33, -15,
					-- layer=2 filter=185 channel=50
					-1, -1, 6, 7, 0, 12, 2, 7, -3,
					-- layer=2 filter=185 channel=51
					-29, -11, -6, -3, -32, -12, -9, -14, -13,
					-- layer=2 filter=185 channel=52
					-6, 15, -22, 17, -27, -18, 22, -53, -29,
					-- layer=2 filter=185 channel=53
					-10, 58, 29, -43, 35, 17, -59, -26, 35,
					-- layer=2 filter=185 channel=54
					-16, -44, 22, -4, -18, -18, 28, -25, -12,
					-- layer=2 filter=185 channel=55
					4, -8, -1, 10, 7, 9, -4, -10, -1,
					-- layer=2 filter=185 channel=56
					-6, -24, 3, -33, -15, -1, 0, -19, 15,
					-- layer=2 filter=185 channel=57
					1, 2, -8, 5, 8, 1, 6, -1, 7,
					-- layer=2 filter=185 channel=58
					-43, -22, 3, 5, 18, 37, -61, -29, -41,
					-- layer=2 filter=185 channel=59
					-19, 25, 23, 0, -27, -3, -66, -9, -16,
					-- layer=2 filter=185 channel=60
					-15, 1, -30, -16, -6, 15, -33, 0, -25,
					-- layer=2 filter=185 channel=61
					-36, 29, -31, -45, -4, -42, -55, 22, -16,
					-- layer=2 filter=185 channel=62
					-34, -6, 8, -13, -52, -6, -28, -22, 4,
					-- layer=2 filter=185 channel=63
					-28, 2, 7, -12, -31, 1, -29, 8, 9,
					-- layer=2 filter=185 channel=64
					26, 3, -1, 0, -7, 2, -13, 16, 7,
					-- layer=2 filter=185 channel=65
					-28, 5, -13, -17, 0, -49, -44, -16, -31,
					-- layer=2 filter=185 channel=66
					13, -5, 17, 30, 52, 12, 28, 24, 6,
					-- layer=2 filter=185 channel=67
					-13, 7, 27, -27, -25, -8, -17, 11, -15,
					-- layer=2 filter=185 channel=68
					9, 5, -3, -3, 8, 5, -2, 8, -3,
					-- layer=2 filter=185 channel=69
					4, -16, -14, 19, 6, 6, 24, 13, -23,
					-- layer=2 filter=185 channel=70
					-25, -17, -14, -24, 22, -1, 4, -26, -1,
					-- layer=2 filter=185 channel=71
					-3, 41, 42, -19, 27, 25, -11, -16, 0,
					-- layer=2 filter=185 channel=72
					0, -22, -19, -20, 2, -31, 11, 14, 3,
					-- layer=2 filter=185 channel=73
					13, -2, 15, -30, 0, 11, 22, 8, 22,
					-- layer=2 filter=185 channel=74
					-38, -19, -16, -50, -29, 0, -18, 2, 10,
					-- layer=2 filter=185 channel=75
					-11, -6, 20, -12, 30, 35, -11, -26, -7,
					-- layer=2 filter=185 channel=76
					-48, 23, 20, -49, -20, 11, -50, -45, 6,
					-- layer=2 filter=185 channel=77
					2, 1, 7, 6, -4, -2, -6, -6, -5,
					-- layer=2 filter=185 channel=78
					1, -3, -16, 2, -26, 2, 10, 17, 15,
					-- layer=2 filter=185 channel=79
					0, 4, 8, 9, 8, -1, -9, -1, -4,
					-- layer=2 filter=185 channel=80
					-1, -10, 10, -6, -25, -9, -4, 10, 5,
					-- layer=2 filter=185 channel=81
					-6, -3, 8, 9, -5, -8, -6, 0, 0,
					-- layer=2 filter=185 channel=82
					-3, 2, -7, -2, -3, -4, -11, 9, 2,
					-- layer=2 filter=185 channel=83
					-9, 8, 31, -2, 19, 6, -46, -25, -9,
					-- layer=2 filter=185 channel=84
					-3, 12, -3, -7, 8, -8, -5, -7, 6,
					-- layer=2 filter=185 channel=85
					3, -6, 9, -3, 2, 0, -1, -1, -2,
					-- layer=2 filter=185 channel=86
					8, 5, -1, 7, 5, 3, -2, -4, -2,
					-- layer=2 filter=185 channel=87
					-21, 6, -35, 0, -41, -10, -13, -13, -7,
					-- layer=2 filter=185 channel=88
					-39, 25, -34, -5, -10, 4, -9, -23, -18,
					-- layer=2 filter=185 channel=89
					-36, -29, -22, 3, 4, 17, -59, -42, -14,
					-- layer=2 filter=185 channel=90
					-7, 12, -1, 9, -7, 10, 3, -4, -5,
					-- layer=2 filter=185 channel=91
					-30, -42, -4, -3, 20, 34, -49, -23, -3,
					-- layer=2 filter=185 channel=92
					-31, -3, 0, 4, -1, 18, -50, -40, -20,
					-- layer=2 filter=185 channel=93
					-11, 22, -8, 30, -7, -36, 21, -2, -19,
					-- layer=2 filter=185 channel=94
					-29, -2, -5, -48, -21, -17, -62, -17, -25,
					-- layer=2 filter=185 channel=95
					4, 6, -6, 3, 7, 0, -3, 10, -2,
					-- layer=2 filter=185 channel=96
					-20, 44, 5, -10, 44, 0, -28, -4, -5,
					-- layer=2 filter=185 channel=97
					35, -15, -4, 19, 11, -5, 9, 4, 1,
					-- layer=2 filter=185 channel=98
					-42, -15, -46, -59, -44, -49, 0, 19, 11,
					-- layer=2 filter=185 channel=99
					47, 39, -3, 18, -3, -3, -26, -10, -9,
					-- layer=2 filter=185 channel=100
					-9, 7, 40, -32, 17, 53, -13, -31, -28,
					-- layer=2 filter=185 channel=101
					-7, 1, 12, 18, 17, 35, 28, -1, -16,
					-- layer=2 filter=185 channel=102
					1, 16, 34, 26, -29, -9, 16, -49, -16,
					-- layer=2 filter=185 channel=103
					-13, -28, -14, -13, -17, -30, 14, 24, -12,
					-- layer=2 filter=185 channel=104
					-1, -24, 17, -9, 27, 19, -35, -49, 15,
					-- layer=2 filter=185 channel=105
					16, -5, -14, -3, -28, -32, 9, 1, -19,
					-- layer=2 filter=185 channel=106
					-43, -27, 3, -4, -7, 14, 4, 3, -16,
					-- layer=2 filter=185 channel=107
					-10, 4, -19, 13, -5, 8, -4, 45, 31,
					-- layer=2 filter=185 channel=108
					5, 34, 43, -20, 6, 24, -7, -23, -20,
					-- layer=2 filter=185 channel=109
					-3, 9, 11, -4, -5, -5, -2, 0, 5,
					-- layer=2 filter=185 channel=110
					2, 32, -30, -1, 32, 8, -47, 13, 25,
					-- layer=2 filter=185 channel=111
					2, -5, 1, 2, 5, -2, 6, -1, -4,
					-- layer=2 filter=185 channel=112
					0, -2, -41, -34, -21, -36, -32, 4, -23,
					-- layer=2 filter=185 channel=113
					0, -8, -40, -22, 5, 5, -30, 2, -27,
					-- layer=2 filter=185 channel=114
					4, -3, -4, -2, -2, 0, -5, -4, 5,
					-- layer=2 filter=185 channel=115
					-2, 2, 10, 6, 10, 0, -7, -5, -8,
					-- layer=2 filter=185 channel=116
					0, -2, -5, 12, -9, 4, -21, -16, -18,
					-- layer=2 filter=185 channel=117
					46, -6, -22, 35, 35, -21, 45, 17, -1,
					-- layer=2 filter=185 channel=118
					-4, 4, -6, 2, 0, -20, -10, 8, 11,
					-- layer=2 filter=185 channel=119
					-16, -44, 7, -51, -24, 10, -3, -11, 24,
					-- layer=2 filter=185 channel=120
					2, 8, 0, -8, 7, -4, 6, 10, -8,
					-- layer=2 filter=185 channel=121
					9, -3, 11, -9, -6, 8, -4, -1, 0,
					-- layer=2 filter=185 channel=122
					7, -7, -4, -7, 2, -4, 0, 6, 2,
					-- layer=2 filter=185 channel=123
					6, -24, -45, -21, -13, -72, -5, -28, -12,
					-- layer=2 filter=185 channel=124
					-12, -14, -3, -4, -6, 10, 16, -1, 37,
					-- layer=2 filter=185 channel=125
					-4, 0, -3, 7, 4, -3, 10, -5, -9,
					-- layer=2 filter=185 channel=126
					-16, 14, -12, -38, 13, -13, -59, -31, -12,
					-- layer=2 filter=185 channel=127
					-41, 5, -13, -35, 6, -1, 5, -19, 4,
					-- layer=2 filter=186 channel=0
					-5, -10, 8, -9, -8, 4, -4, -12, 4,
					-- layer=2 filter=186 channel=1
					1, -1, 0, 6, 8, 3, 5, -10, -1,
					-- layer=2 filter=186 channel=2
					-7, -2, -6, -2, 6, 0, 5, -6, 3,
					-- layer=2 filter=186 channel=3
					5, -1, 5, 4, -7, -7, 1, -13, -3,
					-- layer=2 filter=186 channel=4
					-12, -5, 2, -7, 0, 2, 5, 2, -7,
					-- layer=2 filter=186 channel=5
					-6, 5, -1, 6, -5, -5, -7, -11, -10,
					-- layer=2 filter=186 channel=6
					-9, -5, -2, 2, 4, 1, -9, -2, -9,
					-- layer=2 filter=186 channel=7
					-11, -1, -6, 3, 5, 1, -9, 1, 3,
					-- layer=2 filter=186 channel=8
					5, 1, -9, -6, 8, -3, 8, 9, 4,
					-- layer=2 filter=186 channel=9
					2, -9, -5, -11, -4, -11, -1, -8, -8,
					-- layer=2 filter=186 channel=10
					6, -12, -2, -4, -10, 0, -13, 2, -9,
					-- layer=2 filter=186 channel=11
					0, -2, 0, 4, -8, -10, -4, 1, 3,
					-- layer=2 filter=186 channel=12
					-3, -9, -4, -10, 0, 4, -7, 0, 0,
					-- layer=2 filter=186 channel=13
					-5, 5, 10, 0, -8, 0, -2, 1, 1,
					-- layer=2 filter=186 channel=14
					8, -6, 0, 4, -2, -6, -11, -4, -3,
					-- layer=2 filter=186 channel=15
					7, 2, 7, 4, 3, 6, 6, -2, 2,
					-- layer=2 filter=186 channel=16
					3, -4, -1, -4, -1, 3, 0, 8, -3,
					-- layer=2 filter=186 channel=17
					-9, -2, 9, 10, 8, -4, -6, -7, -1,
					-- layer=2 filter=186 channel=18
					-5, -3, -8, 0, 1, 0, -6, -9, -14,
					-- layer=2 filter=186 channel=19
					2, -9, 8, -10, -7, -6, -2, 7, 3,
					-- layer=2 filter=186 channel=20
					11, 5, 11, 3, -5, -2, -7, -4, -1,
					-- layer=2 filter=186 channel=21
					-1, -4, -2, 0, 6, -1, 3, 0, -7,
					-- layer=2 filter=186 channel=22
					0, 2, 0, -11, -7, -4, 0, 3, 4,
					-- layer=2 filter=186 channel=23
					-4, 7, -1, 6, 7, 0, -7, 6, -8,
					-- layer=2 filter=186 channel=24
					3, 8, 7, 2, 5, -4, -8, 6, -3,
					-- layer=2 filter=186 channel=25
					5, 0, -5, -3, 5, -12, 1, -8, 6,
					-- layer=2 filter=186 channel=26
					1, -1, -3, 6, 3, -9, 8, -9, -1,
					-- layer=2 filter=186 channel=27
					-3, -11, 3, -4, 1, 0, -3, -7, 5,
					-- layer=2 filter=186 channel=28
					-12, 0, -5, -10, -11, 3, 0, -1, -8,
					-- layer=2 filter=186 channel=29
					-9, -8, 6, 4, 6, 0, 4, 9, -4,
					-- layer=2 filter=186 channel=30
					5, -8, -9, 0, 4, -10, 6, 6, -10,
					-- layer=2 filter=186 channel=31
					-3, 9, -9, -9, -7, -10, 0, 7, 0,
					-- layer=2 filter=186 channel=32
					-1, 0, -4, -2, -4, -4, 9, -2, 0,
					-- layer=2 filter=186 channel=33
					-2, -7, 0, -12, 6, -9, 0, 0, 7,
					-- layer=2 filter=186 channel=34
					-5, 0, 5, 5, -5, -4, -9, 7, 6,
					-- layer=2 filter=186 channel=35
					3, -3, 5, -1, 6, -13, -7, 3, -5,
					-- layer=2 filter=186 channel=36
					7, 0, 4, 8, -5, -2, 0, -2, -6,
					-- layer=2 filter=186 channel=37
					7, 0, -8, -3, -1, 2, 0, -11, 7,
					-- layer=2 filter=186 channel=38
					-2, -1, 0, 3, 4, -9, -8, 10, 1,
					-- layer=2 filter=186 channel=39
					3, 6, 6, -1, -8, -9, 8, -9, 9,
					-- layer=2 filter=186 channel=40
					-1, 0, 1, 1, 3, 4, -10, -1, -13,
					-- layer=2 filter=186 channel=41
					6, 0, -6, -9, 1, 0, -5, 6, 0,
					-- layer=2 filter=186 channel=42
					-4, -2, -9, -9, 5, 4, 6, 0, -1,
					-- layer=2 filter=186 channel=43
					6, -3, -6, -2, 5, 2, -7, -3, 1,
					-- layer=2 filter=186 channel=44
					-1, 3, 2, -1, 0, 2, -5, 2, -1,
					-- layer=2 filter=186 channel=45
					4, -3, -7, -4, 4, 2, 4, 1, 7,
					-- layer=2 filter=186 channel=46
					-5, -8, -5, -11, 0, -9, -7, 5, 0,
					-- layer=2 filter=186 channel=47
					-12, -2, -4, 0, 9, 6, -4, -3, 0,
					-- layer=2 filter=186 channel=48
					-4, 0, 1, -5, 7, -5, -8, 10, -1,
					-- layer=2 filter=186 channel=49
					-11, 6, -1, -8, 0, -5, -9, -5, 1,
					-- layer=2 filter=186 channel=50
					1, 1, -2, -4, -4, -3, 2, -6, -4,
					-- layer=2 filter=186 channel=51
					-3, 0, 4, 4, 6, 3, -9, -13, -13,
					-- layer=2 filter=186 channel=52
					-8, -9, -10, 0, -6, -2, -9, -12, -9,
					-- layer=2 filter=186 channel=53
					-3, -2, -5, 0, 2, -2, -5, -11, 7,
					-- layer=2 filter=186 channel=54
					-1, 0, -3, -7, -6, 0, -8, -13, 5,
					-- layer=2 filter=186 channel=55
					7, -7, -7, 3, 8, 3, 4, 0, -2,
					-- layer=2 filter=186 channel=56
					5, -1, -6, 2, -1, 6, 3, -8, -5,
					-- layer=2 filter=186 channel=57
					-3, 10, 0, 6, 6, 8, -7, 6, -3,
					-- layer=2 filter=186 channel=58
					-6, 0, 6, -11, 4, 0, -8, 9, 8,
					-- layer=2 filter=186 channel=59
					-9, -7, -3, 7, 1, 2, -12, 6, -7,
					-- layer=2 filter=186 channel=60
					-11, -3, -8, 1, 6, 2, -1, -1, 10,
					-- layer=2 filter=186 channel=61
					2, -6, 0, -13, -4, 4, -14, 6, -9,
					-- layer=2 filter=186 channel=62
					8, -13, -10, -1, 4, 0, -16, 5, -1,
					-- layer=2 filter=186 channel=63
					-6, -2, 1, 0, 4, -9, 1, -11, -3,
					-- layer=2 filter=186 channel=64
					-2, 0, -2, -10, 7, -8, 7, -3, -7,
					-- layer=2 filter=186 channel=65
					3, 0, 7, -2, -6, -4, 0, -2, -8,
					-- layer=2 filter=186 channel=66
					-8, -8, 6, 4, 9, 5, 10, -4, -2,
					-- layer=2 filter=186 channel=67
					-4, -3, -6, -6, 0, -3, 0, -11, -7,
					-- layer=2 filter=186 channel=68
					5, -6, 0, 1, 8, 6, 3, -7, 5,
					-- layer=2 filter=186 channel=69
					7, -1, 1, -12, -10, -9, -4, 7, -10,
					-- layer=2 filter=186 channel=70
					-5, -7, -10, 4, 0, -13, -3, 3, 2,
					-- layer=2 filter=186 channel=71
					-3, -3, -7, 5, 6, -4, -10, -11, -8,
					-- layer=2 filter=186 channel=72
					-12, 9, -6, -13, -14, -11, 7, 0, -10,
					-- layer=2 filter=186 channel=73
					-8, 1, -5, -10, -9, -2, -7, -18, 2,
					-- layer=2 filter=186 channel=74
					9, 2, -8, -5, 7, -1, -6, 7, -3,
					-- layer=2 filter=186 channel=75
					-8, -1, 8, -7, -4, -6, -2, 0, -3,
					-- layer=2 filter=186 channel=76
					0, -6, -10, 0, -13, -6, -16, -3, -6,
					-- layer=2 filter=186 channel=77
					-6, 3, -4, -8, 3, -6, 6, 9, 9,
					-- layer=2 filter=186 channel=78
					-4, -6, -9, -2, -10, -11, 4, -12, 4,
					-- layer=2 filter=186 channel=79
					7, 5, -1, -5, 5, 10, 9, 8, -4,
					-- layer=2 filter=186 channel=80
					2, -7, -11, 1, -10, -3, -8, -9, 4,
					-- layer=2 filter=186 channel=81
					6, 7, 2, -1, 10, 0, 10, 4, -8,
					-- layer=2 filter=186 channel=82
					8, -5, -9, 8, 2, -6, 0, -2, 3,
					-- layer=2 filter=186 channel=83
					-10, 0, 0, -8, -7, 4, 0, 7, -9,
					-- layer=2 filter=186 channel=84
					5, 3, 5, 0, 9, -6, 0, 0, -1,
					-- layer=2 filter=186 channel=85
					3, 8, -2, -3, -5, 3, 3, 2, 13,
					-- layer=2 filter=186 channel=86
					9, 3, -2, 1, -11, 0, -3, 2, 7,
					-- layer=2 filter=186 channel=87
					1, 2, 5, -7, 4, 5, -7, 0, -10,
					-- layer=2 filter=186 channel=88
					2, 2, 2, -10, -1, -11, -4, 5, 5,
					-- layer=2 filter=186 channel=89
					-14, -9, -9, -5, -8, -6, 3, -14, 3,
					-- layer=2 filter=186 channel=90
					-1, 7, -1, 0, 5, -2, -4, -5, -2,
					-- layer=2 filter=186 channel=91
					5, -5, -18, -5, -15, 13, 3, -10, -3,
					-- layer=2 filter=186 channel=92
					7, 0, -6, -13, 3, 5, -10, -5, 0,
					-- layer=2 filter=186 channel=93
					-4, -1, 0, -3, -3, -7, 1, -1, 7,
					-- layer=2 filter=186 channel=94
					-9, 0, -7, 0, -4, -4, 2, 4, -14,
					-- layer=2 filter=186 channel=95
					-3, 7, 7, -1, 4, 2, -4, -9, -10,
					-- layer=2 filter=186 channel=96
					-2, 3, -6, -1, 0, -8, -5, 6, -4,
					-- layer=2 filter=186 channel=97
					-8, 5, 6, 7, -10, 1, 4, 7, -9,
					-- layer=2 filter=186 channel=98
					6, 6, 4, 8, -10, -11, -9, 3, 0,
					-- layer=2 filter=186 channel=99
					4, 2, -5, 6, 8, 0, 4, -10, -4,
					-- layer=2 filter=186 channel=100
					6, -6, 4, 0, 10, 6, 6, 2, -10,
					-- layer=2 filter=186 channel=101
					-8, 6, 1, -8, 8, -5, -8, 8, 5,
					-- layer=2 filter=186 channel=102
					1, -4, 3, 6, -9, -6, -2, 7, 5,
					-- layer=2 filter=186 channel=103
					-7, -1, -3, 7, -7, 1, 0, 0, 0,
					-- layer=2 filter=186 channel=104
					5, -4, 4, 7, 0, -12, -5, 3, -4,
					-- layer=2 filter=186 channel=105
					6, -12, 0, -10, 4, -3, 6, -7, 5,
					-- layer=2 filter=186 channel=106
					-2, 1, -5, -3, -3, 6, -9, -8, 2,
					-- layer=2 filter=186 channel=107
					-8, 7, 0, -2, 9, 1, -4, -5, 10,
					-- layer=2 filter=186 channel=108
					-1, -1, 0, -9, 6, -4, 1, 1, 2,
					-- layer=2 filter=186 channel=109
					5, 6, 10, 7, 5, -7, 9, 8, -4,
					-- layer=2 filter=186 channel=110
					2, -5, -8, -13, 8, -8, 4, -8, -3,
					-- layer=2 filter=186 channel=111
					8, 0, 4, 0, 0, -7, 6, 3, 3,
					-- layer=2 filter=186 channel=112
					-2, 6, -12, -9, 8, 7, 0, 4, -12,
					-- layer=2 filter=186 channel=113
					-6, 5, -10, -8, 7, -8, -10, 1, -5,
					-- layer=2 filter=186 channel=114
					-4, -4, 11, 8, -3, -5, 7, 4, 5,
					-- layer=2 filter=186 channel=115
					0, 8, 0, 8, -2, 0, -3, -1, 0,
					-- layer=2 filter=186 channel=116
					0, 9, -13, -9, 0, -5, 0, 6, 6,
					-- layer=2 filter=186 channel=117
					2, 0, -6, 0, -12, -1, -10, 4, -8,
					-- layer=2 filter=186 channel=118
					2, -5, -5, -10, 2, 5, 3, 1, -8,
					-- layer=2 filter=186 channel=119
					4, 2, 0, 4, -4, -11, 1, -3, -3,
					-- layer=2 filter=186 channel=120
					-1, 3, 7, 7, -2, 7, -5, -6, 0,
					-- layer=2 filter=186 channel=121
					11, -4, 6, -6, -4, -7, -4, -2, 4,
					-- layer=2 filter=186 channel=122
					8, 1, 6, 5, -10, 4, 3, 0, -6,
					-- layer=2 filter=186 channel=123
					-2, -9, -1, 0, -17, 0, -12, -4, 0,
					-- layer=2 filter=186 channel=124
					-3, -4, -7, 0, 2, 1, 10, -11, 1,
					-- layer=2 filter=186 channel=125
					2, 0, 10, -1, -10, 7, -8, -5, 5,
					-- layer=2 filter=186 channel=126
					3, 10, -1, 9, 1, -7, 8, 7, -8,
					-- layer=2 filter=186 channel=127
					-2, -1, -11, 0, 5, 1, 1, 4, 2,
					-- layer=2 filter=187 channel=0
					3, -29, -9, 12, -14, -21, 0, -21, 17,
					-- layer=2 filter=187 channel=1
					-1, -36, -31, -13, 6, -1, 13, 30, 16,
					-- layer=2 filter=187 channel=2
					3, 6, -2, 2, -7, -4, 11, 0, 1,
					-- layer=2 filter=187 channel=3
					-16, 11, 14, -12, -37, -11, 32, 12, 33,
					-- layer=2 filter=187 channel=4
					-38, 7, 27, 0, 29, 0, -19, 4, -20,
					-- layer=2 filter=187 channel=5
					0, 0, -10, -18, -19, -8, -1, -3, 1,
					-- layer=2 filter=187 channel=6
					51, 28, 6, 29, 56, 19, 48, 36, 2,
					-- layer=2 filter=187 channel=7
					-14, -45, -23, 8, 8, 24, 25, 18, 28,
					-- layer=2 filter=187 channel=8
					-1, 7, 4, -8, 5, 9, 4, 7, -8,
					-- layer=2 filter=187 channel=9
					7, 6, 27, -23, -19, -9, -42, -53, -21,
					-- layer=2 filter=187 channel=10
					-11, -8, -15, 21, -15, 4, 9, -16, 27,
					-- layer=2 filter=187 channel=11
					-12, -16, -16, -25, -20, -21, 1, -26, -9,
					-- layer=2 filter=187 channel=12
					0, -30, -32, -32, 13, 16, 30, 45, 3,
					-- layer=2 filter=187 channel=13
					0, 0, 3, -1, 8, 7, 6, -3, -8,
					-- layer=2 filter=187 channel=14
					-4, -26, -35, -36, -13, 12, 16, 12, -5,
					-- layer=2 filter=187 channel=15
					-7, -10, 10, -30, -21, 8, -34, -18, 33,
					-- layer=2 filter=187 channel=16
					4, 7, 6, 31, 7, 19, -11, -21, -41,
					-- layer=2 filter=187 channel=17
					0, -10, 2, -7, -5, -8, -6, 4, 4,
					-- layer=2 filter=187 channel=18
					-9, 19, 7, 9, 10, -41, -6, -22, -4,
					-- layer=2 filter=187 channel=19
					-7, -23, -1, 12, -15, -13, -12, 20, 17,
					-- layer=2 filter=187 channel=20
					10, -6, -2, 7, -6, -1, -2, -5, -9,
					-- layer=2 filter=187 channel=21
					0, 3, 4, 12, 1, 8, 3, 3, 0,
					-- layer=2 filter=187 channel=22
					-8, -1, -3, 10, -3, 0, 11, -4, -10,
					-- layer=2 filter=187 channel=23
					-15, 5, 15, -25, 6, -5, 7, 0, 8,
					-- layer=2 filter=187 channel=24
					0, 0, -2, 1, -20, -9, -11, -49, -38,
					-- layer=2 filter=187 channel=25
					-47, -27, -19, -13, -41, -4, -49, -38, -49,
					-- layer=2 filter=187 channel=26
					-6, 1, -10, -5, 1, -4, 6, 10, 4,
					-- layer=2 filter=187 channel=27
					6, -12, 10, 18, -8, -10, -16, -33, -20,
					-- layer=2 filter=187 channel=28
					-19, -80, -66, -45, -24, 15, -6, 19, 17,
					-- layer=2 filter=187 channel=29
					8, 0, 0, -5, 11, -6, 2, -6, 0,
					-- layer=2 filter=187 channel=30
					3, 18, 21, -26, -28, 6, -40, 8, -42,
					-- layer=2 filter=187 channel=31
					-1, 35, -29, 18, -7, 5, -53, -31, -3,
					-- layer=2 filter=187 channel=32
					-3, 8, -1, 7, -11, -6, -8, 0, 0,
					-- layer=2 filter=187 channel=33
					-27, -29, -50, -40, -20, 43, 33, 24, 33,
					-- layer=2 filter=187 channel=34
					29, 24, -14, 16, -6, -5, -65, 35, 23,
					-- layer=2 filter=187 channel=35
					-78, -63, -66, -28, -37, -15, 21, 23, 25,
					-- layer=2 filter=187 channel=36
					0, 0, 2, 10, -8, 14, 1, -2, 1,
					-- layer=2 filter=187 channel=37
					0, -4, -8, 0, -20, -4, -6, -8, 2,
					-- layer=2 filter=187 channel=38
					-11, -23, -7, -24, -34, 2, 9, 0, 17,
					-- layer=2 filter=187 channel=39
					9, 33, 10, -8, 7, 39, 17, -36, -8,
					-- layer=2 filter=187 channel=40
					-6, 2, 45, 0, -12, -22, -24, -55, -13,
					-- layer=2 filter=187 channel=41
					-3, 0, 0, 1, 5, 4, -11, 0, -4,
					-- layer=2 filter=187 channel=42
					20, 0, 13, 0, -31, -9, 11, 9, -3,
					-- layer=2 filter=187 channel=43
					-21, -15, 20, 14, -5, -15, 13, 2, 9,
					-- layer=2 filter=187 channel=44
					1, 0, 1, 1, -7, 0, 2, 6, -3,
					-- layer=2 filter=187 channel=45
					33, 15, 0, 54, 38, 40, -30, -24, -15,
					-- layer=2 filter=187 channel=46
					6, 6, 56, 17, 1, 29, 7, -39, -16,
					-- layer=2 filter=187 channel=47
					10, -58, -38, -1, 27, 67, -2, -17, 21,
					-- layer=2 filter=187 channel=48
					0, -1, 3, 1, -2, -6, 1, 4, -4,
					-- layer=2 filter=187 channel=49
					22, 3, 1, 19, 13, -13, 4, -9, -48,
					-- layer=2 filter=187 channel=50
					3, 20, 13, 8, 1, 8, 1, -27, -23,
					-- layer=2 filter=187 channel=51
					-24, -13, -25, -2, -21, -15, -19, -17, -5,
					-- layer=2 filter=187 channel=52
					-21, 5, 16, -4, 5, -15, -4, 37, -9,
					-- layer=2 filter=187 channel=53
					19, -4, 15, 25, 6, -25, 8, -27, 18,
					-- layer=2 filter=187 channel=54
					-5, -26, -39, -5, 9, -5, -2, 14, 5,
					-- layer=2 filter=187 channel=55
					0, 8, -10, 5, 4, -2, -2, -11, 10,
					-- layer=2 filter=187 channel=56
					-12, -9, -4, -18, -16, 9, 5, -22, 8,
					-- layer=2 filter=187 channel=57
					4, 0, -7, 7, 5, 6, 9, -8, 22,
					-- layer=2 filter=187 channel=58
					-18, -25, -33, -43, 14, 13, 57, 42, 32,
					-- layer=2 filter=187 channel=59
					-2, -27, 8, -24, -6, -3, -2, 28, 7,
					-- layer=2 filter=187 channel=60
					-3, -23, -2, -10, 4, 30, 14, 37, 27,
					-- layer=2 filter=187 channel=61
					24, 25, -12, 20, 42, 3, 17, 10, 3,
					-- layer=2 filter=187 channel=62
					48, -2, -22, 35, 24, -24, 20, 14, -48,
					-- layer=2 filter=187 channel=63
					16, 12, -1, 12, 4, 13, -5, -6, -11,
					-- layer=2 filter=187 channel=64
					14, 36, 27, -5, 15, 4, -21, 9, -22,
					-- layer=2 filter=187 channel=65
					11, 12, -3, 12, 26, 9, 17, 15, -6,
					-- layer=2 filter=187 channel=66
					44, -21, 14, -26, -75, 37, 31, -23, 0,
					-- layer=2 filter=187 channel=67
					4, 7, 58, -29, -27, 0, -49, -83, -28,
					-- layer=2 filter=187 channel=68
					6, -6, 2, 0, -4, 6, -1, -6, -9,
					-- layer=2 filter=187 channel=69
					15, 19, 17, 4, 14, 19, 10, -2, -15,
					-- layer=2 filter=187 channel=70
					-35, -38, -50, 5, -16, 35, 30, 27, 38,
					-- layer=2 filter=187 channel=71
					16, 9, 57, 32, 15, -7, -45, -15, -26,
					-- layer=2 filter=187 channel=72
					-13, -53, -36, -26, -61, -8, 6, -12, 19,
					-- layer=2 filter=187 channel=73
					20, 45, 54, 15, 29, 14, -14, -37, 26,
					-- layer=2 filter=187 channel=74
					15, 5, 37, -15, -16, 12, -11, -8, -12,
					-- layer=2 filter=187 channel=75
					-26, -47, -12, 5, 8, 33, 25, 30, 19,
					-- layer=2 filter=187 channel=76
					5, -17, -7, 22, 30, 14, -58, -7, 52,
					-- layer=2 filter=187 channel=77
					7, 5, -2, 1, 0, -2, 4, 3, -6,
					-- layer=2 filter=187 channel=78
					-23, -25, -19, 0, -15, -14, 17, -19, -20,
					-- layer=2 filter=187 channel=79
					2, -5, 2, -5, 1, 1, 7, -5, 0,
					-- layer=2 filter=187 channel=80
					0, 33, 53, 7, -11, 33, -5, -1, -28,
					-- layer=2 filter=187 channel=81
					-2, 8, 4, -8, -7, 0, -1, 1, 0,
					-- layer=2 filter=187 channel=82
					2, -6, -13, 3, -7, 8, -6, -4, -2,
					-- layer=2 filter=187 channel=83
					-1, 16, 26, 4, 32, -2, 8, 33, -46,
					-- layer=2 filter=187 channel=84
					5, 9, 2, -8, -6, -6, -7, 2, -9,
					-- layer=2 filter=187 channel=85
					3, -5, 11, 0, 13, 8, -1, -7, 12,
					-- layer=2 filter=187 channel=86
					6, -22, -15, 4, 0, -11, -4, -8, -17,
					-- layer=2 filter=187 channel=87
					-8, -22, -6, -44, 4, -11, -39, 14, 2,
					-- layer=2 filter=187 channel=88
					15, 22, 31, -9, 27, 3, -22, 1, -26,
					-- layer=2 filter=187 channel=89
					-4, -33, -12, -61, -18, 4, 25, -1, -13,
					-- layer=2 filter=187 channel=90
					7, 0, 10, 4, 0, -3, -6, -8, 3,
					-- layer=2 filter=187 channel=91
					8, -49, 0, -1, -33, 45, 31, -5, 1,
					-- layer=2 filter=187 channel=92
					-1, -32, -38, -19, -11, 16, 21, 8, 2,
					-- layer=2 filter=187 channel=93
					0, 24, 5, 29, 36, 29, 11, -17, 26,
					-- layer=2 filter=187 channel=94
					37, -6, 1, 2, 17, -12, 39, 32, -11,
					-- layer=2 filter=187 channel=95
					4, -5, 4, -5, -11, -18, 12, -16, 7,
					-- layer=2 filter=187 channel=96
					29, 34, 63, 22, 43, 19, 6, 6, 36,
					-- layer=2 filter=187 channel=97
					-28, -24, 30, -50, -26, -3, 4, -20, -6,
					-- layer=2 filter=187 channel=98
					-14, -71, -51, -4, 2, 36, -6, -10, 30,
					-- layer=2 filter=187 channel=99
					34, 54, 27, 2, -12, -5, 5, 7, 0,
					-- layer=2 filter=187 channel=100
					11, -3, 24, -37, -17, 12, -19, 32, -27,
					-- layer=2 filter=187 channel=101
					-26, -39, 27, -36, -49, 18, -25, -50, 0,
					-- layer=2 filter=187 channel=102
					-31, 27, 7, 2, 37, -37, -26, 10, -32,
					-- layer=2 filter=187 channel=103
					35, 2, -28, 4, 27, 43, -8, -17, 33,
					-- layer=2 filter=187 channel=104
					48, 2, 15, 15, 0, -29, 23, -11, -33,
					-- layer=2 filter=187 channel=105
					-2, -20, -37, 1, -46, -48, -21, -30, -28,
					-- layer=2 filter=187 channel=106
					-31, -47, 1, -42, -29, 43, 5, -41, -5,
					-- layer=2 filter=187 channel=107
					-24, -12, -30, -19, 9, -32, 61, -22, 22,
					-- layer=2 filter=187 channel=108
					27, 23, 0, 25, 19, -29, -39, -9, -39,
					-- layer=2 filter=187 channel=109
					-5, 10, -15, -12, 13, 0, -15, 9, 0,
					-- layer=2 filter=187 channel=110
					-9, 16, 11, -17, 24, -9, -37, 13, -4,
					-- layer=2 filter=187 channel=111
					-5, 9, 7, 0, -4, 11, 6, 3, 6,
					-- layer=2 filter=187 channel=112
					2, -14, 21, 4, -20, -2, -3, -27, -2,
					-- layer=2 filter=187 channel=113
					6, -1, 10, -24, -18, 3, 8, 6, -26,
					-- layer=2 filter=187 channel=114
					-8, -9, 0, -6, -6, 6, -17, 1, -2,
					-- layer=2 filter=187 channel=115
					-9, 0, -12, 10, -1, 1, -8, 9, 4,
					-- layer=2 filter=187 channel=116
					-14, -1, -24, -25, 15, 1, -33, -10, 18,
					-- layer=2 filter=187 channel=117
					-21, -21, 8, 23, 8, 7, 30, -1, 12,
					-- layer=2 filter=187 channel=118
					1, 12, 39, 25, -7, -5, 15, 0, 23,
					-- layer=2 filter=187 channel=119
					43, 33, 10, 19, 13, -24, -3, 11, -15,
					-- layer=2 filter=187 channel=120
					7, -2, 3, -10, 0, -9, 2, 10, 9,
					-- layer=2 filter=187 channel=121
					3, 1, -5, 0, -9, 2, -1, -6, 7,
					-- layer=2 filter=187 channel=122
					0, -11, -2, -2, -10, 12, -12, 0, 5,
					-- layer=2 filter=187 channel=123
					-13, -74, -25, -16, -13, 3, 13, 1, 18,
					-- layer=2 filter=187 channel=124
					-41, -47, -8, -62, -13, 18, 9, 20, 36,
					-- layer=2 filter=187 channel=125
					-9, 0, -1, -5, 0, 6, -2, -7, 0,
					-- layer=2 filter=187 channel=126
					36, 65, 17, -25, -14, 17, 43, 43, 78,
					-- layer=2 filter=187 channel=127
					26, 18, -10, -9, -11, -2, -5, 20, -23,
					-- layer=2 filter=188 channel=0
					0, 4, 6, -14, -4, 2, -16, -8, 14,
					-- layer=2 filter=188 channel=1
					11, -41, -12, 13, -1, 4, 35, -17, -8,
					-- layer=2 filter=188 channel=2
					2, -5, 0, 0, -1, -1, -9, -9, 8,
					-- layer=2 filter=188 channel=3
					18, 7, -19, -40, 12, -1, 9, 13, 10,
					-- layer=2 filter=188 channel=4
					-20, -22, 32, 13, -5, 18, -11, 3, -5,
					-- layer=2 filter=188 channel=5
					3, 0, 19, -27, -3, 14, 8, -17, -15,
					-- layer=2 filter=188 channel=6
					-18, -68, -35, 14, -46, -34, 20, 43, -13,
					-- layer=2 filter=188 channel=7
					53, 47, 56, 12, 56, 53, -13, -25, 29,
					-- layer=2 filter=188 channel=8
					7, 11, -9, 3, -1, 7, 6, 0, -3,
					-- layer=2 filter=188 channel=9
					0, -15, -29, -9, 42, 7, 35, 44, 1,
					-- layer=2 filter=188 channel=10
					-2, -5, -11, -15, 1, -4, -15, -1, 10,
					-- layer=2 filter=188 channel=11
					-26, -15, -13, -19, -27, -11, -13, -8, -27,
					-- layer=2 filter=188 channel=12
					4, -13, 22, 26, 27, 12, 12, 9, 3,
					-- layer=2 filter=188 channel=13
					11, 9, -9, 2, -2, 2, -4, 0, -5,
					-- layer=2 filter=188 channel=14
					0, -20, -20, 3, 9, 4, -6, -3, -4,
					-- layer=2 filter=188 channel=15
					1, 14, -44, 27, 0, -53, 27, 36, 1,
					-- layer=2 filter=188 channel=16
					4, 11, -8, 16, 29, 6, -4, 6, -7,
					-- layer=2 filter=188 channel=17
					-1, -2, 6, -6, 1, 5, 8, -2, -7,
					-- layer=2 filter=188 channel=18
					-15, 4, 6, 7, -28, 19, -18, 0, -30,
					-- layer=2 filter=188 channel=19
					3, 14, -1, 21, 0, -15, 41, 22, 2,
					-- layer=2 filter=188 channel=20
					-6, -8, 0, -8, -6, -10, -7, 3, 2,
					-- layer=2 filter=188 channel=21
					-13, -7, -17, 1, -8, -7, 0, -23, -7,
					-- layer=2 filter=188 channel=22
					7, 5, 0, -5, -5, 9, 0, 10, -4,
					-- layer=2 filter=188 channel=23
					7, 21, 19, 48, 4, -11, 39, 17, -10,
					-- layer=2 filter=188 channel=24
					-7, -6, -36, -35, 4, 0, -17, 13, -32,
					-- layer=2 filter=188 channel=25
					-21, 2, -30, -5, 14, -12, -16, 17, -6,
					-- layer=2 filter=188 channel=26
					4, 7, 2, -8, 0, 6, -5, 2, 7,
					-- layer=2 filter=188 channel=27
					-10, -25, -19, 6, 40, 34, -22, 4, 16,
					-- layer=2 filter=188 channel=28
					48, 34, 24, -10, 24, 9, -20, -5, 17,
					-- layer=2 filter=188 channel=29
					0, -9, 2, -4, 6, 0, -8, 5, -4,
					-- layer=2 filter=188 channel=30
					-28, -32, -6, -18, -5, -5, 25, 1, -25,
					-- layer=2 filter=188 channel=31
					39, -18, 15, -40, 48, 3, 35, 78, 38,
					-- layer=2 filter=188 channel=32
					-4, 10, 4, 10, 0, 0, -9, 4, 6,
					-- layer=2 filter=188 channel=33
					15, 15, 7, -6, 25, 36, -32, -22, 49,
					-- layer=2 filter=188 channel=34
					23, 1, -16, 9, -4, -46, 14, -52, -54,
					-- layer=2 filter=188 channel=35
					35, 29, 14, 14, 33, 1, -23, 21, 27,
					-- layer=2 filter=188 channel=36
					9, -6, 8, -1, 12, 0, -5, -7, 2,
					-- layer=2 filter=188 channel=37
					-11, -26, -10, -13, -15, 0, 2, 4, -7,
					-- layer=2 filter=188 channel=38
					16, -26, -21, 7, -2, -4, -27, -10, -23,
					-- layer=2 filter=188 channel=39
					11, -10, -33, -27, 12, 29, -20, -9, -5,
					-- layer=2 filter=188 channel=40
					29, 17, -26, 7, -11, -46, 34, 1, 4,
					-- layer=2 filter=188 channel=41
					-4, 7, 10, 1, -2, 9, 0, 10, -2,
					-- layer=2 filter=188 channel=42
					27, 12, 6, 19, -11, 5, 7, -11, -13,
					-- layer=2 filter=188 channel=43
					8, 39, -33, -10, 17, 16, 10, -3, 7,
					-- layer=2 filter=188 channel=44
					1, 6, -9, -11, 1, -9, 4, 2, 7,
					-- layer=2 filter=188 channel=45
					-21, 4, -5, 14, 42, -8, -45, -14, 17,
					-- layer=2 filter=188 channel=46
					-37, -37, -14, -22, 9, -14, -38, -26, -12,
					-- layer=2 filter=188 channel=47
					38, 33, 32, 43, 58, 9, -2, 5, 12,
					-- layer=2 filter=188 channel=48
					-4, 2, 5, -1, -5, 7, -11, -6, -9,
					-- layer=2 filter=188 channel=49
					-28, -35, 3, 8, -12, -14, 9, 18, -15,
					-- layer=2 filter=188 channel=50
					0, 7, -7, -2, 12, 31, -5, -8, 18,
					-- layer=2 filter=188 channel=51
					-12, -12, -26, -27, -19, -21, -7, -12, -23,
					-- layer=2 filter=188 channel=52
					-12, -15, -38, 0, -46, 15, 26, 10, 0,
					-- layer=2 filter=188 channel=53
					-83, -34, -62, -38, -57, -113, -3, -4, -52,
					-- layer=2 filter=188 channel=54
					8, 28, 29, -2, 6, 2, 2, -12, 16,
					-- layer=2 filter=188 channel=55
					12, 0, 1, 6, -7, 1, -1, -6, -4,
					-- layer=2 filter=188 channel=56
					-40, -26, -11, -39, 2, 1, -7, -17, -9,
					-- layer=2 filter=188 channel=57
					5, 1, -8, 2, -2, -13, 12, -4, 9,
					-- layer=2 filter=188 channel=58
					0, 9, 15, 71, 5, 25, -3, 38, 31,
					-- layer=2 filter=188 channel=59
					46, -12, -56, 21, -3, 8, -8, -5, -5,
					-- layer=2 filter=188 channel=60
					21, 1, -23, 53, 22, -21, -16, -28, -10,
					-- layer=2 filter=188 channel=61
					-14, -23, -28, 10, 6, -22, 6, 12, -24,
					-- layer=2 filter=188 channel=62
					24, -29, 11, 51, -26, -8, 47, 26, -5,
					-- layer=2 filter=188 channel=63
					15, -9, -12, 40, 20, 4, 0, -12, -8,
					-- layer=2 filter=188 channel=64
					-17, -14, -14, -15, 0, 1, 16, 0, -39,
					-- layer=2 filter=188 channel=65
					-25, -68, -3, 27, -11, 3, 0, 0, -11,
					-- layer=2 filter=188 channel=66
					-11, 28, 61, 0, 35, -33, -45, -47, 17,
					-- layer=2 filter=188 channel=67
					-51, -15, -47, -37, 5, -9, 0, 2, -44,
					-- layer=2 filter=188 channel=68
					-2, -5, 3, 8, -6, 0, -1, 9, 1,
					-- layer=2 filter=188 channel=69
					-17, -15, -16, -12, -9, 2, -1, -21, -7,
					-- layer=2 filter=188 channel=70
					9, 12, 12, 16, 30, -10, -16, -1, 17,
					-- layer=2 filter=188 channel=71
					-39, -55, -55, -5, 21, -8, -24, 7, 12,
					-- layer=2 filter=188 channel=72
					7, 25, 40, 1, 25, -10, -8, -37, -4,
					-- layer=2 filter=188 channel=73
					-9, -7, -22, 38, -47, -33, 17, 44, 87,
					-- layer=2 filter=188 channel=74
					11, -6, -14, -15, -30, 7, -18, -19, -11,
					-- layer=2 filter=188 channel=75
					19, 37, 25, 21, 12, 6, 3, -23, 2,
					-- layer=2 filter=188 channel=76
					-24, -50, -47, 59, -107, -54, -46, 41, -16,
					-- layer=2 filter=188 channel=77
					-9, -6, 3, 0, 6, 12, 2, -3, 0,
					-- layer=2 filter=188 channel=78
					-13, -15, 3, -14, -24, -19, 1, 9, -9,
					-- layer=2 filter=188 channel=79
					-9, 4, -2, -7, 0, 9, 5, 3, -8,
					-- layer=2 filter=188 channel=80
					-18, -4, 5, -2, 8, -10, 4, -20, -15,
					-- layer=2 filter=188 channel=81
					17, 6, 4, 16, 7, 2, 7, 9, 10,
					-- layer=2 filter=188 channel=82
					7, 6, 9, -8, -1, 10, 6, 6, 5,
					-- layer=2 filter=188 channel=83
					-21, -18, 2, 16, 8, -4, 16, 5, 4,
					-- layer=2 filter=188 channel=84
					3, -8, 0, -2, 5, -10, -8, 2, -4,
					-- layer=2 filter=188 channel=85
					-3, 0, -9, 3, 7, -4, 15, 4, -5,
					-- layer=2 filter=188 channel=86
					7, -3, -1, 2, 4, 2, -1, -12, 6,
					-- layer=2 filter=188 channel=87
					-7, -16, -31, 25, -41, -39, -50, -53, -17,
					-- layer=2 filter=188 channel=88
					15, -34, -28, 17, -31, 5, 46, 28, 1,
					-- layer=2 filter=188 channel=89
					5, 1, -10, 29, 17, 5, -8, -21, -2,
					-- layer=2 filter=188 channel=90
					8, -1, 0, 0, 0, 0, -3, 1, 6,
					-- layer=2 filter=188 channel=91
					-31, 0, -2, 19, 19, 6, -36, -12, 27,
					-- layer=2 filter=188 channel=92
					-9, -17, -10, 31, 21, 23, 8, -1, 13,
					-- layer=2 filter=188 channel=93
					0, -49, 4, 46, -12, -11, 21, 0, 33,
					-- layer=2 filter=188 channel=94
					-11, -6, -13, 0, -5, -6, 39, 29, 23,
					-- layer=2 filter=188 channel=95
					0, -2, 3, 13, 8, 7, 6, 3, 15,
					-- layer=2 filter=188 channel=96
					13, -25, -49, 52, -14, -52, 21, 29, 30,
					-- layer=2 filter=188 channel=97
					-11, -14, 1, -22, 14, 0, -18, -39, -11,
					-- layer=2 filter=188 channel=98
					33, 32, 30, 11, 51, 10, -23, -11, -13,
					-- layer=2 filter=188 channel=99
					-3, -41, -38, -2, -70, 0, 29, 25, -20,
					-- layer=2 filter=188 channel=100
					25, 1, -10, 14, 22, 4, 7, 20, -14,
					-- layer=2 filter=188 channel=101
					-12, -12, -9, 14, 14, -3, -14, 37, 14,
					-- layer=2 filter=188 channel=102
					-18, -34, -1, 14, -35, -19, 31, 26, 7,
					-- layer=2 filter=188 channel=103
					-15, -12, 14, -39, -29, 16, -12, 9, 35,
					-- layer=2 filter=188 channel=104
					-55, -68, 17, -36, -107, -35, -26, -21, -26,
					-- layer=2 filter=188 channel=105
					42, 21, 3, 51, 7, -24, -46, -5, -18,
					-- layer=2 filter=188 channel=106
					-48, 18, -35, -15, 0, -9, -39, -9, -5,
					-- layer=2 filter=188 channel=107
					-37, 50, -42, 0, 28, 45, -13, -42, -7,
					-- layer=2 filter=188 channel=108
					0, -65, -42, 18, 31, 11, 0, 28, 0,
					-- layer=2 filter=188 channel=109
					0, -1, 0, 6, 4, -7, 12, 5, 15,
					-- layer=2 filter=188 channel=110
					1, -2, -14, 31, 21, 7, 32, -25, -34,
					-- layer=2 filter=188 channel=111
					-2, -2, 5, 3, 7, 9, 8, -4, 1,
					-- layer=2 filter=188 channel=112
					-46, -20, -17, -47, -8, -14, -22, 16, -23,
					-- layer=2 filter=188 channel=113
					-4, -20, 3, 30, -14, -5, 5, -1, -14,
					-- layer=2 filter=188 channel=114
					-11, -2, -7, -4, 12, -1, -9, 9, 2,
					-- layer=2 filter=188 channel=115
					1, -3, 1, -2, -13, 2, 8, 8, 7,
					-- layer=2 filter=188 channel=116
					0, -2, -31, 33, -24, -49, 11, 5, -20,
					-- layer=2 filter=188 channel=117
					-31, -1, 8, -15, 18, 24, -7, -16, -10,
					-- layer=2 filter=188 channel=118
					-1, -14, -18, 20, 12, 0, 29, -6, 31,
					-- layer=2 filter=188 channel=119
					-18, 22, 15, -3, 32, 48, -40, 5, -21,
					-- layer=2 filter=188 channel=120
					-10, 2, 9, 7, -6, 0, -5, -4, 5,
					-- layer=2 filter=188 channel=121
					6, 0, 0, -6, -6, 2, -3, 9, 5,
					-- layer=2 filter=188 channel=122
					-17, -8, -13, -4, -3, 11, -4, -16, -3,
					-- layer=2 filter=188 channel=123
					4, 16, 24, 9, 33, 14, -18, -8, 0,
					-- layer=2 filter=188 channel=124
					0, 0, -23, -4, -63, 4, 20, -43, -43,
					-- layer=2 filter=188 channel=125
					-8, -7, -1, 3, 6, -3, -8, 8, -3,
					-- layer=2 filter=188 channel=126
					-1, 25, -11, 12, 2, -4, -38, 33, 39,
					-- layer=2 filter=188 channel=127
					0, -19, -3, 6, -12, 20, 14, -10, 17,
					-- layer=2 filter=189 channel=0
					7, 0, -17, 5, -2, -18, 4, 25, -1,
					-- layer=2 filter=189 channel=1
					4, 4, -4, 19, -35, -15, 13, -41, -6,
					-- layer=2 filter=189 channel=2
					0, 9, 0, -1, -7, 3, -6, -4, 9,
					-- layer=2 filter=189 channel=3
					4, -10, 4, 13, 9, 5, 2, -2, 0,
					-- layer=2 filter=189 channel=4
					-10, -89, -29, -29, -9, -4, -36, -54, -41,
					-- layer=2 filter=189 channel=5
					0, 17, 5, 3, 1, 5, -1, 46, 28,
					-- layer=2 filter=189 channel=6
					0, -46, 6, 7, -22, 26, 9, 34, 15,
					-- layer=2 filter=189 channel=7
					-30, 7, -16, -8, -40, -10, -8, -45, 46,
					-- layer=2 filter=189 channel=8
					-7, -3, 6, 0, -5, -10, 5, 4, 7,
					-- layer=2 filter=189 channel=9
					-4, -22, -32, -15, -18, 0, -25, -7, -13,
					-- layer=2 filter=189 channel=10
					14, -22, -17, 31, -9, 1, 25, 26, 9,
					-- layer=2 filter=189 channel=11
					11, 9, 28, 5, 24, 35, 17, 22, 27,
					-- layer=2 filter=189 channel=12
					-13, 0, -18, -10, -55, -37, 12, 1, 49,
					-- layer=2 filter=189 channel=13
					4, 0, -3, -6, -1, -9, -9, 6, -6,
					-- layer=2 filter=189 channel=14
					-13, 13, 10, 7, -7, 11, 11, -3, 11,
					-- layer=2 filter=189 channel=15
					50, 15, 2, 31, -13, -13, -9, -45, 19,
					-- layer=2 filter=189 channel=16
					15, -51, -80, 28, -35, -31, -1, -47, 15,
					-- layer=2 filter=189 channel=17
					-6, 10, 0, 0, 2, -8, 2, 5, 2,
					-- layer=2 filter=189 channel=18
					-34, 10, 30, -29, -1, -11, 7, -9, 18,
					-- layer=2 filter=189 channel=19
					0, -36, 8, -23, -36, 18, 8, 20, 22,
					-- layer=2 filter=189 channel=20
					-5, -1, -5, -4, 9, 7, -3, 0, -5,
					-- layer=2 filter=189 channel=21
					13, 16, 24, 15, 12, 8, 4, 8, 16,
					-- layer=2 filter=189 channel=22
					2, 2, -9, 9, 2, 7, -7, -8, -4,
					-- layer=2 filter=189 channel=23
					-7, -38, -66, -5, -51, -10, -8, 32, 5,
					-- layer=2 filter=189 channel=24
					6, -5, -10, 19, 2, 6, 26, 21, -1,
					-- layer=2 filter=189 channel=25
					7, 10, -8, 31, 23, 21, 27, 9, 28,
					-- layer=2 filter=189 channel=26
					-4, 5, 8, -9, 1, -6, -2, -3, -8,
					-- layer=2 filter=189 channel=27
					12, 6, 22, -5, 13, 4, -7, 0, -16,
					-- layer=2 filter=189 channel=28
					-61, -50, 27, -31, -45, -8, -20, -46, -43,
					-- layer=2 filter=189 channel=29
					-6, 4, -9, -3, -9, 0, 6, 7, 6,
					-- layer=2 filter=189 channel=30
					-13, -27, -12, -6, -41, -22, -14, 3, -11,
					-- layer=2 filter=189 channel=31
					10, -32, -39, 42, -35, -69, -32, 32, 13,
					-- layer=2 filter=189 channel=32
					0, 2, -5, 2, -8, -6, 5, -2, 2,
					-- layer=2 filter=189 channel=33
					48, 30, 42, -20, -14, -29, -8, -44, 25,
					-- layer=2 filter=189 channel=34
					29, -14, 9, -8, -33, 33, -10, -26, -2,
					-- layer=2 filter=189 channel=35
					-30, -53, -16, -37, -51, -11, -6, -38, -29,
					-- layer=2 filter=189 channel=36
					-9, 8, 1, 4, 8, -4, 7, 3, 5,
					-- layer=2 filter=189 channel=37
					14, 22, 33, 11, 31, 29, 8, 23, 12,
					-- layer=2 filter=189 channel=38
					7, 0, 15, -20, -10, 8, -58, -9, -15,
					-- layer=2 filter=189 channel=39
					33, -70, -29, 8, -35, -41, 5, -28, 20,
					-- layer=2 filter=189 channel=40
					-37, -13, -9, 63, -12, -41, 9, -26, -10,
					-- layer=2 filter=189 channel=41
					-2, -7, 11, -8, 11, 0, -6, -3, -11,
					-- layer=2 filter=189 channel=42
					-20, -46, -54, -26, -61, -44, 52, -19, 20,
					-- layer=2 filter=189 channel=43
					-1, -14, 16, -14, 13, 0, 5, 5, -12,
					-- layer=2 filter=189 channel=44
					2, 4, 6, 4, 0, 7, -1, 9, -9,
					-- layer=2 filter=189 channel=45
					-22, -8, -10, 11, 29, -27, -82, -59, -24,
					-- layer=2 filter=189 channel=46
					46, -21, -31, -4, -43, -17, -21, -14, -22,
					-- layer=2 filter=189 channel=47
					-91, -50, -8, -65, -37, -47, -34, -83, -13,
					-- layer=2 filter=189 channel=48
					6, 0, -1, 3, 0, 2, -5, -9, 6,
					-- layer=2 filter=189 channel=49
					16, 30, 33, 17, 31, -3, 40, 13, 5,
					-- layer=2 filter=189 channel=50
					13, 21, 9, -7, 1, 2, 1, 13, 7,
					-- layer=2 filter=189 channel=51
					7, 6, 15, 13, 15, 22, 18, 24, 36,
					-- layer=2 filter=189 channel=52
					20, 18, 12, 12, 21, 39, 22, 13, 45,
					-- layer=2 filter=189 channel=53
					5, -23, 19, -30, 24, 5, -33, 28, 38,
					-- layer=2 filter=189 channel=54
					-35, -19, 0, 29, -14, 35, 18, 55, 41,
					-- layer=2 filter=189 channel=55
					8, 6, 1, -12, -2, 1, 3, -6, -9,
					-- layer=2 filter=189 channel=56
					1, 3, 29, -2, 8, 23, 9, 12, 1,
					-- layer=2 filter=189 channel=57
					-5, -11, 1, -5, 0, -8, -4, 10, -6,
					-- layer=2 filter=189 channel=58
					-10, -5, -22, -11, -27, -27, 10, -20, 42,
					-- layer=2 filter=189 channel=59
					16, -7, 4, 9, -11, 32, -21, -29, 24,
					-- layer=2 filter=189 channel=60
					-12, 12, -26, 11, -49, 27, -28, 27, 41,
					-- layer=2 filter=189 channel=61
					-11, 9, -19, 7, -24, -1, 5, 12, -9,
					-- layer=2 filter=189 channel=62
					-18, 10, 14, -19, 4, 28, 9, 29, 44,
					-- layer=2 filter=189 channel=63
					0, -14, -31, 30, -21, -47, 8, 24, -7,
					-- layer=2 filter=189 channel=64
					-45, -62, -55, 20, -24, -47, 36, 8, -12,
					-- layer=2 filter=189 channel=65
					0, -20, -40, 12, -36, 2, 7, 40, 25,
					-- layer=2 filter=189 channel=66
					-19, 6, 25, -23, 5, -45, 12, -6, -2,
					-- layer=2 filter=189 channel=67
					35, 4, -29, -27, -20, -28, -51, -20, -4,
					-- layer=2 filter=189 channel=68
					9, 0, 8, 1, -7, -1, 8, -7, 1,
					-- layer=2 filter=189 channel=69
					-39, -50, -77, 52, -27, -50, 12, -43, -47,
					-- layer=2 filter=189 channel=70
					-60, -9, -5, -32, -49, -6, 24, 10, 13,
					-- layer=2 filter=189 channel=71
					23, 25, 36, 2, 5, 4, -32, -25, -4,
					-- layer=2 filter=189 channel=72
					-46, 19, 38, -12, 34, 20, 10, -5, 27,
					-- layer=2 filter=189 channel=73
					30, -26, 6, 25, 19, 24, -10, -20, -11,
					-- layer=2 filter=189 channel=74
					35, -9, -28, 5, -13, -29, -22, -30, -31,
					-- layer=2 filter=189 channel=75
					-12, 52, 6, -22, -33, -24, 51, -16, 29,
					-- layer=2 filter=189 channel=76
					-19, -23, -4, 24, 17, 35, -50, -14, 5,
					-- layer=2 filter=189 channel=77
					-1, 8, 5, 7, 10, 7, -2, 8, 5,
					-- layer=2 filter=189 channel=78
					10, -1, 18, 21, 32, 16, 22, 33, 39,
					-- layer=2 filter=189 channel=79
					10, 4, 7, -2, 7, 10, 10, 2, 12,
					-- layer=2 filter=189 channel=80
					25, -36, -18, 20, -22, -32, 31, 20, -63,
					-- layer=2 filter=189 channel=81
					0, 17, 12, 10, 3, 14, 1, 2, 15,
					-- layer=2 filter=189 channel=82
					1, -4, 9, 1, 12, 4, 0, 5, 7,
					-- layer=2 filter=189 channel=83
					19, -60, -27, 20, -19, -27, 30, 35, -19,
					-- layer=2 filter=189 channel=84
					0, 1, 8, -8, 2, 10, -8, 6, 0,
					-- layer=2 filter=189 channel=85
					-9, -3, 5, 11, -6, -7, -7, -4, 0,
					-- layer=2 filter=189 channel=86
					1, 0, -8, 5, 12, 4, -6, 7, 1,
					-- layer=2 filter=189 channel=87
					6, 15, 31, -42, -22, 11, -15, -19, 12,
					-- layer=2 filter=189 channel=88
					4, -2, -25, 17, 6, -33, -26, -59, -36,
					-- layer=2 filter=189 channel=89
					-12, 0, 30, -13, -32, 19, 38, -4, 42,
					-- layer=2 filter=189 channel=90
					1, 2, -7, 0, -9, -3, 0, 8, 6,
					-- layer=2 filter=189 channel=91
					-33, 15, -13, -13, -18, 20, -6, 0, 33,
					-- layer=2 filter=189 channel=92
					-4, 21, 5, 1, -42, -15, 10, -7, 6,
					-- layer=2 filter=189 channel=93
					-27, -18, -13, 7, -27, -21, -11, 39, 14,
					-- layer=2 filter=189 channel=94
					-3, -16, -33, 2, -2, -24, -11, 36, -13,
					-- layer=2 filter=189 channel=95
					-1, -11, -7, -15, -4, -22, -3, -5, -7,
					-- layer=2 filter=189 channel=96
					-31, 38, -4, 22, -2, -12, 26, 24, 51,
					-- layer=2 filter=189 channel=97
					-29, -23, -16, -1, -40, -11, -1, 3, -26,
					-- layer=2 filter=189 channel=98
					-49, 19, 28, 0, -7, 9, 11, -19, -8,
					-- layer=2 filter=189 channel=99
					31, 9, -7, 35, 14, 37, 5, 49, 38,
					-- layer=2 filter=189 channel=100
					7, -19, -9, 10, -43, -36, 8, 20, -19,
					-- layer=2 filter=189 channel=101
					16, 18, 2, 13, 7, 16, -5, -26, 12,
					-- layer=2 filter=189 channel=102
					-34, -29, -14, -12, -25, 2, 46, 5, 39,
					-- layer=2 filter=189 channel=103
					-38, 24, -26, 34, -8, 23, 70, -16, 49,
					-- layer=2 filter=189 channel=104
					-4, 18, 38, -2, 22, 8, -12, 28, -5,
					-- layer=2 filter=189 channel=105
					-10, -1, -36, 2, -15, 36, -16, -58, -22,
					-- layer=2 filter=189 channel=106
					5, -5, 3, 25, -20, -3, -1, -12, 15,
					-- layer=2 filter=189 channel=107
					-6, -11, -10, -58, 0, 8, 22, -41, 14,
					-- layer=2 filter=189 channel=108
					16, 14, 23, -3, -10, 0, 13, -9, -6,
					-- layer=2 filter=189 channel=109
					0, 8, -2, 1, 0, 5, 11, 8, 4,
					-- layer=2 filter=189 channel=110
					-20, -11, -35, -18, -24, -44, 9, -2, 11,
					-- layer=2 filter=189 channel=111
					-1, 6, -4, -8, -9, 12, -4, 4, 12,
					-- layer=2 filter=189 channel=112
					-4, -12, -15, -11, -16, -16, 23, 32, 4,
					-- layer=2 filter=189 channel=113
					8, -26, -15, 14, -34, -54, 4, 34, -24,
					-- layer=2 filter=189 channel=114
					-4, 0, -4, -3, -12, -10, 6, 1, -18,
					-- layer=2 filter=189 channel=115
					9, -9, 9, -2, 2, 7, 4, 7, -5,
					-- layer=2 filter=189 channel=116
					0, 25, 0, -35, -44, -11, -4, -50, 18,
					-- layer=2 filter=189 channel=117
					-18, -13, -48, 23, -34, -16, 0, -15, 22,
					-- layer=2 filter=189 channel=118
					13, 0, 14, -13, 15, 7, 5, -2, 6,
					-- layer=2 filter=189 channel=119
					-53, -45, -73, -46, -53, -50, -27, -58, -9,
					-- layer=2 filter=189 channel=120
					-6, 0, -2, 5, -10, -5, 0, 4, -9,
					-- layer=2 filter=189 channel=121
					-3, -7, -1, -3, 9, -3, 7, 0, -2,
					-- layer=2 filter=189 channel=122
					3, -9, -4, -11, 9, 6, 11, 3, 1,
					-- layer=2 filter=189 channel=123
					-44, 11, -12, -15, -9, -18, -20, -33, 36,
					-- layer=2 filter=189 channel=124
					24, -65, -83, 31, -75, 4, -26, -29, 10,
					-- layer=2 filter=189 channel=125
					-1, 0, 5, -9, -5, 7, 5, -6, -9,
					-- layer=2 filter=189 channel=126
					-64, 0, -12, 4, -23, -48, 28, -1, -13,
					-- layer=2 filter=189 channel=127
					29, -51, -40, -16, -40, -66, 10, -25, -22,
					-- layer=2 filter=190 channel=0
					1, 8, 11, -22, 8, -8, -10, 6, -14,
					-- layer=2 filter=190 channel=1
					-2, 1, -10, -4, 31, 27, 48, 6, 14,
					-- layer=2 filter=190 channel=2
					12, -4, -5, 2, 8, 5, 2, -6, 4,
					-- layer=2 filter=190 channel=3
					12, 14, 1, -32, -21, -17, 13, 32, 40,
					-- layer=2 filter=190 channel=4
					24, -12, 11, -2, 24, -10, -27, 7, -23,
					-- layer=2 filter=190 channel=5
					-9, -8, 3, -10, 1, -15, 3, -4, -21,
					-- layer=2 filter=190 channel=6
					16, -4, 13, -10, -33, 34, -1, -47, 7,
					-- layer=2 filter=190 channel=7
					0, 0, -37, 8, 25, -14, 57, 20, 42,
					-- layer=2 filter=190 channel=8
					0, 0, -7, 8, -1, 4, 8, 4, -3,
					-- layer=2 filter=190 channel=9
					6, 26, -8, -39, 15, 1, -45, -56, 2,
					-- layer=2 filter=190 channel=10
					8, 7, 10, -42, 7, -42, 24, 12, -15,
					-- layer=2 filter=190 channel=11
					12, -12, 0, -4, -6, -13, -10, -12, -4,
					-- layer=2 filter=190 channel=12
					-12, 5, 5, 0, 22, 14, 25, 28, -10,
					-- layer=2 filter=190 channel=13
					2, -4, 4, 1, -6, 0, -1, -6, 2,
					-- layer=2 filter=190 channel=14
					7, 0, -19, 5, 17, 4, 13, 19, -3,
					-- layer=2 filter=190 channel=15
					2, -26, -45, -76, 29, 49, -47, 1, 60,
					-- layer=2 filter=190 channel=16
					39, 31, -7, 11, 12, -8, -35, -58, -62,
					-- layer=2 filter=190 channel=17
					0, 1, 8, 1, -8, 6, -2, 7, 7,
					-- layer=2 filter=190 channel=18
					2, -46, -40, -11, -6, 21, -33, -8, 21,
					-- layer=2 filter=190 channel=19
					-8, 4, -1, -3, 5, -7, 49, 17, -1,
					-- layer=2 filter=190 channel=20
					0, -6, -1, 7, 2, -11, -7, 3, -5,
					-- layer=2 filter=190 channel=21
					-6, 3, 13, 9, 5, 14, 5, 15, 5,
					-- layer=2 filter=190 channel=22
					10, 5, 0, 0, 5, 1, -3, -2, 0,
					-- layer=2 filter=190 channel=23
					31, 37, 7, 2, 1, -14, 2, -11, 18,
					-- layer=2 filter=190 channel=24
					15, 18, 18, -15, -27, -16, -17, -30, -21,
					-- layer=2 filter=190 channel=25
					25, 23, 10, 19, -1, -1, -14, -13, -21,
					-- layer=2 filter=190 channel=26
					-4, 8, 4, -3, 0, 2, 9, -4, 6,
					-- layer=2 filter=190 channel=27
					5, 16, 16, 18, 18, -30, 24, 21, 8,
					-- layer=2 filter=190 channel=28
					14, 24, -42, -4, -13, -39, -1, 10, -10,
					-- layer=2 filter=190 channel=29
					-7, -8, -2, -10, 7, 2, -12, 4, -3,
					-- layer=2 filter=190 channel=30
					-23, 20, 19, -21, -14, -5, -35, -47, -33,
					-- layer=2 filter=190 channel=31
					-46, -23, 16, -65, 33, 40, -42, -15, -80,
					-- layer=2 filter=190 channel=32
					4, 5, 3, 7, 2, 0, -6, -6, -7,
					-- layer=2 filter=190 channel=33
					-51, -47, -61, 2, 14, 11, 0, 42, 28,
					-- layer=2 filter=190 channel=34
					-35, -31, 1, -2, -18, 14, -49, -6, 0,
					-- layer=2 filter=190 channel=35
					-15, 18, -10, -17, -40, -41, -13, 18, -6,
					-- layer=2 filter=190 channel=36
					-9, 0, 11, -12, -8, -13, 10, 20, -1,
					-- layer=2 filter=190 channel=37
					1, 12, 3, 4, 0, 0, 0, -13, -21,
					-- layer=2 filter=190 channel=38
					-10, 15, 20, 1, 7, 8, 29, 25, -2,
					-- layer=2 filter=190 channel=39
					-11, 14, 23, -42, 32, 36, 24, -10, -27,
					-- layer=2 filter=190 channel=40
					18, 1, -30, -12, -19, 10, 6, -4, 19,
					-- layer=2 filter=190 channel=41
					11, 3, 0, 1, 4, 9, 10, 0, -8,
					-- layer=2 filter=190 channel=42
					5, 21, -7, 5, 17, -23, 23, 0, -24,
					-- layer=2 filter=190 channel=43
					-20, 8, -41, -55, -28, -11, -42, 14, 34,
					-- layer=2 filter=190 channel=44
					-9, 1, 9, 6, 4, -10, 7, -6, -4,
					-- layer=2 filter=190 channel=45
					21, 26, 8, 29, 30, -10, 28, 32, 4,
					-- layer=2 filter=190 channel=46
					-2, 15, 26, -48, -3, 21, -36, -16, -2,
					-- layer=2 filter=190 channel=47
					30, 13, -29, 45, -6, -24, 4, 33, -2,
					-- layer=2 filter=190 channel=48
					-6, -9, 4, 0, 7, 1, 11, 0, 3,
					-- layer=2 filter=190 channel=49
					34, -6, -50, -49, 1, -20, 16, -35, -3,
					-- layer=2 filter=190 channel=50
					-2, 0, 4, 5, 10, 11, -14, 3, 6,
					-- layer=2 filter=190 channel=51
					-1, 0, -4, -8, -26, -16, -31, -36, -34,
					-- layer=2 filter=190 channel=52
					-5, -2, 19, 7, 18, 13, -12, -10, -3,
					-- layer=2 filter=190 channel=53
					-31, -16, -29, -15, -15, -69, 67, -48, -59,
					-- layer=2 filter=190 channel=54
					34, 2, -31, 20, 14, 16, 23, 11, 31,
					-- layer=2 filter=190 channel=55
					-9, 14, 6, 1, 10, 8, -5, -5, 9,
					-- layer=2 filter=190 channel=56
					28, -25, 4, -6, 14, -8, -27, -39, -23,
					-- layer=2 filter=190 channel=57
					8, 12, -8, 1, -1, -4, 4, -6, -3,
					-- layer=2 filter=190 channel=58
					-20, -2, -11, 20, 21, 35, 41, 42, 3,
					-- layer=2 filter=190 channel=59
					-70, 0, -8, 0, 7, 21, 24, 36, 40,
					-- layer=2 filter=190 channel=60
					-35, -24, 26, -8, 20, 17, 23, -2, -30,
					-- layer=2 filter=190 channel=61
					-61, -16, -26, -27, -60, -20, -16, -54, -30,
					-- layer=2 filter=190 channel=62
					-5, -25, 19, 3, 20, 41, 1, -14, 12,
					-- layer=2 filter=190 channel=63
					-14, 13, -17, -22, 20, -9, -5, -4, -11,
					-- layer=2 filter=190 channel=64
					17, 38, 17, -26, 20, -25, -4, -17, 7,
					-- layer=2 filter=190 channel=65
					-10, -16, -10, -36, -98, -14, -12, -75, -13,
					-- layer=2 filter=190 channel=66
					21, 5, -33, -54, -31, -20, 4, -9, -5,
					-- layer=2 filter=190 channel=67
					-8, 5, -1, -85, -29, 2, -62, -33, 5,
					-- layer=2 filter=190 channel=68
					-1, 5, 5, -7, 0, 7, 1, 8, -7,
					-- layer=2 filter=190 channel=69
					15, 27, 4, -15, 15, -11, -22, -2, -8,
					-- layer=2 filter=190 channel=70
					6, 12, -3, 30, 10, 2, 16, 25, 6,
					-- layer=2 filter=190 channel=71
					-5, 8, -14, 0, 19, -30, 19, 13, -1,
					-- layer=2 filter=190 channel=72
					32, -1, -28, 21, 7, 13, 24, 21, 25,
					-- layer=2 filter=190 channel=73
					-32, 11, -12, -9, -24, -11, -5, -25, -35,
					-- layer=2 filter=190 channel=74
					-3, 23, 8, -45, -32, 1, -65, -20, -12,
					-- layer=2 filter=190 channel=75
					15, -12, 11, 24, 14, -36, 18, -34, -36,
					-- layer=2 filter=190 channel=76
					-44, -34, -22, -29, -32, 31, -13, -12, -4,
					-- layer=2 filter=190 channel=77
					-8, -2, 0, 3, -5, 9, -6, -2, 9,
					-- layer=2 filter=190 channel=78
					18, -29, -15, -8, 8, 17, -37, -33, -28,
					-- layer=2 filter=190 channel=79
					3, 0, 0, -7, 0, 8, 2, -1, -7,
					-- layer=2 filter=190 channel=80
					40, 26, 26, -17, 12, 4, -18, 2, -7,
					-- layer=2 filter=190 channel=81
					19, 16, 15, 0, 10, -1, 13, -7, 4,
					-- layer=2 filter=190 channel=82
					-9, 11, 8, -3, -1, 8, 6, 11, 1,
					-- layer=2 filter=190 channel=83
					0, 28, 6, -3, -7, -6, 7, 7, -44,
					-- layer=2 filter=190 channel=84
					6, -3, -4, 0, -3, 6, 8, 0, 1,
					-- layer=2 filter=190 channel=85
					7, 8, 8, 5, -3, 15, 13, -1, 6,
					-- layer=2 filter=190 channel=86
					-3, -2, 5, 1, -4, 17, 0, -5, -10,
					-- layer=2 filter=190 channel=87
					-53, -57, -18, -15, 1, -20, -48, 0, 37,
					-- layer=2 filter=190 channel=88
					9, 8, 6, -7, 19, 18, -73, 2, -31,
					-- layer=2 filter=190 channel=89
					-6, -5, 3, -3, 31, 20, 29, 5, 13,
					-- layer=2 filter=190 channel=90
					-7, 1, 7, -1, 9, -3, 8, -4, 5,
					-- layer=2 filter=190 channel=91
					-12, 24, 26, 14, 44, 20, 38, 27, -36,
					-- layer=2 filter=190 channel=92
					-15, 16, 2, 2, 16, 27, 27, 12, 8,
					-- layer=2 filter=190 channel=93
					31, -8, -17, -38, 5, -28, 28, -13, -37,
					-- layer=2 filter=190 channel=94
					-40, -38, -19, 10, -2, -12, 54, -49, 7,
					-- layer=2 filter=190 channel=95
					3, -3, 2, -12, -8, -14, 0, -9, -1,
					-- layer=2 filter=190 channel=96
					19, -9, 31, 58, 14, -9, 34, 15, 20,
					-- layer=2 filter=190 channel=97
					17, 37, 0, -12, 4, 11, -42, -11, -22,
					-- layer=2 filter=190 channel=98
					16, 0, -25, 1, -21, -10, -16, 16, 12,
					-- layer=2 filter=190 channel=99
					-34, 1, 8, 2, -21, -22, 13, 5, 0,
					-- layer=2 filter=190 channel=100
					18, 9, 2, -6, -13, -35, 28, 30, 10,
					-- layer=2 filter=190 channel=101
					-18, -8, -13, 5, 13, -48, 3, -4, -13,
					-- layer=2 filter=190 channel=102
					19, -21, 10, 5, -37, -17, 13, -4, -23,
					-- layer=2 filter=190 channel=103
					-19, 64, -9, -5, 18, 21, 2, -13, -70,
					-- layer=2 filter=190 channel=104
					23, -54, -28, -7, 6, 4, 35, -43, -8,
					-- layer=2 filter=190 channel=105
					20, -3, -5, 18, 33, 2, 1, -48, -16,
					-- layer=2 filter=190 channel=106
					-14, 9, -6, 37, 22, 19, -3, 3, -25,
					-- layer=2 filter=190 channel=107
					33, 35, 9, 0, -37, -24, -3, -68, -37,
					-- layer=2 filter=190 channel=108
					13, 12, -8, 3, 3, -8, 47, -5, -17,
					-- layer=2 filter=190 channel=109
					4, -3, -4, -4, 13, -7, 8, -4, -1,
					-- layer=2 filter=190 channel=110
					17, 21, -1, -4, 8, 5, -10, -20, -7,
					-- layer=2 filter=190 channel=111
					9, 8, -11, -7, 2, -9, 3, 0, 4,
					-- layer=2 filter=190 channel=112
					-15, -2, 31, -28, -21, -16, 9, -18, -37,
					-- layer=2 filter=190 channel=113
					2, 13, -6, -39, -40, -18, 1, -26, -38,
					-- layer=2 filter=190 channel=114
					-6, -9, -3, -16, -7, -16, 2, -3, -5,
					-- layer=2 filter=190 channel=115
					-1, -3, -3, -9, 2, 2, -3, -4, -5,
					-- layer=2 filter=190 channel=116
					-19, -44, -22, -8, -28, 2, -48, 17, 23,
					-- layer=2 filter=190 channel=117
					28, -17, -44, -2, -4, -17, 33, 14, -1,
					-- layer=2 filter=190 channel=118
					14, 8, -7, -33, 15, 8, -64, -3, 41,
					-- layer=2 filter=190 channel=119
					52, -23, -31, 25, 12, 1, 0, -5, 3,
					-- layer=2 filter=190 channel=120
					0, -3, -6, -3, 10, 7, 5, 7, 1,
					-- layer=2 filter=190 channel=121
					1, 7, -1, 0, 4, -4, -4, 3, -7,
					-- layer=2 filter=190 channel=122
					5, -2, 10, -3, -3, 4, -16, -4, -6,
					-- layer=2 filter=190 channel=123
					-2, -11, -54, 10, -1, -6, 20, 25, 46,
					-- layer=2 filter=190 channel=124
					-43, -16, -41, -16, 23, 35, -6, 27, 30,
					-- layer=2 filter=190 channel=125
					3, 9, 12, -2, -8, -1, 6, 7, 9,
					-- layer=2 filter=190 channel=126
					-61, 23, 1, -35, 8, -30, 13, -11, 27,
					-- layer=2 filter=190 channel=127
					3, 15, -26, 5, 7, 4, 21, 25, -12,
					-- layer=2 filter=191 channel=0
					-23, 10, 2, -18, 10, 8, 3, -24, -10,
					-- layer=2 filter=191 channel=1
					-12, -27, -5, 36, -18, -22, 5, -4, -6,
					-- layer=2 filter=191 channel=2
					10, 4, -6, -3, 0, -1, 3, -3, 1,
					-- layer=2 filter=191 channel=3
					-28, -2, 0, -15, 2, 2, -16, 0, 12,
					-- layer=2 filter=191 channel=4
					-10, 16, 35, -11, 19, 34, -20, -32, -19,
					-- layer=2 filter=191 channel=5
					-12, -14, -19, -3, -1, -14, 0, 16, 6,
					-- layer=2 filter=191 channel=6
					-12, 0, 42, -9, 3, -7, 33, 6, -5,
					-- layer=2 filter=191 channel=7
					-21, -27, 3, -26, -23, -38, -13, -16, -34,
					-- layer=2 filter=191 channel=8
					4, 8, 8, -8, 7, -7, 0, 4, 3,
					-- layer=2 filter=191 channel=9
					7, 0, 18, 20, 17, 40, 2, 1, 46,
					-- layer=2 filter=191 channel=10
					-23, 10, 4, -29, -8, 17, -8, 1, -1,
					-- layer=2 filter=191 channel=11
					14, -11, -13, 34, -9, -12, 15, 8, -7,
					-- layer=2 filter=191 channel=12
					15, -2, 12, 25, -33, -34, 6, -7, -5,
					-- layer=2 filter=191 channel=13
					5, 9, 2, 6, 10, 6, 3, 0, 9,
					-- layer=2 filter=191 channel=14
					0, -38, -23, 29, 7, -21, 33, 16, 17,
					-- layer=2 filter=191 channel=15
					1, 4, -24, 17, 17, 25, 26, -2, -26,
					-- layer=2 filter=191 channel=16
					-22, -2, 3, 15, 45, 5, -61, -1, -8,
					-- layer=2 filter=191 channel=17
					0, 3, 1, -3, -4, -4, 2, -2, -8,
					-- layer=2 filter=191 channel=18
					43, 47, 22, 71, 51, 2, 43, 46, -8,
					-- layer=2 filter=191 channel=19
					11, -5, 12, -7, 16, 3, -10, -7, -8,
					-- layer=2 filter=191 channel=20
					-8, 9, 0, -5, 8, -7, 1, -9, 4,
					-- layer=2 filter=191 channel=21
					0, 7, 15, -9, -1, -5, 16, 7, 7,
					-- layer=2 filter=191 channel=22
					9, -2, 0, -10, -1, 6, -6, -4, 8,
					-- layer=2 filter=191 channel=23
					-13, 4, 40, -36, 0, 35, -51, -11, 0,
					-- layer=2 filter=191 channel=24
					-16, -9, -23, -20, 0, 16, -5, -10, 10,
					-- layer=2 filter=191 channel=25
					12, -28, -36, 7, -2, -14, 13, -12, -15,
					-- layer=2 filter=191 channel=26
					-6, 8, -9, -8, -10, -2, -5, -5, 0,
					-- layer=2 filter=191 channel=27
					18, -30, -64, 8, -37, -32, 19, -4, -8,
					-- layer=2 filter=191 channel=28
					3, 14, 11, 10, -47, -19, 1, 2, -30,
					-- layer=2 filter=191 channel=29
					4, -5, -6, 6, 0, -1, -3, -3, 3,
					-- layer=2 filter=191 channel=30
					-22, 1, 10, -35, 5, 7, -34, -18, 20,
					-- layer=2 filter=191 channel=31
					-9, -10, 11, -27, -23, 81, -55, -21, 77,
					-- layer=2 filter=191 channel=32
					11, 5, 7, 2, 6, 6, -6, -5, -7,
					-- layer=2 filter=191 channel=33
					25, -3, -28, 27, 32, 32, -2, 3, -40,
					-- layer=2 filter=191 channel=34
					2, 29, -18, 29, -3, -2, 22, 14, -16,
					-- layer=2 filter=191 channel=35
					10, 38, 25, 41, -29, -13, 34, -20, -28,
					-- layer=2 filter=191 channel=36
					-7, 15, 10, -6, 10, -1, 1, -3, -2,
					-- layer=2 filter=191 channel=37
					27, -23, -30, 28, -2, -15, 25, 28, 2,
					-- layer=2 filter=191 channel=38
					-21, -19, -31, 21, -18, 3, 22, -1, 18,
					-- layer=2 filter=191 channel=39
					-1, 0, 13, -11, 22, 2, -28, -37, 0,
					-- layer=2 filter=191 channel=40
					-12, -12, -36, 5, 0, 32, -38, 2, 22,
					-- layer=2 filter=191 channel=41
					3, 11, 6, -1, 0, -7, 4, -6, -2,
					-- layer=2 filter=191 channel=42
					17, 19, 3, -10, 3, 0, -8, 4, 12,
					-- layer=2 filter=191 channel=43
					8, 11, 17, 12, -10, -34, -9, 9, -30,
					-- layer=2 filter=191 channel=44
					-7, -4, 9, 2, -4, -2, 2, -4, 6,
					-- layer=2 filter=191 channel=45
					40, 29, -18, 9, 2, 13, 30, -10, 32,
					-- layer=2 filter=191 channel=46
					-5, 9, 24, 4, 1, 9, -24, -11, 2,
					-- layer=2 filter=191 channel=47
					-23, -22, -14, 27, -6, 28, -21, -3, -10,
					-- layer=2 filter=191 channel=48
					-5, -6, -9, -1, 4, 5, 2, 4, 7,
					-- layer=2 filter=191 channel=49
					-5, 19, 10, 12, 42, -6, 20, 7, -12,
					-- layer=2 filter=191 channel=50
					-7, 0, -8, -6, -3, -2, 8, -2, 7,
					-- layer=2 filter=191 channel=51
					5, -16, -14, 20, -15, -12, 21, -6, 0,
					-- layer=2 filter=191 channel=52
					-18, -13, -21, 6, -18, -25, -20, -31, 0,
					-- layer=2 filter=191 channel=53
					-45, -19, -16, 36, -41, -38, 21, -10, 22,
					-- layer=2 filter=191 channel=54
					-13, -12, -21, 9, -11, 2, 13, -14, -7,
					-- layer=2 filter=191 channel=55
					12, -2, 5, -2, 6, -2, 14, 1, -9,
					-- layer=2 filter=191 channel=56
					4, -12, -16, 19, -5, -18, 25, 17, 8,
					-- layer=2 filter=191 channel=57
					6, 11, -2, 12, 16, 10, -2, 12, -2,
					-- layer=2 filter=191 channel=58
					34, 8, 21, 9, -9, -43, 7, -35, -39,
					-- layer=2 filter=191 channel=59
					-1, -13, 19, 35, 11, 13, 10, 0, -27,
					-- layer=2 filter=191 channel=60
					-8, -2, -5, 3, 2, -4, 44, 18, -18,
					-- layer=2 filter=191 channel=61
					28, -23, 34, -49, 41, -15, 7, 20, 5,
					-- layer=2 filter=191 channel=62
					13, 8, 29, 57, 2, -10, 35, 6, -41,
					-- layer=2 filter=191 channel=63
					0, -6, 15, -35, 27, 19, -39, 6, -11,
					-- layer=2 filter=191 channel=64
					-32, -2, 14, -34, 36, 28, -42, -7, 21,
					-- layer=2 filter=191 channel=65
					14, 16, 35, -30, 9, 11, 6, 38, 5,
					-- layer=2 filter=191 channel=66
					-7, -16, -17, -9, -2, 9, 35, 5, -52,
					-- layer=2 filter=191 channel=67
					-2, 10, 13, -11, -13, 25, -28, -27, 12,
					-- layer=2 filter=191 channel=68
					-4, 3, 8, -2, -1, 0, -3, -2, 7,
					-- layer=2 filter=191 channel=69
					-21, -10, 2, 12, 29, 13, -16, 27, 21,
					-- layer=2 filter=191 channel=70
					8, 2, -8, 0, -10, 4, 12, -11, -37,
					-- layer=2 filter=191 channel=71
					47, -29, -29, 18, -13, -16, 16, -5, -25,
					-- layer=2 filter=191 channel=72
					30, -14, 0, 6, -15, 2, 1, 41, 5,
					-- layer=2 filter=191 channel=73
					-43, 3, 9, -51, 0, 8, -13, -21, 13,
					-- layer=2 filter=191 channel=74
					-17, 15, 6, -27, 6, 31, -62, -17, 3,
					-- layer=2 filter=191 channel=75
					-13, -35, -39, 28, 3, -34, -20, 0, -67,
					-- layer=2 filter=191 channel=76
					17, -30, -20, -5, -14, -44, 7, 14, -11,
					-- layer=2 filter=191 channel=77
					-3, -7, -8, -6, -7, 7, 5, -3, 5,
					-- layer=2 filter=191 channel=78
					-4, -10, 5, 15, -3, -29, 20, -8, -11,
					-- layer=2 filter=191 channel=79
					-8, -8, -6, 8, -3, -4, -5, -7, -8,
					-- layer=2 filter=191 channel=80
					-12, 4, 25, -43, -1, 16, -46, -7, -13,
					-- layer=2 filter=191 channel=81
					5, 9, 9, -5, -5, -8, 2, 9, -6,
					-- layer=2 filter=191 channel=82
					-3, 7, -7, -4, 5, 0, -10, 0, -1,
					-- layer=2 filter=191 channel=83
					12, -8, 21, -38, 4, 14, -54, -27, -11,
					-- layer=2 filter=191 channel=84
					0, 0, -3, 2, 4, 7, 10, -6, 3,
					-- layer=2 filter=191 channel=85
					-5, -1, -5, 0, -17, -13, -3, -12, -6,
					-- layer=2 filter=191 channel=86
					-5, 8, -10, -10, 7, 9, 6, -2, 0,
					-- layer=2 filter=191 channel=87
					13, 35, 25, 23, -20, -21, 10, -14, -51,
					-- layer=2 filter=191 channel=88
					-24, -4, 15, -9, 3, 37, -55, -13, 14,
					-- layer=2 filter=191 channel=89
					3, -23, -7, 29, -8, -40, 21, 5, 0,
					-- layer=2 filter=191 channel=90
					-9, 3, 6, -2, 0, -3, 4, -6, 0,
					-- layer=2 filter=191 channel=91
					73, 0, 3, 19, -26, -54, 27, -12, -33,
					-- layer=2 filter=191 channel=92
					31, -24, -1, 29, -43, -31, 23, 15, 0,
					-- layer=2 filter=191 channel=93
					3, 22, 50, 34, 19, 10, 38, 0, -31,
					-- layer=2 filter=191 channel=94
					-24, -15, 9, -23, 6, 6, -1, 37, -27,
					-- layer=2 filter=191 channel=95
					-13, 6, 0, -6, 2, -10, -2, 6, -5,
					-- layer=2 filter=191 channel=96
					-74, -17, 29, -28, -27, 21, -24, -18, -10,
					-- layer=2 filter=191 channel=97
					8, -10, -20, 17, 68, 25, -24, -19, 30,
					-- layer=2 filter=191 channel=98
					-12, 9, -15, 14, -52, -7, 7, 15, 0,
					-- layer=2 filter=191 channel=99
					2, -41, -6, 23, 23, -2, -5, -22, 35,
					-- layer=2 filter=191 channel=100
					-4, 6, -18, -33, -47, -6, -20, -24, -26,
					-- layer=2 filter=191 channel=101
					49, 2, -35, 21, -8, -21, 51, -7, 4,
					-- layer=2 filter=191 channel=102
					2, 40, 0, 18, 21, 10, 17, -9, 8,
					-- layer=2 filter=191 channel=103
					12, -8, -9, 17, -22, 9, 17, 39, -7,
					-- layer=2 filter=191 channel=104
					22, 32, 32, 19, 4, 4, 36, 8, -1,
					-- layer=2 filter=191 channel=105
					21, 16, -7, -16, -50, -32, -14, 39, -28,
					-- layer=2 filter=191 channel=106
					21, -10, 0, 24, -16, -11, 44, -9, -5,
					-- layer=2 filter=191 channel=107
					-35, -29, 32, -37, -15, 22, 40, -5, 22,
					-- layer=2 filter=191 channel=108
					-8, -12, -52, 0, -24, -44, 31, -26, -21,
					-- layer=2 filter=191 channel=109
					1, 4, 15, -4, -2, -2, -7, -6, 8,
					-- layer=2 filter=191 channel=110
					-12, 0, 16, -22, -18, 27, -49, -14, 13,
					-- layer=2 filter=191 channel=111
					3, 0, -9, 0, 8, -11, 0, -8, 6,
					-- layer=2 filter=191 channel=112
					32, -7, -4, -17, 5, -1, 11, -10, 3,
					-- layer=2 filter=191 channel=113
					1, 0, 12, -22, -8, 16, -48, -9, 37,
					-- layer=2 filter=191 channel=114
					10, 3, 8, 1, 4, 7, -16, -1, -6,
					-- layer=2 filter=191 channel=115
					4, 0, 4, 13, 4, 5, -1, 3, -2,
					-- layer=2 filter=191 channel=116
					-3, 19, 34, 19, -11, -11, 7, 0, -54,
					-- layer=2 filter=191 channel=117
					-14, 15, 0, -29, 0, 11, -12, -1, 27,
					-- layer=2 filter=191 channel=118
					11, 27, 30, -9, 1, -7, -1, 4, -34,
					-- layer=2 filter=191 channel=119
					7, 0, 4, 34, 35, 22, 10, 21, -26,
					-- layer=2 filter=191 channel=120
					3, -4, 2, -10, -4, 3, 3, 1, 4,
					-- layer=2 filter=191 channel=121
					1, 7, -8, 0, 8, 10, -3, 2, -7,
					-- layer=2 filter=191 channel=122
					-1, 17, 6, 7, 10, 13, 7, -9, 11,
					-- layer=2 filter=191 channel=123
					-19, -17, 30, 0, -10, -3, -16, 14, 3,
					-- layer=2 filter=191 channel=124
					-17, -18, 8, 0, -16, -6, -8, -38, -12,
					-- layer=2 filter=191 channel=125
					2, -9, 5, -6, 0, 6, 1, -7, 5,
					-- layer=2 filter=191 channel=126
					61, -53, -10, 64, -11, -2, 27, 11, -21,
					-- layer=2 filter=191 channel=127
					-11, 5, 10, -23, 28, 0, 2, 9, 23,
					-- layer=2 filter=192 channel=0
					19, 22, -16, -8, -30, -51, 26, 19, -2,
					-- layer=2 filter=192 channel=1
					-40, -9, 5, 16, -5, 19, 4, 33, 30,
					-- layer=2 filter=192 channel=2
					2, -1, 10, -8, 5, -3, 6, 8, 1,
					-- layer=2 filter=192 channel=3
					8, 10, -21, 15, 2, -20, 36, 8, 18,
					-- layer=2 filter=192 channel=4
					-2, 26, 2, 2, 9, 7, -20, -27, -7,
					-- layer=2 filter=192 channel=5
					20, 20, -1, 18, -28, -67, 39, 0, -9,
					-- layer=2 filter=192 channel=6
					16, 20, -3, 13, -12, -33, 6, -30, 21,
					-- layer=2 filter=192 channel=7
					15, 33, 15, -11, 39, 26, 4, 22, 4,
					-- layer=2 filter=192 channel=8
					0, -11, -3, -5, -4, 8, 9, -4, -2,
					-- layer=2 filter=192 channel=9
					-5, 0, 22, -45, -45, -24, -10, -66, -10,
					-- layer=2 filter=192 channel=10
					7, -3, -19, 0, -21, -37, 49, 19, 6,
					-- layer=2 filter=192 channel=11
					18, -2, -18, 23, -15, -28, 13, -29, -42,
					-- layer=2 filter=192 channel=12
					-10, 12, 9, 5, 14, -8, -1, 34, -7,
					-- layer=2 filter=192 channel=13
					4, 3, 6, 8, 9, 9, 8, -3, 2,
					-- layer=2 filter=192 channel=14
					-35, -11, 3, 10, -9, -34, -39, -6, -60,
					-- layer=2 filter=192 channel=15
					17, -23, -3, 45, -12, 6, -16, -9, 13,
					-- layer=2 filter=192 channel=16
					-51, -2, 28, -95, -28, -23, -99, -44, -28,
					-- layer=2 filter=192 channel=17
					-7, -7, -9, -3, -3, -10, -4, 9, 1,
					-- layer=2 filter=192 channel=18
					21, -16, -6, 31, -23, 23, 1, 15, 18,
					-- layer=2 filter=192 channel=19
					2, 3, 10, 14, 38, -5, 12, 17, 13,
					-- layer=2 filter=192 channel=20
					-10, 3, 10, 1, 6, 11, -6, 4, 0,
					-- layer=2 filter=192 channel=21
					3, 6, 0, 0, 0, 14, 12, 8, 20,
					-- layer=2 filter=192 channel=22
					-5, 7, -2, -4, 1, 4, -8, -10, 9,
					-- layer=2 filter=192 channel=23
					-5, -9, -2, -23, 21, 8, -68, -20, -3,
					-- layer=2 filter=192 channel=24
					3, 24, 32, -10, 14, -14, 19, 1, -5,
					-- layer=2 filter=192 channel=25
					23, 40, 29, 7, 15, -12, 25, -6, -48,
					-- layer=2 filter=192 channel=26
					5, -6, -11, 1, 0, 9, -3, 0, -8,
					-- layer=2 filter=192 channel=27
					-24, 12, 8, 29, 0, -62, -3, -49, -87,
					-- layer=2 filter=192 channel=28
					5, 9, 6, -1, -10, -26, 19, 3, 11,
					-- layer=2 filter=192 channel=29
					0, 2, -10, 5, 0, 2, 0, 0, -8,
					-- layer=2 filter=192 channel=30
					5, -19, -1, -40, -62, -7, 4, -44, 37,
					-- layer=2 filter=192 channel=31
					-8, -45, 8, 43, 15, 17, -43, -49, -47,
					-- layer=2 filter=192 channel=32
					-8, 1, -11, 3, -9, 7, -7, -5, 5,
					-- layer=2 filter=192 channel=33
					-23, 0, -45, 36, 33, 22, 6, 37, -10,
					-- layer=2 filter=192 channel=34
					36, 27, 6, 19, 45, -8, 4, 35, 2,
					-- layer=2 filter=192 channel=35
					9, 10, 10, 40, 0, -4, 33, -4, 8,
					-- layer=2 filter=192 channel=36
					8, -4, -3, -10, 4, 5, 5, -7, -4,
					-- layer=2 filter=192 channel=37
					19, -6, -12, 35, 13, -32, 2, -14, -46,
					-- layer=2 filter=192 channel=38
					-5, 30, -7, 41, -28, -2, -10, -17, -27,
					-- layer=2 filter=192 channel=39
					-5, 37, 61, 17, 52, 15, -17, -38, -6,
					-- layer=2 filter=192 channel=40
					6, 16, -73, 21, -26, -33, -32, 31, -4,
					-- layer=2 filter=192 channel=41
					8, 6, -1, -1, 7, -2, 1, 0, -1,
					-- layer=2 filter=192 channel=42
					5, -4, 35, -35, 28, 43, -69, -6, 14,
					-- layer=2 filter=192 channel=43
					-6, 25, -74, 46, -17, -72, 29, 41, 27,
					-- layer=2 filter=192 channel=44
					5, -8, -8, 3, 5, 13, 6, 3, -1,
					-- layer=2 filter=192 channel=45
					-15, 11, 21, 5, -32, -92, -9, -37, -28,
					-- layer=2 filter=192 channel=46
					18, -28, -2, 13, -33, -31, 18, 7, 12,
					-- layer=2 filter=192 channel=47
					-51, -13, -40, -70, -19, 3, -34, 28, 14,
					-- layer=2 filter=192 channel=48
					-6, 0, 8, 0, 5, 4, -8, 5, 2,
					-- layer=2 filter=192 channel=49
					0, -16, 5, -9, -11, 35, 4, -6, -6,
					-- layer=2 filter=192 channel=50
					-18, 0, -2, 18, -7, -4, 13, 12, -4,
					-- layer=2 filter=192 channel=51
					-9, -4, -38, 17, -26, -14, 16, -18, -32,
					-- layer=2 filter=192 channel=52
					0, -14, -12, 43, -28, 7, -15, -38, -14,
					-- layer=2 filter=192 channel=53
					-24, 4, -22, 25, -16, -17, 21, -36, -53,
					-- layer=2 filter=192 channel=54
					14, 8, -10, 15, 21, 20, 23, 22, 21,
					-- layer=2 filter=192 channel=55
					-7, 0, 11, -1, 5, 4, 10, 0, 10,
					-- layer=2 filter=192 channel=56
					14, 1, 4, 12, -3, -43, 0, -28, -46,
					-- layer=2 filter=192 channel=57
					0, 14, 1, -10, -4, 7, -4, -15, 0,
					-- layer=2 filter=192 channel=58
					4, 28, 38, 3, 37, 21, -5, 58, 24,
					-- layer=2 filter=192 channel=59
					-38, 36, 9, 40, 53, -5, 1, 34, -31,
					-- layer=2 filter=192 channel=60
					13, 22, -7, 30, 23, 29, 34, 51, 30,
					-- layer=2 filter=192 channel=61
					16, -14, 6, -37, -16, 0, 3, -8, 22,
					-- layer=2 filter=192 channel=62
					15, -35, -27, 7, -6, -7, 42, 0, 14,
					-- layer=2 filter=192 channel=63
					-11, 7, 12, -25, 0, 14, 8, 34, -19,
					-- layer=2 filter=192 channel=64
					-8, -12, 38, -55, 19, 24, -72, -3, 14,
					-- layer=2 filter=192 channel=65
					17, -29, -32, 16, -15, -16, 11, -23, 15,
					-- layer=2 filter=192 channel=66
					-27, -45, -19, -40, -7, -6, 14, 8, 40,
					-- layer=2 filter=192 channel=67
					3, 2, 2, 11, -66, -37, 32, 2, -4,
					-- layer=2 filter=192 channel=68
					7, -3, 7, -3, -9, 7, -5, -6, -8,
					-- layer=2 filter=192 channel=69
					-31, -3, 27, -29, 45, 59, -75, 12, 48,
					-- layer=2 filter=192 channel=70
					37, 9, 11, 28, 11, 18, 34, 25, -5,
					-- layer=2 filter=192 channel=71
					-5, 27, -1, 36, 5, -41, 5, -25, -71,
					-- layer=2 filter=192 channel=72
					-7, 17, 12, -9, 5, 5, 27, 24, -11,
					-- layer=2 filter=192 channel=73
					-3, 32, 20, -19, 29, 21, -35, -10, 7,
					-- layer=2 filter=192 channel=74
					-11, 9, 13, 11, 8, 14, -4, 21, -14,
					-- layer=2 filter=192 channel=75
					-74, -86, -5, -32, -10, -16, 23, -6, 0,
					-- layer=2 filter=192 channel=76
					10, -63, -32, -26, -11, -13, 11, -75, -27,
					-- layer=2 filter=192 channel=77
					-2, -6, 7, -9, 5, 4, -10, 8, 0,
					-- layer=2 filter=192 channel=78
					13, -20, -11, 18, -21, -9, 15, -20, -5,
					-- layer=2 filter=192 channel=79
					-8, 1, -4, 1, -1, -9, 0, -5, 2,
					-- layer=2 filter=192 channel=80
					-18, -12, -11, -44, -12, -25, -54, -44, -58,
					-- layer=2 filter=192 channel=81
					19, 18, 18, 23, 3, 26, 7, 17, 14,
					-- layer=2 filter=192 channel=82
					9, 2, -10, -3, 8, 2, 1, 3, 5,
					-- layer=2 filter=192 channel=83
					-16, 8, 30, -16, -26, 10, 2, -4, 0,
					-- layer=2 filter=192 channel=84
					4, -2, -1, 4, -3, -10, 4, 0, 3,
					-- layer=2 filter=192 channel=85
					0, 4, -4, 3, 0, 6, -3, 3, 9,
					-- layer=2 filter=192 channel=86
					0, -6, 1, 16, -1, 6, 2, 1, -9,
					-- layer=2 filter=192 channel=87
					36, 3, -12, 51, -9, 20, 26, 21, 40,
					-- layer=2 filter=192 channel=88
					-10, -12, 21, -17, -28, 22, -20, 3, -6,
					-- layer=2 filter=192 channel=89
					-35, 11, 5, 23, 7, 0, -23, 12, -12,
					-- layer=2 filter=192 channel=90
					1, 7, -7, 0, 9, 7, 0, 0, -6,
					-- layer=2 filter=192 channel=91
					6, 10, 33, 9, 44, 13, 29, 32, 0,
					-- layer=2 filter=192 channel=92
					-21, 23, 29, 19, -6, 10, -23, 23, 4,
					-- layer=2 filter=192 channel=93
					17, -1, -41, 21, 0, -42, 9, -13, 20,
					-- layer=2 filter=192 channel=94
					-39, -37, -15, -34, -23, -13, -16, -11, 13,
					-- layer=2 filter=192 channel=95
					14, 13, 0, 10, -6, -4, -5, -3, 6,
					-- layer=2 filter=192 channel=96
					-24, -24, -2, -40, -11, -17, -61, -33, -12,
					-- layer=2 filter=192 channel=97
					4, -18, 6, -21, -5, -14, -22, -6, -21,
					-- layer=2 filter=192 channel=98
					-10, -27, -10, -39, -7, 0, 17, 8, 16,
					-- layer=2 filter=192 channel=99
					15, 1, 22, 45, 50, -4, 12, -29, -4,
					-- layer=2 filter=192 channel=100
					2, 24, 2, -10, 13, -23, 23, 45, 11,
					-- layer=2 filter=192 channel=101
					24, 10, -5, 7, 4, -33, -1, -12, -61,
					-- layer=2 filter=192 channel=102
					20, -22, 4, 11, -8, -13, -13, -11, 5,
					-- layer=2 filter=192 channel=103
					7, -3, -11, 9, -41, 5, 51, 15, -24,
					-- layer=2 filter=192 channel=104
					16, 0, -32, 7, -12, 24, 3, -20, 0,
					-- layer=2 filter=192 channel=105
					3, 20, 11, -7, -28, 23, 23, 2, -36,
					-- layer=2 filter=192 channel=106
					11, 22, 20, 6, 7, -24, 34, 1, -37,
					-- layer=2 filter=192 channel=107
					-3, -53, 46, -11, -15, 37, 25, -1, 12,
					-- layer=2 filter=192 channel=108
					-18, 25, -3, 8, -8, -39, 10, -46, -33,
					-- layer=2 filter=192 channel=109
					-12, 4, -17, 0, 0, -3, 3, 2, 11,
					-- layer=2 filter=192 channel=110
					11, 16, 54, -33, 14, 49, -69, 7, 14,
					-- layer=2 filter=192 channel=111
					4, -5, -4, 1, 0, 7, 9, -9, 3,
					-- layer=2 filter=192 channel=112
					33, 10, -17, 18, -1, -8, 28, 6, -2,
					-- layer=2 filter=192 channel=113
					6, -16, 14, -16, -24, 20, -21, -32, 14,
					-- layer=2 filter=192 channel=114
					2, -4, 0, -8, -4, -5, -15, -4, -2,
					-- layer=2 filter=192 channel=115
					1, -3, -7, -3, 2, 8, 3, 4, 2,
					-- layer=2 filter=192 channel=116
					16, -19, -33, 51, -42, 9, 9, 14, 32,
					-- layer=2 filter=192 channel=117
					-11, -4, 14, -34, 9, -1, 10, -8, 18,
					-- layer=2 filter=192 channel=118
					5, 0, -30, -21, -15, -37, 12, 22, 17,
					-- layer=2 filter=192 channel=119
					21, -2, -18, 23, 11, -9, -14, -9, -3,
					-- layer=2 filter=192 channel=120
					-10, 0, -3, 10, 0, 10, -6, 4, 9,
					-- layer=2 filter=192 channel=121
					-6, -8, 11, 0, 2, 0, 7, 9, 3,
					-- layer=2 filter=192 channel=122
					3, 15, 0, 7, -13, 1, -9, -15, 5,
					-- layer=2 filter=192 channel=123
					2, 33, -4, -29, 10, 3, 31, 13, 21,
					-- layer=2 filter=192 channel=124
					-4, -47, -19, 7, -16, -4, -31, -1, 61,
					-- layer=2 filter=192 channel=125
					2, 2, -1, -10, 3, 11, 0, 0, 0,
					-- layer=2 filter=192 channel=126
					27, 27, -2, 22, -54, -22, 0, 2, -2,
					-- layer=2 filter=192 channel=127
					-11, 8, -3, -14, 14, 22, 6, 17, 28,
					-- layer=2 filter=193 channel=0
					-32, 1, -6, -16, -10, -20, -4, -12, -6,
					-- layer=2 filter=193 channel=1
					12, 2, -10, 1, -3, -12, 5, -43, -23,
					-- layer=2 filter=193 channel=2
					1, 7, -1, 1, 9, -2, -4, 4, -7,
					-- layer=2 filter=193 channel=3
					-17, -4, -4, 27, 27, 10, 60, 33, 38,
					-- layer=2 filter=193 channel=4
					-42, -9, 2, -6, 10, 5, -29, -38, -24,
					-- layer=2 filter=193 channel=5
					2, 12, 6, -36, -29, -24, -17, -13, -19,
					-- layer=2 filter=193 channel=6
					-82, -69, -62, -98, -137, -13, 3, -44, 25,
					-- layer=2 filter=193 channel=7
					7, 13, 43, 98, 44, 32, 7, 10, 11,
					-- layer=2 filter=193 channel=8
					1, -8, 8, -3, -4, 8, -8, -8, 9,
					-- layer=2 filter=193 channel=9
					18, 23, 24, 14, 22, 13, 4, 7, -4,
					-- layer=2 filter=193 channel=10
					-40, -10, -3, -10, 8, 10, 19, 25, 18,
					-- layer=2 filter=193 channel=11
					35, 32, 14, -23, -36, -15, -5, 16, -21,
					-- layer=2 filter=193 channel=12
					48, 8, 10, 24, 23, 38, -34, -84, -4,
					-- layer=2 filter=193 channel=13
					-9, 7, -3, -3, 10, 0, 0, 5, 6,
					-- layer=2 filter=193 channel=14
					24, 19, 0, -4, 7, 10, -25, -53, -28,
					-- layer=2 filter=193 channel=15
					30, 12, 6, 30, -5, -6, -18, 18, -22,
					-- layer=2 filter=193 channel=16
					-30, -33, -14, 22, -1, -7, 22, 42, 26,
					-- layer=2 filter=193 channel=17
					-1, -10, 3, 4, -4, -9, -4, -5, 7,
					-- layer=2 filter=193 channel=18
					26, 25, -33, -43, -14, 14, -57, -19, 29,
					-- layer=2 filter=193 channel=19
					-16, -20, -12, -14, -56, -21, -5, -29, -8,
					-- layer=2 filter=193 channel=20
					0, -2, -2, -8, -3, 6, -5, 8, 2,
					-- layer=2 filter=193 channel=21
					18, 22, -8, -4, -14, -9, 7, -3, 6,
					-- layer=2 filter=193 channel=22
					4, -9, 8, -6, -4, 4, 3, 3, 1,
					-- layer=2 filter=193 channel=23
					-2, 6, -14, 21, -10, 24, 11, -9, 6,
					-- layer=2 filter=193 channel=24
					-4, -15, -15, 29, 34, 18, 39, 32, 20,
					-- layer=2 filter=193 channel=25
					-5, -20, -20, 1, 6, -24, 33, 21, -12,
					-- layer=2 filter=193 channel=26
					-7, -2, 8, -8, -7, 0, 6, 0, -10,
					-- layer=2 filter=193 channel=27
					9, 26, 60, 16, 14, 7, 18, -3, -14,
					-- layer=2 filter=193 channel=28
					22, 29, 16, 1, -24, -38, 29, 12, -5,
					-- layer=2 filter=193 channel=29
					1, 3, -9, -1, 6, 9, 4, 5, 3,
					-- layer=2 filter=193 channel=30
					0, -7, 1, -12, -15, -12, 1, 13, 27,
					-- layer=2 filter=193 channel=31
					-74, 44, 51, 22, 13, 59, -14, -55, -47,
					-- layer=2 filter=193 channel=32
					9, -1, -8, -6, 0, 10, 7, -3, 8,
					-- layer=2 filter=193 channel=33
					-24, 14, 30, 33, 40, 2, 13, 6, 11,
					-- layer=2 filter=193 channel=34
					-30, -39, -69, -30, -55, -57, -11, -10, 34,
					-- layer=2 filter=193 channel=35
					29, 11, 1, 2, -7, -38, 11, 16, 3,
					-- layer=2 filter=193 channel=36
					4, 4, 11, 3, 10, -4, -5, 8, -5,
					-- layer=2 filter=193 channel=37
					11, 13, 20, -10, -17, -16, 0, 13, -1,
					-- layer=2 filter=193 channel=38
					30, 33, 26, -16, 6, 17, -17, -23, -10,
					-- layer=2 filter=193 channel=39
					0, -7, -1, 34, 6, 17, 5, 22, 0,
					-- layer=2 filter=193 channel=40
					17, 37, 15, 32, -26, 41, -8, -41, 28,
					-- layer=2 filter=193 channel=41
					5, 6, -2, -3, -9, 0, -12, 0, 12,
					-- layer=2 filter=193 channel=42
					34, 0, 2, 43, 13, 17, 24, -4, 28,
					-- layer=2 filter=193 channel=43
					19, 19, 2, -21, -10, 1, 15, 9, 6,
					-- layer=2 filter=193 channel=44
					10, -2, 9, -6, 9, -7, 8, 10, 5,
					-- layer=2 filter=193 channel=45
					-53, -26, 20, 20, -9, -7, 40, 34, 48,
					-- layer=2 filter=193 channel=46
					-56, -47, -10, -12, -13, -29, -33, -18, -18,
					-- layer=2 filter=193 channel=47
					-27, -9, 17, 34, -8, 1, 29, 11, 9,
					-- layer=2 filter=193 channel=48
					6, -2, -2, -4, 0, -1, -7, -2, -7,
					-- layer=2 filter=193 channel=49
					12, 26, 27, -26, 2, 41, 11, 68, 82,
					-- layer=2 filter=193 channel=50
					-1, -12, -15, 9, 21, 16, 10, 0, 2,
					-- layer=2 filter=193 channel=51
					21, 30, 24, -36, -31, -40, -7, -15, -16,
					-- layer=2 filter=193 channel=52
					5, 26, -16, -35, -60, -29, -21, -20, -11,
					-- layer=2 filter=193 channel=53
					3, -24, 25, -41, -43, 18, -12, -66, -10,
					-- layer=2 filter=193 channel=54
					-14, -32, -1, 18, -33, -7, 14, 11, 41,
					-- layer=2 filter=193 channel=55
					6, 12, 2, 10, 6, 11, -4, 9, 0,
					-- layer=2 filter=193 channel=56
					40, 44, 37, -11, -2, -14, 3, 7, -23,
					-- layer=2 filter=193 channel=57
					-1, -1, -11, 0, -5, 0, -3, -6, -3,
					-- layer=2 filter=193 channel=58
					42, 24, -9, 9, 28, 47, -28, -31, -32,
					-- layer=2 filter=193 channel=59
					19, 8, -28, -10, -26, -11, -62, -27, -57,
					-- layer=2 filter=193 channel=60
					-28, -5, -18, -14, -64, -35, -48, -29, -48,
					-- layer=2 filter=193 channel=61
					-27, 5, -23, -29, -48, -38, -23, 35, -10,
					-- layer=2 filter=193 channel=62
					-21, -37, 1, -77, -99, -9, -33, -5, 11,
					-- layer=2 filter=193 channel=63
					6, -13, -11, 3, -9, -17, -2, 3, -13,
					-- layer=2 filter=193 channel=64
					-16, -2, -1, 14, 0, 13, 36, 37, 37,
					-- layer=2 filter=193 channel=65
					-72, -34, -67, -108, -61, -38, -70, -50, -27,
					-- layer=2 filter=193 channel=66
					2, 4, -30, 23, 38, 44, 54, -2, 1,
					-- layer=2 filter=193 channel=67
					-20, -10, -18, -2, -21, -24, -16, -7, -34,
					-- layer=2 filter=193 channel=68
					5, 4, -9, 4, 7, -3, 6, -2, 3,
					-- layer=2 filter=193 channel=69
					-12, -8, 8, 18, 7, 28, 36, 28, 27,
					-- layer=2 filter=193 channel=70
					-15, -2, 9, -30, -29, -17, 15, -3, -15,
					-- layer=2 filter=193 channel=71
					26, 22, 41, 19, 25, 17, 4, -15, -38,
					-- layer=2 filter=193 channel=72
					28, 29, 21, 16, 1, -2, -10, -5, 10,
					-- layer=2 filter=193 channel=73
					4, 46, 84, 39, 19, 35, 61, 54, 17,
					-- layer=2 filter=193 channel=74
					17, 3, 7, -10, -4, 4, -15, -6, -24,
					-- layer=2 filter=193 channel=75
					18, 7, 6, 15, 31, 29, -42, -50, -69,
					-- layer=2 filter=193 channel=76
					0, -47, -9, -16, 14, -4, -5, -34, 19,
					-- layer=2 filter=193 channel=77
					-10, -9, 8, -5, 2, -2, -2, -3, 0,
					-- layer=2 filter=193 channel=78
					-4, 15, -7, -20, -8, 3, 18, 54, 33,
					-- layer=2 filter=193 channel=79
					3, 6, 4, -1, 11, 4, 11, -5, -1,
					-- layer=2 filter=193 channel=80
					-16, -17, 0, 37, 18, 14, 13, 17, 17,
					-- layer=2 filter=193 channel=81
					-8, -11, -4, -6, -10, -5, -1, -8, 8,
					-- layer=2 filter=193 channel=82
					-7, -8, -6, -6, 1, -5, -4, 8, 0,
					-- layer=2 filter=193 channel=83
					-6, -31, -20, 14, 10, 19, 5, -8, -22,
					-- layer=2 filter=193 channel=84
					9, 7, -6, 3, -2, 0, -5, 10, -3,
					-- layer=2 filter=193 channel=85
					13, 9, 15, 15, 4, -8, -8, -5, -10,
					-- layer=2 filter=193 channel=86
					5, -4, -4, 19, 6, -8, -8, 12, -14,
					-- layer=2 filter=193 channel=87
					16, 10, -67, -98, -90, -45, -34, -3, 47,
					-- layer=2 filter=193 channel=88
					3, -9, -15, -30, -7, -8, -11, -5, -9,
					-- layer=2 filter=193 channel=89
					46, 19, -22, 23, 10, 15, -22, -10, -46,
					-- layer=2 filter=193 channel=90
					7, -9, 0, 5, 10, 8, -8, 10, -3,
					-- layer=2 filter=193 channel=91
					29, -1, 0, 26, 22, 19, -12, -47, -46,
					-- layer=2 filter=193 channel=92
					28, 15, 3, 13, 12, 23, -2, -56, -29,
					-- layer=2 filter=193 channel=93
					-57, 29, 1, -46, -7, -4, 29, 22, -4,
					-- layer=2 filter=193 channel=94
					-54, -39, -18, -33, -143, -45, -50, -20, 1,
					-- layer=2 filter=193 channel=95
					-16, -19, -9, -9, 3, -16, 11, -16, -4,
					-- layer=2 filter=193 channel=96
					-7, -38, -25, -37, -87, -55, -23, -19, 26,
					-- layer=2 filter=193 channel=97
					13, -18, -1, 45, 32, 12, -5, 4, 10,
					-- layer=2 filter=193 channel=98
					-6, 14, 25, 4, -30, -30, 19, 20, 12,
					-- layer=2 filter=193 channel=99
					35, 15, 24, -46, -36, -24, 4, -11, -10,
					-- layer=2 filter=193 channel=100
					3, -6, 5, 31, 9, 18, -30, -25, -44,
					-- layer=2 filter=193 channel=101
					23, -24, -1, -10, 16, -14, -15, -62, -76,
					-- layer=2 filter=193 channel=102
					-17, -47, -46, -92, -101, -18, -52, -10, 70,
					-- layer=2 filter=193 channel=103
					-17, 8, 17, 11, 6, 28, 15, -9, 15,
					-- layer=2 filter=193 channel=104
					-20, 10, 16, -66, -62, 11, -33, -7, 42,
					-- layer=2 filter=193 channel=105
					-13, 2, 13, -26, -20, -18, -37, 24, -12,
					-- layer=2 filter=193 channel=106
					-4, -15, -4, 3, -8, -9, -28, -33, -55,
					-- layer=2 filter=193 channel=107
					-17, -12, -3, 47, -34, -30, 6, -60, -4,
					-- layer=2 filter=193 channel=108
					15, 3, 26, 37, 29, -5, 23, 19, 11,
					-- layer=2 filter=193 channel=109
					-2, 6, -2, 11, 7, 2, -7, 2, 4,
					-- layer=2 filter=193 channel=110
					-10, -1, -7, 40, 11, 6, 36, 25, 10,
					-- layer=2 filter=193 channel=111
					-9, -6, 8, -10, 9, 5, 1, 0, -6,
					-- layer=2 filter=193 channel=112
					-58, 8, -2, -38, -41, -34, -39, -9, -31,
					-- layer=2 filter=193 channel=113
					-17, 21, 8, -1, -27, -1, -3, 13, -17,
					-- layer=2 filter=193 channel=114
					16, 6, 7, 4, 12, -5, 7, 1, -13,
					-- layer=2 filter=193 channel=115
					-6, 0, -2, 10, 6, -1, -5, -4, -3,
					-- layer=2 filter=193 channel=116
					4, 46, -84, -84, -102, -52, -45, -16, 48,
					-- layer=2 filter=193 channel=117
					0, 0, 41, 65, -18, -16, 21, -2, 23,
					-- layer=2 filter=193 channel=118
					-29, -25, -19, 0, 7, 20, 28, 37, 43,
					-- layer=2 filter=193 channel=119
					-12, -19, -9, -21, 2, 3, -19, -24, -8,
					-- layer=2 filter=193 channel=120
					0, 7, -2, -3, 2, -6, -1, -2, 3,
					-- layer=2 filter=193 channel=121
					4, -9, 5, 3, 0, -4, -1, 4, -7,
					-- layer=2 filter=193 channel=122
					5, -7, 4, -2, 1, 7, -6, 7, -4,
					-- layer=2 filter=193 channel=123
					-2, -3, 23, 24, -21, 2, 3, 9, 22,
					-- layer=2 filter=193 channel=124
					30, -26, 19, 25, 13, -6, -11, -36, -11,
					-- layer=2 filter=193 channel=125
					-8, 1, 9, 0, 8, -2, -8, 2, -3,
					-- layer=2 filter=193 channel=126
					-8, -5, -31, 83, -30, 0, -30, -61, -20,
					-- layer=2 filter=193 channel=127
					-6, -1, -19, -31, -29, -21, -49, -42, -53,
					-- layer=2 filter=194 channel=0
					13, 9, 13, -3, 15, 10, 13, 10, 12,
					-- layer=2 filter=194 channel=1
					-5, -13, -26, -14, -19, 0, 68, 17, -46,
					-- layer=2 filter=194 channel=2
					0, 1, 4, -7, 5, 0, -3, -5, 7,
					-- layer=2 filter=194 channel=3
					7, 26, 18, -10, 15, -16, 0, -6, -15,
					-- layer=2 filter=194 channel=4
					11, -13, 12, 17, -28, 22, -1, 4, 11,
					-- layer=2 filter=194 channel=5
					20, 33, -8, 20, 13, 13, 25, 13, 0,
					-- layer=2 filter=194 channel=6
					9, -69, -37, -145, -98, -87, -41, -56, -37,
					-- layer=2 filter=194 channel=7
					33, -5, 19, 10, 15, 35, 18, 7, 11,
					-- layer=2 filter=194 channel=8
					-6, -8, -8, -9, -8, 5, -5, -4, 7,
					-- layer=2 filter=194 channel=9
					13, 38, 21, -33, -27, 6, -1, -9, -17,
					-- layer=2 filter=194 channel=10
					26, 5, 19, 11, 18, 20, 4, 8, 18,
					-- layer=2 filter=194 channel=11
					30, 14, 7, 27, 29, 9, 5, 29, -4,
					-- layer=2 filter=194 channel=12
					28, 7, 11, 30, 1, 7, 63, 16, -35,
					-- layer=2 filter=194 channel=13
					0, -3, -5, 11, -1, 1, -4, -3, -2,
					-- layer=2 filter=194 channel=14
					20, 13, -11, -12, -7, -10, 44, 9, -21,
					-- layer=2 filter=194 channel=15
					-7, 5, -3, 17, 12, 2, 9, 7, 19,
					-- layer=2 filter=194 channel=16
					-18, -25, -7, -39, -12, 28, -18, 13, 28,
					-- layer=2 filter=194 channel=17
					0, 7, 11, 4, 6, 3, 5, 11, 0,
					-- layer=2 filter=194 channel=18
					-53, -50, -10, -30, -56, -8, 9, 7, -44,
					-- layer=2 filter=194 channel=19
					-31, -57, -26, 15, -18, -26, 43, 23, 0,
					-- layer=2 filter=194 channel=20
					-3, -2, -11, 8, -2, 6, -4, 5, 1,
					-- layer=2 filter=194 channel=21
					-3, 3, -14, -21, -4, 0, -17, 5, 18,
					-- layer=2 filter=194 channel=22
					-3, 5, 4, 8, 0, -2, 3, 0, 4,
					-- layer=2 filter=194 channel=23
					-24, -18, 17, 10, -29, 32, 9, 11, 26,
					-- layer=2 filter=194 channel=24
					17, 18, 10, -10, 13, -17, -15, -20, -12,
					-- layer=2 filter=194 channel=25
					10, -2, -15, -2, -17, -16, -10, -25, -13,
					-- layer=2 filter=194 channel=26
					8, 0, 8, 8, -8, -9, 0, -9, 1,
					-- layer=2 filter=194 channel=27
					-12, 10, -5, 23, 24, 23, 2, 28, 20,
					-- layer=2 filter=194 channel=28
					29, -25, -6, 20, 2, 27, 6, -3, 19,
					-- layer=2 filter=194 channel=29
					-5, 1, 6, -2, -5, -5, -9, -6, -10,
					-- layer=2 filter=194 channel=30
					-12, 5, -6, 0, -28, -25, -6, 4, 22,
					-- layer=2 filter=194 channel=31
					8, 42, 28, 12, 57, 57, -36, -61, -1,
					-- layer=2 filter=194 channel=32
					0, -11, -2, -4, 6, 7, 3, -11, 5,
					-- layer=2 filter=194 channel=33
					15, 11, 11, 23, 33, 21, 5, 30, -3,
					-- layer=2 filter=194 channel=34
					1, -18, -65, 39, -22, -80, -13, -9, 12,
					-- layer=2 filter=194 channel=35
					10, -22, -41, 10, 1, 5, -16, -10, 3,
					-- layer=2 filter=194 channel=36
					5, -5, 0, 9, -7, 7, 19, -1, 1,
					-- layer=2 filter=194 channel=37
					23, 8, 5, 9, 19, 15, 6, 18, 14,
					-- layer=2 filter=194 channel=38
					20, 25, 22, 10, 12, 16, 3, -2, 2,
					-- layer=2 filter=194 channel=39
					6, 8, 24, 24, 19, 29, 23, 40, 19,
					-- layer=2 filter=194 channel=40
					1, -22, 1, -57, -55, 17, 7, 46, -2,
					-- layer=2 filter=194 channel=41
					8, 6, -1, 10, 8, 4, 11, 2, -8,
					-- layer=2 filter=194 channel=42
					15, -16, 8, -8, -11, 37, 18, 11, 26,
					-- layer=2 filter=194 channel=43
					-7, 0, -4, -15, 22, 8, -22, 10, -20,
					-- layer=2 filter=194 channel=44
					-5, 8, 8, -3, -7, 8, 3, -5, 12,
					-- layer=2 filter=194 channel=45
					-24, -30, -28, 18, 13, 35, -8, -14, 28,
					-- layer=2 filter=194 channel=46
					-21, -10, 28, 14, -12, -4, 11, -2, 28,
					-- layer=2 filter=194 channel=47
					16, 7, 2, 18, 0, 43, 2, 0, 31,
					-- layer=2 filter=194 channel=48
					7, 7, 9, 7, 4, 3, -7, -9, 3,
					-- layer=2 filter=194 channel=49
					-58, -6, 17, -65, -63, -19, 27, -11, 26,
					-- layer=2 filter=194 channel=50
					-4, 8, 5, 7, -3, 11, 20, 25, 11,
					-- layer=2 filter=194 channel=51
					25, 26, 10, 15, 23, -4, 12, 10, 15,
					-- layer=2 filter=194 channel=52
					-13, -19, 17, 26, -19, -22, -2, 44, -11,
					-- layer=2 filter=194 channel=53
					8, -69, -40, -32, 31, -116, 36, -75, -50,
					-- layer=2 filter=194 channel=54
					19, -3, -17, 11, -27, 0, 48, -6, 0,
					-- layer=2 filter=194 channel=55
					-1, 13, 10, -1, 5, 4, -2, 4, 0,
					-- layer=2 filter=194 channel=56
					41, 26, 6, 14, 25, 6, 1, 12, 9,
					-- layer=2 filter=194 channel=57
					-5, -6, -8, -14, -8, -16, 2, -1, 2,
					-- layer=2 filter=194 channel=58
					28, 15, 0, 40, 16, 25, 50, 20, -7,
					-- layer=2 filter=194 channel=59
					-19, -16, -10, 43, 15, -25, 38, 16, -2,
					-- layer=2 filter=194 channel=60
					-14, 2, -12, 25, 15, 13, 26, 14, 20,
					-- layer=2 filter=194 channel=61
					-55, -26, -41, -32, -16, -43, -35, 15, -10,
					-- layer=2 filter=194 channel=62
					-27, -26, -17, -39, -80, -28, 18, 10, 1,
					-- layer=2 filter=194 channel=63
					-1, 4, 26, 16, -10, 16, 21, 11, 6,
					-- layer=2 filter=194 channel=64
					5, 5, 23, -11, -13, 8, 24, 29, 23,
					-- layer=2 filter=194 channel=65
					-40, -64, -39, -44, -69, -41, -32, -42, -43,
					-- layer=2 filter=194 channel=66
					-3, -54, 59, 50, 25, 21, 16, -4, 63,
					-- layer=2 filter=194 channel=67
					15, 8, 20, -5, -23, -11, -6, -18, 4,
					-- layer=2 filter=194 channel=68
					9, 9, -2, -3, -6, -1, -9, 1, 8,
					-- layer=2 filter=194 channel=69
					-7, 20, 14, -9, -15, 40, 9, 31, 41,
					-- layer=2 filter=194 channel=70
					5, -21, -15, 24, 14, 9, 14, -6, 7,
					-- layer=2 filter=194 channel=71
					9, 25, -21, 0, 14, 9, 0, 10, 21,
					-- layer=2 filter=194 channel=72
					25, -2, 26, 14, 30, 22, 47, 28, 20,
					-- layer=2 filter=194 channel=73
					50, 48, 76, 59, 79, 82, 43, 9, 49,
					-- layer=2 filter=194 channel=74
					2, 14, 26, 17, 7, -5, 17, 13, 0,
					-- layer=2 filter=194 channel=75
					24, -39, -20, -3, -8, 13, 6, -26, -45,
					-- layer=2 filter=194 channel=76
					9, -55, -33, -23, -8, 28, -31, -80, -46,
					-- layer=2 filter=194 channel=77
					8, -11, 0, -5, -6, -8, 4, 10, -3,
					-- layer=2 filter=194 channel=78
					31, 12, -10, -5, -11, -9, 28, 12, -19,
					-- layer=2 filter=194 channel=79
					-1, -4, -8, -1, 8, -6, -5, 1, -3,
					-- layer=2 filter=194 channel=80
					12, 8, 23, 20, 4, 22, 0, 6, 8,
					-- layer=2 filter=194 channel=81
					8, 5, 10, 10, 24, 6, 16, 8, 9,
					-- layer=2 filter=194 channel=82
					0, -6, 2, 5, -3, -1, 4, 3, 0,
					-- layer=2 filter=194 channel=83
					-17, -32, -21, 7, -26, -21, -10, -4, 13,
					-- layer=2 filter=194 channel=84
					4, 4, -1, 7, -7, 10, 4, 4, -8,
					-- layer=2 filter=194 channel=85
					16, 9, 0, 0, 13, -2, 14, 13, 10,
					-- layer=2 filter=194 channel=86
					2, -5, 6, -4, -6, 14, 16, -16, 2,
					-- layer=2 filter=194 channel=87
					13, -27, -41, -22, -78, -29, -56, -30, -21,
					-- layer=2 filter=194 channel=88
					17, 10, 12, -6, -33, -10, 6, 7, -23,
					-- layer=2 filter=194 channel=89
					-2, -25, -9, 5, -14, -8, 63, -5, -21,
					-- layer=2 filter=194 channel=90
					2, 9, 4, 2, -3, 0, 0, 9, -2,
					-- layer=2 filter=194 channel=91
					11, -5, 16, 15, 11, 33, 20, -7, -1,
					-- layer=2 filter=194 channel=92
					22, 16, 7, 13, -20, 20, 69, 31, -30,
					-- layer=2 filter=194 channel=93
					19, -38, 30, -6, -41, 8, 14, 51, -10,
					-- layer=2 filter=194 channel=94
					-81, -69, -43, -44, -89, -68, -2, 2, -32,
					-- layer=2 filter=194 channel=95
					-4, -10, -1, 2, -15, -7, 0, -7, -17,
					-- layer=2 filter=194 channel=96
					-89, -51, -64, -36, -66, -77, -30, -69, -13,
					-- layer=2 filter=194 channel=97
					22, 20, 3, 11, -14, -4, -1, -16, -3,
					-- layer=2 filter=194 channel=98
					9, -3, 6, 30, 26, 20, 2, 22, 32,
					-- layer=2 filter=194 channel=99
					15, -11, -30, 49, 5, 33, 53, 28, 32,
					-- layer=2 filter=194 channel=100
					10, 7, 3, -15, 11, 14, -5, 2, -20,
					-- layer=2 filter=194 channel=101
					16, 16, -29, 7, 6, -3, -20, -7, 11,
					-- layer=2 filter=194 channel=102
					-59, -60, -80, -70, -104, -50, -30, -73, 1,
					-- layer=2 filter=194 channel=103
					-29, -13, 4, -56, -58, -14, 16, 26, 9,
					-- layer=2 filter=194 channel=104
					-46, -30, -9, -64, -38, -46, 2, 4, -21,
					-- layer=2 filter=194 channel=105
					-38, -72, -23, -2, -22, 34, -48, -3, -12,
					-- layer=2 filter=194 channel=106
					32, -26, -13, 4, 11, -12, -2, -21, -8,
					-- layer=2 filter=194 channel=107
					16, 14, 66, 5, 20, 9, -52, 6, 12,
					-- layer=2 filter=194 channel=108
					-1, 6, -30, 1, -10, 8, 11, -13, 16,
					-- layer=2 filter=194 channel=109
					14, 19, 3, -12, 4, -2, 7, -8, -1,
					-- layer=2 filter=194 channel=110
					-25, -21, -31, -6, -21, 0, -23, -3, -11,
					-- layer=2 filter=194 channel=111
					2, 3, 6, -1, 11, 4, -3, -8, -11,
					-- layer=2 filter=194 channel=112
					21, -3, -1, -9, 13, 3, -16, 16, 12,
					-- layer=2 filter=194 channel=113
					-35, 0, -27, 25, -8, -28, -38, 33, 36,
					-- layer=2 filter=194 channel=114
					0, 6, 8, -12, -1, -10, 1, -14, 3,
					-- layer=2 filter=194 channel=115
					-5, 9, 2, -4, 2, 6, -2, 9, -7,
					-- layer=2 filter=194 channel=116
					-10, -5, -46, 5, -63, -6, -45, 0, -14,
					-- layer=2 filter=194 channel=117
					24, -13, -12, -9, 1, 36, 42, 0, 13,
					-- layer=2 filter=194 channel=118
					7, 8, 23, 8, 8, 9, -3, 3, -22,
					-- layer=2 filter=194 channel=119
					-14, 8, 29, -24, -23, 40, 4, -13, 0,
					-- layer=2 filter=194 channel=120
					-6, 4, -6, -6, -2, -6, 1, 6, 5,
					-- layer=2 filter=194 channel=121
					6, -4, 0, -6, -3, -5, -7, -1, 1,
					-- layer=2 filter=194 channel=122
					5, -1, -9, -5, 10, 0, 1, -1, -3,
					-- layer=2 filter=194 channel=123
					-13, -12, 20, 2, 2, 16, 18, 11, 33,
					-- layer=2 filter=194 channel=124
					9, -35, -4, -2, -20, -5, 32, -24, -20,
					-- layer=2 filter=194 channel=125
					-9, -6, 12, -4, 3, 8, 7, 8, 5,
					-- layer=2 filter=194 channel=126
					-7, 0, -33, 31, 12, 11, -31, -8, 30,
					-- layer=2 filter=194 channel=127
					2, 20, 2, -11, -32, -9, 0, -9, -1,
					-- layer=2 filter=195 channel=0
					10, 12, 30, 17, 14, -9, 8, 7, 18,
					-- layer=2 filter=195 channel=1
					5, 23, 3, 9, 36, 5, -12, 9, -15,
					-- layer=2 filter=195 channel=2
					-8, 3, -7, 6, 9, -2, -6, 11, 6,
					-- layer=2 filter=195 channel=3
					14, -3, -10, 15, -6, 3, 2, 10, 6,
					-- layer=2 filter=195 channel=4
					-1, 16, -2, -6, -1, -7, -19, 9, -20,
					-- layer=2 filter=195 channel=5
					11, -25, 6, 0, 7, -8, -14, 3, 3,
					-- layer=2 filter=195 channel=6
					-5, 29, -52, 20, 1, 27, 24, 45, -38,
					-- layer=2 filter=195 channel=7
					42, 30, 24, 50, 46, 19, 26, 48, -27,
					-- layer=2 filter=195 channel=8
					-2, 6, -9, 8, -3, -1, 10, 4, -6,
					-- layer=2 filter=195 channel=9
					2, -4, -25, -2, -9, -9, 41, 49, 18,
					-- layer=2 filter=195 channel=10
					19, 36, 11, 6, 0, -14, 18, -9, -13,
					-- layer=2 filter=195 channel=11
					-20, -10, -40, 17, 17, -8, 0, 6, -16,
					-- layer=2 filter=195 channel=12
					14, -2, -8, 21, 22, 25, -32, -22, 7,
					-- layer=2 filter=195 channel=13
					-3, -5, 5, 2, -3, -2, -5, -6, 3,
					-- layer=2 filter=195 channel=14
					24, 17, -6, 5, 22, 29, -39, -11, 0,
					-- layer=2 filter=195 channel=15
					-45, 1, -6, -51, -1, -35, -36, -32, -10,
					-- layer=2 filter=195 channel=16
					-18, 2, 0, -14, -8, 26, -44, -1, -2,
					-- layer=2 filter=195 channel=17
					-1, -5, -11, -2, 6, 9, -2, 2, -6,
					-- layer=2 filter=195 channel=18
					-19, -5, -8, -40, -10, -27, -54, -65, -6,
					-- layer=2 filter=195 channel=19
					-3, -11, 7, 10, 59, 20, 21, 7, 10,
					-- layer=2 filter=195 channel=20
					0, 6, -9, -2, 10, 2, 5, 6, 3,
					-- layer=2 filter=195 channel=21
					5, -3, -22, -14, -4, -13, -17, -14, -7,
					-- layer=2 filter=195 channel=22
					-2, -2, 3, 10, 2, -5, -5, -9, 4,
					-- layer=2 filter=195 channel=23
					-29, -1, -2, -10, 17, 2, 10, 7, -14,
					-- layer=2 filter=195 channel=24
					-7, 0, -17, -6, -15, -2, 2, -9, -1,
					-- layer=2 filter=195 channel=25
					1, -9, -23, -5, -5, 23, 8, 18, 17,
					-- layer=2 filter=195 channel=26
					-5, -6, 7, -9, 9, -1, -6, 1, 6,
					-- layer=2 filter=195 channel=27
					-36, -7, 34, 5, 3, 29, 18, -11, -9,
					-- layer=2 filter=195 channel=28
					8, 18, 18, 26, 25, 24, -47, -39, -25,
					-- layer=2 filter=195 channel=29
					-2, 0, 8, 3, -5, 9, -7, 3, 1,
					-- layer=2 filter=195 channel=30
					-9, 13, -2, -21, -2, -17, 26, -3, 28,
					-- layer=2 filter=195 channel=31
					-69, -34, 31, -9, 76, -44, 17, -14, -6,
					-- layer=2 filter=195 channel=32
					-6, -9, 3, -10, -6, 1, 4, 9, 5,
					-- layer=2 filter=195 channel=33
					23, 20, 8, -6, -34, -63, -50, -16, 22,
					-- layer=2 filter=195 channel=34
					9, -50, -72, -62, -58, 32, -27, -25, 20,
					-- layer=2 filter=195 channel=35
					8, 16, 9, 22, 48, 30, -35, 6, -11,
					-- layer=2 filter=195 channel=36
					5, 11, 4, -10, 3, 15, 13, 6, 16,
					-- layer=2 filter=195 channel=37
					-10, -21, -14, -6, -6, -2, 5, 4, 1,
					-- layer=2 filter=195 channel=38
					22, 23, 15, 21, -3, 6, 8, 7, -6,
					-- layer=2 filter=195 channel=39
					-18, 14, 6, -5, 27, -4, -11, 49, -19,
					-- layer=2 filter=195 channel=40
					-38, 39, 39, -40, 44, -25, -46, -31, -26,
					-- layer=2 filter=195 channel=41
					9, 5, -3, 4, -2, -4, -3, -9, 6,
					-- layer=2 filter=195 channel=42
					-29, 10, -28, -20, 23, -20, -24, -1, -16,
					-- layer=2 filter=195 channel=43
					-4, -45, -85, -17, -32, -55, 31, -38, 13,
					-- layer=2 filter=195 channel=44
					0, 7, 4, 3, 0, 7, -8, -10, 0,
					-- layer=2 filter=195 channel=45
					-64, 18, 36, -20, -1, 61, 15, -1, 4,
					-- layer=2 filter=195 channel=46
					18, 20, -5, 13, -15, -49, 42, 22, -17,
					-- layer=2 filter=195 channel=47
					-7, 45, 34, 21, 24, 9, -37, -29, -36,
					-- layer=2 filter=195 channel=48
					6, -8, 2, -8, -4, -6, 0, 0, -5,
					-- layer=2 filter=195 channel=49
					-26, -4, -12, -28, -38, 12, -39, -22, -24,
					-- layer=2 filter=195 channel=50
					16, 22, 3, 9, 16, 0, -2, -4, -1,
					-- layer=2 filter=195 channel=51
					-5, -20, -8, 0, 7, 12, 6, 11, -2,
					-- layer=2 filter=195 channel=52
					-19, -42, 5, 14, 5, 11, 0, 3, 6,
					-- layer=2 filter=195 channel=53
					27, 16, -5, 19, 35, 3, 0, -41, -54,
					-- layer=2 filter=195 channel=54
					-1, 2, -1, -1, 11, 4, -20, 28, -29,
					-- layer=2 filter=195 channel=55
					5, -1, -11, -1, 7, 6, -3, 7, -6,
					-- layer=2 filter=195 channel=56
					1, -23, -35, 4, 12, -13, 5, 17, 9,
					-- layer=2 filter=195 channel=57
					4, 0, -1, 7, -1, -13, 6, -9, -14,
					-- layer=2 filter=195 channel=58
					24, 16, -33, 5, 15, 16, 9, -10, 6,
					-- layer=2 filter=195 channel=59
					20, 15, -2, 43, 18, 12, 16, -12, -24,
					-- layer=2 filter=195 channel=60
					11, -5, -45, 25, -14, -16, -13, -26, -27,
					-- layer=2 filter=195 channel=61
					-37, 28, 38, 7, 9, 34, -20, -19, -76,
					-- layer=2 filter=195 channel=62
					-4, -4, -21, -35, 5, 12, 0, 4, 4,
					-- layer=2 filter=195 channel=63
					20, 30, -12, -13, -6, 1, -3, 10, -33,
					-- layer=2 filter=195 channel=64
					-24, -8, -22, 9, -3, 0, 2, 14, -5,
					-- layer=2 filter=195 channel=65
					-8, 35, 29, 6, 18, 34, -3, 22, -34,
					-- layer=2 filter=195 channel=66
					39, -30, 32, -37, -36, -47, -7, -38, 20,
					-- layer=2 filter=195 channel=67
					10, -33, -45, 30, 1, -38, 54, 46, 24,
					-- layer=2 filter=195 channel=68
					4, -7, -5, -5, 3, -5, 5, 5, 2,
					-- layer=2 filter=195 channel=69
					-20, -18, -37, -4, 3, 5, -3, -14, -15,
					-- layer=2 filter=195 channel=70
					20, -1, 36, 12, 19, 10, -24, -6, -9,
					-- layer=2 filter=195 channel=71
					-21, -38, -8, 3, 16, 23, 17, 11, 0,
					-- layer=2 filter=195 channel=72
					19, 28, 0, 31, 5, 0, 9, 28, -7,
					-- layer=2 filter=195 channel=73
					3, -7, -17, 46, 9, -49, 13, -44, -70,
					-- layer=2 filter=195 channel=74
					13, 21, 13, 32, 21, -20, 26, 6, 1,
					-- layer=2 filter=195 channel=75
					-37, -29, -53, 25, 65, 11, 3, -16, 0,
					-- layer=2 filter=195 channel=76
					40, -58, -33, 42, 26, -4, 47, -11, -26,
					-- layer=2 filter=195 channel=77
					-6, -3, 0, -8, -6, -3, -9, 5, 1,
					-- layer=2 filter=195 channel=78
					-36, -39, -44, -21, 12, 18, -13, -3, -14,
					-- layer=2 filter=195 channel=79
					-8, 0, 2, -1, -2, -2, 3, 7, 9,
					-- layer=2 filter=195 channel=80
					-11, -8, -24, -5, 4, -25, 0, 0, -15,
					-- layer=2 filter=195 channel=81
					-14, -3, -23, -24, -22, -4, -6, -5, -12,
					-- layer=2 filter=195 channel=82
					2, 2, 10, -2, -2, -8, -5, 9, 7,
					-- layer=2 filter=195 channel=83
					-37, 30, 5, -25, 28, 40, -19, -15, -31,
					-- layer=2 filter=195 channel=84
					3, -7, 4, 8, -3, 5, 4, -10, -4,
					-- layer=2 filter=195 channel=85
					-22, 4, -1, -16, -13, -14, -11, -2, -7,
					-- layer=2 filter=195 channel=86
					-16, -2, 26, 0, 3, -4, 1, -15, -6,
					-- layer=2 filter=195 channel=87
					8, -15, -57, 29, 26, -49, 1, 17, -5,
					-- layer=2 filter=195 channel=88
					6, 37, 14, 2, 6, -4, 0, 12, 10,
					-- layer=2 filter=195 channel=89
					9, -4, -44, 20, 24, 6, 0, 8, 1,
					-- layer=2 filter=195 channel=90
					12, -10, 7, -7, 5, 6, -5, -11, -6,
					-- layer=2 filter=195 channel=91
					0, -6, -61, 8, 11, -15, -25, 11, 3,
					-- layer=2 filter=195 channel=92
					-10, 26, -7, 0, 35, 9, -6, 7, -17,
					-- layer=2 filter=195 channel=93
					8, 44, -36, -35, 14, -50, 18, -27, -15,
					-- layer=2 filter=195 channel=94
					-24, -33, -31, 6, -8, 23, 29, 8, -20,
					-- layer=2 filter=195 channel=95
					3, 5, 2, -9, -11, 16, 2, 12, -1,
					-- layer=2 filter=195 channel=96
					53, 9, 4, 66, -22, -5, 19, 28, 13,
					-- layer=2 filter=195 channel=97
					-5, 2, -12, 27, -9, 12, 14, -6, 19,
					-- layer=2 filter=195 channel=98
					-10, 27, 23, 14, 29, 17, -24, -57, -51,
					-- layer=2 filter=195 channel=99
					10, -31, -6, 45, 26, 7, 33, -28, -5,
					-- layer=2 filter=195 channel=100
					32, 7, 9, -3, 42, -6, -10, -13, 13,
					-- layer=2 filter=195 channel=101
					-14, -24, -14, 7, -9, 20, 10, 21, 17,
					-- layer=2 filter=195 channel=102
					-1, -18, -6, 16, -11, 21, 15, -21, -35,
					-- layer=2 filter=195 channel=103
					-46, -1, -15, -59, -23, -19, -59, -60, 19,
					-- layer=2 filter=195 channel=104
					24, -24, -8, -5, -53, 17, -21, -28, -15,
					-- layer=2 filter=195 channel=105
					14, -12, 38, 28, 8, -9, 26, 9, -31,
					-- layer=2 filter=195 channel=106
					2, -6, -30, 17, -9, 17, 24, -5, 13,
					-- layer=2 filter=195 channel=107
					-37, 9, -16, -4, -29, 4, 38, 36, 50,
					-- layer=2 filter=195 channel=108
					-38, 5, 37, 12, 21, 37, 15, -38, -8,
					-- layer=2 filter=195 channel=109
					29, 1, -15, 6, 10, 0, 17, 16, -5,
					-- layer=2 filter=195 channel=110
					3, 8, 14, 5, 11, 22, 9, 42, -11,
					-- layer=2 filter=195 channel=111
					6, 1, 12, 0, 1, -6, -12, 1, 6,
					-- layer=2 filter=195 channel=112
					-14, 15, -5, 5, 2, 1, -25, -3, -10,
					-- layer=2 filter=195 channel=113
					37, 49, 34, -14, 8, -1, 6, -24, -24,
					-- layer=2 filter=195 channel=114
					7, 8, 19, -3, 15, 12, -2, 0, -3,
					-- layer=2 filter=195 channel=115
					0, -8, 0, -2, -9, 1, 2, -12, 4,
					-- layer=2 filter=195 channel=116
					11, -7, -40, -2, 4, -35, -19, -1, -23,
					-- layer=2 filter=195 channel=117
					-7, -8, -11, 1, 65, 1, 37, 29, -15,
					-- layer=2 filter=195 channel=118
					10, -3, -34, -20, -14, 9, -3, 1, 6,
					-- layer=2 filter=195 channel=119
					2, -15, -10, -28, 21, -25, -19, -33, -17,
					-- layer=2 filter=195 channel=120
					-7, 8, -4, -8, 8, -10, 10, -8, 1,
					-- layer=2 filter=195 channel=121
					0, 8, -1, -2, 6, -9, -10, -10, -2,
					-- layer=2 filter=195 channel=122
					-9, -12, 0, 9, 7, 6, 2, -11, 3,
					-- layer=2 filter=195 channel=123
					24, 19, 5, 54, 22, -7, 23, 1, -46,
					-- layer=2 filter=195 channel=124
					-13, -6, -35, -48, 17, -26, -6, 20, -1,
					-- layer=2 filter=195 channel=125
					0, 7, -11, 7, 5, -6, 3, -7, -5,
					-- layer=2 filter=195 channel=126
					55, -3, -13, 15, -48, -3, -7, 40, 22,
					-- layer=2 filter=195 channel=127
					0, 37, 46, 0, -16, 18, 0, -9, -6,
					-- layer=2 filter=196 channel=0
					6, -1, -6, 2, -4, 6, 0, -6, -10,
					-- layer=2 filter=196 channel=1
					-1, -7, 3, 3, -16, 0, -9, -8, -1,
					-- layer=2 filter=196 channel=2
					-10, 8, -2, -5, 0, 6, 3, -7, 1,
					-- layer=2 filter=196 channel=3
					-9, 1, -5, 9, 6, -6, 1, 7, -2,
					-- layer=2 filter=196 channel=4
					0, 6, -13, 9, 0, 3, -7, -3, -6,
					-- layer=2 filter=196 channel=5
					-6, 0, -9, 6, -1, -4, -9, -1, -1,
					-- layer=2 filter=196 channel=6
					-14, 0, -6, 3, 6, -9, -7, 0, -5,
					-- layer=2 filter=196 channel=7
					-18, -14, -16, 7, -16, -10, 4, -2, 7,
					-- layer=2 filter=196 channel=8
					-1, -4, 3, 10, 1, 0, -11, -2, -3,
					-- layer=2 filter=196 channel=9
					-5, 1, 2, -5, 4, -7, 1, 9, -1,
					-- layer=2 filter=196 channel=10
					-1, -5, -9, -4, 7, 4, 4, -9, 2,
					-- layer=2 filter=196 channel=11
					-8, -2, 0, 0, -4, 2, -12, -10, -3,
					-- layer=2 filter=196 channel=12
					0, 4, 12, -8, 0, -15, -9, -1, -14,
					-- layer=2 filter=196 channel=13
					-3, 6, -7, 2, -8, 4, 4, -8, -1,
					-- layer=2 filter=196 channel=14
					-8, 4, -6, -2, -6, -9, 1, -2, 3,
					-- layer=2 filter=196 channel=15
					-3, 3, 1, -3, -6, -2, 0, 6, 0,
					-- layer=2 filter=196 channel=16
					0, -9, -4, -8, 7, 6, -9, -6, 0,
					-- layer=2 filter=196 channel=17
					-9, -5, 6, -8, 4, 0, -6, 2, 3,
					-- layer=2 filter=196 channel=18
					16, 1, -22, -7, 3, -10, 4, 3, 0,
					-- layer=2 filter=196 channel=19
					1, 8, 0, -1, -9, -10, 4, 3, 8,
					-- layer=2 filter=196 channel=20
					-6, -6, 1, -10, -4, 8, 2, -8, 2,
					-- layer=2 filter=196 channel=21
					-7, -6, -1, -1, 4, 0, -4, 4, -6,
					-- layer=2 filter=196 channel=22
					5, -9, -6, -1, -5, 10, 10, -4, 9,
					-- layer=2 filter=196 channel=23
					2, 0, -10, -6, -2, -13, -2, -11, 2,
					-- layer=2 filter=196 channel=24
					6, 1, -5, -9, 8, -9, 6, -7, -9,
					-- layer=2 filter=196 channel=25
					-5, 1, 7, -21, -8, -16, -1, -8, -13,
					-- layer=2 filter=196 channel=26
					0, 4, -7, 10, 10, 7, 4, 8, 2,
					-- layer=2 filter=196 channel=27
					-3, 6, -5, 0, -9, -7, -8, -7, -2,
					-- layer=2 filter=196 channel=28
					-1, -10, -8, -4, -4, 4, 0, 1, -10,
					-- layer=2 filter=196 channel=29
					3, -6, -4, 8, 6, -5, 1, -1, -5,
					-- layer=2 filter=196 channel=30
					3, 7, -1, 1, -6, 2, 0, -8, -7,
					-- layer=2 filter=196 channel=31
					1, -9, 2, 2, -6, 9, -2, -8, 9,
					-- layer=2 filter=196 channel=32
					9, 1, -11, -9, 3, 7, -10, 0, 5,
					-- layer=2 filter=196 channel=33
					-9, -1, -7, 1, -5, -11, 0, -6, -6,
					-- layer=2 filter=196 channel=34
					3, -6, -5, -1, -3, 6, -10, -3, 1,
					-- layer=2 filter=196 channel=35
					-9, -14, -4, -11, 8, -6, -8, -16, -19,
					-- layer=2 filter=196 channel=36
					-1, -1, 2, 1, 0, -4, 2, -4, 1,
					-- layer=2 filter=196 channel=37
					-1, -13, 5, 6, -2, -12, -1, -12, -4,
					-- layer=2 filter=196 channel=38
					0, -1, -14, -1, 0, -9, -10, -5, 7,
					-- layer=2 filter=196 channel=39
					3, -12, 0, -5, -11, -1, 0, -5, -6,
					-- layer=2 filter=196 channel=40
					4, 6, -8, 6, -2, 3, 4, -4, -11,
					-- layer=2 filter=196 channel=41
					3, 1, -7, -7, -7, 9, 5, -3, -10,
					-- layer=2 filter=196 channel=42
					7, -9, -4, -12, 4, 0, 5, 0, -1,
					-- layer=2 filter=196 channel=43
					2, -3, -10, 2, 8, -6, 0, -9, 4,
					-- layer=2 filter=196 channel=44
					0, -1, 6, 0, 6, 2, -11, -10, 0,
					-- layer=2 filter=196 channel=45
					-8, -6, 8, 0, 2, -4, -1, 0, -2,
					-- layer=2 filter=196 channel=46
					-9, -9, -11, -9, -7, -3, 6, 7, 1,
					-- layer=2 filter=196 channel=47
					-12, -15, 0, -2, -5, 11, -12, 3, 7,
					-- layer=2 filter=196 channel=48
					-9, 7, 1, -1, -1, 5, -4, -8, -4,
					-- layer=2 filter=196 channel=49
					-6, -13, 0, 1, -5, -8, 4, -4, -8,
					-- layer=2 filter=196 channel=50
					10, 0, 6, 6, 5, 6, 4, 4, -5,
					-- layer=2 filter=196 channel=51
					-12, 0, -8, -9, -5, -11, -1, 4, 6,
					-- layer=2 filter=196 channel=52
					-13, -2, 2, 1, 1, 5, 3, 3, -2,
					-- layer=2 filter=196 channel=53
					-4, 1, 6, -10, -2, 4, 7, 5, 7,
					-- layer=2 filter=196 channel=54
					0, 0, -3, -5, -15, -13, -5, -15, -7,
					-- layer=2 filter=196 channel=55
					0, 2, -4, -9, -4, -2, 3, -12, 0,
					-- layer=2 filter=196 channel=56
					-8, -9, 5, -7, -11, -9, -9, -4, 4,
					-- layer=2 filter=196 channel=57
					8, -4, -2, -1, 12, 10, 1, 10, -2,
					-- layer=2 filter=196 channel=58
					0, -4, 8, 3, 0, 0, -10, -15, 1,
					-- layer=2 filter=196 channel=59
					5, 8, 5, 2, -4, -12, -4, 2, -7,
					-- layer=2 filter=196 channel=60
					-3, -1, -10, -19, -1, -7, 5, -1, -14,
					-- layer=2 filter=196 channel=61
					-9, 11, 2, 6, 1, -11, -9, -14, -8,
					-- layer=2 filter=196 channel=62
					-4, 2, -20, 7, 2, -3, 0, -8, -6,
					-- layer=2 filter=196 channel=63
					1, 9, -4, -9, -5, -14, 3, -7, 1,
					-- layer=2 filter=196 channel=64
					-10, -4, 3, -5, -4, 0, -2, 2, 9,
					-- layer=2 filter=196 channel=65
					4, 1, 1, 0, -3, -9, -5, 2, 0,
					-- layer=2 filter=196 channel=66
					1, 12, 4, 4, -3, -7, -10, 5, 1,
					-- layer=2 filter=196 channel=67
					6, 7, 0, 9, 4, -1, -1, 7, 5,
					-- layer=2 filter=196 channel=68
					5, -10, -4, -5, 9, 6, -10, 7, -7,
					-- layer=2 filter=196 channel=69
					-2, 1, 3, -13, -16, -10, 0, -8, 3,
					-- layer=2 filter=196 channel=70
					9, 1, -6, -2, -9, 3, -1, -11, -17,
					-- layer=2 filter=196 channel=71
					-4, -6, 0, 10, 10, -3, 3, 2, -5,
					-- layer=2 filter=196 channel=72
					-12, 3, -15, -6, 0, 8, -5, 7, 5,
					-- layer=2 filter=196 channel=73
					-5, -12, 14, -10, -5, -6, -3, -7, 1,
					-- layer=2 filter=196 channel=74
					4, -11, -12, 5, 10, -2, -3, -9, -4,
					-- layer=2 filter=196 channel=75
					11, -7, 1, -8, -1, 12, 0, 0, 0,
					-- layer=2 filter=196 channel=76
					5, 7, -10, 3, -4, -9, 9, 0, 11,
					-- layer=2 filter=196 channel=77
					7, -9, -4, 2, 0, 0, 4, -4, -2,
					-- layer=2 filter=196 channel=78
					-13, -2, 6, -7, -4, 3, -12, -1, -2,
					-- layer=2 filter=196 channel=79
					-4, 7, 6, -6, 8, 9, 6, 6, 0,
					-- layer=2 filter=196 channel=80
					-10, -2, -5, -5, -9, 3, 0, -3, -11,
					-- layer=2 filter=196 channel=81
					3, 3, 4, 2, 10, -3, -7, 3, 7,
					-- layer=2 filter=196 channel=82
					-2, -5, 8, 6, -2, -2, -8, -4, 5,
					-- layer=2 filter=196 channel=83
					-7, 0, 4, -8, -10, 8, -10, -7, -11,
					-- layer=2 filter=196 channel=84
					-2, -8, 4, 9, -5, 0, 8, 3, -4,
					-- layer=2 filter=196 channel=85
					-10, 0, 2, 5, 4, 6, 4, 2, 0,
					-- layer=2 filter=196 channel=86
					-12, -9, 8, -1, 4, -4, -7, -5, 3,
					-- layer=2 filter=196 channel=87
					-11, 1, 3, 2, 7, 0, 7, 0, -7,
					-- layer=2 filter=196 channel=88
					-4, 4, -12, 6, 0, -11, 2, -5, -5,
					-- layer=2 filter=196 channel=89
					3, -5, -7, -10, 2, -2, -9, 3, -2,
					-- layer=2 filter=196 channel=90
					8, 7, 8, -5, -2, -10, 9, 9, 5,
					-- layer=2 filter=196 channel=91
					-4, -8, 5, -8, -11, -7, -3, -5, -13,
					-- layer=2 filter=196 channel=92
					-9, -8, 10, -4, -1, 0, 8, -4, -6,
					-- layer=2 filter=196 channel=93
					2, -8, 0, -4, 3, -8, -6, 3, 8,
					-- layer=2 filter=196 channel=94
					-8, 0, 3, -3, 3, -3, 7, -4, -6,
					-- layer=2 filter=196 channel=95
					-11, -11, -2, -7, 0, 1, -3, -1, -10,
					-- layer=2 filter=196 channel=96
					0, -5, -7, -5, 3, -2, 5, -9, -10,
					-- layer=2 filter=196 channel=97
					-4, -3, 7, 7, -8, -6, -9, 4, 2,
					-- layer=2 filter=196 channel=98
					0, -13, -1, -3, -4, 12, -3, -2, 6,
					-- layer=2 filter=196 channel=99
					-9, 1, -16, -7, -7, 1, 8, 4, 11,
					-- layer=2 filter=196 channel=100
					7, 1, -5, 4, -8, -2, -2, 5, -9,
					-- layer=2 filter=196 channel=101
					4, -9, 1, -12, -3, -4, -12, 1, -10,
					-- layer=2 filter=196 channel=102
					6, -1, -7, -13, 2, -11, -1, 6, 5,
					-- layer=2 filter=196 channel=103
					6, 1, -3, -5, -1, 7, 8, -7, -7,
					-- layer=2 filter=196 channel=104
					-9, 4, -10, 7, -5, 2, 7, 7, -5,
					-- layer=2 filter=196 channel=105
					-7, -11, -3, 6, 6, -2, 0, 1, 0,
					-- layer=2 filter=196 channel=106
					7, 3, 2, -5, -1, -4, -8, 0, -7,
					-- layer=2 filter=196 channel=107
					-7, 0, 7, -1, 1, 9, 0, -3, 4,
					-- layer=2 filter=196 channel=108
					-14, 5, -9, 2, 0, -3, 11, -3, -7,
					-- layer=2 filter=196 channel=109
					2, -9, 1, -1, -3, 8, 3, 9, -9,
					-- layer=2 filter=196 channel=110
					-11, 3, -1, -19, -10, 5, -6, -11, -4,
					-- layer=2 filter=196 channel=111
					-4, 9, 4, 3, 7, -11, -5, -11, -10,
					-- layer=2 filter=196 channel=112
					-3, -2, -9, -7, -6, 7, -3, -1, -8,
					-- layer=2 filter=196 channel=113
					6, -9, 1, 0, -7, -5, -9, -9, 0,
					-- layer=2 filter=196 channel=114
					4, 9, -2, 6, -4, -9, -8, 8, 5,
					-- layer=2 filter=196 channel=115
					4, -4, 6, 2, -10, 2, -4, 1, 5,
					-- layer=2 filter=196 channel=116
					-7, -1, -9, -4, -12, -7, -6, -6, -14,
					-- layer=2 filter=196 channel=117
					-13, -14, -4, -2, -3, -3, -13, -7, 5,
					-- layer=2 filter=196 channel=118
					-2, 4, 0, 5, -2, -1, -8, -1, -5,
					-- layer=2 filter=196 channel=119
					11, -4, -10, -1, -15, -4, 0, 0, -17,
					-- layer=2 filter=196 channel=120
					-2, -5, -7, 6, -5, 8, -1, 6, 3,
					-- layer=2 filter=196 channel=121
					0, 3, -5, 11, 11, 8, -1, -2, 6,
					-- layer=2 filter=196 channel=122
					0, -2, -8, 8, -11, 1, -5, 9, -7,
					-- layer=2 filter=196 channel=123
					-3, -12, 5, -3, -9, -6, -7, -2, 10,
					-- layer=2 filter=196 channel=124
					-6, 0, 10, -2, -13, -14, -6, -7, -3,
					-- layer=2 filter=196 channel=125
					0, 3, 0, 8, -11, 2, -5, 0, -5,
					-- layer=2 filter=196 channel=126
					7, 2, 7, 4, 7, 2, -10, 8, -4,
					-- layer=2 filter=196 channel=127
					0, 1, -3, -13, 0, -15, -5, -6, -8,
					-- layer=2 filter=197 channel=0
					-13, -1, -19, -20, -9, -7, -16, -22, -14,
					-- layer=2 filter=197 channel=1
					11, 5, 8, 11, 0, -4, -10, 0, -17,
					-- layer=2 filter=197 channel=2
					7, -4, -4, -8, 0, -9, 1, 4, 0,
					-- layer=2 filter=197 channel=3
					-17, -6, -17, -12, -5, -13, -20, -16, -3,
					-- layer=2 filter=197 channel=4
					-17, -23, -18, -6, -16, -19, -10, -6, -8,
					-- layer=2 filter=197 channel=5
					-11, -21, -11, -24, -10, -18, -15, -18, -7,
					-- layer=2 filter=197 channel=6
					-14, 16, 14, -37, -14, 6, -15, -13, -5,
					-- layer=2 filter=197 channel=7
					-14, -14, -5, -2, -1, -10, 0, -14, 7,
					-- layer=2 filter=197 channel=8
					-10, 4, 6, -6, 10, -6, -6, -4, 6,
					-- layer=2 filter=197 channel=9
					-28, -2, -3, -26, -25, -31, -10, -9, -27,
					-- layer=2 filter=197 channel=10
					-17, -23, -20, -12, -20, -11, -11, -18, -13,
					-- layer=2 filter=197 channel=11
					-6, -19, -14, -15, -15, -3, -17, -19, -5,
					-- layer=2 filter=197 channel=12
					-8, -14, -15, -13, -22, -21, -14, -8, -21,
					-- layer=2 filter=197 channel=13
					0, -8, 5, 0, 7, -1, -7, 7, -9,
					-- layer=2 filter=197 channel=14
					-2, 1, -1, -3, -12, -17, -7, -19, -15,
					-- layer=2 filter=197 channel=15
					1, -6, -6, 7, -14, -17, -17, -10, -1,
					-- layer=2 filter=197 channel=16
					0, -1, 8, 12, 4, 8, 5, 18, 5,
					-- layer=2 filter=197 channel=17
					2, 3, 10, 8, 1, -3, -7, -10, -8,
					-- layer=2 filter=197 channel=18
					-21, -16, 2, 3, -30, -19, -5, -17, -16,
					-- layer=2 filter=197 channel=19
					5, 6, 7, -19, -1, -4, -9, -8, -5,
					-- layer=2 filter=197 channel=20
					4, -10, -3, 4, -9, 6, 10, -9, -2,
					-- layer=2 filter=197 channel=21
					8, -7, -9, -5, 2, 1, 5, -5, 3,
					-- layer=2 filter=197 channel=22
					0, 8, -1, 4, -9, -1, 0, -2, -9,
					-- layer=2 filter=197 channel=23
					-7, -12, -15, -1, 1, -2, -8, 4, 0,
					-- layer=2 filter=197 channel=24
					-20, -5, -20, -22, -15, -11, -24, -16, -19,
					-- layer=2 filter=197 channel=25
					-10, 2, 0, -6, -8, -2, -14, 0, 0,
					-- layer=2 filter=197 channel=26
					-7, -4, -2, 7, -6, 0, 2, 10, 2,
					-- layer=2 filter=197 channel=27
					-20, -4, 4, -2, -8, 1, -11, -15, -35,
					-- layer=2 filter=197 channel=28
					-16, -4, 2, -3, 8, 5, -8, -6, -1,
					-- layer=2 filter=197 channel=29
					-10, 8, 1, -9, 6, 8, -2, -2, -2,
					-- layer=2 filter=197 channel=30
					-3, -16, -17, 5, -2, -23, 3, -5, -12,
					-- layer=2 filter=197 channel=31
					7, -17, 7, -1, -22, 13, -17, -4, 32,
					-- layer=2 filter=197 channel=32
					7, -9, 0, -6, -1, 9, -8, -8, 8,
					-- layer=2 filter=197 channel=33
					-25, 0, 4, 0, -10, -8, -21, -17, -6,
					-- layer=2 filter=197 channel=34
					-9, -18, -1, 24, -7, -5, 15, -40, 0,
					-- layer=2 filter=197 channel=35
					-10, -6, -12, 9, 12, 0, -2, -5, -16,
					-- layer=2 filter=197 channel=36
					8, 10, 4, -1, 0, 2, -8, -2, -3,
					-- layer=2 filter=197 channel=37
					-14, -15, -9, -4, -15, -14, -17, -8, -7,
					-- layer=2 filter=197 channel=38
					-3, -15, -13, -16, 0, -14, -10, -9, -24,
					-- layer=2 filter=197 channel=39
					-9, 0, -7, 1, 3, -16, -1, 16, 6,
					-- layer=2 filter=197 channel=40
					-6, 18, 0, 8, -26, 2, -28, -15, -14,
					-- layer=2 filter=197 channel=41
					7, 1, 8, 7, 4, -4, -7, 5, 6,
					-- layer=2 filter=197 channel=42
					-5, 0, 3, -4, 2, 13, -2, -5, 0,
					-- layer=2 filter=197 channel=43
					-17, -12, -2, -17, -8, -17, -10, -22, -7,
					-- layer=2 filter=197 channel=44
					-5, 0, -6, 9, -5, 5, -1, 5, 9,
					-- layer=2 filter=197 channel=45
					9, 3, 2, -12, -17, -19, -9, -1, 2,
					-- layer=2 filter=197 channel=46
					-13, -16, -15, -7, -4, -9, -18, -12, -19,
					-- layer=2 filter=197 channel=47
					-4, 5, -16, -26, -9, -22, -5, -3, -10,
					-- layer=2 filter=197 channel=48
					-1, 0, 8, -3, -4, -7, 2, -1, -3,
					-- layer=2 filter=197 channel=49
					-18, -31, 6, -3, -31, 1, 7, -21, -6,
					-- layer=2 filter=197 channel=50
					8, -3, 3, -9, -5, 9, 9, -6, -9,
					-- layer=2 filter=197 channel=51
					-16, -10, -9, -11, -15, -8, -24, -14, -18,
					-- layer=2 filter=197 channel=52
					2, -10, -20, -8, -19, -10, 0, -20, -13,
					-- layer=2 filter=197 channel=53
					-16, -9, 3, 0, -6, -4, 5, -11, -3,
					-- layer=2 filter=197 channel=54
					-15, -18, -3, -9, -16, -14, 0, -12, -18,
					-- layer=2 filter=197 channel=55
					-5, 7, -9, 0, -1, 3, -4, -9, -9,
					-- layer=2 filter=197 channel=56
					-8, -8, -6, -14, -9, -21, -9, -10, -21,
					-- layer=2 filter=197 channel=57
					0, -10, 1, -5, -5, 1, 9, 8, 8,
					-- layer=2 filter=197 channel=58
					-2, -5, -22, -1, -20, -11, -8, 0, -13,
					-- layer=2 filter=197 channel=59
					1, -1, -13, 0, -12, -6, -12, -11, -8,
					-- layer=2 filter=197 channel=60
					-4, -16, -24, -7, -16, -9, -10, -27, -9,
					-- layer=2 filter=197 channel=61
					-9, 7, -3, -14, -10, -21, -15, -8, -13,
					-- layer=2 filter=197 channel=62
					1, -15, 2, 6, -5, 7, -15, -23, -14,
					-- layer=2 filter=197 channel=63
					-9, 2, -14, -15, 0, -17, -7, 2, -8,
					-- layer=2 filter=197 channel=64
					-13, -1, -16, -7, -15, 8, -9, -4, 5,
					-- layer=2 filter=197 channel=65
					2, 0, -9, -15, -9, 1, -24, -7, 6,
					-- layer=2 filter=197 channel=66
					21, 12, -3, 4, 6, 15, 0, 11, -9,
					-- layer=2 filter=197 channel=67
					-17, -10, -24, -29, -11, -28, -15, -17, -20,
					-- layer=2 filter=197 channel=68
					6, 0, -2, 10, 4, 5, 9, -8, -4,
					-- layer=2 filter=197 channel=69
					0, -2, -11, 8, -13, -3, -2, 0, 10,
					-- layer=2 filter=197 channel=70
					-2, -10, -9, -15, 6, -9, -17, -13, -15,
					-- layer=2 filter=197 channel=71
					-11, -4, -3, -10, 5, -6, -6, -7, -3,
					-- layer=2 filter=197 channel=72
					2, 13, 5, 3, -12, -20, -19, -1, -15,
					-- layer=2 filter=197 channel=73
					1, 14, 3, -24, -24, -6, -22, -13, -13,
					-- layer=2 filter=197 channel=74
					-11, -15, -1, -6, -13, -8, -18, -1, -17,
					-- layer=2 filter=197 channel=75
					-7, 10, 20, -5, 6, 17, -15, -7, -7,
					-- layer=2 filter=197 channel=76
					-6, -5, -2, -12, -5, 5, -7, -15, -6,
					-- layer=2 filter=197 channel=77
					5, 2, -11, -4, -5, -2, -4, 2, 5,
					-- layer=2 filter=197 channel=78
					-16, -15, 4, -14, -22, -14, -4, -7, -19,
					-- layer=2 filter=197 channel=79
					5, 8, -2, 1, -5, -6, -6, -10, -5,
					-- layer=2 filter=197 channel=80
					-6, -13, -21, -9, -2, 4, -3, 4, -10,
					-- layer=2 filter=197 channel=81
					5, -9, 0, -4, -1, -2, 6, 0, -11,
					-- layer=2 filter=197 channel=82
					1, 10, 9, -9, 7, 0, 4, 8, 3,
					-- layer=2 filter=197 channel=83
					8, -1, -1, 8, -2, 3, 0, -2, 10,
					-- layer=2 filter=197 channel=84
					-5, -11, -6, 2, -4, -11, -10, -5, 0,
					-- layer=2 filter=197 channel=85
					-1, 6, -9, -3, 4, 6, -3, 8, 0,
					-- layer=2 filter=197 channel=86
					1, 0, 2, 8, -8, 5, 4, 1, -2,
					-- layer=2 filter=197 channel=87
					-7, -10, -7, 9, 11, 9, -7, -22, 0,
					-- layer=2 filter=197 channel=88
					-5, -3, -9, -9, 0, -13, -4, 6, -9,
					-- layer=2 filter=197 channel=89
					6, -2, -7, 19, -1, -9, -1, 5, -22,
					-- layer=2 filter=197 channel=90
					-6, 7, 3, 9, 1, 1, 3, -10, -2,
					-- layer=2 filter=197 channel=91
					-9, -11, -4, -5, -5, -8, -6, 8, -23,
					-- layer=2 filter=197 channel=92
					-12, 6, -2, 8, -6, -20, -6, -10, -8,
					-- layer=2 filter=197 channel=93
					13, 10, 11, -2, -8, 18, -2, -20, 17,
					-- layer=2 filter=197 channel=94
					-37, 9, 2, -16, -4, -8, -26, -6, -16,
					-- layer=2 filter=197 channel=95
					-7, 8, -6, -9, -3, -10, 4, -3, -8,
					-- layer=2 filter=197 channel=96
					-11, -22, 0, -3, -6, -8, -8, -7, 3,
					-- layer=2 filter=197 channel=97
					-27, -16, -13, -13, -19, -14, -18, -21, -13,
					-- layer=2 filter=197 channel=98
					-9, 1, -17, -3, 6, -8, -15, -3, -12,
					-- layer=2 filter=197 channel=99
					-4, -14, -4, -12, -13, -14, -15, -10, -15,
					-- layer=2 filter=197 channel=100
					0, -11, -7, -6, -2, 6, -7, 6, -2,
					-- layer=2 filter=197 channel=101
					-23, -12, 11, 0, -13, -12, 0, -15, 2,
					-- layer=2 filter=197 channel=102
					-10, -20, 2, 14, -4, -13, 12, -14, -5,
					-- layer=2 filter=197 channel=103
					-25, -19, -27, 22, 3, -4, -2, -6, -1,
					-- layer=2 filter=197 channel=104
					-18, -7, 11, 8, -25, 4, -5, -16, -5,
					-- layer=2 filter=197 channel=105
					-23, 11, 3, -5, 12, -1, -14, -16, -18,
					-- layer=2 filter=197 channel=106
					-22, -30, -12, -12, -2, -21, -25, -2, -25,
					-- layer=2 filter=197 channel=107
					-13, 12, 21, -5, -6, -14, -4, 2, 2,
					-- layer=2 filter=197 channel=108
					-11, -10, 3, -3, -15, -1, -5, -9, -8,
					-- layer=2 filter=197 channel=109
					-8, -2, 7, -1, 0, 8, -5, 0, -7,
					-- layer=2 filter=197 channel=110
					-2, -2, -15, 5, 2, 9, -5, -1, 12,
					-- layer=2 filter=197 channel=111
					5, 4, -4, 1, 2, -5, 7, 3, 9,
					-- layer=2 filter=197 channel=112
					-23, -20, -9, -6, -9, -20, -19, -4, -16,
					-- layer=2 filter=197 channel=113
					0, -13, -7, -12, 8, -16, 1, 10, -11,
					-- layer=2 filter=197 channel=114
					4, 4, 4, -6, -9, 5, -2, -8, -6,
					-- layer=2 filter=197 channel=115
					-10, -1, -4, 8, -3, -9, 1, 7, 0,
					-- layer=2 filter=197 channel=116
					-5, -4, -8, 14, -1, -14, -14, -27, -10,
					-- layer=2 filter=197 channel=117
					-24, -12, 2, -15, -13, 0, 11, 0, -14,
					-- layer=2 filter=197 channel=118
					-25, -23, -6, -13, -6, -3, -18, -24, -13,
					-- layer=2 filter=197 channel=119
					-6, -16, -9, -8, -30, -11, 0, 0, 2,
					-- layer=2 filter=197 channel=120
					-8, -1, 6, 4, 0, 5, 4, -7, 0,
					-- layer=2 filter=197 channel=121
					-8, 2, 7, 4, -4, 2, -10, 10, 7,
					-- layer=2 filter=197 channel=122
					8, 6, 11, -6, -3, 0, -2, -2, -1,
					-- layer=2 filter=197 channel=123
					-24, 4, -3, 3, -10, -19, -11, -16, -8,
					-- layer=2 filter=197 channel=124
					-8, 6, 11, -6, -13, -3, -1, -20, -1,
					-- layer=2 filter=197 channel=125
					-1, -10, -7, 4, -3, -5, -1, 10, 1,
					-- layer=2 filter=197 channel=126
					-18, 0, 1, -8, -20, -19, 0, -3, -9,
					-- layer=2 filter=197 channel=127
					-5, 0, -4, 1, -20, -7, -1, -11, -11,
					-- layer=2 filter=198 channel=0
					10, 24, 6, 9, 13, 11, -11, -13, 9,
					-- layer=2 filter=198 channel=1
					6, -13, 22, 2, 27, 7, -28, -27, -15,
					-- layer=2 filter=198 channel=2
					11, 11, 8, -4, 0, 3, 11, 7, 1,
					-- layer=2 filter=198 channel=3
					19, 25, -23, -39, -20, -14, -11, 1, -17,
					-- layer=2 filter=198 channel=4
					15, -22, 17, 0, 0, -24, -49, -5, 4,
					-- layer=2 filter=198 channel=5
					7, -7, 21, 1, 16, 28, -12, 0, 15,
					-- layer=2 filter=198 channel=6
					14, -2, -13, 2, 16, -23, 32, -20, -15,
					-- layer=2 filter=198 channel=7
					-2, 17, -1, -7, -29, -25, -33, 18, -24,
					-- layer=2 filter=198 channel=8
					5, -2, -2, 1, -1, 3, -5, -9, -7,
					-- layer=2 filter=198 channel=9
					24, -10, -24, -20, -9, -18, -46, 0, -16,
					-- layer=2 filter=198 channel=10
					-5, 23, -2, -28, -1, 24, -29, -29, -15,
					-- layer=2 filter=198 channel=11
					-8, 38, 8, 17, 15, -1, -15, 11, -21,
					-- layer=2 filter=198 channel=12
					20, 4, 10, 34, 30, 2, -13, -30, -4,
					-- layer=2 filter=198 channel=13
					-2, 9, -8, -4, 1, 11, 5, -5, 0,
					-- layer=2 filter=198 channel=14
					48, -9, 7, 15, 42, 4, 12, -27, -28,
					-- layer=2 filter=198 channel=15
					-37, 8, -43, -18, 25, -27, -9, 2, -64,
					-- layer=2 filter=198 channel=16
					-57, -27, -9, -41, -14, -11, -5, 14, 32,
					-- layer=2 filter=198 channel=17
					2, -3, 9, -6, -12, -8, 8, -7, -10,
					-- layer=2 filter=198 channel=18
					27, 18, 10, 24, 53, -18, 5, 34, -5,
					-- layer=2 filter=198 channel=19
					-31, -31, -7, 31, 59, 32, -45, -10, -50,
					-- layer=2 filter=198 channel=20
					10, 9, -5, 6, 4, 1, 5, -4, -6,
					-- layer=2 filter=198 channel=21
					0, -15, 1, -16, -16, 1, -7, -18, -11,
					-- layer=2 filter=198 channel=22
					-11, -8, 2, -3, 9, 3, -2, -2, -7,
					-- layer=2 filter=198 channel=23
					25, -28, -24, 22, -43, -34, 45, 15, -9,
					-- layer=2 filter=198 channel=24
					17, 4, -2, 12, 38, 26, 51, 61, 39,
					-- layer=2 filter=198 channel=25
					-16, -12, 7, -1, -3, -4, -8, 26, 34,
					-- layer=2 filter=198 channel=26
					10, 7, -2, 9, 3, 3, 4, 0, -12,
					-- layer=2 filter=198 channel=27
					-26, 4, 5, 1, 14, 53, -8, 42, 56,
					-- layer=2 filter=198 channel=28
					-6, -14, -20, -10, 10, -16, -7, -78, -98,
					-- layer=2 filter=198 channel=29
					3, -2, 7, -5, 9, 6, -8, -5, -2,
					-- layer=2 filter=198 channel=30
					18, 18, -6, -46, 0, 23, 0, -4, -29,
					-- layer=2 filter=198 channel=31
					5, -6, 13, 57, 21, 1, -20, 45, 43,
					-- layer=2 filter=198 channel=32
					7, 11, 11, 7, 0, -6, -5, 8, 0,
					-- layer=2 filter=198 channel=33
					10, 7, -40, 27, -10, 4, 11, -6, -25,
					-- layer=2 filter=198 channel=34
					-26, -7, -13, 0, 10, -6, 66, 6, -47,
					-- layer=2 filter=198 channel=35
					-14, -1, -25, 13, -8, -6, 0, -25, -14,
					-- layer=2 filter=198 channel=36
					-1, 6, 16, -1, 9, 9, 1, -10, -1,
					-- layer=2 filter=198 channel=37
					0, 25, 5, 5, 14, 8, 2, 17, 1,
					-- layer=2 filter=198 channel=38
					-7, -5, 16, -30, 9, 28, -33, 3, 27,
					-- layer=2 filter=198 channel=39
					19, 16, -12, 8, 3, -13, 5, 60, 52,
					-- layer=2 filter=198 channel=40
					12, 14, -92, -6, 30, 28, -25, 44, 1,
					-- layer=2 filter=198 channel=41
					-5, 5, 1, 1, 0, 9, 0, -6, -10,
					-- layer=2 filter=198 channel=42
					-8, -10, -3, -8, 0, -8, 39, 21, 2,
					-- layer=2 filter=198 channel=43
					7, -8, -9, -22, -12, -62, -19, -19, -51,
					-- layer=2 filter=198 channel=44
					9, -8, -2, 1, -9, -10, -4, 3, -3,
					-- layer=2 filter=198 channel=45
					13, -5, 34, 21, -1, 24, -3, 23, 26,
					-- layer=2 filter=198 channel=46
					-21, 16, -18, -36, 3, 9, -55, -13, -35,
					-- layer=2 filter=198 channel=47
					19, -2, 0, 9, 24, 6, -20, -28, -49,
					-- layer=2 filter=198 channel=48
					-4, 2, -6, -1, 7, 7, 0, -11, 0,
					-- layer=2 filter=198 channel=49
					5, 2, 28, 57, 22, -7, 0, 7, 6,
					-- layer=2 filter=198 channel=50
					17, -14, 1, -20, 0, 12, 14, 0, -8,
					-- layer=2 filter=198 channel=51
					15, 35, 32, -11, 17, 3, -16, 16, 6,
					-- layer=2 filter=198 channel=52
					-3, 16, 1, -23, -5, 16, -16, 7, 6,
					-- layer=2 filter=198 channel=53
					28, 7, 1, -28, -17, 21, -24, -23, -18,
					-- layer=2 filter=198 channel=54
					-10, -33, -13, -10, -32, -46, 28, -9, -37,
					-- layer=2 filter=198 channel=55
					-3, -6, -5, -9, 8, -5, -3, -11, 0,
					-- layer=2 filter=198 channel=56
					-3, 34, 28, 5, 18, 14, -10, 24, 5,
					-- layer=2 filter=198 channel=57
					3, 7, -2, 0, -3, -4, 10, 8, 2,
					-- layer=2 filter=198 channel=58
					13, 30, 19, 48, -2, 6, 11, -34, -10,
					-- layer=2 filter=198 channel=59
					-11, 22, -6, 29, 3, 34, -25, -12, 26,
					-- layer=2 filter=198 channel=60
					9, 5, 37, -7, 4, 31, -13, -40, -2,
					-- layer=2 filter=198 channel=61
					17, 72, 63, 17, 79, 55, -7, 38, 54,
					-- layer=2 filter=198 channel=62
					-19, -7, -3, -12, 12, -24, -7, -27, -76,
					-- layer=2 filter=198 channel=63
					43, 6, 0, 14, -10, -19, 1, -14, 3,
					-- layer=2 filter=198 channel=64
					29, -11, -27, 29, 6, -14, 61, 30, 13,
					-- layer=2 filter=198 channel=65
					9, 33, 55, 9, 69, 16, -12, 44, 6,
					-- layer=2 filter=198 channel=66
					-48, 19, 26, -20, -27, -51, -1, -23, 40,
					-- layer=2 filter=198 channel=67
					-10, -10, -25, -33, -7, 13, -33, -27, -56,
					-- layer=2 filter=198 channel=68
					0, -5, -6, -5, -2, 11, 6, -1, 7,
					-- layer=2 filter=198 channel=69
					29, -22, -28, 12, -7, -17, 55, 18, 17,
					-- layer=2 filter=198 channel=70
					-5, -12, -2, 16, 18, -8, -9, -57, -61,
					-- layer=2 filter=198 channel=71
					-36, -15, -7, 33, 22, 18, 12, 16, 6,
					-- layer=2 filter=198 channel=72
					-2, -10, -14, 27, 35, 6, 26, 24, -14,
					-- layer=2 filter=198 channel=73
					-4, -14, -21, 31, -50, 25, 54, -18, -33,
					-- layer=2 filter=198 channel=74
					31, 33, -31, 6, -17, -6, -29, -31, 9,
					-- layer=2 filter=198 channel=75
					-33, 23, 0, -7, 22, -3, -61, -76, -94,
					-- layer=2 filter=198 channel=76
					-6, 10, 3, -80, -26, 2, 13, 7, -10,
					-- layer=2 filter=198 channel=77
					-3, -2, 6, 7, 0, -8, 2, -3, -1,
					-- layer=2 filter=198 channel=78
					-14, 0, 36, 31, 21, -21, -4, -8, -17,
					-- layer=2 filter=198 channel=79
					0, -7, -1, 9, -7, -3, -7, 10, -7,
					-- layer=2 filter=198 channel=80
					20, 1, -15, -24, -22, -34, -9, 9, 19,
					-- layer=2 filter=198 channel=81
					-10, 8, -6, -2, 3, 7, -12, -2, -1,
					-- layer=2 filter=198 channel=82
					-6, -4, 10, 1, -9, -3, -1, -8, -10,
					-- layer=2 filter=198 channel=83
					21, -24, 5, 12, -5, -12, -18, 8, -38,
					-- layer=2 filter=198 channel=84
					3, 8, 9, 7, 7, -4, -7, 3, -6,
					-- layer=2 filter=198 channel=85
					7, -1, -14, -17, 0, 0, 6, 2, 10,
					-- layer=2 filter=198 channel=86
					-1, -13, -7, 2, 6, -15, -11, 0, 2,
					-- layer=2 filter=198 channel=87
					14, -35, 0, -8, 10, -37, 25, 9, -35,
					-- layer=2 filter=198 channel=88
					43, 3, -16, -19, 8, -29, -12, -6, -7,
					-- layer=2 filter=198 channel=89
					3, -21, -13, 43, 41, 2, 26, -27, -36,
					-- layer=2 filter=198 channel=90
					-8, 6, -5, -5, -6, 9, -5, 0, -8,
					-- layer=2 filter=198 channel=91
					-1, -9, -9, 5, 17, 24, 0, -49, 14,
					-- layer=2 filter=198 channel=92
					18, -30, 23, 13, 47, 20, -3, -5, 15,
					-- layer=2 filter=198 channel=93
					28, -6, 21, 35, 48, 39, 2, 10, -23,
					-- layer=2 filter=198 channel=94
					4, -24, 8, -19, 20, 8, -43, 0, -5,
					-- layer=2 filter=198 channel=95
					1, 12, 21, 12, -1, 18, 18, 18, 26,
					-- layer=2 filter=198 channel=96
					22, -19, 20, 8, -26, -23, 36, 13, -9,
					-- layer=2 filter=198 channel=97
					15, -15, -44, 16, 21, -5, -21, -4, -14,
					-- layer=2 filter=198 channel=98
					-2, 19, 4, 27, 15, 4, -16, -31, -34,
					-- layer=2 filter=198 channel=99
					-10, -24, -21, -14, 17, 18, -36, -26, 25,
					-- layer=2 filter=198 channel=100
					24, -22, -15, -24, 5, 42, -17, -14, 0,
					-- layer=2 filter=198 channel=101
					-6, 9, -15, 30, 1, 14, -16, -11, -5,
					-- layer=2 filter=198 channel=102
					12, -21, 12, 31, 8, -3, -29, -6, 17,
					-- layer=2 filter=198 channel=103
					-24, -63, -18, -35, 21, 15, -26, 16, 1,
					-- layer=2 filter=198 channel=104
					-28, -16, 15, 22, 8, 19, -12, 1, -46,
					-- layer=2 filter=198 channel=105
					-77, -13, 0, -24, 26, 21, -31, -1, -23,
					-- layer=2 filter=198 channel=106
					-11, -11, -8, -8, 22, -1, -42, 0, 0,
					-- layer=2 filter=198 channel=107
					27, -72, -5, -40, -31, -9, -44, -10, -48,
					-- layer=2 filter=198 channel=108
					-10, -19, 15, 6, 13, -6, -36, -19, -14,
					-- layer=2 filter=198 channel=109
					0, 4, 0, 10, 12, -1, 4, 4, 2,
					-- layer=2 filter=198 channel=110
					0, -23, 10, 38, 10, 25, 91, 75, 50,
					-- layer=2 filter=198 channel=111
					-2, 4, 4, -7, 9, -2, -2, 8, 5,
					-- layer=2 filter=198 channel=112
					-3, 41, 16, 7, 19, 31, -48, 14, -17,
					-- layer=2 filter=198 channel=113
					-10, 13, 47, 1, 16, 23, 13, 22, -40,
					-- layer=2 filter=198 channel=114
					12, 10, 0, -1, -12, 0, 5, 3, -1,
					-- layer=2 filter=198 channel=115
					-7, 2, 8, -9, -4, -9, 2, 5, 7,
					-- layer=2 filter=198 channel=116
					-10, -28, -10, -13, -10, -67, -22, 0, -43,
					-- layer=2 filter=198 channel=117
					-20, -11, -2, -32, 8, 5, 5, 7, -77,
					-- layer=2 filter=198 channel=118
					4, -3, 0, 7, -1, -40, 7, -6, -7,
					-- layer=2 filter=198 channel=119
					-11, -5, 14, -27, 25, -10, 24, -7, 11,
					-- layer=2 filter=198 channel=120
					5, -2, -5, 6, -8, -4, 0, 2, 0,
					-- layer=2 filter=198 channel=121
					4, -7, -3, -6, 1, -10, 5, 5, 3,
					-- layer=2 filter=198 channel=122
					-13, 5, -5, 5, 2, -3, 15, 3, 6,
					-- layer=2 filter=198 channel=123
					30, -20, -6, -7, -6, -14, 0, -8, -69,
					-- layer=2 filter=198 channel=124
					-11, -17, -20, -18, 13, -38, 37, 8, -65,
					-- layer=2 filter=198 channel=125
					-6, 2, -10, -8, -5, 10, -8, 0, -8,
					-- layer=2 filter=198 channel=126
					6, 17, -2, -25, 48, -10, 38, -9, -17,
					-- layer=2 filter=198 channel=127
					27, -16, 18, 0, 11, 9, -11, -13, 6,
					-- layer=2 filter=199 channel=0
					-7, -2, -9, 8, -7, 7, -3, -1, -3,
					-- layer=2 filter=199 channel=1
					1, -4, -7, 0, -6, -1, -10, -9, -10,
					-- layer=2 filter=199 channel=2
					-5, 1, 5, 4, 1, -6, 0, -7, 5,
					-- layer=2 filter=199 channel=3
					-3, 6, -5, -8, 0, -7, 0, -14, -8,
					-- layer=2 filter=199 channel=4
					2, 0, -8, 2, -8, -2, -7, 3, 8,
					-- layer=2 filter=199 channel=5
					0, -4, -12, -2, 3, 5, 7, -10, 2,
					-- layer=2 filter=199 channel=6
					6, 13, -10, -10, 7, 0, 6, -1, 7,
					-- layer=2 filter=199 channel=7
					6, -2, -4, 6, 7, -8, 1, -3, -4,
					-- layer=2 filter=199 channel=8
					-5, -3, 10, 8, -5, 10, -8, -8, 6,
					-- layer=2 filter=199 channel=9
					-3, -9, 0, -5, -9, 3, -11, 0, -3,
					-- layer=2 filter=199 channel=10
					-10, 7, 5, -6, -8, -9, -7, 5, 1,
					-- layer=2 filter=199 channel=11
					-5, -9, 1, 1, -6, -5, -11, -12, -3,
					-- layer=2 filter=199 channel=12
					-12, -5, 3, -6, 3, 0, -15, 9, 5,
					-- layer=2 filter=199 channel=13
					8, 8, -2, -7, -1, -5, -6, 3, 5,
					-- layer=2 filter=199 channel=14
					0, -4, -10, -13, 2, -10, -9, -2, 2,
					-- layer=2 filter=199 channel=15
					-14, 0, 6, -6, -7, -5, 0, -9, 0,
					-- layer=2 filter=199 channel=16
					5, -9, 6, 7, -5, -10, -3, 5, -6,
					-- layer=2 filter=199 channel=17
					10, 5, -8, -6, -2, -6, 7, 7, 10,
					-- layer=2 filter=199 channel=18
					-12, 3, 0, -8, 4, 6, 0, 2, -3,
					-- layer=2 filter=199 channel=19
					-1, 6, 13, 0, 1, -2, 3, -11, -14,
					-- layer=2 filter=199 channel=20
					2, 8, -1, -1, -8, -3, 7, -4, -4,
					-- layer=2 filter=199 channel=21
					4, -3, -2, -11, -11, 6, 0, -10, 0,
					-- layer=2 filter=199 channel=22
					3, 3, -5, 0, 4, 5, -8, -10, -3,
					-- layer=2 filter=199 channel=23
					-11, -4, 1, -7, -11, 7, -13, -11, -11,
					-- layer=2 filter=199 channel=24
					-5, -17, 1, -13, 0, -12, -5, -5, -7,
					-- layer=2 filter=199 channel=25
					-1, 0, 6, -9, 3, -5, -13, 4, 0,
					-- layer=2 filter=199 channel=26
					-10, 2, -1, -1, -7, -6, 0, -3, 7,
					-- layer=2 filter=199 channel=27
					-3, -7, 10, 5, 0, 1, -2, -10, -8,
					-- layer=2 filter=199 channel=28
					0, -5, -6, -3, -11, -6, 1, -8, 0,
					-- layer=2 filter=199 channel=29
					1, 5, -4, -5, 3, -3, -4, -10, 6,
					-- layer=2 filter=199 channel=30
					-14, -11, 0, -2, -4, 7, -10, 6, -11,
					-- layer=2 filter=199 channel=31
					-10, -1, -8, 6, 0, 2, 8, -3, 2,
					-- layer=2 filter=199 channel=32
					-10, -6, -8, 0, 9, -7, 3, -5, -8,
					-- layer=2 filter=199 channel=33
					-7, -1, 9, -4, 4, 5, -11, -10, -4,
					-- layer=2 filter=199 channel=34
					-4, -2, -7, -2, 5, -5, 0, 6, -7,
					-- layer=2 filter=199 channel=35
					0, -7, -5, 2, -1, 2, 5, -10, 4,
					-- layer=2 filter=199 channel=36
					-9, -4, 0, -7, 5, -4, 8, -6, 7,
					-- layer=2 filter=199 channel=37
					-15, 0, 5, -12, 0, 4, 5, -12, 1,
					-- layer=2 filter=199 channel=38
					0, -3, -9, 7, 3, -10, 0, -1, 5,
					-- layer=2 filter=199 channel=39
					3, -5, 0, -4, 7, 5, -1, -1, -4,
					-- layer=2 filter=199 channel=40
					-11, 3, -8, 2, -10, 2, -3, -5, 3,
					-- layer=2 filter=199 channel=41
					9, -2, -2, -11, 5, -9, -2, -7, -1,
					-- layer=2 filter=199 channel=42
					-3, 0, -9, 1, 0, 2, -11, 0, -6,
					-- layer=2 filter=199 channel=43
					-3, -9, -10, 4, -9, 3, -10, -3, 3,
					-- layer=2 filter=199 channel=44
					8, 0, 2, -6, -4, 9, -8, 3, -1,
					-- layer=2 filter=199 channel=45
					-10, -6, -10, 6, 5, -3, -7, 7, 3,
					-- layer=2 filter=199 channel=46
					-7, 1, 0, -11, -1, 0, -10, 2, -11,
					-- layer=2 filter=199 channel=47
					-5, -2, -7, -12, -7, 0, 0, -15, 4,
					-- layer=2 filter=199 channel=48
					8, -7, 3, 1, 6, 0, -4, 11, 5,
					-- layer=2 filter=199 channel=49
					2, 0, 3, -2, 1, 0, -5, -6, 3,
					-- layer=2 filter=199 channel=50
					-3, 4, -6, -9, 10, -5, -5, -5, 4,
					-- layer=2 filter=199 channel=51
					-15, -9, -9, -11, 5, -13, -11, -13, -13,
					-- layer=2 filter=199 channel=52
					-16, -2, -6, 5, 4, -10, -1, -5, -3,
					-- layer=2 filter=199 channel=53
					8, -7, -3, 1, -1, 10, 3, 3, 9,
					-- layer=2 filter=199 channel=54
					-2, -5, -16, -12, 6, -2, 0, -5, -4,
					-- layer=2 filter=199 channel=55
					6, -4, 3, -9, -7, 0, -9, 5, -6,
					-- layer=2 filter=199 channel=56
					-11, 0, -7, -8, -3, -10, -3, -1, 0,
					-- layer=2 filter=199 channel=57
					4, 4, -9, 8, -9, 0, 8, -2, -8,
					-- layer=2 filter=199 channel=58
					-13, -4, 3, -11, -8, 4, -5, 12, -3,
					-- layer=2 filter=199 channel=59
					-4, 9, -6, 0, 1, 4, 1, 2, -3,
					-- layer=2 filter=199 channel=60
					-1, -5, 2, -9, -10, -13, 0, 0, 0,
					-- layer=2 filter=199 channel=61
					-2, 0, 4, 1, 5, -2, -12, -8, -14,
					-- layer=2 filter=199 channel=62
					-6, -13, -2, -5, -9, -5, -7, -5, 1,
					-- layer=2 filter=199 channel=63
					-10, 4, 2, -4, -9, 2, -8, 0, 5,
					-- layer=2 filter=199 channel=64
					4, -3, 0, 0, 1, -11, -13, -4, 1,
					-- layer=2 filter=199 channel=65
					0, 0, -10, -9, -10, -7, -13, 8, 6,
					-- layer=2 filter=199 channel=66
					3, 7, -5, 3, 8, 4, -6, 8, -1,
					-- layer=2 filter=199 channel=67
					-9, -6, -12, 0, 1, -8, 0, 3, 2,
					-- layer=2 filter=199 channel=68
					7, -1, -3, 0, 2, -9, -7, -9, 0,
					-- layer=2 filter=199 channel=69
					-2, 6, -10, -5, -14, 0, 1, -3, 4,
					-- layer=2 filter=199 channel=70
					5, 1, -10, 4, 7, 3, 0, 1, -1,
					-- layer=2 filter=199 channel=71
					2, 7, 0, 5, -8, 7, -7, -2, -1,
					-- layer=2 filter=199 channel=72
					0, 5, -6, -8, 1, -4, 5, -10, -13,
					-- layer=2 filter=199 channel=73
					-13, 8, -2, -2, -3, -1, -1, 6, 8,
					-- layer=2 filter=199 channel=74
					4, 0, -11, -6, 1, -3, -1, -1, -8,
					-- layer=2 filter=199 channel=75
					1, 4, 0, 6, 0, 9, -5, 8, -3,
					-- layer=2 filter=199 channel=76
					0, 10, -13, -6, -1, 10, 0, 0, 0,
					-- layer=2 filter=199 channel=77
					-10, 0, -4, -7, -2, -8, 0, -4, 0,
					-- layer=2 filter=199 channel=78
					2, -1, 3, 4, -4, -6, -5, 4, -8,
					-- layer=2 filter=199 channel=79
					-10, 7, 5, 5, -7, 7, -1, -11, 9,
					-- layer=2 filter=199 channel=80
					-11, 5, 4, -4, 3, -6, 1, -5, -3,
					-- layer=2 filter=199 channel=81
					-10, 7, -9, -9, 3, -1, -5, -8, -6,
					-- layer=2 filter=199 channel=82
					5, -10, -8, 5, -11, -6, 1, 4, 2,
					-- layer=2 filter=199 channel=83
					3, -9, 3, -6, -6, 3, -10, 6, 1,
					-- layer=2 filter=199 channel=84
					-4, 2, -3, 8, 6, 0, -1, 6, 0,
					-- layer=2 filter=199 channel=85
					4, 5, 1, -7, 5, 4, -8, -1, -2,
					-- layer=2 filter=199 channel=86
					-1, -10, 0, -5, -11, 3, -4, -11, -6,
					-- layer=2 filter=199 channel=87
					-15, -9, -4, -5, -11, 4, 2, -4, -10,
					-- layer=2 filter=199 channel=88
					-12, -10, -11, 7, 7, 5, -5, -8, -8,
					-- layer=2 filter=199 channel=89
					3, 7, 2, -12, -5, -9, 5, -13, -3,
					-- layer=2 filter=199 channel=90
					10, 2, 5, -6, -4, -3, 4, -1, -5,
					-- layer=2 filter=199 channel=91
					-8, -3, -2, 6, -2, -2, 5, -9, -4,
					-- layer=2 filter=199 channel=92
					0, 6, -9, 0, -10, -2, -6, -8, 4,
					-- layer=2 filter=199 channel=93
					-2, -2, -13, -6, -2, -2, -4, 4, -11,
					-- layer=2 filter=199 channel=94
					13, 4, 6, 6, -6, 12, 4, 10, -7,
					-- layer=2 filter=199 channel=95
					-8, -2, 9, -1, -4, -11, 8, 9, -4,
					-- layer=2 filter=199 channel=96
					-6, -5, -3, 0, -7, -1, -8, -7, 7,
					-- layer=2 filter=199 channel=97
					-1, -3, -14, -7, 5, -4, -2, -9, -4,
					-- layer=2 filter=199 channel=98
					0, -2, 2, -10, 6, -1, -9, -9, -8,
					-- layer=2 filter=199 channel=99
					1, -3, 8, -3, -3, 3, -6, -5, 7,
					-- layer=2 filter=199 channel=100
					2, 7, -11, -8, -10, 3, -1, 3, -11,
					-- layer=2 filter=199 channel=101
					0, 0, -10, -10, -2, -3, 4, -9, -5,
					-- layer=2 filter=199 channel=102
					-10, 0, 4, -7, 7, 0, -8, -10, 2,
					-- layer=2 filter=199 channel=103
					-1, 0, -11, 8, 0, -6, 3, -2, -7,
					-- layer=2 filter=199 channel=104
					-8, -13, 0, 4, -10, -11, 0, 4, 2,
					-- layer=2 filter=199 channel=105
					4, 3, -3, 1, -12, 5, -10, 6, 0,
					-- layer=2 filter=199 channel=106
					-14, -3, 2, -11, 0, 0, 11, -2, 6,
					-- layer=2 filter=199 channel=107
					-2, 1, -3, -5, 7, -9, -3, 4, 7,
					-- layer=2 filter=199 channel=108
					3, -13, 6, -14, 5, 5, 0, 5, 1,
					-- layer=2 filter=199 channel=109
					9, -7, 7, 3, -8, -7, -3, 0, 4,
					-- layer=2 filter=199 channel=110
					0, -4, 2, -2, 7, -9, 0, -4, -5,
					-- layer=2 filter=199 channel=111
					1, 6, -4, -10, 7, -5, 5, 2, 2,
					-- layer=2 filter=199 channel=112
					4, -7, -4, 0, 3, 0, -9, 3, -2,
					-- layer=2 filter=199 channel=113
					-11, 3, -11, -13, -5, -10, -7, 0, -11,
					-- layer=2 filter=199 channel=114
					-9, 4, 3, -9, 5, 1, 10, -3, -9,
					-- layer=2 filter=199 channel=115
					-3, 0, 8, 0, -9, -4, -7, 1, -5,
					-- layer=2 filter=199 channel=116
					-4, 0, -10, 6, 5, -8, -8, 3, 4,
					-- layer=2 filter=199 channel=117
					0, -6, -5, 4, 5, -8, -13, -1, -2,
					-- layer=2 filter=199 channel=118
					-2, -4, -8, -2, -2, 6, 0, -6, -10,
					-- layer=2 filter=199 channel=119
					3, -4, -11, -13, 8, -9, 6, 4, 2,
					-- layer=2 filter=199 channel=120
					3, 7, 10, 7, 9, -9, 9, -4, 0,
					-- layer=2 filter=199 channel=121
					1, 2, 5, -6, 1, -3, -5, -9, 7,
					-- layer=2 filter=199 channel=122
					3, 8, -8, 7, 4, 0, -4, 10, 1,
					-- layer=2 filter=199 channel=123
					-4, -1, -5, -1, -1, 3, 2, 0, -11,
					-- layer=2 filter=199 channel=124
					-2, -3, 3, 0, -7, 6, 0, 1, 1,
					-- layer=2 filter=199 channel=125
					6, -4, -6, 6, 10, 1, 3, 3, 5,
					-- layer=2 filter=199 channel=126
					-1, 5, 7, -11, -4, -9, 1, -1, 4,
					-- layer=2 filter=199 channel=127
					-3, 7, -6, -1, 2, 8, -12, -11, -9,
					-- layer=2 filter=200 channel=0
					-10, -20, -13, -26, -17, -3, 1, 8, -2,
					-- layer=2 filter=200 channel=1
					-32, 2, -16, 10, 0, 8, 3, 9, -3,
					-- layer=2 filter=200 channel=2
					6, -1, -11, 0, 4, 11, 11, -5, 12,
					-- layer=2 filter=200 channel=3
					-5, -47, -35, -27, -24, -16, 31, 32, 4,
					-- layer=2 filter=200 channel=4
					-31, -10, 20, 10, 4, -25, -24, 20, 14,
					-- layer=2 filter=200 channel=5
					-36, -25, -25, -24, -18, -36, 2, -2, 11,
					-- layer=2 filter=200 channel=6
					29, 42, -4, 3, 54, 46, -7, 5, 10,
					-- layer=2 filter=200 channel=7
					25, -27, 8, 21, -22, -13, -38, -1, -8,
					-- layer=2 filter=200 channel=8
					2, 8, 5, 3, -7, 7, 8, 0, 8,
					-- layer=2 filter=200 channel=9
					-1, 0, 0, -33, -26, -34, -9, -6, 0,
					-- layer=2 filter=200 channel=10
					0, -16, -8, -37, -24, -31, -9, -19, 0,
					-- layer=2 filter=200 channel=11
					-8, -18, -36, 0, -26, -10, -20, -18, -2,
					-- layer=2 filter=200 channel=12
					8, 14, 5, -31, -13, -25, 5, 25, -17,
					-- layer=2 filter=200 channel=13
					-13, 5, 6, 10, 10, -1, -6, -7, 3,
					-- layer=2 filter=200 channel=14
					-1, 7, 9, 1, -9, -34, 10, 16, 0,
					-- layer=2 filter=200 channel=15
					-16, -25, -7, 3, -40, -18, -54, 10, -50,
					-- layer=2 filter=200 channel=16
					-47, -25, 9, -14, -13, -7, 1, 5, 20,
					-- layer=2 filter=200 channel=17
					7, -6, 1, -4, 9, -2, 0, 4, -4,
					-- layer=2 filter=200 channel=18
					32, 17, 8, 42, -17, 24, 34, 17, 34,
					-- layer=2 filter=200 channel=19
					-39, 20, -30, -10, -15, 26, 7, 34, 8,
					-- layer=2 filter=200 channel=20
					-7, -1, 5, -5, 7, 8, -3, -8, 4,
					-- layer=2 filter=200 channel=21
					-20, 13, 7, -15, 11, -5, -12, 12, 12,
					-- layer=2 filter=200 channel=22
					3, -11, -7, 5, 3, -1, 10, -9, 5,
					-- layer=2 filter=200 channel=23
					-10, -4, 11, -30, -21, -18, -30, -27, -34,
					-- layer=2 filter=200 channel=24
					23, -44, -1, 18, -38, -11, 16, -6, -9,
					-- layer=2 filter=200 channel=25
					-12, -77, -35, -15, -70, -3, -31, -13, -14,
					-- layer=2 filter=200 channel=26
					-5, -6, -2, 3, 4, -9, 5, -10, -8,
					-- layer=2 filter=200 channel=27
					-44, -63, -71, -8, 5, -2, 5, 38, 8,
					-- layer=2 filter=200 channel=28
					-1, -16, 24, 14, -5, -18, 6, 19, 2,
					-- layer=2 filter=200 channel=29
					9, -4, 2, 1, -9, -8, 1, 2, -8,
					-- layer=2 filter=200 channel=30
					-22, -34, 11, 5, 21, -6, 10, -11, 48,
					-- layer=2 filter=200 channel=31
					32, 51, 4, 62, -26, 56, -51, -41, -49,
					-- layer=2 filter=200 channel=32
					-8, -3, 1, 3, 1, -7, -2, -4, 0,
					-- layer=2 filter=200 channel=33
					-32, 4, 26, 26, 20, 12, 0, 36, -8,
					-- layer=2 filter=200 channel=34
					9, -15, 36, 47, 4, 41, 21, -6, -5,
					-- layer=2 filter=200 channel=35
					-14, -36, -24, 0, -29, -5, 39, 21, 18,
					-- layer=2 filter=200 channel=36
					4, 4, -1, -10, 6, 0, 8, 0, 3,
					-- layer=2 filter=200 channel=37
					-24, -16, -54, -9, -5, -7, -20, -3, -8,
					-- layer=2 filter=200 channel=38
					-39, -6, -23, -8, 22, 9, 31, 40, 21,
					-- layer=2 filter=200 channel=39
					-23, 17, 50, -13, 7, -16, -8, -35, 11,
					-- layer=2 filter=200 channel=40
					-1, -53, 0, 15, -24, -29, -18, -5, -53,
					-- layer=2 filter=200 channel=41
					7, 0, 10, -2, -4, 7, -10, -6, 4,
					-- layer=2 filter=200 channel=42
					-10, 13, 5, -16, 8, -13, -51, 5, -29,
					-- layer=2 filter=200 channel=43
					-39, -76, -70, -12, -44, -19, 34, -14, 3,
					-- layer=2 filter=200 channel=44
					5, -4, -6, -4, 1, 2, -3, 7, 8,
					-- layer=2 filter=200 channel=45
					2, -51, -42, 26, 5, -13, 3, 46, 16,
					-- layer=2 filter=200 channel=46
					-48, 16, 0, -14, 15, 7, 0, -6, 0,
					-- layer=2 filter=200 channel=47
					-5, -26, 15, 10, -26, -20, 22, 50, 18,
					-- layer=2 filter=200 channel=48
					5, 3, 5, 0, -2, 6, 6, 3, 1,
					-- layer=2 filter=200 channel=49
					23, -7, -18, 30, -5, -24, -38, -3, -7,
					-- layer=2 filter=200 channel=50
					10, 11, -11, 0, 25, 15, 2, -5, 3,
					-- layer=2 filter=200 channel=51
					-30, -42, -38, -3, 0, -3, -27, -3, -2,
					-- layer=2 filter=200 channel=52
					-16, 19, 22, 26, 52, 18, -25, 23, 1,
					-- layer=2 filter=200 channel=53
					15, -48, -64, 37, -48, -10, -16, 2, -2,
					-- layer=2 filter=200 channel=54
					-3, 25, 15, -23, -19, -8, -9, 14, 8,
					-- layer=2 filter=200 channel=55
					13, 0, 8, 11, -4, -3, 8, 0, 7,
					-- layer=2 filter=200 channel=56
					-19, -31, -43, 1, -30, -36, -29, -25, -8,
					-- layer=2 filter=200 channel=57
					-10, 0, -2, 1, -1, 8, -1, 5, 2,
					-- layer=2 filter=200 channel=58
					-29, 20, 20, 0, -9, 11, 14, 35, 7,
					-- layer=2 filter=200 channel=59
					-23, -39, 0, -17, -2, 53, 23, 29, 14,
					-- layer=2 filter=200 channel=60
					-12, -16, -1, -10, 4, 36, 15, 0, 30,
					-- layer=2 filter=200 channel=61
					44, -32, -10, -17, -9, 6, 0, -29, 10,
					-- layer=2 filter=200 channel=62
					19, 30, -9, 23, 9, 6, -33, -18, -11,
					-- layer=2 filter=200 channel=63
					1, 13, 21, -16, -14, 14, -12, -12, -3,
					-- layer=2 filter=200 channel=64
					17, 10, 18, 12, 17, 26, -28, -22, -9,
					-- layer=2 filter=200 channel=65
					21, 43, -36, 1, 23, 30, -16, -8, 1,
					-- layer=2 filter=200 channel=66
					-4, -15, -16, -10, 40, -29, -32, -32, 10,
					-- layer=2 filter=200 channel=67
					-50, 6, 24, -44, -29, -37, -29, 0, -20,
					-- layer=2 filter=200 channel=68
					3, 2, -8, 0, -7, -1, 7, 8, 5,
					-- layer=2 filter=200 channel=69
					5, -11, 8, 6, 18, -1, -24, -16, 9,
					-- layer=2 filter=200 channel=70
					13, -13, 13, -17, -24, -9, 13, 12, 3,
					-- layer=2 filter=200 channel=71
					-19, -57, -70, -3, 0, -21, 0, 16, 0,
					-- layer=2 filter=200 channel=72
					48, 60, 74, 9, -60, 14, -14, 33, -18,
					-- layer=2 filter=200 channel=73
					4, -15, -23, 21, -25, 13, 16, -26, -2,
					-- layer=2 filter=200 channel=74
					-4, 16, 23, -7, -4, 11, 9, 42, 3,
					-- layer=2 filter=200 channel=75
					48, -17, 54, -42, -26, 4, 68, 86, 15,
					-- layer=2 filter=200 channel=76
					-8, 20, -50, 14, -29, 0, -20, -42, 5,
					-- layer=2 filter=200 channel=77
					-4, 1, 10, 4, -5, 1, 5, 10, 9,
					-- layer=2 filter=200 channel=78
					15, -21, -43, 8, -16, -12, 5, -38, 9,
					-- layer=2 filter=200 channel=79
					5, 6, 2, -5, 11, 5, 7, 9, -4,
					-- layer=2 filter=200 channel=80
					-51, -23, -2, -22, 3, -2, -5, 15, 0,
					-- layer=2 filter=200 channel=81
					-14, -1, -15, 0, 5, -2, 5, 0, -3,
					-- layer=2 filter=200 channel=82
					-3, 3, -3, 1, -2, 10, -1, 6, 8,
					-- layer=2 filter=200 channel=83
					-4, -41, 4, -51, -31, 2, 15, 11, -9,
					-- layer=2 filter=200 channel=84
					3, 6, 1, -5, 10, -2, 8, 6, 9,
					-- layer=2 filter=200 channel=85
					8, -12, 5, -3, 5, -3, -5, 0, -4,
					-- layer=2 filter=200 channel=86
					3, -3, -6, 16, 0, 1, 5, -5, -9,
					-- layer=2 filter=200 channel=87
					-20, -24, -17, 50, -17, 26, -38, 37, 7,
					-- layer=2 filter=200 channel=88
					9, 2, 25, -16, 14, -20, -6, 4, -13,
					-- layer=2 filter=200 channel=89
					-9, 17, 12, -36, -37, -17, 0, 29, -17,
					-- layer=2 filter=200 channel=90
					1, -9, 7, -9, 7, -9, 7, 4, 7,
					-- layer=2 filter=200 channel=91
					-15, 0, -7, -64, -18, 1, 3, 11, 23,
					-- layer=2 filter=200 channel=92
					-5, 33, 1, -17, -50, -14, 1, 2, -12,
					-- layer=2 filter=200 channel=93
					-46, 30, -30, -8, 23, 40, -4, -39, -18,
					-- layer=2 filter=200 channel=94
					-7, -22, -11, 4, 17, 4, 11, 17, 2,
					-- layer=2 filter=200 channel=95
					5, -20, 15, -20, -8, -9, 8, -9, -1,
					-- layer=2 filter=200 channel=96
					-16, 71, 15, 16, 35, 65, -7, 30, 37,
					-- layer=2 filter=200 channel=97
					7, -35, -10, -14, -8, -36, 13, 9, 11,
					-- layer=2 filter=200 channel=98
					9, -16, 10, 1, -44, -38, 6, 20, 4,
					-- layer=2 filter=200 channel=99
					33, 6, -22, 0, 38, 0, 8, 1, 11,
					-- layer=2 filter=200 channel=100
					-36, -41, -14, -47, -2, 7, 10, 49, 11,
					-- layer=2 filter=200 channel=101
					-49, -88, -9, -29, -36, -21, 17, -8, -45,
					-- layer=2 filter=200 channel=102
					26, 49, -7, 40, 63, 25, -16, 29, 15,
					-- layer=2 filter=200 channel=103
					42, 49, -8, 9, -18, 34, 31, -2, 24,
					-- layer=2 filter=200 channel=104
					0, -6, -16, 37, -13, -24, -20, 22, 0,
					-- layer=2 filter=200 channel=105
					-4, 15, 40, 18, -44, 37, -6, -13, 28,
					-- layer=2 filter=200 channel=106
					-36, -48, -5, -40, -18, -11, -28, -14, -4,
					-- layer=2 filter=200 channel=107
					2, 16, 13, 15, -31, 2, 1, -14, 11,
					-- layer=2 filter=200 channel=108
					-5, -11, -39, -12, -7, -5, -2, 3, 6,
					-- layer=2 filter=200 channel=109
					-2, 0, 12, 12, -18, -29, 2, -2, 16,
					-- layer=2 filter=200 channel=110
					-5, 0, 17, -3, -12, -16, -19, 9, -13,
					-- layer=2 filter=200 channel=111
					0, -10, 10, 2, 0, -7, 4, -2, -9,
					-- layer=2 filter=200 channel=112
					-4, -70, -8, -20, -35, 1, -29, -62, 1,
					-- layer=2 filter=200 channel=113
					-3, -22, 20, 15, 19, 12, 37, -20, 58,
					-- layer=2 filter=200 channel=114
					5, 7, 11, 9, -1, 0, 6, -3, -1,
					-- layer=2 filter=200 channel=115
					-6, -9, 9, -1, 1, -8, -4, 10, 9,
					-- layer=2 filter=200 channel=116
					-15, -11, 7, 32, -16, 33, -33, 19, 16,
					-- layer=2 filter=200 channel=117
					-28, -23, 27, 39, -32, 0, -14, 29, -10,
					-- layer=2 filter=200 channel=118
					-25, -27, -68, -19, -27, -27, 0, -25, 8,
					-- layer=2 filter=200 channel=119
					13, 7, -15, 12, -4, 1, 11, 2, 14,
					-- layer=2 filter=200 channel=120
					0, -1, 2, -6, 5, -7, -2, -6, 5,
					-- layer=2 filter=200 channel=121
					11, -10, 8, -6, -9, 1, 8, 0, -11,
					-- layer=2 filter=200 channel=122
					-11, 0, 4, 0, 4, 0, 17, -2, -3,
					-- layer=2 filter=200 channel=123
					-18, 20, 28, 6, -10, 38, 5, 29, -7,
					-- layer=2 filter=200 channel=124
					-31, 2, -15, 19, 6, 15, -22, -14, 34,
					-- layer=2 filter=200 channel=125
					7, -5, 3, -4, 6, 9, -5, -7, -2,
					-- layer=2 filter=200 channel=126
					-6, 1, -10, 60, -20, 31, 18, 26, 4,
					-- layer=2 filter=200 channel=127
					7, 9, 41, 12, 20, 24, 23, 11, 23,
					-- layer=2 filter=201 channel=0
					-27, -3, 20, -32, 2, -3, -4, 0, -4,
					-- layer=2 filter=201 channel=1
					-13, -3, -12, -11, 0, 4, 38, -9, 6,
					-- layer=2 filter=201 channel=2
					9, -6, 4, 5, -9, -1, -4, 5, 4,
					-- layer=2 filter=201 channel=3
					16, 17, -27, 0, 30, 25, 24, -9, -2,
					-- layer=2 filter=201 channel=4
					15, -9, 27, 34, 8, -24, 9, -4, -16,
					-- layer=2 filter=201 channel=5
					-41, -28, -7, 9, 5, 17, 0, 18, 4,
					-- layer=2 filter=201 channel=6
					40, 19, 15, 5, 5, 41, -23, 34, 40,
					-- layer=2 filter=201 channel=7
					34, 7, 11, 23, 7, 19, 38, 33, 40,
					-- layer=2 filter=201 channel=8
					10, -11, 4, -1, 2, -1, 7, -2, -11,
					-- layer=2 filter=201 channel=9
					27, 35, 34, -29, -16, 12, -15, -41, -32,
					-- layer=2 filter=201 channel=10
					2, 4, -3, -25, 6, -14, 7, -22, -16,
					-- layer=2 filter=201 channel=11
					-39, -27, -24, -13, 12, -9, -11, 0, 13,
					-- layer=2 filter=201 channel=12
					-15, 6, 5, 14, 3, 5, 29, 19, 39,
					-- layer=2 filter=201 channel=13
					-10, 4, 0, 8, -6, 7, 8, 8, 5,
					-- layer=2 filter=201 channel=14
					1, 0, 27, 28, 0, 7, 16, -12, 12,
					-- layer=2 filter=201 channel=15
					-2, -34, -40, -32, 30, -5, -13, 58, 6,
					-- layer=2 filter=201 channel=16
					23, 5, 33, 3, -5, -32, -27, -63, -46,
					-- layer=2 filter=201 channel=17
					4, 5, -2, 2, -9, 6, 5, -4, -7,
					-- layer=2 filter=201 channel=18
					24, -26, -48, -6, -7, -22, 28, 21, 14,
					-- layer=2 filter=201 channel=19
					-36, -47, -23, -8, -24, 0, 32, 5, 17,
					-- layer=2 filter=201 channel=20
					2, -8, 1, 7, -11, -5, 0, -7, -7,
					-- layer=2 filter=201 channel=21
					-11, -5, 2, -6, -9, 0, -19, -11, -21,
					-- layer=2 filter=201 channel=22
					1, -15, -3, 8, 9, -11, -4, -6, -4,
					-- layer=2 filter=201 channel=23
					46, 5, -4, 24, -46, -28, 16, -24, -46,
					-- layer=2 filter=201 channel=24
					21, 6, -1, 9, 39, 8, 8, 14, -20,
					-- layer=2 filter=201 channel=25
					-37, 12, -21, 13, 32, 6, 11, 29, -5,
					-- layer=2 filter=201 channel=26
					9, 0, -6, -4, 2, 0, -1, 8, -1,
					-- layer=2 filter=201 channel=27
					-25, -35, 15, 25, 11, 8, 50, 44, 13,
					-- layer=2 filter=201 channel=28
					4, -26, 3, -36, -3, -44, 34, -37, -17,
					-- layer=2 filter=201 channel=29
					7, 3, -7, -5, -1, 10, -7, -9, -7,
					-- layer=2 filter=201 channel=30
					4, 26, -2, -21, -9, 7, 0, -5, -33,
					-- layer=2 filter=201 channel=31
					-61, -68, -56, -130, -47, -42, -24, -35, -41,
					-- layer=2 filter=201 channel=32
					7, -4, -6, 0, 7, 9, -9, -1, -8,
					-- layer=2 filter=201 channel=33
					17, -10, 0, 43, 35, 11, 12, 29, -11,
					-- layer=2 filter=201 channel=34
					-37, 0, -15, 0, -2, 5, -37, 5, 21,
					-- layer=2 filter=201 channel=35
					-29, -26, -54, -29, -31, -49, 18, -13, -21,
					-- layer=2 filter=201 channel=36
					2, -3, 5, 11, 2, -6, 9, -4, -6,
					-- layer=2 filter=201 channel=37
					-14, -36, -14, -4, 19, 25, 2, 28, 34,
					-- layer=2 filter=201 channel=38
					-60, -24, -1, -14, 0, -7, 0, 42, 8,
					-- layer=2 filter=201 channel=39
					27, 15, 11, 17, -19, 8, 2, -30, -65,
					-- layer=2 filter=201 channel=40
					-3, -1, -21, 3, 36, 11, 43, 13, -5,
					-- layer=2 filter=201 channel=41
					-6, -10, 5, 2, -9, 0, 1, 0, 3,
					-- layer=2 filter=201 channel=42
					23, 16, -3, -31, 10, -33, -6, -52, -30,
					-- layer=2 filter=201 channel=43
					-17, -4, -35, -78, -7, -50, 2, 9, 33,
					-- layer=2 filter=201 channel=44
					-6, -4, 5, 3, -8, -10, 10, -2, -5,
					-- layer=2 filter=201 channel=45
					2, 2, 71, 51, 47, -5, 21, 13, -17,
					-- layer=2 filter=201 channel=46
					9, 21, 12, -23, 21, 19, -35, -30, -40,
					-- layer=2 filter=201 channel=47
					3, -2, 32, 47, 45, -1, -2, -15, 56,
					-- layer=2 filter=201 channel=48
					-10, 0, 6, -4, -6, 8, 1, 4, -5,
					-- layer=2 filter=201 channel=49
					31, -9, -30, -51, -4, -15, 21, 15, -5,
					-- layer=2 filter=201 channel=50
					-14, -15, -1, -3, 27, 17, 24, 10, -4,
					-- layer=2 filter=201 channel=51
					-37, -15, -37, -36, -19, 1, -25, -1, -9,
					-- layer=2 filter=201 channel=52
					-18, -23, -26, 49, -2, 32, 43, 18, 42,
					-- layer=2 filter=201 channel=53
					-3, -25, -26, -6, -12, -34, -7, 32, -20,
					-- layer=2 filter=201 channel=54
					-2, -8, -25, -14, 3, -5, 35, 2, 3,
					-- layer=2 filter=201 channel=55
					-6, 9, 0, 9, -1, 2, 0, 1, 1,
					-- layer=2 filter=201 channel=56
					-6, -34, -3, 0, 22, 15, 6, -3, 33,
					-- layer=2 filter=201 channel=57
					0, -5, -12, -2, -10, -2, 7, -9, -7,
					-- layer=2 filter=201 channel=58
					-41, -5, -28, 45, -7, 0, 30, 12, 8,
					-- layer=2 filter=201 channel=59
					-52, 3, -41, 11, 49, 0, 22, 23, 26,
					-- layer=2 filter=201 channel=60
					-51, -8, -8, -24, 6, 10, 26, 22, 14,
					-- layer=2 filter=201 channel=61
					-7, 13, -15, -40, -54, 23, -34, 4, 2,
					-- layer=2 filter=201 channel=62
					-3, -32, -1, -18, 0, 6, -7, 19, 12,
					-- layer=2 filter=201 channel=63
					16, 19, 3, 4, -30, -18, 7, -17, -33,
					-- layer=2 filter=201 channel=64
					27, 39, 31, 23, -7, -9, 0, -15, -66,
					-- layer=2 filter=201 channel=65
					-4, -5, -37, -35, -35, 22, -53, 4, 44,
					-- layer=2 filter=201 channel=66
					27, 29, 21, 3, 29, 2, 4, 30, 44,
					-- layer=2 filter=201 channel=67
					21, 8, 38, -50, -22, 24, -21, -9, -19,
					-- layer=2 filter=201 channel=68
					6, -3, -4, -7, 0, 3, 7, -1, -2,
					-- layer=2 filter=201 channel=69
					37, 18, 36, -4, -6, 2, 17, -32, -33,
					-- layer=2 filter=201 channel=70
					-23, -19, -40, -1, 0, -18, 15, -17, 9,
					-- layer=2 filter=201 channel=71
					-36, -37, 9, 4, -16, -14, 38, 13, 0,
					-- layer=2 filter=201 channel=72
					28, -16, -1, 2, 10, 18, 1, -21, 18,
					-- layer=2 filter=201 channel=73
					-88, -51, -29, -62, -43, -21, -38, -30, -17,
					-- layer=2 filter=201 channel=74
					-4, -4, 18, -37, 0, 14, -12, -27, -19,
					-- layer=2 filter=201 channel=75
					20, 26, 16, 21, 37, 33, 14, 9, 16,
					-- layer=2 filter=201 channel=76
					-36, -11, -49, 34, -5, -34, -37, 4, -45,
					-- layer=2 filter=201 channel=77
					6, 3, -6, -6, -9, -3, 4, -8, 3,
					-- layer=2 filter=201 channel=78
					-28, 6, -41, -30, 18, 8, -1, -1, 2,
					-- layer=2 filter=201 channel=79
					-5, 8, -1, -4, 3, 0, -9, 2, 2,
					-- layer=2 filter=201 channel=80
					10, 9, 34, 5, -6, 24, -10, -26, 17,
					-- layer=2 filter=201 channel=81
					-10, 2, -5, 0, -6, 2, 12, 5, 15,
					-- layer=2 filter=201 channel=82
					0, 3, 7, 0, -2, 0, 10, 5, -2,
					-- layer=2 filter=201 channel=83
					-4, 6, 9, 0, -53, 10, 36, -28, -26,
					-- layer=2 filter=201 channel=84
					2, 0, 5, 4, 4, -7, -2, -5, 5,
					-- layer=2 filter=201 channel=85
					5, 0, 0, 14, 13, -6, 1, 2, 1,
					-- layer=2 filter=201 channel=86
					1, -18, 6, 25, 5, 10, 5, 11, -12,
					-- layer=2 filter=201 channel=87
					0, -5, -23, 7, -7, -33, -5, 47, -4,
					-- layer=2 filter=201 channel=88
					46, 9, 19, 8, -29, -4, -19, -23, -32,
					-- layer=2 filter=201 channel=89
					-50, -19, -10, 9, 13, 35, 12, 12, 30,
					-- layer=2 filter=201 channel=90
					5, -9, -9, 1, 8, -8, -5, -9, 8,
					-- layer=2 filter=201 channel=91
					-39, 3, -16, -11, 32, 26, 22, 24, 39,
					-- layer=2 filter=201 channel=92
					-23, 3, 7, 0, 6, 24, 26, 6, 35,
					-- layer=2 filter=201 channel=93
					-37, -24, -5, 30, 30, 71, 3, 17, 56,
					-- layer=2 filter=201 channel=94
					0, -35, -8, -54, -6, 12, 7, 13, -2,
					-- layer=2 filter=201 channel=95
					13, -4, 5, 3, 2, 10, -5, 0, 6,
					-- layer=2 filter=201 channel=96
					5, -24, 8, 41, 8, 22, -36, 50, 25,
					-- layer=2 filter=201 channel=97
					5, 6, 23, -2, -8, 31, -10, -8, -24,
					-- layer=2 filter=201 channel=98
					-1, -16, 8, -5, 2, 7, 24, -25, 35,
					-- layer=2 filter=201 channel=99
					-36, -42, -29, 18, -31, 4, -10, 0, 32,
					-- layer=2 filter=201 channel=100
					-17, -17, -31, -26, 5, -12, 6, 30, 16,
					-- layer=2 filter=201 channel=101
					-19, -5, -47, 36, 4, -39, 1, -24, -26,
					-- layer=2 filter=201 channel=102
					-4, -8, -49, -12, -8, 0, -29, 18, 25,
					-- layer=2 filter=201 channel=103
					35, -1, 2, 29, 40, 59, 17, -29, 20,
					-- layer=2 filter=201 channel=104
					3, -73, -41, -23, -9, 0, 18, 5, -6,
					-- layer=2 filter=201 channel=105
					28, -24, 6, -8, -31, -42, -1, -51, -27,
					-- layer=2 filter=201 channel=106
					-33, 16, -13, 4, 39, -12, -3, -10, -11,
					-- layer=2 filter=201 channel=107
					-1, 3, 7, -7, 25, 18, -33, -11, 36,
					-- layer=2 filter=201 channel=108
					-22, -61, -5, 11, -26, 14, 16, 27, 9,
					-- layer=2 filter=201 channel=109
					11, -2, 11, -4, -7, 5, 2, 3, 2,
					-- layer=2 filter=201 channel=110
					31, 7, 5, 23, -6, -2, -3, -33, -25,
					-- layer=2 filter=201 channel=111
					3, 9, 6, -2, 4, -2, 3, -10, 10,
					-- layer=2 filter=201 channel=112
					-19, -8, -14, -67, 15, 19, 8, -1, 0,
					-- layer=2 filter=201 channel=113
					4, 32, -5, -14, -29, 11, 25, -32, -8,
					-- layer=2 filter=201 channel=114
					1, -7, 3, -4, -6, -13, 8, 2, 0,
					-- layer=2 filter=201 channel=115
					-4, 9, -4, 1, -9, 2, -5, 8, 0,
					-- layer=2 filter=201 channel=116
					16, -21, -23, 40, 7, -2, 3, 34, 7,
					-- layer=2 filter=201 channel=117
					-11, -33, -8, 14, -28, -30, 20, -4, 17,
					-- layer=2 filter=201 channel=118
					26, 14, -14, -8, 7, -15, -29, 17, 15,
					-- layer=2 filter=201 channel=119
					23, 7, -42, 15, 2, -32, 34, -24, -32,
					-- layer=2 filter=201 channel=120
					-10, -10, 7, -4, 6, 10, 7, -4, -9,
					-- layer=2 filter=201 channel=121
					9, -10, -5, 12, -1, -1, -3, 0, 0,
					-- layer=2 filter=201 channel=122
					-14, 2, -7, 7, 0, -6, -14, -10, 10,
					-- layer=2 filter=201 channel=123
					45, 4, 2, 15, -32, -8, -6, 15, 38,
					-- layer=2 filter=201 channel=124
					-47, 8, -29, 10, 13, -6, -38, 20, -26,
					-- layer=2 filter=201 channel=125
					9, -11, 0, 0, 11, 12, 9, -3, 0,
					-- layer=2 filter=201 channel=126
					13, -18, -2, -14, -15, 4, 11, -51, 16,
					-- layer=2 filter=201 channel=127
					-2, 11, 11, 16, -31, -9, 5, -22, -18,
					-- layer=2 filter=202 channel=0
					-10, 8, 3, 2, 6, 13, 23, 13, 3,
					-- layer=2 filter=202 channel=1
					4, 4, -7, 22, 22, -2, -4, -2, 15,
					-- layer=2 filter=202 channel=2
					-4, -2, -11, 0, 0, -3, 7, 8, 6,
					-- layer=2 filter=202 channel=3
					-23, -30, 26, 6, -41, 9, 3, -31, -21,
					-- layer=2 filter=202 channel=4
					-54, -2, -32, -49, 0, 5, -33, 30, -2,
					-- layer=2 filter=202 channel=5
					-4, -11, 26, -13, 20, 24, -24, -23, 12,
					-- layer=2 filter=202 channel=6
					16, -4, -27, -8, -5, 38, -47, -39, 37,
					-- layer=2 filter=202 channel=7
					-24, 11, 9, 18, -29, -13, -37, 32, 25,
					-- layer=2 filter=202 channel=8
					-5, 6, -10, -1, -6, -10, 2, -5, 0,
					-- layer=2 filter=202 channel=9
					-3, -11, -11, -19, -10, -20, -8, -7, 1,
					-- layer=2 filter=202 channel=10
					-2, -10, 28, 7, -5, -6, 28, 21, 31,
					-- layer=2 filter=202 channel=11
					2, -4, 5, 0, 2, 15, -19, -4, -7,
					-- layer=2 filter=202 channel=12
					-6, 11, -1, 3, -15, -13, -9, -1, 24,
					-- layer=2 filter=202 channel=13
					2, 0, 4, -5, 0, -2, -3, 7, -4,
					-- layer=2 filter=202 channel=14
					-14, 4, -3, 3, 12, -29, -10, 2, 9,
					-- layer=2 filter=202 channel=15
					-20, -26, -2, -14, -43, -23, -4, -33, 10,
					-- layer=2 filter=202 channel=16
					-29, -42, -20, -9, -24, -43, -20, -22, -14,
					-- layer=2 filter=202 channel=17
					0, 2, -3, 3, -4, 7, 3, 8, 0,
					-- layer=2 filter=202 channel=18
					-17, -15, -17, -30, 19, -26, -26, -2, -8,
					-- layer=2 filter=202 channel=19
					0, -21, -4, 11, -2, 4, 0, 7, 11,
					-- layer=2 filter=202 channel=20
					0, -11, -6, -10, 6, -6, -3, 0, 0,
					-- layer=2 filter=202 channel=21
					10, 1, -12, -11, -6, -2, 0, 2, -5,
					-- layer=2 filter=202 channel=22
					-1, -6, 8, -10, 7, -7, -3, -1, -7,
					-- layer=2 filter=202 channel=23
					-41, -19, -15, -18, -37, -17, -30, 0, 0,
					-- layer=2 filter=202 channel=24
					-8, 11, 17, -5, -33, -21, -1, -19, -24,
					-- layer=2 filter=202 channel=25
					-18, -15, -10, 0, -26, -12, -14, -29, -16,
					-- layer=2 filter=202 channel=26
					-8, 9, 0, 10, 3, 7, -5, 1, -1,
					-- layer=2 filter=202 channel=27
					10, 0, -1, 6, -6, -2, 6, -20, -7,
					-- layer=2 filter=202 channel=28
					-47, -31, 15, -62, -32, -21, 8, 8, 0,
					-- layer=2 filter=202 channel=29
					-4, 8, -5, -1, -12, -1, 0, -8, 1,
					-- layer=2 filter=202 channel=30
					31, -35, -10, 27, -13, -12, 19, -3, -21,
					-- layer=2 filter=202 channel=31
					-32, -14, -38, -31, 12, 3, -17, -23, -7,
					-- layer=2 filter=202 channel=32
					-9, 6, -7, -9, 8, 0, -7, -9, 7,
					-- layer=2 filter=202 channel=33
					-42, 7, 1, 4, -31, 9, 0, -11, 0,
					-- layer=2 filter=202 channel=34
					12, -25, 26, 18, 19, -15, -21, -16, -2,
					-- layer=2 filter=202 channel=35
					-25, -34, 23, -64, -18, -17, 13, 17, -5,
					-- layer=2 filter=202 channel=36
					-3, -7, 6, -4, 1, -11, -10, -4, -2,
					-- layer=2 filter=202 channel=37
					0, -10, 0, 7, 11, 15, -17, -16, 10,
					-- layer=2 filter=202 channel=38
					23, 7, 0, 25, -25, -13, -12, -23, 3,
					-- layer=2 filter=202 channel=39
					-13, -24, -26, -12, -34, -24, -40, -31, -22,
					-- layer=2 filter=202 channel=40
					-35, -1, 2, -41, -12, 22, 17, -35, -1,
					-- layer=2 filter=202 channel=41
					6, -10, 1, -6, -7, -6, -4, 2, -3,
					-- layer=2 filter=202 channel=42
					-30, -18, -22, -16, -14, -32, -49, -21, 13,
					-- layer=2 filter=202 channel=43
					-14, 0, -14, -29, -17, -37, -25, -20, -45,
					-- layer=2 filter=202 channel=44
					0, 1, 9, 2, -5, 0, 10, -4, -9,
					-- layer=2 filter=202 channel=45
					4, -21, -47, 4, 1, 8, 0, 0, 0,
					-- layer=2 filter=202 channel=46
					10, -54, -12, 7, 6, 14, 20, 2, -4,
					-- layer=2 filter=202 channel=47
					-71, -14, -37, -43, -17, -25, 0, 30, 14,
					-- layer=2 filter=202 channel=48
					-3, 1, -10, 0, 0, 1, -10, -3, 4,
					-- layer=2 filter=202 channel=49
					-10, -33, -26, -5, 35, -14, -31, -13, 10,
					-- layer=2 filter=202 channel=50
					-2, 6, 11, 9, 0, -4, 17, 14, 1,
					-- layer=2 filter=202 channel=51
					-3, 16, 1, 5, 20, 0, -3, -9, 12,
					-- layer=2 filter=202 channel=52
					3, 19, -26, 3, 8, -28, 27, 20, 27,
					-- layer=2 filter=202 channel=53
					4, -66, -31, -7, 9, 3, 6, -5, 54,
					-- layer=2 filter=202 channel=54
					-42, -35, 7, -17, -9, 21, 2, 16, 10,
					-- layer=2 filter=202 channel=55
					-2, -3, 7, 0, -6, 10, 4, -7, -1,
					-- layer=2 filter=202 channel=56
					-13, -16, -1, -40, -28, -2, -37, -3, -19,
					-- layer=2 filter=202 channel=57
					-4, 3, 12, -5, 0, -3, 8, 6, 11,
					-- layer=2 filter=202 channel=58
					-19, 7, 5, 19, -25, -4, -16, -14, -11,
					-- layer=2 filter=202 channel=59
					-9, 28, -10, 11, -18, 6, 0, 0, -22,
					-- layer=2 filter=202 channel=60
					7, -2, -8, 9, -17, -13, -18, 19, -5,
					-- layer=2 filter=202 channel=61
					-10, 2, 1, 17, 11, -11, -29, 27, -1,
					-- layer=2 filter=202 channel=62
					5, -2, -31, 9, 5, 26, -56, 5, 7,
					-- layer=2 filter=202 channel=63
					-4, -5, -39, -19, 2, -48, -54, 30, -51,
					-- layer=2 filter=202 channel=64
					31, -11, -39, 16, -2, -32, -13, -51, -4,
					-- layer=2 filter=202 channel=65
					23, 9, -19, 32, -19, 7, -23, -6, 20,
					-- layer=2 filter=202 channel=66
					17, -25, -65, 10, -55, 4, 13, -28, 0,
					-- layer=2 filter=202 channel=67
					27, -38, -12, 7, -37, -13, -9, -19, 19,
					-- layer=2 filter=202 channel=68
					-10, 7, 2, 8, 7, -4, 2, -2, 3,
					-- layer=2 filter=202 channel=69
					-3, -20, -45, -1, -42, -18, -63, -60, -15,
					-- layer=2 filter=202 channel=70
					-47, -66, 29, -60, 4, 7, 21, 12, 2,
					-- layer=2 filter=202 channel=71
					0, -14, 16, -14, -19, -3, -10, -27, -7,
					-- layer=2 filter=202 channel=72
					8, 33, 4, 9, -29, -9, -32, 13, 0,
					-- layer=2 filter=202 channel=73
					-20, -40, 3, 4, 8, -20, -7, 12, 12,
					-- layer=2 filter=202 channel=74
					22, -8, -8, 7, -21, -16, -11, -13, 15,
					-- layer=2 filter=202 channel=75
					-23, -4, 1, -20, -35, -5, -19, 4, -13,
					-- layer=2 filter=202 channel=76
					-20, -19, -37, -23, 19, 44, 13, 9, 38,
					-- layer=2 filter=202 channel=77
					5, 0, -9, -12, 0, -10, 4, 4, 0,
					-- layer=2 filter=202 channel=78
					1, -1, -8, 4, -8, 1, -28, 13, 1,
					-- layer=2 filter=202 channel=79
					-9, -9, 7, 1, 8, -4, 5, -8, -5,
					-- layer=2 filter=202 channel=80
					-16, -38, -4, -36, -48, 0, -16, -16, -33,
					-- layer=2 filter=202 channel=81
					0, 5, 1, 2, 8, -5, 5, -2, -11,
					-- layer=2 filter=202 channel=82
					6, -8, 3, 0, 7, 6, 0, 7, -9,
					-- layer=2 filter=202 channel=83
					-25, -31, -12, -4, -48, 13, 7, 9, 3,
					-- layer=2 filter=202 channel=84
					-1, 9, 6, -6, 5, -1, 5, 0, -10,
					-- layer=2 filter=202 channel=85
					-5, -11, 4, 7, 1, 0, 3, -7, 6,
					-- layer=2 filter=202 channel=86
					2, 8, -1, 0, 0, -4, -10, -4, -1,
					-- layer=2 filter=202 channel=87
					-29, -10, -42, -37, -2, -26, -2, 29, 18,
					-- layer=2 filter=202 channel=88
					0, -13, -47, 0, -18, -35, -39, -41, -1,
					-- layer=2 filter=202 channel=89
					-8, 22, -24, 2, 5, 30, -6, 18, 15,
					-- layer=2 filter=202 channel=90
					8, -3, 4, 2, 3, 10, 7, -4, -3,
					-- layer=2 filter=202 channel=91
					-13, 29, -11, -12, -28, -11, -8, -2, 6,
					-- layer=2 filter=202 channel=92
					0, 15, -26, 2, 6, 8, -19, 3, 24,
					-- layer=2 filter=202 channel=93
					13, -21, -46, 15, -12, -12, -54, -7, 31,
					-- layer=2 filter=202 channel=94
					14, -33, -45, 31, -19, 5, -34, 32, 18,
					-- layer=2 filter=202 channel=95
					2, 0, -10, -4, 6, -7, 2, 4, -8,
					-- layer=2 filter=202 channel=96
					-26, -16, 14, -46, 48, 25, 11, 38, 4,
					-- layer=2 filter=202 channel=97
					-6, -15, -29, -27, -9, -9, -40, 26, -20,
					-- layer=2 filter=202 channel=98
					-75, -14, -24, -16, -28, 0, 2, 40, 1,
					-- layer=2 filter=202 channel=99
					-20, 9, -16, 28, 24, 15, 3, 29, 16,
					-- layer=2 filter=202 channel=100
					35, -23, 6, -10, -22, -33, -26, -3, -19,
					-- layer=2 filter=202 channel=101
					-24, -6, 16, -44, -5, 4, -26, -25, -8,
					-- layer=2 filter=202 channel=102
					-35, -11, -15, -5, 56, -26, 4, 16, -8,
					-- layer=2 filter=202 channel=103
					-24, 27, 5, -3, 28, 3, 46, 36, 45,
					-- layer=2 filter=202 channel=104
					-8, -27, -17, -14, -4, 36, -1, 32, 11,
					-- layer=2 filter=202 channel=105
					-25, 18, -60, 0, -5, -18, -9, 20, -7,
					-- layer=2 filter=202 channel=106
					-23, 5, -20, -44, -49, -16, -16, -32, -11,
					-- layer=2 filter=202 channel=107
					-10, -15, -6, 24, 24, -27, 3, 10, 4,
					-- layer=2 filter=202 channel=108
					9, -7, -10, -1, 22, -24, -8, 0, 4,
					-- layer=2 filter=202 channel=109
					1, -2, 0, -11, 1, -11, 0, 8, -11,
					-- layer=2 filter=202 channel=110
					8, -24, 4, -9, -7, -32, -13, -27, -39,
					-- layer=2 filter=202 channel=111
					6, 1, 3, 7, 4, -3, -11, -1, 3,
					-- layer=2 filter=202 channel=112
					-9, 4, -19, -7, -15, -13, -2, 6, -3,
					-- layer=2 filter=202 channel=113
					15, -8, -15, -2, -29, -5, -7, 2, -46,
					-- layer=2 filter=202 channel=114
					0, 5, -6, 1, -4, -10, -8, -1, 5,
					-- layer=2 filter=202 channel=115
					6, 4, 7, -6, -14, 0, 2, 8, 1,
					-- layer=2 filter=202 channel=116
					-22, -32, -27, -25, 22, -38, -3, 9, 22,
					-- layer=2 filter=202 channel=117
					-44, -32, 10, 4, -23, -23, -34, 29, 27,
					-- layer=2 filter=202 channel=118
					-30, -14, 5, 5, -14, -1, -6, 2, -11,
					-- layer=2 filter=202 channel=119
					-29, -27, -29, -26, -8, -48, -19, -17, -39,
					-- layer=2 filter=202 channel=120
					-4, 4, 6, 6, 2, -2, 0, 6, -10,
					-- layer=2 filter=202 channel=121
					-4, 2, -8, 4, -10, 6, 2, 8, -2,
					-- layer=2 filter=202 channel=122
					2, -8, 7, 4, 4, -3, 0, -5, -1,
					-- layer=2 filter=202 channel=123
					-33, 34, -14, 7, -42, 4, 1, 40, 6,
					-- layer=2 filter=202 channel=124
					-30, 14, -19, -17, -31, -1, -19, -21, -6,
					-- layer=2 filter=202 channel=125
					8, 4, -5, -5, -3, 0, 6, 5, 0,
					-- layer=2 filter=202 channel=126
					9, -7, 8, -10, 28, -31, -23, 11, -12,
					-- layer=2 filter=202 channel=127
					-6, -22, -10, -21, 2, -22, -27, -18, -22,
					-- layer=2 filter=203 channel=0
					2, -2, -5, -15, -14, -8, -10, -2, 6,
					-- layer=2 filter=203 channel=1
					-14, -13, -11, -7, 6, 1, -1, 4, -8,
					-- layer=2 filter=203 channel=2
					-2, 3, 5, 3, -3, 0, -9, -5, 11,
					-- layer=2 filter=203 channel=3
					1, -2, -8, -14, -7, 5, 1, -8, -2,
					-- layer=2 filter=203 channel=4
					0, 5, -7, -10, 1, 2, -7, -3, -7,
					-- layer=2 filter=203 channel=5
					-8, 2, -6, -7, -6, 0, 0, -4, -3,
					-- layer=2 filter=203 channel=6
					-8, -20, -8, -8, -12, -9, -13, -11, 2,
					-- layer=2 filter=203 channel=7
					0, 7, -8, 3, 9, -7, -10, -7, -3,
					-- layer=2 filter=203 channel=8
					4, 1, -10, 0, 4, 0, 7, 2, -8,
					-- layer=2 filter=203 channel=9
					-10, 0, 0, -11, -7, 0, -12, -8, 6,
					-- layer=2 filter=203 channel=10
					-3, 3, -14, -9, -10, -9, -9, -9, 2,
					-- layer=2 filter=203 channel=11
					-9, 3, -4, 1, -13, -3, 2, -8, 3,
					-- layer=2 filter=203 channel=12
					-11, 5, -6, 2, 4, -15, 0, 2, -10,
					-- layer=2 filter=203 channel=13
					-1, 4, -1, 6, 6, -8, -5, 0, -8,
					-- layer=2 filter=203 channel=14
					0, 3, -11, -7, 2, 4, -1, -12, -10,
					-- layer=2 filter=203 channel=15
					-18, -10, -11, -5, -6, 4, -9, -7, 4,
					-- layer=2 filter=203 channel=16
					-13, 5, -6, -14, -8, -12, -11, -9, -3,
					-- layer=2 filter=203 channel=17
					9, 5, -3, -4, 1, -4, -8, 0, -7,
					-- layer=2 filter=203 channel=18
					8, -6, -12, -9, -4, -18, -16, -1, -6,
					-- layer=2 filter=203 channel=19
					5, 6, -7, 2, 1, -12, -2, -18, -7,
					-- layer=2 filter=203 channel=20
					11, 8, -4, 2, -9, -8, 6, 6, -1,
					-- layer=2 filter=203 channel=21
					9, -1, -8, 1, 3, -7, -6, -8, 7,
					-- layer=2 filter=203 channel=22
					3, 2, 5, 0, -3, 9, -2, -4, -2,
					-- layer=2 filter=203 channel=23
					0, -15, -4, -9, -11, 4, -9, -12, 4,
					-- layer=2 filter=203 channel=24
					2, 5, 0, 0, 0, 8, 0, 0, 2,
					-- layer=2 filter=203 channel=25
					8, 7, 0, -15, 6, -2, 5, 0, 3,
					-- layer=2 filter=203 channel=26
					8, 8, -8, 0, -5, 4, -9, -4, 8,
					-- layer=2 filter=203 channel=27
					5, 2, -14, 1, -6, -15, 1, -9, -11,
					-- layer=2 filter=203 channel=28
					-5, 10, -3, -13, -5, 1, -5, 4, -9,
					-- layer=2 filter=203 channel=29
					-6, 1, -6, 3, 9, -6, 0, -8, 7,
					-- layer=2 filter=203 channel=30
					-14, -6, -8, 4, -7, 6, 0, -7, -13,
					-- layer=2 filter=203 channel=31
					2, -9, 6, 5, -6, -7, 4, -9, 0,
					-- layer=2 filter=203 channel=32
					-4, 1, 6, -11, 4, 5, 9, 9, -11,
					-- layer=2 filter=203 channel=33
					-11, -11, -1, -7, 4, 1, 0, -8, -11,
					-- layer=2 filter=203 channel=34
					-10, -6, -13, -13, -16, -12, -17, -9, -14,
					-- layer=2 filter=203 channel=35
					0, -6, -11, -15, 7, 0, -9, 0, 0,
					-- layer=2 filter=203 channel=36
					-10, 8, -7, 3, -9, -2, -10, 3, -5,
					-- layer=2 filter=203 channel=37
					5, 3, -11, -7, 1, 3, -4, 0, -7,
					-- layer=2 filter=203 channel=38
					-1, -1, -12, 2, -14, -15, 0, -9, -16,
					-- layer=2 filter=203 channel=39
					3, -9, -3, -2, -5, 0, -4, -12, 1,
					-- layer=2 filter=203 channel=40
					-8, -2, 0, -14, 4, -8, -5, -2, 4,
					-- layer=2 filter=203 channel=41
					1, -11, 6, 11, -9, 8, -8, -4, -1,
					-- layer=2 filter=203 channel=42
					1, 4, -10, 4, 4, 10, -4, -16, -6,
					-- layer=2 filter=203 channel=43
					1, 0, -4, 1, -10, -1, -12, -10, -13,
					-- layer=2 filter=203 channel=44
					1, 0, 1, -6, 1, -9, -11, 4, -3,
					-- layer=2 filter=203 channel=45
					-10, -6, -7, -3, -4, 5, -5, -3, -8,
					-- layer=2 filter=203 channel=46
					0, 3, -13, 2, 5, -2, -14, 0, 0,
					-- layer=2 filter=203 channel=47
					-7, -3, -6, -6, 2, -2, 3, -13, -4,
					-- layer=2 filter=203 channel=48
					3, -1, -6, 1, 7, -2, 8, 6, 0,
					-- layer=2 filter=203 channel=49
					-7, -5, -8, -5, -5, -5, -4, -5, -7,
					-- layer=2 filter=203 channel=50
					11, -1, -4, 0, -1, 5, -6, -5, 4,
					-- layer=2 filter=203 channel=51
					-14, 0, -14, 4, 0, -2, 0, -11, 0,
					-- layer=2 filter=203 channel=52
					-5, -13, 3, -10, -14, 2, -17, -1, -14,
					-- layer=2 filter=203 channel=53
					0, -19, 3, 10, -5, 0, 4, -2, 0,
					-- layer=2 filter=203 channel=54
					-7, -18, 3, -23, 4, -4, 1, -10, 8,
					-- layer=2 filter=203 channel=55
					6, 2, -4, -3, -6, -7, -10, 1, 4,
					-- layer=2 filter=203 channel=56
					3, 0, 5, -12, -8, -2, 2, 6, -10,
					-- layer=2 filter=203 channel=57
					7, 11, 0, 0, 5, 9, -4, 6, -1,
					-- layer=2 filter=203 channel=58
					-5, 9, -2, -12, -9, -10, -6, -9, -1,
					-- layer=2 filter=203 channel=59
					-10, -11, -15, 4, -12, -9, -11, -15, 4,
					-- layer=2 filter=203 channel=60
					0, -6, 3, 3, -1, -11, -8, -1, -1,
					-- layer=2 filter=203 channel=61
					-9, 11, 9, -11, -7, 1, 11, -18, 5,
					-- layer=2 filter=203 channel=62
					-14, -7, 5, -10, -3, 0, -3, -6, -9,
					-- layer=2 filter=203 channel=63
					5, 0, -8, -12, 0, 6, -1, -11, -6,
					-- layer=2 filter=203 channel=64
					-5, -10, -7, 7, -10, 7, -14, -13, -14,
					-- layer=2 filter=203 channel=65
					3, -2, 0, -1, -1, -9, -9, -7, 9,
					-- layer=2 filter=203 channel=66
					6, 8, -6, -9, -4, 3, -6, -4, 8,
					-- layer=2 filter=203 channel=67
					-10, -5, -4, -4, -11, -11, -13, 0, -2,
					-- layer=2 filter=203 channel=68
					3, 9, -1, 1, -3, -8, -9, -5, -7,
					-- layer=2 filter=203 channel=69
					4, -7, -1, 4, -8, -12, -18, 5, -7,
					-- layer=2 filter=203 channel=70
					0, -3, -3, -4, -8, -9, -6, -3, -7,
					-- layer=2 filter=203 channel=71
					-8, -9, -6, 2, -2, -11, -10, -1, -2,
					-- layer=2 filter=203 channel=72
					0, 6, 0, 3, 14, 7, 1, -7, -1,
					-- layer=2 filter=203 channel=73
					-3, -2, 0, -13, -2, 1, 12, -15, 8,
					-- layer=2 filter=203 channel=74
					-7, -4, 1, 4, -9, -11, 0, -5, -11,
					-- layer=2 filter=203 channel=75
					4, 11, -7, -10, -7, 9, 5, 4, 3,
					-- layer=2 filter=203 channel=76
					-5, -2, -5, 11, -14, 3, -4, -17, 11,
					-- layer=2 filter=203 channel=77
					6, 7, -7, -9, 3, 4, -11, -5, 8,
					-- layer=2 filter=203 channel=78
					3, -1, -6, -18, 0, -15, -1, 3, -4,
					-- layer=2 filter=203 channel=79
					-7, 8, 8, -1, 0, -7, 11, -5, -3,
					-- layer=2 filter=203 channel=80
					1, 5, -5, -7, -12, 5, 1, -8, -5,
					-- layer=2 filter=203 channel=81
					0, 2, 3, -10, 0, -4, 5, 0, 0,
					-- layer=2 filter=203 channel=82
					8, 2, -8, 0, -6, -6, -6, -6, -2,
					-- layer=2 filter=203 channel=83
					-13, -9, 2, -8, 0, -4, -8, 7, 0,
					-- layer=2 filter=203 channel=84
					-1, -3, 1, 4, -6, -8, 2, -8, 3,
					-- layer=2 filter=203 channel=85
					4, 3, -5, 6, 8, -8, 7, 2, -7,
					-- layer=2 filter=203 channel=86
					-3, -3, -3, -7, 1, -10, -1, 3, -5,
					-- layer=2 filter=203 channel=87
					3, -8, 5, -6, 1, -16, -12, -15, 3,
					-- layer=2 filter=203 channel=88
					-8, -4, -16, -6, -11, 5, -16, -7, -7,
					-- layer=2 filter=203 channel=89
					0, -6, 0, -2, 10, -4, -17, -1, -10,
					-- layer=2 filter=203 channel=90
					-5, -9, -8, 7, 6, -9, -7, 5, -8,
					-- layer=2 filter=203 channel=91
					-1, 10, 6, 4, -4, 7, 1, -5, 2,
					-- layer=2 filter=203 channel=92
					0, 0, -13, -6, 5, 0, -18, -3, 0,
					-- layer=2 filter=203 channel=93
					-4, -10, -11, 0, 6, -14, 4, 5, -5,
					-- layer=2 filter=203 channel=94
					6, -9, 5, -3, -18, -9, 3, -12, 9,
					-- layer=2 filter=203 channel=95
					-8, -1, 2, 7, -9, 6, 1, -5, -1,
					-- layer=2 filter=203 channel=96
					0, -15, -17, 12, 7, 4, 0, 2, -7,
					-- layer=2 filter=203 channel=97
					-3, -4, 6, 3, 9, 0, -6, -7, 0,
					-- layer=2 filter=203 channel=98
					12, 6, -5, -7, 4, 0, 5, -4, -9,
					-- layer=2 filter=203 channel=99
					-2, 0, -7, 3, -12, 3, 3, -4, 0,
					-- layer=2 filter=203 channel=100
					-15, -12, -8, -12, -6, -6, -6, -2, 5,
					-- layer=2 filter=203 channel=101
					-9, -3, 2, -5, -8, 3, 0, -7, -7,
					-- layer=2 filter=203 channel=102
					2, -10, 1, 11, -5, 4, 1, -2, -13,
					-- layer=2 filter=203 channel=103
					4, -9, -3, 7, -8, 3, 4, -7, 7,
					-- layer=2 filter=203 channel=104
					5, -7, -8, -14, -8, 1, -16, -5, 4,
					-- layer=2 filter=203 channel=105
					-3, -6, 4, 0, 4, -2, 0, 2, -5,
					-- layer=2 filter=203 channel=106
					0, -10, 0, -3, 3, -14, 5, 6, -6,
					-- layer=2 filter=203 channel=107
					-4, 1, -3, -5, -8, 6, -2, 2, -2,
					-- layer=2 filter=203 channel=108
					-8, 0, 0, -5, -8, -5, -2, -2, 0,
					-- layer=2 filter=203 channel=109
					3, 8, -4, -6, -5, -7, -4, 4, 0,
					-- layer=2 filter=203 channel=110
					0, 1, -13, -3, 7, -4, -9, -2, -6,
					-- layer=2 filter=203 channel=111
					-2, -2, 6, 8, -9, 3, -10, -2, 3,
					-- layer=2 filter=203 channel=112
					-9, -8, -5, -16, 5, -7, 5, -4, 3,
					-- layer=2 filter=203 channel=113
					3, -1, -8, -13, -2, -9, -2, -11, 4,
					-- layer=2 filter=203 channel=114
					-10, -9, 2, 8, 8, 3, 3, -6, 8,
					-- layer=2 filter=203 channel=115
					-4, 0, 0, 3, 8, 7, -6, 8, -6,
					-- layer=2 filter=203 channel=116
					-2, -2, -9, -6, 8, -15, -20, 9, -12,
					-- layer=2 filter=203 channel=117
					-7, -9, -17, -13, 5, 9, 0, -7, -17,
					-- layer=2 filter=203 channel=118
					-9, -6, -3, -8, 0, -8, -7, 1, -13,
					-- layer=2 filter=203 channel=119
					-3, -9, -8, -13, 3, -16, -14, -12, -8,
					-- layer=2 filter=203 channel=120
					4, 3, -10, -5, 3, -2, -3, 9, -1,
					-- layer=2 filter=203 channel=121
					-4, 8, 7, -1, 5, 5, 3, 5, -8,
					-- layer=2 filter=203 channel=122
					-3, -3, 2, 1, -7, -4, -9, 9, 4,
					-- layer=2 filter=203 channel=123
					7, -4, -3, 9, 10, 1, -17, -8, -2,
					-- layer=2 filter=203 channel=124
					-8, -14, -5, 8, 8, 2, -18, -16, -2,
					-- layer=2 filter=203 channel=125
					5, 3, -5, -7, 11, -8, 6, -11, -5,
					-- layer=2 filter=203 channel=126
					0, 2, 1, 0, -9, 5, 9, -10, 0,
					-- layer=2 filter=203 channel=127
					-1, -11, -6, -4, -8, -2, -13, -9, 5,
					-- layer=2 filter=204 channel=0
					-10, -11, -20, -9, -27, -20, 10, -9, -22,
					-- layer=2 filter=204 channel=1
					20, 14, 31, -10, -3, 12, -26, 3, 14,
					-- layer=2 filter=204 channel=2
					-7, 2, -8, -2, -2, 13, 3, 4, 6,
					-- layer=2 filter=204 channel=3
					31, 0, -28, 12, -1, 0, 8, 10, -6,
					-- layer=2 filter=204 channel=4
					-31, -41, -33, 8, -21, -46, -14, -28, -24,
					-- layer=2 filter=204 channel=5
					-8, -10, 9, 5, 2, 10, 12, 12, 0,
					-- layer=2 filter=204 channel=6
					-40, -2, -14, 10, 33, 16, -30, -29, -24,
					-- layer=2 filter=204 channel=7
					20, 0, -43, 29, 27, -11, 13, 46, 0,
					-- layer=2 filter=204 channel=8
					-11, -7, 5, 0, 7, -1, -6, 10, -10,
					-- layer=2 filter=204 channel=9
					9, 8, -26, 19, 10, -24, 8, 21, -14,
					-- layer=2 filter=204 channel=10
					29, 20, -33, 5, 0, -24, 23, 8, -14,
					-- layer=2 filter=204 channel=11
					-8, -4, -10, 5, 12, -9, -27, 5, -12,
					-- layer=2 filter=204 channel=12
					16, 24, 17, -11, -36, -15, -16, -7, 8,
					-- layer=2 filter=204 channel=13
					4, 0, 0, -3, 3, 2, -5, 9, -7,
					-- layer=2 filter=204 channel=14
					15, 31, 16, -23, -13, 7, -15, -11, -23,
					-- layer=2 filter=204 channel=15
					22, 33, 0, 10, 43, 21, 9, -3, 7,
					-- layer=2 filter=204 channel=16
					8, -29, -56, 14, 1, -62, 0, -13, -11,
					-- layer=2 filter=204 channel=17
					2, 11, 7, -8, 7, 0, 4, 7, 1,
					-- layer=2 filter=204 channel=18
					-26, 0, 3, 29, 11, 29, 31, -9, 34,
					-- layer=2 filter=204 channel=19
					-16, 3, 15, -7, 35, 1, -10, 49, 35,
					-- layer=2 filter=204 channel=20
					-4, -3, -4, 8, 8, 8, 9, -5, 8,
					-- layer=2 filter=204 channel=21
					-3, 0, 0, -5, 3, 3, 0, -6, -16,
					-- layer=2 filter=204 channel=22
					-7, 0, -2, -7, 2, 11, -8, -8, -2,
					-- layer=2 filter=204 channel=23
					8, -17, -6, 36, -28, -15, 5, -1, -41,
					-- layer=2 filter=204 channel=24
					54, 1, -38, 16, -45, -5, 5, -23, -7,
					-- layer=2 filter=204 channel=25
					-28, -51, -19, -26, -47, -15, -50, -47, -25,
					-- layer=2 filter=204 channel=26
					-5, 9, 10, 6, 5, -7, -3, 1, 7,
					-- layer=2 filter=204 channel=27
					-18, 10, 12, -4, 1, 0, -2, 8, 12,
					-- layer=2 filter=204 channel=28
					6, -24, -52, 35, -17, -36, 31, 16, -8,
					-- layer=2 filter=204 channel=29
					7, 7, 2, 9, 6, -4, 2, 8, 9,
					-- layer=2 filter=204 channel=30
					4, 6, -18, 7, 19, -17, 10, -6, -11,
					-- layer=2 filter=204 channel=31
					58, 34, -57, 74, -34, -29, -24, 17, -33,
					-- layer=2 filter=204 channel=32
					5, 0, -10, 2, 7, 2, 1, 8, -2,
					-- layer=2 filter=204 channel=33
					67, 59, 38, 1, 7, -29, 14, -17, -47,
					-- layer=2 filter=204 channel=34
					-12, -51, -31, 28, 42, 7, -6, -5, -12,
					-- layer=2 filter=204 channel=35
					-12, -4, -2, -12, -12, -19, 2, 11, 10,
					-- layer=2 filter=204 channel=36
					-5, 11, -2, 0, 0, -7, 12, -1, -8,
					-- layer=2 filter=204 channel=37
					-6, 14, 9, -6, 11, 16, -8, 0, 1,
					-- layer=2 filter=204 channel=38
					0, 8, -6, -13, 2, 17, -15, -9, -39,
					-- layer=2 filter=204 channel=39
					11, 1, -37, 4, -16, -39, 34, 22, -15,
					-- layer=2 filter=204 channel=40
					29, -27, 12, -4, -16, 43, -42, -33, 45,
					-- layer=2 filter=204 channel=41
					10, 5, 6, 8, -1, -10, -2, 3, -2,
					-- layer=2 filter=204 channel=42
					17, 30, 13, 33, -12, 15, 20, -7, -10,
					-- layer=2 filter=204 channel=43
					27, -8, -18, -5, 5, 30, 45, 21, 28,
					-- layer=2 filter=204 channel=44
					4, 4, -7, 3, 1, -4, 2, -5, 1,
					-- layer=2 filter=204 channel=45
					-19, -23, -12, 10, -7, -1, 7, 14, 26,
					-- layer=2 filter=204 channel=46
					8, 15, -20, -30, 16, -62, 15, 13, -20,
					-- layer=2 filter=204 channel=47
					6, -20, 10, -4, -9, -50, -13, -33, -48,
					-- layer=2 filter=204 channel=48
					-10, -1, -10, 9, -7, -6, 0, 3, -10,
					-- layer=2 filter=204 channel=49
					-31, 44, 42, 21, 16, 40, 40, -19, 6,
					-- layer=2 filter=204 channel=50
					27, 29, 21, -1, -1, 4, -9, -11, 12,
					-- layer=2 filter=204 channel=51
					-10, 1, 4, -6, 16, 24, -18, -4, -19,
					-- layer=2 filter=204 channel=52
					-40, 5, 22, -11, 10, 11, -11, -3, 0,
					-- layer=2 filter=204 channel=53
					-17, 41, 37, 3, 51, -8, 13, 3, -51,
					-- layer=2 filter=204 channel=54
					0, -28, -27, -4, -10, -9, -10, -24, -15,
					-- layer=2 filter=204 channel=55
					8, 5, -11, -2, 4, -5, 0, 7, -10,
					-- layer=2 filter=204 channel=56
					2, -2, 9, 20, 24, -2, -17, -5, -13,
					-- layer=2 filter=204 channel=57
					-3, 0, -11, -11, -10, -2, -11, -7, 3,
					-- layer=2 filter=204 channel=58
					28, 22, 12, 20, -10, -22, -30, 16, 17,
					-- layer=2 filter=204 channel=59
					18, -9, 49, 26, -5, 5, 0, 5, 6,
					-- layer=2 filter=204 channel=60
					4, -13, 23, 3, 16, 55, -8, 6, 11,
					-- layer=2 filter=204 channel=61
					-13, 18, 54, 17, 48, 60, 3, 5, 52,
					-- layer=2 filter=204 channel=62
					-50, -25, -9, -4, 4, 3, -47, -34, -20,
					-- layer=2 filter=204 channel=63
					17, -14, -7, 19, -22, -47, 37, 17, -42,
					-- layer=2 filter=204 channel=64
					21, 1, -18, 50, 0, -6, 12, -8, -13,
					-- layer=2 filter=204 channel=65
					-1, 50, 22, 19, 55, 52, -13, 11, 32,
					-- layer=2 filter=204 channel=66
					-23, 39, 16, 18, 2, -41, 9, -26, 1,
					-- layer=2 filter=204 channel=67
					19, 19, -18, 36, 43, -44, 17, 8, -28,
					-- layer=2 filter=204 channel=68
					0, 6, 7, 3, -8, -6, 6, -9, -5,
					-- layer=2 filter=204 channel=69
					-4, 0, -5, 6, -5, -6, 0, -9, -17,
					-- layer=2 filter=204 channel=70
					-32, -23, -7, -9, -13, -23, -17, 7, 8,
					-- layer=2 filter=204 channel=71
					-17, -12, 19, 2, 30, 2, -6, 20, 8,
					-- layer=2 filter=204 channel=72
					29, -1, -23, -33, 13, -1, 33, 24, 2,
					-- layer=2 filter=204 channel=73
					29, 18, -63, -16, 53, 17, 19, 56, 3,
					-- layer=2 filter=204 channel=74
					18, -10, -27, 9, 6, -39, 4, 21, -2,
					-- layer=2 filter=204 channel=75
					-23, 5, 10, 0, -16, -21, 48, -49, -46,
					-- layer=2 filter=204 channel=76
					-34, -2, -12, 7, -28, -29, -30, 6, -1,
					-- layer=2 filter=204 channel=77
					8, -9, -4, -4, -5, 2, 3, 7, -10,
					-- layer=2 filter=204 channel=78
					-22, -22, -30, 4, -17, -12, -12, -23, -16,
					-- layer=2 filter=204 channel=79
					-5, 2, 7, -2, -5, 0, 2, -3, -5,
					-- layer=2 filter=204 channel=80
					23, -36, -66, 24, -17, -42, 37, 35, 14,
					-- layer=2 filter=204 channel=81
					-1, 7, -10, 4, -8, 0, -9, -3, -7,
					-- layer=2 filter=204 channel=82
					0, -10, 8, 0, 3, 3, -1, 4, 0,
					-- layer=2 filter=204 channel=83
					4, -2, -9, -20, -32, -45, -1, -14, -17,
					-- layer=2 filter=204 channel=84
					1, 1, -7, -7, 5, 0, 2, -1, -2,
					-- layer=2 filter=204 channel=85
					-2, -5, -8, 8, 0, 4, 5, -3, -4,
					-- layer=2 filter=204 channel=86
					-9, 5, 25, 8, 19, 16, 8, 25, -2,
					-- layer=2 filter=204 channel=87
					-37, -15, -18, 26, -11, 22, -23, -45, 11,
					-- layer=2 filter=204 channel=88
					31, 13, 4, 6, -13, -18, 5, -6, -7,
					-- layer=2 filter=204 channel=89
					-16, -17, -7, -12, -25, -22, 16, -2, 9,
					-- layer=2 filter=204 channel=90
					3, 0, 1, -5, 9, -4, 6, 4, 6,
					-- layer=2 filter=204 channel=91
					-23, -8, 16, -15, -30, -19, 0, -9, 7,
					-- layer=2 filter=204 channel=92
					5, 5, 31, -26, -25, 0, -27, -2, 12,
					-- layer=2 filter=204 channel=93
					-34, 14, -1, 2, 2, 19, -31, 8, 2,
					-- layer=2 filter=204 channel=94
					4, 8, 35, 32, 30, 40, -1, 29, 1,
					-- layer=2 filter=204 channel=95
					3, 2, -5, 6, -1, -8, 14, -1, -3,
					-- layer=2 filter=204 channel=96
					-26, -10, 23, -8, -13, 20, -4, -16, -39,
					-- layer=2 filter=204 channel=97
					53, -1, -17, 17, -7, -43, 25, -38, -47,
					-- layer=2 filter=204 channel=98
					0, -38, -28, -1, -20, -34, -29, -10, -6,
					-- layer=2 filter=204 channel=99
					-24, -8, 49, 22, 31, 18, -22, 9, 0,
					-- layer=2 filter=204 channel=100
					-5, -49, -51, 5, -36, -13, 5, 15, 1,
					-- layer=2 filter=204 channel=101
					-7, -15, 13, 2, 13, 10, -34, 15, -1,
					-- layer=2 filter=204 channel=102
					-43, 14, 7, -10, 0, 61, -24, -14, 22,
					-- layer=2 filter=204 channel=103
					14, 35, 4, 7, -33, 38, -76, 19, -12,
					-- layer=2 filter=204 channel=104
					-17, 29, 53, 5, 41, 37, 39, 20, 5,
					-- layer=2 filter=204 channel=105
					-5, -55, 7, 16, -51, -28, 9, 24, 8,
					-- layer=2 filter=204 channel=106
					20, 19, -4, 6, -4, -18, -17, -23, -64,
					-- layer=2 filter=204 channel=107
					16, 14, -10, -1, -31, 24, 4, -6, -39,
					-- layer=2 filter=204 channel=108
					-24, 26, 11, -11, 29, 11, -9, -23, -5,
					-- layer=2 filter=204 channel=109
					-10, 4, 14, -17, 9, -6, 4, -1, -11,
					-- layer=2 filter=204 channel=110
					20, -32, 19, 25, -30, -11, 3, 12, 27,
					-- layer=2 filter=204 channel=111
					0, -8, -4, 0, 7, 1, -3, -12, -5,
					-- layer=2 filter=204 channel=112
					-4, 32, 46, -15, 5, 13, -27, -9, 0,
					-- layer=2 filter=204 channel=113
					-3, 16, 38, 0, 17, 0, 10, 7, -7,
					-- layer=2 filter=204 channel=114
					-2, 19, -6, 8, 7, 13, 0, 4, 1,
					-- layer=2 filter=204 channel=115
					4, -10, 12, 6, 2, 8, 9, -10, 0,
					-- layer=2 filter=204 channel=116
					-56, 8, 4, 20, 20, 34, -13, -36, -2,
					-- layer=2 filter=204 channel=117
					-18, 20, -14, -22, 4, -11, -9, 25, -37,
					-- layer=2 filter=204 channel=118
					13, -24, -18, 20, 5, -1, 19, -13, 21,
					-- layer=2 filter=204 channel=119
					-15, -55, -24, 22, -21, -15, 8, -23, 16,
					-- layer=2 filter=204 channel=120
					5, 8, -7, -3, 2, 10, -2, -6, -8,
					-- layer=2 filter=204 channel=121
					-6, -6, -2, -8, 7, -5, -10, -1, 5,
					-- layer=2 filter=204 channel=122
					-14, 7, 0, 8, 4, -9, 3, 3, -15,
					-- layer=2 filter=204 channel=123
					26, -36, -5, 3, 40, -20, 29, 28, -7,
					-- layer=2 filter=204 channel=124
					26, 6, -7, 32, 25, 21, -2, -29, -1,
					-- layer=2 filter=204 channel=125
					-6, -10, -7, -2, -1, -12, -5, -7, 8,
					-- layer=2 filter=204 channel=126
					6, -59, 32, -18, 21, 15, 0, 41, -10,
					-- layer=2 filter=204 channel=127
					25, 18, -14, -28, -15, -3, 5, 3, -32,
					-- layer=2 filter=205 channel=0
					18, -10, 21, 20, 0, -38, 67, -23, -9,
					-- layer=2 filter=205 channel=1
					-15, 23, -6, -10, 13, 35, -53, -16, 41,
					-- layer=2 filter=205 channel=2
					-2, 2, -6, 2, -2, 3, -1, -6, 7,
					-- layer=2 filter=205 channel=3
					18, -16, -21, 36, 1, -45, 31, 27, -40,
					-- layer=2 filter=205 channel=4
					-8, 11, 12, -66, 24, 24, -18, 17, 20,
					-- layer=2 filter=205 channel=5
					-17, -2, -10, 12, -50, -43, 35, 13, -40,
					-- layer=2 filter=205 channel=6
					-17, -24, -74, -50, -47, -38, -37, -42, -21,
					-- layer=2 filter=205 channel=7
					-9, -32, -32, -21, 22, 4, 21, 12, 18,
					-- layer=2 filter=205 channel=8
					6, -7, 6, 1, 7, 2, -3, -5, -3,
					-- layer=2 filter=205 channel=9
					-28, 12, 46, -20, 1, 10, 22, -19, -21,
					-- layer=2 filter=205 channel=10
					-2, -13, 5, 33, 3, -17, 32, -21, -31,
					-- layer=2 filter=205 channel=11
					14, -8, -12, 27, -4, -14, 26, 9, 0,
					-- layer=2 filter=205 channel=12
					-2, 21, -14, -11, 12, 3, -49, 13, 31,
					-- layer=2 filter=205 channel=13
					8, 4, -4, -9, 6, 5, -4, 10, -9,
					-- layer=2 filter=205 channel=14
					-3, 17, -4, -25, 0, -4, -31, -11, 30,
					-- layer=2 filter=205 channel=15
					-5, -25, -76, 0, -4, -28, 28, -21, 50,
					-- layer=2 filter=205 channel=16
					-11, 15, 47, -55, -5, 42, -54, 6, 23,
					-- layer=2 filter=205 channel=17
					-3, -8, 1, -7, 6, 1, 2, 3, -5,
					-- layer=2 filter=205 channel=18
					8, 32, -26, -8, -5, -18, -15, 53, 16,
					-- layer=2 filter=205 channel=19
					3, 15, 4, -16, 39, 45, -35, 8, 20,
					-- layer=2 filter=205 channel=20
					0, -4, -10, -5, 0, 1, -1, -1, 4,
					-- layer=2 filter=205 channel=21
					18, 15, 17, 22, 6, -8, 14, 14, 0,
					-- layer=2 filter=205 channel=22
					-2, 7, -6, -2, 3, 9, -10, 5, -6,
					-- layer=2 filter=205 channel=23
					4, 4, 56, -76, -22, 25, -57, -45, 4,
					-- layer=2 filter=205 channel=24
					2, -22, -8, 47, -11, -12, 47, 5, -59,
					-- layer=2 filter=205 channel=25
					39, -18, -36, 56, -25, -13, 61, 9, -40,
					-- layer=2 filter=205 channel=26
					-8, -9, -12, -4, -1, -10, -6, 1, -3,
					-- layer=2 filter=205 channel=27
					-14, 12, 38, -22, 4, 21, 0, -7, -1,
					-- layer=2 filter=205 channel=28
					-12, 12, 30, -33, -39, -46, 18, 38, 28,
					-- layer=2 filter=205 channel=29
					1, 0, -10, -4, -4, 4, 1, 5, -5,
					-- layer=2 filter=205 channel=30
					-14, 32, 14, -49, -23, 9, -45, 7, -2,
					-- layer=2 filter=205 channel=31
					-72, 2, 63, -24, 36, 21, 0, -45, 49,
					-- layer=2 filter=205 channel=32
					4, -8, 8, -2, -7, 0, 13, 6, 0,
					-- layer=2 filter=205 channel=33
					20, -34, -39, 9, -16, -14, -22, 25, 27,
					-- layer=2 filter=205 channel=34
					-35, 3, 1, -27, 0, -65, -91, -20, -38,
					-- layer=2 filter=205 channel=35
					-7, 21, 17, -26, -49, -55, 1, 39, 23,
					-- layer=2 filter=205 channel=36
					7, -6, -19, 10, 17, -13, 0, -13, 0,
					-- layer=2 filter=205 channel=37
					-8, 2, 9, 2, -20, -8, 7, -12, -7,
					-- layer=2 filter=205 channel=38
					-31, 1, -2, -16, -56, -9, -21, -2, -11,
					-- layer=2 filter=205 channel=39
					-22, -5, 6, -67, -12, 37, -64, -24, 4,
					-- layer=2 filter=205 channel=40
					-13, -10, -29, -32, -67, -6, 0, 18, 26,
					-- layer=2 filter=205 channel=41
					-1, 6, -7, -6, 0, -7, -6, 10, 4,
					-- layer=2 filter=205 channel=42
					4, 29, 27, -51, 6, 12, -75, -9, 31,
					-- layer=2 filter=205 channel=43
					0, 11, -21, -35, -25, -58, 1, 3, -16,
					-- layer=2 filter=205 channel=44
					8, -8, 4, 11, -9, 3, 10, -7, -8,
					-- layer=2 filter=205 channel=45
					-18, 23, 41, -21, 25, 26, -14, -21, 54,
					-- layer=2 filter=205 channel=46
					-36, -13, 10, -27, -11, 32, -38, 1, -19,
					-- layer=2 filter=205 channel=47
					-6, 1, 38, -19, 26, -4, 14, 37, 54,
					-- layer=2 filter=205 channel=48
					2, -5, -3, 5, 4, 2, -11, -3, -8,
					-- layer=2 filter=205 channel=49
					16, 45, -7, 0, 21, 13, 3, 13, 25,
					-- layer=2 filter=205 channel=50
					21, 16, 27, 19, 32, 8, -11, -13, -18,
					-- layer=2 filter=205 channel=51
					37, 7, -18, 40, -17, -31, 31, -1, -22,
					-- layer=2 filter=205 channel=52
					8, -14, -32, -59, -17, -52, -26, -2, 18,
					-- layer=2 filter=205 channel=53
					9, -21, -34, 2, 27, 12, 35, -2, -16,
					-- layer=2 filter=205 channel=54
					-3, 4, -8, -18, 11, 1, -19, 27, 16,
					-- layer=2 filter=205 channel=55
					-2, 3, -10, 3, 2, -8, 10, 11, -4,
					-- layer=2 filter=205 channel=56
					9, -11, -14, 9, -23, -23, 59, 18, -3,
					-- layer=2 filter=205 channel=57
					-5, -2, -3, 2, -2, -7, -2, -6, -3,
					-- layer=2 filter=205 channel=58
					1, 3, -30, -24, 19, 2, -42, 2, 37,
					-- layer=2 filter=205 channel=59
					-15, -13, 0, -40, -27, 11, -40, -59, 41,
					-- layer=2 filter=205 channel=60
					-9, -10, -11, 19, -1, -8, -22, 12, -28,
					-- layer=2 filter=205 channel=61
					-19, -18, 9, 5, 18, 23, 28, 1, 11,
					-- layer=2 filter=205 channel=62
					14, 29, -26, -16, -13, -20, -74, -6, 4,
					-- layer=2 filter=205 channel=63
					-50, -14, 34, -60, -15, 39, -43, -41, -3,
					-- layer=2 filter=205 channel=64
					-54, 8, 4, -82, -23, 2, -72, -40, -5,
					-- layer=2 filter=205 channel=65
					-35, -13, -25, -15, -6, -25, -6, -63, 10,
					-- layer=2 filter=205 channel=66
					20, -14, 4, -1, -25, 43, 34, 33, 41,
					-- layer=2 filter=205 channel=67
					-20, 4, 17, -30, -43, 11, 23, 42, -15,
					-- layer=2 filter=205 channel=68
					-3, 2, -4, 9, -4, 0, -1, -1, -2,
					-- layer=2 filter=205 channel=69
					-28, 1, 7, -48, 6, 27, -88, -45, 20,
					-- layer=2 filter=205 channel=70
					-21, -5, 11, -36, -40, -44, 13, 37, 15,
					-- layer=2 filter=205 channel=71
					-12, 25, 8, -2, 8, 12, -7, -26, 2,
					-- layer=2 filter=205 channel=72
					35, 7, -12, -28, 7, 11, -18, 37, 8,
					-- layer=2 filter=205 channel=73
					19, -14, 0, 52, 31, 20, 57, 8, 40,
					-- layer=2 filter=205 channel=74
					-26, 8, -9, -36, -3, 42, -54, -25, 17,
					-- layer=2 filter=205 channel=75
					-72, 21, 6, -53, -5, 51, -9, -27, 51,
					-- layer=2 filter=205 channel=76
					12, -14, 14, 1, 58, -18, 61, -28, 1,
					-- layer=2 filter=205 channel=77
					3, 9, 5, -10, 9, -3, -10, -3, 11,
					-- layer=2 filter=205 channel=78
					58, -4, -11, 14, -13, 2, 0, -26, 8,
					-- layer=2 filter=205 channel=79
					-9, -1, -7, 0, 0, -5, -6, -6, -8,
					-- layer=2 filter=205 channel=80
					-40, 12, 4, -50, -41, 22, -32, -32, 2,
					-- layer=2 filter=205 channel=81
					0, 0, 20, 4, -9, 2, -18, -8, 1,
					-- layer=2 filter=205 channel=82
					8, 9, 4, -3, 0, -9, -12, -11, 0,
					-- layer=2 filter=205 channel=83
					-14, 3, 38, -46, 31, 55, -62, -25, 31,
					-- layer=2 filter=205 channel=84
					-10, 0, -9, -6, -9, 2, 0, -1, -6,
					-- layer=2 filter=205 channel=85
					21, 4, 0, -2, 4, 5, 15, 4, -8,
					-- layer=2 filter=205 channel=86
					-6, -6, -4, 10, -2, 7, -1, 13, 21,
					-- layer=2 filter=205 channel=87
					-30, -10, -45, -38, -28, -71, 43, 15, 14,
					-- layer=2 filter=205 channel=88
					-31, -4, 24, -38, -22, 21, -51, -16, 8,
					-- layer=2 filter=205 channel=89
					28, 24, -14, -44, 25, 24, -24, -50, 48,
					-- layer=2 filter=205 channel=90
					-10, -6, 9, -1, -7, -3, 6, -2, 3,
					-- layer=2 filter=205 channel=91
					-11, 0, -12, -19, 8, -19, -32, 3, 50,
					-- layer=2 filter=205 channel=92
					0, 44, 13, -23, 22, 31, -57, 30, 50,
					-- layer=2 filter=205 channel=93
					17, 14, -13, -70, -29, -31, -78, -44, -45,
					-- layer=2 filter=205 channel=94
					6, -2, -41, -6, 11, 45, 7, 36, 18,
					-- layer=2 filter=205 channel=95
					-4, -4, 0, -18, -20, -17, -18, 3, 0,
					-- layer=2 filter=205 channel=96
					-32, -31, 21, -50, -18, -30, -15, -36, 2,
					-- layer=2 filter=205 channel=97
					-28, -16, -4, -6, -13, 49, -20, -60, 1,
					-- layer=2 filter=205 channel=98
					-34, 27, 21, -37, -7, -31, 22, 18, 16,
					-- layer=2 filter=205 channel=99
					28, -7, 1, 22, 17, -20, 47, -28, 22,
					-- layer=2 filter=205 channel=100
					-44, 0, 28, -26, 5, 6, -65, -51, 10,
					-- layer=2 filter=205 channel=101
					27, 7, -17, 11, -2, -35, 39, -3, -6,
					-- layer=2 filter=205 channel=102
					-13, 18, 12, -58, 33, 9, -24, 36, 37,
					-- layer=2 filter=205 channel=103
					-16, -2, 9, -2, -42, -49, -2, 19, 4,
					-- layer=2 filter=205 channel=104
					13, 23, -47, -12, -5, -17, -8, 21, 27,
					-- layer=2 filter=205 channel=105
					14, 39, 5, 30, 50, 4, 52, -14, 13,
					-- layer=2 filter=205 channel=106
					24, -9, -15, 17, -41, -71, 52, 28, -49,
					-- layer=2 filter=205 channel=107
					-24, 19, 44, 48, -18, -12, -6, 45, 38,
					-- layer=2 filter=205 channel=108
					-12, 48, 32, -52, 28, 7, -23, -35, 15,
					-- layer=2 filter=205 channel=109
					14, 0, 7, 2, 10, -26, -2, 5, -1,
					-- layer=2 filter=205 channel=110
					8, 8, 16, -66, -1, -1, -47, -27, 20,
					-- layer=2 filter=205 channel=111
					0, 0, 4, -9, 5, -3, -5, 2, -9,
					-- layer=2 filter=205 channel=112
					13, 23, 18, 72, 0, -19, 77, 30, 18,
					-- layer=2 filter=205 channel=113
					-26, 46, 28, -59, 3, 1, -15, -27, 7,
					-- layer=2 filter=205 channel=114
					-11, -5, 0, 4, -14, -17, -4, -4, -2,
					-- layer=2 filter=205 channel=115
					-9, -7, 9, 5, -3, 5, -8, 1, -8,
					-- layer=2 filter=205 channel=116
					-30, -18, -38, -55, -53, -64, -13, 37, -8,
					-- layer=2 filter=205 channel=117
					-6, 3, -19, 28, 35, 14, 11, 37, 16,
					-- layer=2 filter=205 channel=118
					-11, -23, -18, 0, -30, -24, -4, -25, -13,
					-- layer=2 filter=205 channel=119
					-5, 15, 40, -38, 16, 30, -40, 54, 65,
					-- layer=2 filter=205 channel=120
					5, 8, 2, 6, -3, -2, -2, 10, -3,
					-- layer=2 filter=205 channel=121
					-9, -10, 1, 10, -8, -1, -3, -9, 9,
					-- layer=2 filter=205 channel=122
					-7, -14, -6, -5, 8, -3, 12, 6, -11,
					-- layer=2 filter=205 channel=123
					-8, 1, -10, -8, 29, 17, 17, 13, 10,
					-- layer=2 filter=205 channel=124
					6, -12, -40, 15, 14, -13, 16, 0, 32,
					-- layer=2 filter=205 channel=125
					10, 10, -9, -5, 0, -9, -10, 3, 6,
					-- layer=2 filter=205 channel=126
					10, 38, 48, -43, -7, 1, -76, -36, 31,
					-- layer=2 filter=205 channel=127
					-10, 8, 52, -25, -3, 37, -33, 12, 67,
					-- layer=2 filter=206 channel=0
					-19, -12, 8, 9, 0, -2, -6, 18, 17,
					-- layer=2 filter=206 channel=1
					-18, -18, 15, -48, -32, -7, -12, 4, 25,
					-- layer=2 filter=206 channel=2
					11, 2, -7, -7, -3, 3, -8, 11, 9,
					-- layer=2 filter=206 channel=3
					6, -12, -5, 3, 7, -14, 19, 12, 12,
					-- layer=2 filter=206 channel=4
					-8, 6, -6, 4, 19, 14, 41, 38, 44,
					-- layer=2 filter=206 channel=5
					-28, 6, -8, 3, -8, 4, -7, 19, 29,
					-- layer=2 filter=206 channel=6
					-19, -21, -52, -38, -17, -21, -15, -8, -4,
					-- layer=2 filter=206 channel=7
					-66, -49, -8, -52, -93, -49, -23, -13, 0,
					-- layer=2 filter=206 channel=8
					-4, -4, 6, -2, 8, 7, -4, -1, -7,
					-- layer=2 filter=206 channel=9
					16, -7, -24, 20, 23, -22, 18, -15, 0,
					-- layer=2 filter=206 channel=10
					10, 2, -18, 11, 12, 1, 15, 19, 28,
					-- layer=2 filter=206 channel=11
					0, 11, 11, -21, -1, 5, -10, -3, 15,
					-- layer=2 filter=206 channel=12
					-41, -57, -13, -74, -70, -23, -44, -7, -14,
					-- layer=2 filter=206 channel=13
					-2, -4, 6, 0, 10, -10, 2, -3, 2,
					-- layer=2 filter=206 channel=14
					-33, -13, 28, -59, -50, 1, -14, -50, -28,
					-- layer=2 filter=206 channel=15
					0, -2, 1, -63, 38, 13, -42, -7, 0,
					-- layer=2 filter=206 channel=16
					-24, -27, 7, 4, 8, 7, 26, 16, 11,
					-- layer=2 filter=206 channel=17
					4, -9, -12, -3, 0, 5, 8, 6, -7,
					-- layer=2 filter=206 channel=18
					-8, -1, 0, -52, -14, 7, -27, -8, -7,
					-- layer=2 filter=206 channel=19
					-21, -13, -30, -23, 0, 8, -32, -18, 14,
					-- layer=2 filter=206 channel=20
					-3, 8, -4, 3, -8, 2, -2, 7, 7,
					-- layer=2 filter=206 channel=21
					-14, -4, 3, -3, -13, -8, -2, -16, -3,
					-- layer=2 filter=206 channel=22
					-8, -8, -3, -7, 3, -7, -5, -9, 4,
					-- layer=2 filter=206 channel=23
					-9, 6, -6, 22, 11, -7, 14, 41, 12,
					-- layer=2 filter=206 channel=24
					-5, 1, 36, -7, 8, -11, 6, 16, 20,
					-- layer=2 filter=206 channel=25
					-21, 0, 15, -3, 1, -3, 12, 14, 3,
					-- layer=2 filter=206 channel=26
					-10, -5, 6, 5, -5, -1, 2, 0, 11,
					-- layer=2 filter=206 channel=27
					-6, -28, -30, -10, -7, 44, -10, 1, 52,
					-- layer=2 filter=206 channel=28
					-92, -30, -34, -41, -14, -3, -32, 19, -15,
					-- layer=2 filter=206 channel=29
					-4, -8, 2, -8, -10, 0, 2, -7, 4,
					-- layer=2 filter=206 channel=30
					10, -13, 11, 17, 2, 21, 23, 0, 15,
					-- layer=2 filter=206 channel=31
					34, 67, 29, -13, 49, 26, -35, 19, 33,
					-- layer=2 filter=206 channel=32
					-8, 0, -5, 0, 0, 5, -4, 0, 5,
					-- layer=2 filter=206 channel=33
					-28, -35, 42, -93, -15, 2, -45, 12, 59,
					-- layer=2 filter=206 channel=34
					36, -45, 28, -38, -22, 52, 16, 16, -23,
					-- layer=2 filter=206 channel=35
					-49, -2, -12, -15, 13, 1, -29, -12, -32,
					-- layer=2 filter=206 channel=36
					4, 7, 0, -6, 5, -12, 1, -4, -9,
					-- layer=2 filter=206 channel=37
					6, 5, -10, 2, -3, 6, -5, 11, 27,
					-- layer=2 filter=206 channel=38
					-34, -31, -1, -26, 5, 21, -34, 14, 34,
					-- layer=2 filter=206 channel=39
					-31, -11, -21, 11, 7, -22, 7, 0, -13,
					-- layer=2 filter=206 channel=40
					2, -14, 2, -29, 33, -25, -15, -14, -44,
					-- layer=2 filter=206 channel=41
					-7, 2, 1, 1, 10, -8, -8, 6, 7,
					-- layer=2 filter=206 channel=42
					-8, 3, -12, 3, 2, -33, 16, 13, 0,
					-- layer=2 filter=206 channel=43
					14, -15, -47, 22, 4, 25, -2, 14, 7,
					-- layer=2 filter=206 channel=44
					-6, 8, 2, 3, 5, -6, -3, 0, -2,
					-- layer=2 filter=206 channel=45
					14, 5, -15, -22, 54, 62, -23, 0, 34,
					-- layer=2 filter=206 channel=46
					-15, -20, -13, 2, 8, 0, 18, 21, 39,
					-- layer=2 filter=206 channel=47
					-57, -30, 27, -52, -18, -23, 10, -4, 3,
					-- layer=2 filter=206 channel=48
					0, -4, -6, 8, 7, -9, 1, -6, -6,
					-- layer=2 filter=206 channel=49
					25, 24, 41, -6, 10, -16, 8, -24, 10,
					-- layer=2 filter=206 channel=50
					-18, 6, 11, 3, -13, 8, -13, -1, -2,
					-- layer=2 filter=206 channel=51
					-2, 12, 23, 3, 10, 11, -13, -10, 5,
					-- layer=2 filter=206 channel=52
					19, 9, 1, -26, -25, -18, -6, -5, -2,
					-- layer=2 filter=206 channel=53
					18, 34, -29, -3, 40, -8, -47, -7, 6,
					-- layer=2 filter=206 channel=54
					-57, -17, -3, -29, -19, -7, -8, 37, 35,
					-- layer=2 filter=206 channel=55
					-8, 1, -2, -2, -2, -10, 6, 0, -1,
					-- layer=2 filter=206 channel=56
					-9, 6, -16, 4, -1, 9, -22, -14, 10,
					-- layer=2 filter=206 channel=57
					0, -4, 1, 8, 3, -4, -9, -8, -6,
					-- layer=2 filter=206 channel=58
					-69, -23, -18, -56, -47, -42, -66, -8, -2,
					-- layer=2 filter=206 channel=59
					-24, -36, 13, -61, -13, 14, -69, 12, 45,
					-- layer=2 filter=206 channel=60
					-15, -15, 3, -24, -9, 44, -3, 0, -5,
					-- layer=2 filter=206 channel=61
					-12, -6, -2, -11, 7, 12, -13, -11, 21,
					-- layer=2 filter=206 channel=62
					15, 15, -9, -37, 36, 4, 39, 9, -3,
					-- layer=2 filter=206 channel=63
					-22, -1, -26, 10, -5, -16, 17, 41, -2,
					-- layer=2 filter=206 channel=64
					12, -20, 12, 8, -13, -2, 40, 16, 0,
					-- layer=2 filter=206 channel=65
					25, -42, -4, -7, -8, 8, -18, -3, 12,
					-- layer=2 filter=206 channel=66
					-7, -3, 0, -21, -17, -21, 0, -11, 9,
					-- layer=2 filter=206 channel=67
					3, -1, -18, 7, 23, -9, -1, 3, 16,
					-- layer=2 filter=206 channel=68
					3, -1, 3, -7, 10, 7, 9, -5, -9,
					-- layer=2 filter=206 channel=69
					-11, -15, -1, -4, 3, -7, 42, 21, 0,
					-- layer=2 filter=206 channel=70
					-38, -21, -25, -10, 3, 18, -19, -2, -12,
					-- layer=2 filter=206 channel=71
					40, -4, 0, -11, 2, 37, -14, -19, 18,
					-- layer=2 filter=206 channel=72
					-76, -28, -10, -77, -59, 19, -54, -27, 5,
					-- layer=2 filter=206 channel=73
					7, 69, -45, 24, 34, 32, 28, 45, 6,
					-- layer=2 filter=206 channel=74
					-23, -25, -35, 7, 12, -15, 21, 29, -20,
					-- layer=2 filter=206 channel=75
					-49, -45, -33, -57, 6, 20, -19, -48, -43,
					-- layer=2 filter=206 channel=76
					-16, 1, -19, -30, 58, -9, 44, -15, 30,
					-- layer=2 filter=206 channel=77
					0, 8, -5, -5, 5, 10, -4, -8, 9,
					-- layer=2 filter=206 channel=78
					-1, -1, 0, 7, 12, 2, 16, 3, 5,
					-- layer=2 filter=206 channel=79
					10, -7, 9, -1, -4, 0, -6, -3, 11,
					-- layer=2 filter=206 channel=80
					7, 0, -16, 23, 20, 6, 45, 12, 35,
					-- layer=2 filter=206 channel=81
					4, 0, -2, 0, 10, -3, 9, 4, 3,
					-- layer=2 filter=206 channel=82
					-9, -6, 6, 2, 3, 5, 1, 0, 9,
					-- layer=2 filter=206 channel=83
					-9, -2, 16, 20, 4, 51, 11, 30, 34,
					-- layer=2 filter=206 channel=84
					-3, -1, -8, 0, 11, 6, 11, 9, -9,
					-- layer=2 filter=206 channel=85
					-12, 7, -16, 11, -8, 2, -5, -8, 6,
					-- layer=2 filter=206 channel=86
					4, 8, 26, -3, -10, 0, -6, -11, -2,
					-- layer=2 filter=206 channel=87
					-12, 12, 21, -59, 38, 22, -25, 38, 63,
					-- layer=2 filter=206 channel=88
					1, -21, 22, -2, 26, 15, 3, 24, 10,
					-- layer=2 filter=206 channel=89
					-28, -26, 12, -63, -14, 0, -35, -25, 11,
					-- layer=2 filter=206 channel=90
					-8, -3, 1, 4, -6, -5, 6, -8, -9,
					-- layer=2 filter=206 channel=91
					-62, -45, -43, -79, -29, -25, -28, 13, -2,
					-- layer=2 filter=206 channel=92
					-41, -25, -20, -75, -41, -43, -59, -11, -22,
					-- layer=2 filter=206 channel=93
					32, -7, -54, -9, -9, 5, 1, 8, -58,
					-- layer=2 filter=206 channel=94
					-30, 12, -25, -20, 23, 15, -1, -18, -19,
					-- layer=2 filter=206 channel=95
					-23, 0, -8, -5, 0, -5, -2, 1, 0,
					-- layer=2 filter=206 channel=96
					-14, 44, 22, -16, -12, 11, -21, -10, -6,
					-- layer=2 filter=206 channel=97
					0, -20, 2, 2, -18, -21, 30, -8, 22,
					-- layer=2 filter=206 channel=98
					-42, -63, -2, -39, -4, -39, 16, 13, -7,
					-- layer=2 filter=206 channel=99
					49, 0, 19, -1, 1, -2, -5, -34, 12,
					-- layer=2 filter=206 channel=100
					-15, -12, -36, -9, 12, 9, -17, 26, 45,
					-- layer=2 filter=206 channel=101
					42, 31, 16, -1, 1, -15, -6, -27, -21,
					-- layer=2 filter=206 channel=102
					24, 23, 13, -19, 1, 8, -11, -31, 4,
					-- layer=2 filter=206 channel=103
					27, -10, 7, -30, 22, 25, -37, -9, 9,
					-- layer=2 filter=206 channel=104
					12, 42, 9, -28, 65, -8, -32, -9, -11,
					-- layer=2 filter=206 channel=105
					-60, -7, 11, -58, 15, -39, 40, -29, 33,
					-- layer=2 filter=206 channel=106
					-34, -13, 3, -16, -24, 0, -14, 0, 20,
					-- layer=2 filter=206 channel=107
					-16, 5, 35, -26, 30, 6, -8, 23, -31,
					-- layer=2 filter=206 channel=108
					18, 7, 9, -11, -7, 35, -14, -18, 14,
					-- layer=2 filter=206 channel=109
					13, -7, -12, 12, -5, -2, -4, 4, 6,
					-- layer=2 filter=206 channel=110
					-15, -26, 3, 2, -15, 15, -7, 15, 22,
					-- layer=2 filter=206 channel=111
					-1, 4, -4, -12, 2, 7, -9, 6, 6,
					-- layer=2 filter=206 channel=112
					27, 2, 2, -4, 9, 0, -10, 6, 13,
					-- layer=2 filter=206 channel=113
					3, -24, 8, 10, -2, 2, 24, -8, -19,
					-- layer=2 filter=206 channel=114
					-3, 0, 5, -8, -8, -20, -6, -10, -17,
					-- layer=2 filter=206 channel=115
					-9, -3, -8, -2, -6, 3, -8, -1, 1,
					-- layer=2 filter=206 channel=116
					13, -1, -6, -61, -15, 25, -44, 29, 41,
					-- layer=2 filter=206 channel=117
					28, 19, 23, -18, -35, -17, -4, 14, 14,
					-- layer=2 filter=206 channel=118
					27, -9, -30, 21, 3, -12, 51, 21, 37,
					-- layer=2 filter=206 channel=119
					-22, -7, -11, -25, 0, 24, 32, 23, 19,
					-- layer=2 filter=206 channel=120
					-7, 3, 5, -3, -3, -6, -1, -10, 5,
					-- layer=2 filter=206 channel=121
					0, 9, -4, 4, 8, -2, 9, -8, 6,
					-- layer=2 filter=206 channel=122
					3, 3, 3, -6, 9, 13, 1, 13, 1,
					-- layer=2 filter=206 channel=123
					-54, -24, 15, -65, -28, -28, -9, -6, 7,
					-- layer=2 filter=206 channel=124
					-33, 7, 25, -73, 15, 8, -7, -20, 46,
					-- layer=2 filter=206 channel=125
					-1, 6, 6, 1, 5, 2, -3, 1, -6,
					-- layer=2 filter=206 channel=126
					-60, 38, -51, 0, -26, 14, -11, -1, -59,
					-- layer=2 filter=206 channel=127
					-11, -20, 20, -6, -10, 20, 15, 33, 13,
					-- layer=2 filter=207 channel=0
					1, -4, 0, -5, 3, -7, -12, -7, -4,
					-- layer=2 filter=207 channel=1
					-7, -13, -12, -13, -10, -7, 4, 2, -4,
					-- layer=2 filter=207 channel=2
					-2, 8, -1, -5, 9, -3, 1, 6, 8,
					-- layer=2 filter=207 channel=3
					-7, 8, 8, -6, -3, -7, 3, 7, 8,
					-- layer=2 filter=207 channel=4
					-13, -20, -1, -10, -8, -8, -6, 1, -9,
					-- layer=2 filter=207 channel=5
					2, -2, -3, -4, 1, 2, -16, -2, -4,
					-- layer=2 filter=207 channel=6
					-8, 0, 6, -11, -4, 0, 0, -11, -4,
					-- layer=2 filter=207 channel=7
					1, -1, -15, -21, -3, 3, 13, 11, -5,
					-- layer=2 filter=207 channel=8
					0, -1, -1, 11, -7, 2, 11, -7, -1,
					-- layer=2 filter=207 channel=9
					0, -4, -1, -11, -14, -6, -8, -15, -10,
					-- layer=2 filter=207 channel=10
					4, -8, -5, -3, -5, 4, -16, -1, -9,
					-- layer=2 filter=207 channel=11
					-6, -3, -14, 3, -5, -10, -8, 0, -3,
					-- layer=2 filter=207 channel=12
					-3, -3, -6, -14, -27, -11, -11, -9, -1,
					-- layer=2 filter=207 channel=13
					-9, 2, -4, -11, 8, 3, -11, 3, -8,
					-- layer=2 filter=207 channel=14
					0, -10, -14, -14, -26, -19, -18, 2, -10,
					-- layer=2 filter=207 channel=15
					-7, -14, -1, -11, 2, -12, -13, 0, -11,
					-- layer=2 filter=207 channel=16
					-4, 10, -3, 0, 1, 3, -8, -7, -3,
					-- layer=2 filter=207 channel=17
					9, -8, -4, 0, -1, 1, 1, 10, 6,
					-- layer=2 filter=207 channel=18
					-2, -16, -15, 1, 17, -13, -9, 0, 4,
					-- layer=2 filter=207 channel=19
					-2, -2, -4, -6, -12, -4, 8, 1, 0,
					-- layer=2 filter=207 channel=20
					-1, -11, 3, 4, -7, -4, 3, 0, -7,
					-- layer=2 filter=207 channel=21
					-1, 0, 4, -4, -9, -11, -1, -7, 5,
					-- layer=2 filter=207 channel=22
					-6, 8, -6, 0, 7, 8, 1, -9, 4,
					-- layer=2 filter=207 channel=23
					-10, -7, -14, 1, -13, -6, -9, 8, -7,
					-- layer=2 filter=207 channel=24
					-1, -15, -10, -16, -18, -7, -10, -14, -16,
					-- layer=2 filter=207 channel=25
					-3, -7, -8, 7, -2, -9, -8, -3, 7,
					-- layer=2 filter=207 channel=26
					0, -8, -8, 6, -6, -1, -8, 3, -7,
					-- layer=2 filter=207 channel=27
					-16, -11, 2, -10, 2, -9, 6, -3, 2,
					-- layer=2 filter=207 channel=28
					3, -6, -2, 2, 6, 8, 0, -2, 7,
					-- layer=2 filter=207 channel=29
					-3, 3, 0, 0, -1, -7, 6, 0, 4,
					-- layer=2 filter=207 channel=30
					-11, 0, -8, -8, 0, -14, -13, 2, -3,
					-- layer=2 filter=207 channel=31
					6, -11, -6, -15, -12, -6, 0, -10, 0,
					-- layer=2 filter=207 channel=32
					-2, -9, -6, -2, -10, 7, 0, 4, -3,
					-- layer=2 filter=207 channel=33
					-11, -7, -11, -22, -11, -8, -1, 2, -1,
					-- layer=2 filter=207 channel=34
					5, -18, -2, -6, -1, -5, 9, 0, 3,
					-- layer=2 filter=207 channel=35
					-2, -22, -19, 4, 2, 5, -4, 1, 4,
					-- layer=2 filter=207 channel=36
					3, -2, -4, 0, 0, 0, 2, -7, -3,
					-- layer=2 filter=207 channel=37
					-9, -18, -15, -4, 5, -15, 8, 0, -16,
					-- layer=2 filter=207 channel=38
					-8, -17, -11, 6, -11, -7, -13, 3, 7,
					-- layer=2 filter=207 channel=39
					-16, -14, -7, 0, -8, 0, -10, -6, -7,
					-- layer=2 filter=207 channel=40
					-16, -9, -14, -9, -17, 8, -15, -8, -14,
					-- layer=2 filter=207 channel=41
					0, 3, -7, -9, -9, -7, 0, 3, 8,
					-- layer=2 filter=207 channel=42
					1, 2, -11, -15, -17, -18, -15, -9, -12,
					-- layer=2 filter=207 channel=43
					-7, -16, 2, 4, 1, -2, -1, -2, -8,
					-- layer=2 filter=207 channel=44
					2, -3, -9, -4, -8, -11, 5, -9, 0,
					-- layer=2 filter=207 channel=45
					3, -2, 1, -8, 1, -13, 0, 6, 0,
					-- layer=2 filter=207 channel=46
					-1, -14, -13, 4, -3, -19, -3, -9, -2,
					-- layer=2 filter=207 channel=47
					-13, -4, 0, 3, 2, -2, -5, -14, 1,
					-- layer=2 filter=207 channel=48
					-6, 4, 0, -10, 5, 7, 8, -7, 0,
					-- layer=2 filter=207 channel=49
					4, -16, 12, -2, 7, 11, 2, 13, 6,
					-- layer=2 filter=207 channel=50
					-9, -5, -4, 5, -5, -9, 0, 5, -1,
					-- layer=2 filter=207 channel=51
					2, -10, 1, 6, -3, 0, 0, -9, -3,
					-- layer=2 filter=207 channel=52
					-17, 4, -11, -7, -8, -12, -1, -1, -13,
					-- layer=2 filter=207 channel=53
					-10, -14, -2, -6, -10, -6, -4, -6, 11,
					-- layer=2 filter=207 channel=54
					-6, -8, -7, -10, -17, 1, 5, 0, 0,
					-- layer=2 filter=207 channel=55
					4, -2, 0, -11, -3, 0, -4, 0, 7,
					-- layer=2 filter=207 channel=56
					-8, -7, -18, -3, 4, -7, -13, 0, -14,
					-- layer=2 filter=207 channel=57
					-11, 0, -6, 3, -2, -6, 0, 6, -2,
					-- layer=2 filter=207 channel=58
					-5, -2, -3, -26, -22, -10, -7, -7, -7,
					-- layer=2 filter=207 channel=59
					-4, 0, -6, 0, 0, 2, 1, -14, 1,
					-- layer=2 filter=207 channel=60
					2, -11, -4, -5, -12, -5, 0, 3, -5,
					-- layer=2 filter=207 channel=61
					-13, 6, 1, 1, -7, -3, 4, -11, -5,
					-- layer=2 filter=207 channel=62
					-9, -12, 0, 5, -7, -2, 3, 0, -1,
					-- layer=2 filter=207 channel=63
					-6, -13, 0, -7, 1, -8, 0, 0, -3,
					-- layer=2 filter=207 channel=64
					2, 1, -13, 0, -15, -6, -11, 4, -10,
					-- layer=2 filter=207 channel=65
					4, -9, 4, -8, 0, -8, 13, -10, 10,
					-- layer=2 filter=207 channel=66
					-1, -6, -1, 7, 4, -3, -5, 6, -6,
					-- layer=2 filter=207 channel=67
					-3, -19, -12, -8, -7, -5, -10, -17, -14,
					-- layer=2 filter=207 channel=68
					-8, 8, -6, -5, 6, -1, -3, -2, 4,
					-- layer=2 filter=207 channel=69
					2, 1, -5, -8, -25, -4, -2, -10, -10,
					-- layer=2 filter=207 channel=70
					-2, -20, -13, 7, 13, 15, 3, -6, -9,
					-- layer=2 filter=207 channel=71
					-17, -6, 0, 4, -6, -7, 4, 2, -19,
					-- layer=2 filter=207 channel=72
					-1, -6, -1, -13, -9, -10, 12, -8, -7,
					-- layer=2 filter=207 channel=73
					-7, -1, 4, -8, -12, -3, -14, -8, -12,
					-- layer=2 filter=207 channel=74
					1, -5, -15, 4, 0, -7, -3, -16, -4,
					-- layer=2 filter=207 channel=75
					5, -22, 10, 1, 2, -15, -17, -12, 3,
					-- layer=2 filter=207 channel=76
					-4, -18, 10, -9, -15, 1, 3, 1, 4,
					-- layer=2 filter=207 channel=77
					-4, -1, 1, -3, 3, -5, 9, 8, -10,
					-- layer=2 filter=207 channel=78
					-2, -17, -8, -15, -10, -8, -14, -9, -11,
					-- layer=2 filter=207 channel=79
					4, 3, -2, -2, -7, -6, -7, 6, 6,
					-- layer=2 filter=207 channel=80
					-2, -12, -3, 0, -5, -18, -13, 0, -18,
					-- layer=2 filter=207 channel=81
					4, -4, 0, -14, -5, -6, -14, 1, -2,
					-- layer=2 filter=207 channel=82
					2, -7, -2, -12, -8, -11, 8, 3, -11,
					-- layer=2 filter=207 channel=83
					-8, 3, -10, -10, -9, -1, 0, 4, -10,
					-- layer=2 filter=207 channel=84
					-2, 6, -2, -8, -1, 11, -7, 9, -1,
					-- layer=2 filter=207 channel=85
					-4, 6, 4, -8, 7, -12, -3, -10, -5,
					-- layer=2 filter=207 channel=86
					-1, -4, 6, 6, 9, 7, 5, 6, -4,
					-- layer=2 filter=207 channel=87
					-4, -13, 1, 0, -4, -3, -17, 1, -4,
					-- layer=2 filter=207 channel=88
					0, 0, -17, -12, -13, -7, -5, 0, 0,
					-- layer=2 filter=207 channel=89
					5, -4, -2, -27, -25, -16, -15, -9, -6,
					-- layer=2 filter=207 channel=90
					2, 7, -5, 2, 0, 2, -5, -1, -4,
					-- layer=2 filter=207 channel=91
					0, -8, -12, -28, -15, -5, -4, 6, 1,
					-- layer=2 filter=207 channel=92
					-5, -3, 2, -29, -24, -22, -11, -1, -14,
					-- layer=2 filter=207 channel=93
					-8, -14, -4, -5, -3, -4, 2, -3, -7,
					-- layer=2 filter=207 channel=94
					0, -5, 5, 13, 3, 0, 2, -6, 2,
					-- layer=2 filter=207 channel=95
					4, 6, -9, -2, 0, 9, 8, 5, 2,
					-- layer=2 filter=207 channel=96
					-1, -7, 10, -1, 2, -4, -13, 10, 4,
					-- layer=2 filter=207 channel=97
					-7, -8, -4, -18, -11, -4, -16, -17, -15,
					-- layer=2 filter=207 channel=98
					-12, -4, -5, -6, 3, 10, 2, -12, 0,
					-- layer=2 filter=207 channel=99
					-11, -4, 11, -2, 0, 2, 13, 4, -5,
					-- layer=2 filter=207 channel=100
					4, -11, 1, -13, 0, -13, -15, 0, 0,
					-- layer=2 filter=207 channel=101
					2, 2, -15, 7, -2, -4, -2, -5, -19,
					-- layer=2 filter=207 channel=102
					3, -1, -5, 0, 3, 0, -13, 12, 1,
					-- layer=2 filter=207 channel=103
					-9, -7, -9, -11, 6, -11, 4, -9, 3,
					-- layer=2 filter=207 channel=104
					-17, -16, 9, 6, -5, -7, -6, 10, -2,
					-- layer=2 filter=207 channel=105
					6, 0, 1, -3, -4, -6, -18, -2, -7,
					-- layer=2 filter=207 channel=106
					7, -20, -3, -12, -17, -8, -13, -5, -9,
					-- layer=2 filter=207 channel=107
					-10, -5, -17, -18, -8, -10, -2, -1, 1,
					-- layer=2 filter=207 channel=108
					-10, 2, 2, 0, 9, -18, -13, -8, -7,
					-- layer=2 filter=207 channel=109
					-5, 7, -7, 3, -10, 7, 6, 6, -10,
					-- layer=2 filter=207 channel=110
					2, -6, -18, -2, -22, -14, -11, 0, -6,
					-- layer=2 filter=207 channel=111
					7, 4, 8, 2, 1, -5, 0, -4, 1,
					-- layer=2 filter=207 channel=112
					1, -15, -3, -2, -1, -7, -8, -1, -17,
					-- layer=2 filter=207 channel=113
					-10, -10, -20, 4, -4, -9, -5, -17, -6,
					-- layer=2 filter=207 channel=114
					-5, 7, -1, 5, 6, -5, -6, -5, -4,
					-- layer=2 filter=207 channel=115
					-10, 7, 0, -7, -5, 5, -7, 7, -2,
					-- layer=2 filter=207 channel=116
					1, -10, 10, 9, 1, -5, 4, 15, 13,
					-- layer=2 filter=207 channel=117
					3, 4, -2, -9, -17, -1, -3, 0, -3,
					-- layer=2 filter=207 channel=118
					-16, -14, -5, -3, -1, -9, -4, -10, 0,
					-- layer=2 filter=207 channel=119
					7, -8, 4, -10, -12, -9, -6, -4, -2,
					-- layer=2 filter=207 channel=120
					3, 2, 9, -8, 0, -7, -4, -8, -3,
					-- layer=2 filter=207 channel=121
					-4, 0, -1, -6, 4, 1, -1, -8, 4,
					-- layer=2 filter=207 channel=122
					1, 5, -4, 6, -5, 5, 2, 8, 5,
					-- layer=2 filter=207 channel=123
					5, -6, -7, -16, -15, 0, 14, 7, 1,
					-- layer=2 filter=207 channel=124
					-4, -10, -11, -10, -13, 9, -3, 0, 2,
					-- layer=2 filter=207 channel=125
					-1, -10, 4, 0, 9, 0, -3, -2, 9,
					-- layer=2 filter=207 channel=126
					4, 6, 2, -3, -1, -7, 1, 4, -11,
					-- layer=2 filter=207 channel=127
					-5, 9, -15, -6, -3, -20, 0, 7, 6,
					-- layer=2 filter=208 channel=0
					1, 16, 15, -13, 14, 17, -17, 10, 14,
					-- layer=2 filter=208 channel=1
					-23, -20, -1, -38, -20, -7, -34, -24, -8,
					-- layer=2 filter=208 channel=2
					2, 8, 0, 2, -2, 0, 0, -5, -3,
					-- layer=2 filter=208 channel=3
					4, 25, 26, 19, -3, -5, -19, -20, -3,
					-- layer=2 filter=208 channel=4
					3, -36, -2, -3, -20, 1, 2, -18, -2,
					-- layer=2 filter=208 channel=5
					7, 24, 11, 0, 19, 10, 2, 2, 19,
					-- layer=2 filter=208 channel=6
					27, -1, -21, -21, 39, -4, 8, 2, -3,
					-- layer=2 filter=208 channel=7
					12, 4, -4, 7, -43, 3, -14, -49, -25,
					-- layer=2 filter=208 channel=8
					9, -5, 4, -10, 1, 4, 4, 10, 9,
					-- layer=2 filter=208 channel=9
					3, 27, 13, 17, -2, 23, -11, 7, -15,
					-- layer=2 filter=208 channel=10
					3, 19, 28, 14, 17, 28, -3, -10, -8,
					-- layer=2 filter=208 channel=11
					10, 23, -1, 9, 4, 3, 14, 33, 9,
					-- layer=2 filter=208 channel=12
					4, -56, -3, -23, -6, -25, -20, -18, -28,
					-- layer=2 filter=208 channel=13
					-2, -7, -3, -4, -5, 9, 3, 4, 11,
					-- layer=2 filter=208 channel=14
					-10, -27, -7, 12, -4, 19, 20, -8, -6,
					-- layer=2 filter=208 channel=15
					17, 7, 16, -24, -5, -34, 25, 32, -4,
					-- layer=2 filter=208 channel=16
					-4, -7, 18, -7, 4, -1, -18, -41, -19,
					-- layer=2 filter=208 channel=17
					1, 0, 9, 6, 0, 5, -9, -10, 5,
					-- layer=2 filter=208 channel=18
					35, 49, 33, 10, 15, -3, 7, 31, 12,
					-- layer=2 filter=208 channel=19
					5, -6, 6, -6, -18, -19, -38, -35, -38,
					-- layer=2 filter=208 channel=20
					-1, -7, 4, 10, -2, 9, -8, 7, -7,
					-- layer=2 filter=208 channel=21
					-1, -8, -3, -4, 0, -7, 3, -12, 9,
					-- layer=2 filter=208 channel=22
					-5, 1, 5, -5, 6, -9, -6, 8, -6,
					-- layer=2 filter=208 channel=23
					-2, -22, 11, -11, -46, -25, -21, -11, -20,
					-- layer=2 filter=208 channel=24
					24, 1, 18, 19, 11, 13, 9, -8, -12,
					-- layer=2 filter=208 channel=25
					5, -5, 0, -1, 5, -11, 0, 8, -4,
					-- layer=2 filter=208 channel=26
					12, -8, -7, -1, 7, -5, 10, -5, -1,
					-- layer=2 filter=208 channel=27
					-12, 7, 9, 9, 19, 40, 0, 20, 45,
					-- layer=2 filter=208 channel=28
					-15, -14, -43, 22, 10, -8, 1, 28, 1,
					-- layer=2 filter=208 channel=29
					-8, 9, -1, 1, 2, -5, 1, 2, -6,
					-- layer=2 filter=208 channel=30
					-11, 23, 30, -13, -25, -7, -20, -14, -22,
					-- layer=2 filter=208 channel=31
					13, 4, 29, -39, 47, -19, 23, 21, -7,
					-- layer=2 filter=208 channel=32
					-9, 5, 6, -5, 2, 4, -2, -12, -5,
					-- layer=2 filter=208 channel=33
					0, -46, -57, 33, 10, 17, -2, -21, -19,
					-- layer=2 filter=208 channel=34
					-18, 5, -19, -10, 27, 2, -40, 8, 31,
					-- layer=2 filter=208 channel=35
					7, -10, -8, 18, 16, -1, -12, 1, 16,
					-- layer=2 filter=208 channel=36
					9, -12, -6, 1, 4, -12, -9, 6, 9,
					-- layer=2 filter=208 channel=37
					7, 12, -10, -14, 25, -1, 2, 19, 13,
					-- layer=2 filter=208 channel=38
					-13, 9, -18, -29, 18, -11, 16, -12, 26,
					-- layer=2 filter=208 channel=39
					0, -15, -15, -10, -45, 8, -38, -32, -35,
					-- layer=2 filter=208 channel=40
					19, -1, -7, -35, -12, 48, -23, 48, -13,
					-- layer=2 filter=208 channel=41
					8, -2, -6, 6, 8, -9, 7, 1, -5,
					-- layer=2 filter=208 channel=42
					26, -19, 9, -6, -32, -18, 2, 9, -18,
					-- layer=2 filter=208 channel=43
					28, 18, 33, -20, 21, -42, -28, -29, 1,
					-- layer=2 filter=208 channel=44
					-9, 0, -5, -3, -1, -6, 6, -8, -2,
					-- layer=2 filter=208 channel=45
					40, 7, 7, 14, -23, -18, 21, -40, -4,
					-- layer=2 filter=208 channel=46
					-17, 16, 22, -10, 18, 12, -21, -21, -25,
					-- layer=2 filter=208 channel=47
					-5, -29, -53, 14, -11, -6, 24, -13, -45,
					-- layer=2 filter=208 channel=48
					6, 2, -5, 0, -4, 1, 3, 3, -1,
					-- layer=2 filter=208 channel=49
					27, 44, 61, -2, 36, 19, -5, 18, -8,
					-- layer=2 filter=208 channel=50
					13, 12, -12, 7, 3, 15, -14, 17, 14,
					-- layer=2 filter=208 channel=51
					3, 16, -15, -11, 14, 1, 1, 23, 29,
					-- layer=2 filter=208 channel=52
					7, 2, -32, -15, -26, 26, 4, 16, -3,
					-- layer=2 filter=208 channel=53
					22, 4, 27, -8, -18, 0, -21, -15, 1,
					-- layer=2 filter=208 channel=54
					-21, -14, -30, 0, -1, -14, 18, 26, 9,
					-- layer=2 filter=208 channel=55
					-10, -6, -2, 2, -5, -8, 11, -7, 4,
					-- layer=2 filter=208 channel=56
					8, 16, 2, 11, 16, 15, 0, 12, 21,
					-- layer=2 filter=208 channel=57
					9, 8, -4, 2, -7, 4, 7, 4, 3,
					-- layer=2 filter=208 channel=58
					30, -41, -13, -24, -11, -27, 18, -24, -24,
					-- layer=2 filter=208 channel=59
					19, -1, -35, -22, -19, 13, -9, 1, -21,
					-- layer=2 filter=208 channel=60
					-47, -18, -31, -69, 4, -4, -3, -3, -6,
					-- layer=2 filter=208 channel=61
					17, 30, 35, -10, 36, 0, -24, 23, 11,
					-- layer=2 filter=208 channel=62
					-29, -8, -35, -13, 10, -36, -24, 16, 19,
					-- layer=2 filter=208 channel=63
					-17, -24, 4, -42, -31, -21, -22, 2, -20,
					-- layer=2 filter=208 channel=64
					21, 1, 24, 32, -1, -2, 5, -20, 9,
					-- layer=2 filter=208 channel=65
					0, 11, 10, 11, 36, 31, 16, 15, 27,
					-- layer=2 filter=208 channel=66
					17, -59, -31, -5, -4, -8, 16, 3, -12,
					-- layer=2 filter=208 channel=67
					-25, -12, 16, -42, 3, 10, -33, -31, -25,
					-- layer=2 filter=208 channel=68
					-4, -5, -1, -5, 2, 4, 2, -4, 6,
					-- layer=2 filter=208 channel=69
					-1, -3, 6, 25, 19, 14, 8, -15, 1,
					-- layer=2 filter=208 channel=70
					5, -2, -24, 13, 0, 29, 10, 4, 22,
					-- layer=2 filter=208 channel=71
					-13, 1, 0, -1, 13, 29, -12, 0, 9,
					-- layer=2 filter=208 channel=72
					-20, -35, -31, 42, 11, -1, 24, 18, 3,
					-- layer=2 filter=208 channel=73
					39, 58, 32, 5, 44, -8, 10, -11, -8,
					-- layer=2 filter=208 channel=74
					-25, -19, 10, -26, -10, -11, -9, -23, -12,
					-- layer=2 filter=208 channel=75
					10, -60, -73, -35, -53, -13, -12, -41, -44,
					-- layer=2 filter=208 channel=76
					52, 21, 24, -47, 9, -39, -29, 4, -36,
					-- layer=2 filter=208 channel=77
					-4, 9, 6, 7, 7, 1, 3, 9, 0,
					-- layer=2 filter=208 channel=78
					4, 8, -17, 5, 5, -16, 4, 13, 1,
					-- layer=2 filter=208 channel=79
					5, 1, -9, -5, 1, 2, 4, 9, -5,
					-- layer=2 filter=208 channel=80
					12, 9, 18, 3, 0, -4, -29, -25, -13,
					-- layer=2 filter=208 channel=81
					-3, 0, -10, -9, -3, 7, 0, -8, -2,
					-- layer=2 filter=208 channel=82
					-8, 3, 2, 5, 3, 10, 0, -2, -8,
					-- layer=2 filter=208 channel=83
					-11, -26, 15, 0, -29, 0, -9, -28, -14,
					-- layer=2 filter=208 channel=84
					2, 10, 6, 2, 4, 5, 3, 11, -3,
					-- layer=2 filter=208 channel=85
					3, 11, -6, -2, 6, -2, -12, 5, 4,
					-- layer=2 filter=208 channel=86
					-15, -2, 4, -12, -12, -5, -6, -8, -6,
					-- layer=2 filter=208 channel=87
					48, -16, -10, 1, 7, 42, -18, 47, 16,
					-- layer=2 filter=208 channel=88
					-25, -40, 8, -2, 6, -21, -15, -7, 6,
					-- layer=2 filter=208 channel=89
					16, -34, -34, 0, -5, -19, 0, -10, -26,
					-- layer=2 filter=208 channel=90
					0, 7, 4, 1, -11, 0, -6, 6, -2,
					-- layer=2 filter=208 channel=91
					-8, -46, -74, -18, -40, -32, -15, -45, -39,
					-- layer=2 filter=208 channel=92
					-23, -32, -19, -4, -1, 4, -28, -6, 3,
					-- layer=2 filter=208 channel=93
					30, 0, 27, 0, -10, 0, -47, -52, -35,
					-- layer=2 filter=208 channel=94
					14, 16, 32, -40, -13, -2, -57, -7, -33,
					-- layer=2 filter=208 channel=95
					8, -3, -7, 0, 9, -3, -4, 7, 7,
					-- layer=2 filter=208 channel=96
					-33, 2, 5, -10, 30, 23, 13, 26, 5,
					-- layer=2 filter=208 channel=97
					4, 5, 18, 25, 12, -1, 28, 16, -5,
					-- layer=2 filter=208 channel=98
					12, -12, -8, 36, -3, 20, 17, 35, -2,
					-- layer=2 filter=208 channel=99
					-6, -2, -6, -15, -14, 2, -10, -2, -29,
					-- layer=2 filter=208 channel=100
					2, -10, 10, -33, 16, 17, 17, -15, -15,
					-- layer=2 filter=208 channel=101
					-14, -12, 10, 18, -3, 18, -8, -8, -40,
					-- layer=2 filter=208 channel=102
					-2, 21, 17, 5, 20, 23, 7, 13, -8,
					-- layer=2 filter=208 channel=103
					18, -21, -55, -68, 6, 44, -5, -5, -13,
					-- layer=2 filter=208 channel=104
					13, 24, 19, 17, 15, 30, -39, 24, 18,
					-- layer=2 filter=208 channel=105
					-5, 43, 11, -8, -20, -5, 10, -20, -33,
					-- layer=2 filter=208 channel=106
					4, -18, 11, 10, -4, -9, 9, -4, -24,
					-- layer=2 filter=208 channel=107
					7, 16, 11, -23, 29, -9, -37, 6, 41,
					-- layer=2 filter=208 channel=108
					-35, -6, 22, -14, 10, 12, -15, -18, -12,
					-- layer=2 filter=208 channel=109
					1, -12, 12, 4, 1, 1, -2, -2, -16,
					-- layer=2 filter=208 channel=110
					-4, -29, 7, 10, -5, -20, 2, -10, -24,
					-- layer=2 filter=208 channel=111
					-2, -8, -10, -4, -6, -7, -1, 9, -6,
					-- layer=2 filter=208 channel=112
					20, 13, 17, 0, 28, 11, -19, 14, 26,
					-- layer=2 filter=208 channel=113
					2, 6, 35, 8, -18, 18, -29, 0, 12,
					-- layer=2 filter=208 channel=114
					-10, -11, -3, -13, -9, -14, -10, -13, -3,
					-- layer=2 filter=208 channel=115
					0, 10, -8, -2, -11, -5, 1, 1, 4,
					-- layer=2 filter=208 channel=116
					11, 11, -5, -10, -3, 0, -31, 36, 4,
					-- layer=2 filter=208 channel=117
					16, 34, 31, -6, -28, -4, -26, -32, -7,
					-- layer=2 filter=208 channel=118
					16, 25, 25, -3, 5, -2, -12, 14, -13,
					-- layer=2 filter=208 channel=119
					12, -2, -6, -11, 7, -11, 12, -11, 23,
					-- layer=2 filter=208 channel=120
					0, -1, 3, -1, -4, 2, 0, -1, 8,
					-- layer=2 filter=208 channel=121
					-9, 0, 7, 3, 2, -11, 5, -5, 5,
					-- layer=2 filter=208 channel=122
					5, 0, -2, -6, -4, 11, 4, 6, -6,
					-- layer=2 filter=208 channel=123
					6, -37, -41, 10, -35, -8, -4, -16, -22,
					-- layer=2 filter=208 channel=124
					35, -21, 25, 8, 16, -45, 6, 10, -28,
					-- layer=2 filter=208 channel=125
					6, -10, 1, -12, -3, 2, 10, -2, 6,
					-- layer=2 filter=208 channel=126
					-44, 12, 8, -29, -21, -56, -20, 4, -24,
					-- layer=2 filter=208 channel=127
					-2, -29, -2, -1, -8, -9, -39, -18, 11,
					-- layer=2 filter=209 channel=0
					-10, 5, 0, 0, -4, 6, -4, 8, -7,
					-- layer=2 filter=209 channel=1
					-15, -6, 8, -9, -11, -6, -7, -16, -20,
					-- layer=2 filter=209 channel=2
					5, -1, -9, -3, 6, 3, 4, 5, -11,
					-- layer=2 filter=209 channel=3
					5, 3, -9, 0, -11, 0, -4, 0, 0,
					-- layer=2 filter=209 channel=4
					-12, -7, -6, 0, -14, -3, -3, 0, 2,
					-- layer=2 filter=209 channel=5
					-2, -3, -10, 5, -2, -4, -5, -4, 0,
					-- layer=2 filter=209 channel=6
					1, 7, -7, -13, -3, 0, 3, -6, -2,
					-- layer=2 filter=209 channel=7
					-3, 4, 7, 1, 6, -13, 1, -6, 0,
					-- layer=2 filter=209 channel=8
					-5, 0, 2, -2, 2, 8, -7, -4, -3,
					-- layer=2 filter=209 channel=9
					1, 2, -2, 3, -4, 7, 1, -9, -7,
					-- layer=2 filter=209 channel=10
					-6, -4, 0, 0, -3, 6, 0, -11, -1,
					-- layer=2 filter=209 channel=11
					2, -18, -2, 1, -15, 0, -17, -5, -18,
					-- layer=2 filter=209 channel=12
					-5, 4, 0, -5, -4, -13, -7, -7, -11,
					-- layer=2 filter=209 channel=13
					0, 0, 8, -10, 8, -4, 8, 3, -2,
					-- layer=2 filter=209 channel=14
					-8, -8, 4, -9, -8, 0, -6, -9, 1,
					-- layer=2 filter=209 channel=15
					3, -12, 0, -9, -13, -2, -4, -12, 0,
					-- layer=2 filter=209 channel=16
					-9, -10, -4, -3, -1, -6, 4, -1, -2,
					-- layer=2 filter=209 channel=17
					4, -9, 3, 8, 4, 7, -7, -3, -4,
					-- layer=2 filter=209 channel=18
					1, -1, -7, 10, 5, 7, -1, -5, -12,
					-- layer=2 filter=209 channel=19
					-10, -1, -11, 0, 3, -12, -17, -4, -1,
					-- layer=2 filter=209 channel=20
					8, -5, 7, -11, 0, -11, 4, -3, 6,
					-- layer=2 filter=209 channel=21
					7, 1, -10, -4, -9, 1, 4, 6, -7,
					-- layer=2 filter=209 channel=22
					4, -9, -9, -7, -9, 2, 1, -8, 7,
					-- layer=2 filter=209 channel=23
					-2, 0, -7, -14, -15, -12, -1, -3, 0,
					-- layer=2 filter=209 channel=24
					3, -4, -9, 0, -11, -3, -2, 4, -12,
					-- layer=2 filter=209 channel=25
					-6, -10, -11, -4, 0, -12, 4, 0, -3,
					-- layer=2 filter=209 channel=26
					-3, 0, 6, 10, 4, -5, -9, 8, -1,
					-- layer=2 filter=209 channel=27
					-7, 7, 4, -8, -4, -3, -15, -7, 2,
					-- layer=2 filter=209 channel=28
					-11, -4, -5, -11, 2, 2, 2, -11, -10,
					-- layer=2 filter=209 channel=29
					-12, -4, 3, -3, -10, 2, -9, -2, 5,
					-- layer=2 filter=209 channel=30
					-3, -9, -17, 8, -10, -6, -2, 0, 7,
					-- layer=2 filter=209 channel=31
					-7, -8, 0, 1, 0, -2, 1, 0, -11,
					-- layer=2 filter=209 channel=32
					0, -4, 6, -10, -9, 7, 4, 1, 2,
					-- layer=2 filter=209 channel=33
					-14, -9, 8, -14, -12, -2, -13, -6, -6,
					-- layer=2 filter=209 channel=34
					-3, 2, -14, -4, -8, -1, -1, -12, -12,
					-- layer=2 filter=209 channel=35
					-8, -9, -9, 2, -12, 4, -12, 0, 3,
					-- layer=2 filter=209 channel=36
					-3, -1, -11, 8, -4, -8, 7, -4, 8,
					-- layer=2 filter=209 channel=37
					-8, 4, -2, -3, -12, -12, -1, -5, -14,
					-- layer=2 filter=209 channel=38
					-1, 10, -10, -6, 10, -1, -15, -6, 0,
					-- layer=2 filter=209 channel=39
					-2, -1, 2, -10, 0, -2, -7, 0, -4,
					-- layer=2 filter=209 channel=40
					-14, -6, 0, -11, 4, -11, -9, -11, 0,
					-- layer=2 filter=209 channel=41
					4, 8, -8, -10, 4, 3, 7, -3, 7,
					-- layer=2 filter=209 channel=42
					0, -1, 7, -11, -5, 9, 2, -14, -5,
					-- layer=2 filter=209 channel=43
					1, -12, 6, -8, -10, -4, 5, -13, -2,
					-- layer=2 filter=209 channel=44
					2, 3, 9, 4, 0, -5, 1, -5, 2,
					-- layer=2 filter=209 channel=45
					-3, -6, -10, 3, -3, -11, -14, -7, 5,
					-- layer=2 filter=209 channel=46
					9, 5, -8, 2, -4, 0, -7, 8, -11,
					-- layer=2 filter=209 channel=47
					-11, 0, 0, -10, -1, 4, -11, -1, 1,
					-- layer=2 filter=209 channel=48
					10, 1, 0, 0, 5, 4, -4, 4, -3,
					-- layer=2 filter=209 channel=49
					-4, -13, -9, -2, 2, 10, 6, -3, -12,
					-- layer=2 filter=209 channel=50
					-1, -2, 0, 9, -8, 7, -9, 9, -8,
					-- layer=2 filter=209 channel=51
					-6, -12, -13, -3, 3, 3, 2, -12, -9,
					-- layer=2 filter=209 channel=52
					-15, -6, -21, -14, -5, 1, 0, -2, -14,
					-- layer=2 filter=209 channel=53
					-6, 4, -13, -2, 5, -5, 6, -2, 0,
					-- layer=2 filter=209 channel=54
					0, -6, -8, -3, -9, 3, -4, -3, -20,
					-- layer=2 filter=209 channel=55
					-9, 3, 7, -2, 1, -1, -9, 0, 3,
					-- layer=2 filter=209 channel=56
					-14, -5, -11, -15, -3, -10, -2, -9, -12,
					-- layer=2 filter=209 channel=57
					-10, 4, -8, 2, 1, -8, -11, -6, -5,
					-- layer=2 filter=209 channel=58
					4, -14, 3, -5, -5, -7, -17, -16, -16,
					-- layer=2 filter=209 channel=59
					2, -11, -9, -5, 1, -8, -6, -9, -3,
					-- layer=2 filter=209 channel=60
					-13, 14, -10, -10, 3, -19, -13, -5, -11,
					-- layer=2 filter=209 channel=61
					-9, 8, -13, -11, 2, -11, -15, 4, 4,
					-- layer=2 filter=209 channel=62
					0, 5, -8, 5, 6, -2, -4, 0, -2,
					-- layer=2 filter=209 channel=63
					-1, 3, 1, -9, 0, -4, -8, 1, 2,
					-- layer=2 filter=209 channel=64
					0, 3, -13, -6, -5, 4, -8, -3, -12,
					-- layer=2 filter=209 channel=65
					-1, -2, -3, 0, -8, -12, -8, -4, -13,
					-- layer=2 filter=209 channel=66
					-10, -9, 0, 0, 5, -1, -5, 5, 8,
					-- layer=2 filter=209 channel=67
					0, -8, 1, 10, -4, 0, -1, 3, 6,
					-- layer=2 filter=209 channel=68
					4, 3, -11, 0, 7, -4, -5, -11, 5,
					-- layer=2 filter=209 channel=69
					4, -2, -2, -5, 1, -3, 5, -3, 5,
					-- layer=2 filter=209 channel=70
					0, -12, -9, -6, -2, 3, 7, -7, -6,
					-- layer=2 filter=209 channel=71
					-14, 16, 0, -3, -6, 0, -6, -2, -13,
					-- layer=2 filter=209 channel=72
					-1, 6, 0, 3, -12, -5, -8, -13, -1,
					-- layer=2 filter=209 channel=73
					-11, -7, -16, -16, 4, 0, -13, 0, 6,
					-- layer=2 filter=209 channel=74
					-3, 4, -1, -1, -10, -8, 6, 0, -2,
					-- layer=2 filter=209 channel=75
					-9, -13, -10, -3, -12, -7, 0, 1, -5,
					-- layer=2 filter=209 channel=76
					-3, -8, -16, 0, -10, -16, 5, 0, 5,
					-- layer=2 filter=209 channel=77
					5, 8, 6, -12, 1, 0, 4, 3, -11,
					-- layer=2 filter=209 channel=78
					-2, 0, -4, -4, -8, -6, 7, 3, -9,
					-- layer=2 filter=209 channel=79
					0, 4, -5, 7, 0, 0, -7, -2, -6,
					-- layer=2 filter=209 channel=80
					5, -12, -6, 1, -7, 5, 8, -11, -2,
					-- layer=2 filter=209 channel=81
					-2, -1, -12, -2, 6, -7, 0, -6, 5,
					-- layer=2 filter=209 channel=82
					-8, 2, -3, 8, -3, 4, 3, -7, 3,
					-- layer=2 filter=209 channel=83
					-6, -10, -7, -7, 3, -2, -2, -7, 0,
					-- layer=2 filter=209 channel=84
					-4, 3, 5, 4, 6, -8, -6, 3, 8,
					-- layer=2 filter=209 channel=85
					-6, 10, 0, 3, -6, -9, 9, 5, 10,
					-- layer=2 filter=209 channel=86
					-2, 8, 4, 1, 10, -2, 0, -1, -9,
					-- layer=2 filter=209 channel=87
					-3, -15, 0, 0, 2, -6, -10, 1, -6,
					-- layer=2 filter=209 channel=88
					-10, -19, -15, 1, 7, -12, -11, 3, 2,
					-- layer=2 filter=209 channel=89
					-8, -2, -2, -1, -22, -6, -18, -10, -12,
					-- layer=2 filter=209 channel=90
					-7, 7, 7, 4, -10, 5, 3, 10, 0,
					-- layer=2 filter=209 channel=91
					-3, -12, -4, -17, -7, -4, -2, -11, -6,
					-- layer=2 filter=209 channel=92
					-11, 3, -1, -6, -20, -5, -12, -1, -3,
					-- layer=2 filter=209 channel=93
					-15, 5, 2, -13, 10, -15, -6, 10, -16,
					-- layer=2 filter=209 channel=94
					-6, 4, 2, -19, -12, -5, -7, -12, -13,
					-- layer=2 filter=209 channel=95
					5, -9, 5, -4, -1, -10, 6, -1, -2,
					-- layer=2 filter=209 channel=96
					-14, 1, 5, -9, -8, -18, 0, -4, -3,
					-- layer=2 filter=209 channel=97
					3, -8, -6, -5, -3, 1, 7, -9, -4,
					-- layer=2 filter=209 channel=98
					-17, -11, -7, -1, -3, -3, -7, -15, -3,
					-- layer=2 filter=209 channel=99
					-12, -6, -17, 0, -7, -12, -21, -7, -3,
					-- layer=2 filter=209 channel=100
					2, 3, -3, 0, 1, -9, 8, 5, -12,
					-- layer=2 filter=209 channel=101
					-14, 6, -4, 0, 1, 0, 0, 0, -5,
					-- layer=2 filter=209 channel=102
					-20, -12, 3, -7, 1, -17, 0, -15, 10,
					-- layer=2 filter=209 channel=103
					2, 6, 5, 7, -10, -8, 6, 3, -7,
					-- layer=2 filter=209 channel=104
					-1, -1, -5, -11, 0, -2, 10, -12, 1,
					-- layer=2 filter=209 channel=105
					-7, -4, 4, -15, -8, 13, 7, -4, 0,
					-- layer=2 filter=209 channel=106
					0, -10, 0, -6, -10, -4, -13, -8, 0,
					-- layer=2 filter=209 channel=107
					-4, 9, 5, 8, -8, 8, 0, 5, -2,
					-- layer=2 filter=209 channel=108
					-1, 4, -6, 2, 0, 0, -8, -5, -12,
					-- layer=2 filter=209 channel=109
					0, -5, -3, -6, -10, -12, -8, 5, -5,
					-- layer=2 filter=209 channel=110
					-5, 2, 0, -16, 3, 2, -11, -10, -6,
					-- layer=2 filter=209 channel=111
					-6, -7, 0, -4, -11, -5, -11, 8, 3,
					-- layer=2 filter=209 channel=112
					-15, 6, -4, -5, 7, -3, -7, -6, -9,
					-- layer=2 filter=209 channel=113
					-7, 0, -4, -3, -8, -1, 6, 4, 0,
					-- layer=2 filter=209 channel=114
					-1, 10, -7, 8, -2, -7, 0, 2, -6,
					-- layer=2 filter=209 channel=115
					-5, 9, -2, -8, -9, 1, 0, 1, -8,
					-- layer=2 filter=209 channel=116
					-7, 0, -13, 4, -2, 4, -13, -16, -2,
					-- layer=2 filter=209 channel=117
					-10, -3, -5, -14, -5, -3, -14, -19, -1,
					-- layer=2 filter=209 channel=118
					4, -15, 0, 1, 0, 7, -9, -2, -12,
					-- layer=2 filter=209 channel=119
					-7, -10, -5, -12, -9, -6, -11, -4, -10,
					-- layer=2 filter=209 channel=120
					-3, -8, 6, 9, 0, -8, -3, -10, 7,
					-- layer=2 filter=209 channel=121
					-6, 0, -3, -8, -9, 0, -2, 7, -5,
					-- layer=2 filter=209 channel=122
					2, -2, 6, -7, -6, -9, 4, -1, 0,
					-- layer=2 filter=209 channel=123
					-10, -11, -3, 0, -15, -12, -7, -3, 9,
					-- layer=2 filter=209 channel=124
					-15, -11, -8, 0, -5, -13, -12, -15, -9,
					-- layer=2 filter=209 channel=125
					-2, -9, 8, 2, 6, -10, -7, 8, -8,
					-- layer=2 filter=209 channel=126
					-9, 2, 5, 5, -1, 7, -10, -9, -3,
					-- layer=2 filter=209 channel=127
					-7, -10, 6, -12, 0, 0, 1, -9, -17,
					-- layer=2 filter=210 channel=0
					-31, -18, -19, -69, -59, -25, -48, -47, -61,
					-- layer=2 filter=210 channel=1
					11, 12, -5, 29, -1, -48, -11, 4, -26,
					-- layer=2 filter=210 channel=2
					1, -8, 7, 8, -9, 6, -9, -5, -3,
					-- layer=2 filter=210 channel=3
					-37, -45, -8, -58, -73, -11, -20, 10, 6,
					-- layer=2 filter=210 channel=4
					17, -50, 9, 39, -16, -30, 7, 1, -15,
					-- layer=2 filter=210 channel=5
					-7, -10, -30, -47, -45, -16, -27, -30, -30,
					-- layer=2 filter=210 channel=6
					-67, 17, -8, 5, 35, -64, -20, 26, 35,
					-- layer=2 filter=210 channel=7
					-89, -19, -11, 37, -22, 32, -23, 9, 36,
					-- layer=2 filter=210 channel=8
					-6, -2, 8, 7, 1, -1, 1, 1, 5,
					-- layer=2 filter=210 channel=9
					-7, -37, -58, -40, -56, -4, -55, 6, -10,
					-- layer=2 filter=210 channel=10
					-17, -51, -9, -63, -59, -18, -58, -40, -21,
					-- layer=2 filter=210 channel=11
					-5, -41, -25, -24, -1, -12, -13, 7, -11,
					-- layer=2 filter=210 channel=12
					15, 20, -5, -8, -30, -70, 2, -8, -25,
					-- layer=2 filter=210 channel=13
					-2, 0, 1, 4, 5, 2, 3, 1, 2,
					-- layer=2 filter=210 channel=14
					-3, -15, -8, 1, -19, -41, -11, -9, -32,
					-- layer=2 filter=210 channel=15
					29, 27, 29, 25, 56, 23, 14, 27, 25,
					-- layer=2 filter=210 channel=16
					-107, -81, -31, 23, 1, 55, -10, 8, 18,
					-- layer=2 filter=210 channel=17
					7, -6, 5, -9, 5, -5, 9, 0, -2,
					-- layer=2 filter=210 channel=18
					-11, -77, 34, -7, -5, -3, 18, 36, 3,
					-- layer=2 filter=210 channel=19
					29, 27, 23, 47, 30, -22, 20, 4, -15,
					-- layer=2 filter=210 channel=20
					9, -4, 7, -4, -3, -1, 9, 7, -3,
					-- layer=2 filter=210 channel=21
					-29, -1, -6, -21, -9, -2, -14, -9, -9,
					-- layer=2 filter=210 channel=22
					11, 3, 6, 6, 0, -3, 5, 7, -4,
					-- layer=2 filter=210 channel=23
					-40, -59, -14, -16, 0, -7, 8, 52, 44,
					-- layer=2 filter=210 channel=24
					-67, -65, -28, -74, -27, 1, -38, -1, 36,
					-- layer=2 filter=210 channel=25
					-55, -20, -15, 0, -8, -6, -5, 20, 12,
					-- layer=2 filter=210 channel=26
					10, 0, 9, 4, -7, -5, -5, 1, -2,
					-- layer=2 filter=210 channel=27
					44, 42, -1, 34, -5, -50, 13, -23, -30,
					-- layer=2 filter=210 channel=28
					-45, -43, 32, -10, -18, 19, -23, -11, -76,
					-- layer=2 filter=210 channel=29
					3, -4, 1, 3, 7, -1, 6, 4, -3,
					-- layer=2 filter=210 channel=30
					33, -13, -32, -1, -17, -28, -20, -33, 2,
					-- layer=2 filter=210 channel=31
					26, 2, 22, 0, 18, 35, 15, -6, 49,
					-- layer=2 filter=210 channel=32
					6, 9, 5, 1, 8, -9, -1, -1, -1,
					-- layer=2 filter=210 channel=33
					-33, -7, 12, 7, -24, 5, 33, -47, 3,
					-- layer=2 filter=210 channel=34
					-14, -48, 29, 15, 17, 32, -5, -5, -18,
					-- layer=2 filter=210 channel=35
					12, 7, 18, 3, 9, 18, 33, -14, -17,
					-- layer=2 filter=210 channel=36
					-9, 1, -1, 6, -1, 4, 3, 6, -3,
					-- layer=2 filter=210 channel=37
					14, 2, -23, -6, 0, -29, -3, -6, -11,
					-- layer=2 filter=210 channel=38
					35, 8, -11, 5, -30, -34, -22, -22, -31,
					-- layer=2 filter=210 channel=39
					-55, -2, -56, -10, 17, -5, 17, 2, 62,
					-- layer=2 filter=210 channel=40
					19, 31, 17, 42, 5, 74, 11, 68, -12,
					-- layer=2 filter=210 channel=41
					4, -2, -1, -4, 7, 9, 6, 1, 1,
					-- layer=2 filter=210 channel=42
					-41, -30, -29, 0, -17, -12, -21, -28, 29,
					-- layer=2 filter=210 channel=43
					-4, -32, 5, -23, -17, -4, -8, -12, -2,
					-- layer=2 filter=210 channel=44
					-7, 9, 0, 7, 4, -2, 0, 0, -4,
					-- layer=2 filter=210 channel=45
					61, 49, 3, 57, -9, 9, 35, -45, -14,
					-- layer=2 filter=210 channel=46
					25, -19, -80, 14, -8, -54, -34, -29, -32,
					-- layer=2 filter=210 channel=47
					-23, 17, -28, 12, -25, 17, -5, -21, -73,
					-- layer=2 filter=210 channel=48
					0, 5, 8, 7, -7, 4, -5, 7, 9,
					-- layer=2 filter=210 channel=49
					-65, -62, 0, -8, 7, -15, -47, 33, -3,
					-- layer=2 filter=210 channel=50
					-3, -4, 9, 1, 6, 7, 7, 1, 2,
					-- layer=2 filter=210 channel=51
					-16, -47, -40, -36, -19, -18, -32, -6, -9,
					-- layer=2 filter=210 channel=52
					13, -3, -16, -13, -24, -8, 13, 7, -34,
					-- layer=2 filter=210 channel=53
					-15, -5, -24, 15, 17, -41, -2, 45, 14,
					-- layer=2 filter=210 channel=54
					-6, 10, 3, -16, -8, 9, -16, -13, 20,
					-- layer=2 filter=210 channel=55
					1, 4, -1, -6, -9, -10, 3, -3, 3,
					-- layer=2 filter=210 channel=56
					-5, -51, -13, -32, -22, -7, -16, -12, -20,
					-- layer=2 filter=210 channel=57
					-2, -1, 7, -1, 5, 10, -8, -10, 3,
					-- layer=2 filter=210 channel=58
					15, 32, 2, -7, 7, -87, 49, -6, 1,
					-- layer=2 filter=210 channel=59
					28, 24, 6, -13, -1, -14, 33, 6, -31,
					-- layer=2 filter=210 channel=60
					0, 28, 5, 6, -3, 10, -23, 24, -41,
					-- layer=2 filter=210 channel=61
					-77, 8, -45, -37, 16, -20, 18, 16, 26,
					-- layer=2 filter=210 channel=62
					-32, 1, 10, 19, 30, -31, -59, 31, 20,
					-- layer=2 filter=210 channel=63
					-25, -25, -42, -42, -15, 22, 17, 17, 8,
					-- layer=2 filter=210 channel=64
					-97, -57, -19, -54, -24, 17, 11, 19, 37,
					-- layer=2 filter=210 channel=65
					-45, -19, -53, -9, 0, -70, -18, 21, 30,
					-- layer=2 filter=210 channel=66
					0, -10, -22, 20, 25, 0, 45, -8, -7,
					-- layer=2 filter=210 channel=67
					-13, 7, -68, -28, -15, -37, 9, -4, -1,
					-- layer=2 filter=210 channel=68
					-5, -2, -8, 4, -5, -11, -7, 7, -4,
					-- layer=2 filter=210 channel=69
					-31, -25, -26, -1, 13, -2, -14, 19, -18,
					-- layer=2 filter=210 channel=70
					43, 17, 27, -7, -7, -1, 4, -47, -47,
					-- layer=2 filter=210 channel=71
					19, 24, -10, 17, 2, -43, 20, 9, 1,
					-- layer=2 filter=210 channel=72
					-63, -27, -34, 38, -13, -4, -35, -24, 22,
					-- layer=2 filter=210 channel=73
					-4, 19, 18, 11, -3, 20, 17, 41, 58,
					-- layer=2 filter=210 channel=74
					-1, -9, -15, 0, -37, 22, 20, 13, -30,
					-- layer=2 filter=210 channel=75
					54, 8, -6, -17, -21, -3, 29, -27, -78,
					-- layer=2 filter=210 channel=76
					-2, 2, -7, 15, 63, 1, 16, 53, 30,
					-- layer=2 filter=210 channel=77
					2, -7, 1, 8, -11, 0, -1, -2, -6,
					-- layer=2 filter=210 channel=78
					-22, -48, -6, 14, 13, -10, -3, 15, 26,
					-- layer=2 filter=210 channel=79
					2, -5, 6, 7, 0, 5, 0, 0, -5,
					-- layer=2 filter=210 channel=80
					-19, -29, -4, -8, -60, -28, -39, -22, 4,
					-- layer=2 filter=210 channel=81
					6, 9, 5, 6, 0, 3, 7, -5, -3,
					-- layer=2 filter=210 channel=82
					5, 1, -5, 9, -8, 2, -1, 2, 7,
					-- layer=2 filter=210 channel=83
					58, 26, 9, 22, 7, -55, 48, -11, -19,
					-- layer=2 filter=210 channel=84
					-11, 6, 5, -11, -9, 0, 3, -11, -7,
					-- layer=2 filter=210 channel=85
					8, -4, 0, -5, 7, 5, 7, 0, 8,
					-- layer=2 filter=210 channel=86
					3, 1, -1, 8, -1, 9, -2, -3, -6,
					-- layer=2 filter=210 channel=87
					-5, 38, -5, -3, 12, 7, -16, 22, -15,
					-- layer=2 filter=210 channel=88
					2, -14, -65, -26, -36, -3, 41, -33, -18,
					-- layer=2 filter=210 channel=89
					15, 8, 25, 16, 4, -21, 3, 15, -32,
					-- layer=2 filter=210 channel=90
					8, 6, -10, -2, -3, -7, -3, -4, -6,
					-- layer=2 filter=210 channel=91
					14, 36, 13, 16, 10, -2, 60, 34, -34,
					-- layer=2 filter=210 channel=92
					-11, 3, -13, 7, 4, -57, 7, 10, 12,
					-- layer=2 filter=210 channel=93
					-35, -12, -22, 32, 25, -38, -31, 40, 34,
					-- layer=2 filter=210 channel=94
					-50, 30, -16, -4, 6, -42, -26, 2, -9,
					-- layer=2 filter=210 channel=95
					10, 5, -16, 19, 2, -13, 8, 3, -4,
					-- layer=2 filter=210 channel=96
					-50, -47, -6, -24, -30, -30, 24, 60, -58,
					-- layer=2 filter=210 channel=97
					-6, -15, -64, -42, -14, -9, -63, -43, 7,
					-- layer=2 filter=210 channel=98
					-53, -14, 16, 15, 2, 13, -10, -43, -54,
					-- layer=2 filter=210 channel=99
					33, 25, 19, 22, 38, 1, 13, 11, -24,
					-- layer=2 filter=210 channel=100
					45, 27, -3, -10, -11, -42, 13, -7, -8,
					-- layer=2 filter=210 channel=101
					-19, -20, -15, 13, -2, 6, 43, 14, 12,
					-- layer=2 filter=210 channel=102
					-22, -79, 9, 16, -39, -6, 5, 39, 1,
					-- layer=2 filter=210 channel=103
					-39, -44, -4, -9, -39, -17, -16, -31, 0,
					-- layer=2 filter=210 channel=104
					-55, -41, -9, -15, -12, -23, -16, 24, -11,
					-- layer=2 filter=210 channel=105
					-12, 38, 28, 40, 88, 21, -11, -20, 0,
					-- layer=2 filter=210 channel=106
					0, -11, 9, 2, 18, -32, 0, -10, -19,
					-- layer=2 filter=210 channel=107
					-31, -39, 20, 7, -30, 11, 10, -63, 16,
					-- layer=2 filter=210 channel=108
					44, 8, -3, -1, -4, -36, 2, -15, -21,
					-- layer=2 filter=210 channel=109
					-1, 0, -5, -8, -12, -9, -8, 7, 8,
					-- layer=2 filter=210 channel=110
					-61, -42, -29, 16, -27, 10, 5, 15, -5,
					-- layer=2 filter=210 channel=111
					3, 6, 1, 3, 10, 10, -6, -1, 3,
					-- layer=2 filter=210 channel=112
					-53, -31, -70, -54, 0, 16, -16, -14, -1,
					-- layer=2 filter=210 channel=113
					14, -63, -2, -32, -50, -4, 13, -5, -7,
					-- layer=2 filter=210 channel=114
					11, 0, 3, 2, 2, -10, 5, -9, -12,
					-- layer=2 filter=210 channel=115
					5, 9, -6, 7, 1, 9, -2, -2, -2,
					-- layer=2 filter=210 channel=116
					-1, 20, 0, 10, -10, 0, -9, 28, -36,
					-- layer=2 filter=210 channel=117
					-39, 9, -13, 47, -36, 50, 0, -28, 15,
					-- layer=2 filter=210 channel=118
					-23, -29, -6, -13, 2, -21, -42, -41, 14,
					-- layer=2 filter=210 channel=119
					-3, -55, 15, 3, 2, -3, 17, -9, -41,
					-- layer=2 filter=210 channel=120
					-6, -5, 1, 5, 4, 1, -3, -2, -4,
					-- layer=2 filter=210 channel=121
					-9, -7, 0, 11, -9, -9, -3, 5, -1,
					-- layer=2 filter=210 channel=122
					4, 0, 0, 12, 8, 2, 1, 9, 1,
					-- layer=2 filter=210 channel=123
					-59, -23, -14, -3, 2, -14, 2, 7, 29,
					-- layer=2 filter=210 channel=124
					12, -6, 13, 12, 18, 1, 2, 3, 51,
					-- layer=2 filter=210 channel=125
					11, 0, -8, 3, 0, 9, -10, 0, 0,
					-- layer=2 filter=210 channel=126
					-66, 7, -8, -9, -23, -56, 40, 51, -9,
					-- layer=2 filter=210 channel=127
					41, 11, -16, 15, -20, -21, -19, 2, 1,
					-- layer=2 filter=211 channel=0
					12, 6, 0, 3, 28, 28, -7, 16, 0,
					-- layer=2 filter=211 channel=1
					-15, -66, -40, -46, -26, -24, 27, 32, 21,
					-- layer=2 filter=211 channel=2
					4, 3, 5, 6, 0, -9, -6, -8, 7,
					-- layer=2 filter=211 channel=3
					33, 49, 36, 8, 11, 23, -31, -1, -35,
					-- layer=2 filter=211 channel=4
					6, 16, -18, 0, 7, 8, 25, -47, 30,
					-- layer=2 filter=211 channel=5
					9, -43, -5, 33, 27, 14, -4, 19, 31,
					-- layer=2 filter=211 channel=6
					4, -37, 17, 51, -29, 15, 18, -29, -4,
					-- layer=2 filter=211 channel=7
					-11, -20, -28, 5, 10, 20, 22, 12, 31,
					-- layer=2 filter=211 channel=8
					6, -6, -4, 3, -4, 10, 5, 4, 4,
					-- layer=2 filter=211 channel=9
					6, 33, 18, -9, 5, 3, -65, -17, -20,
					-- layer=2 filter=211 channel=10
					21, 34, 32, 9, 18, 28, -25, 27, -9,
					-- layer=2 filter=211 channel=11
					-1, -26, -11, 6, -6, -2, 26, 10, 9,
					-- layer=2 filter=211 channel=12
					14, -52, -57, 21, 2, -34, 21, 50, 60,
					-- layer=2 filter=211 channel=13
					-6, -7, 5, 5, -4, 1, 1, 6, 3,
					-- layer=2 filter=211 channel=14
					-40, -52, -43, -3, 3, -48, 17, 21, 33,
					-- layer=2 filter=211 channel=15
					-43, -17, 21, -5, 33, 39, 13, 36, 0,
					-- layer=2 filter=211 channel=16
					-3, -19, -42, -29, -36, 10, -29, -27, 4,
					-- layer=2 filter=211 channel=17
					-9, 1, -2, 3, -6, 1, 9, 9, 0,
					-- layer=2 filter=211 channel=18
					-14, -36, -43, -18, -5, -13, 8, -3, -4,
					-- layer=2 filter=211 channel=19
					-24, -19, -27, -5, -47, -14, 7, -34, 4,
					-- layer=2 filter=211 channel=20
					-1, -8, -9, 1, 1, -3, 8, -4, -2,
					-- layer=2 filter=211 channel=21
					-7, 8, -1, 9, -5, 2, -9, 4, -6,
					-- layer=2 filter=211 channel=22
					-10, -9, -3, 2, 3, 8, -5, -4, -5,
					-- layer=2 filter=211 channel=23
					4, -21, -30, -38, -62, -20, -27, -54, 1,
					-- layer=2 filter=211 channel=24
					33, 72, 38, 21, 34, 3, -69, -41, -66,
					-- layer=2 filter=211 channel=25
					14, 40, 16, 16, 4, 3, -34, -14, -27,
					-- layer=2 filter=211 channel=26
					-5, 0, -10, 2, -8, -2, 4, 0, 3,
					-- layer=2 filter=211 channel=27
					-78, -88, -92, 25, 14, 16, 28, 37, 42,
					-- layer=2 filter=211 channel=28
					-78, -23, -9, 0, 35, 5, 15, 69, 31,
					-- layer=2 filter=211 channel=29
					-3, -2, -9, -12, 4, 2, -8, 6, 8,
					-- layer=2 filter=211 channel=30
					15, -22, 12, -30, -25, 2, -7, -26, -14,
					-- layer=2 filter=211 channel=31
					21, -20, -3, -31, 4, 28, 26, 36, -60,
					-- layer=2 filter=211 channel=32
					-2, -1, -5, 0, -6, 1, -8, 6, 6,
					-- layer=2 filter=211 channel=33
					-17, -13, -56, 0, 31, 35, -10, 40, 27,
					-- layer=2 filter=211 channel=34
					-46, 12, -34, -11, 23, -12, 10, -9, -44,
					-- layer=2 filter=211 channel=35
					-39, -17, -48, -9, 11, -6, 25, 28, -5,
					-- layer=2 filter=211 channel=36
					-1, -8, 14, 6, 0, 0, -4, 11, -1,
					-- layer=2 filter=211 channel=37
					-22, -42, -18, 7, -12, 13, 22, 11, 26,
					-- layer=2 filter=211 channel=38
					-37, -57, -67, 3, 10, -2, 7, 7, 29,
					-- layer=2 filter=211 channel=39
					11, -34, -33, 6, -9, 5, -73, -68, -31,
					-- layer=2 filter=211 channel=40
					-34, -4, -6, 9, 5, 0, 42, 28, 10,
					-- layer=2 filter=211 channel=41
					1, -3, -4, 11, -8, 2, -12, -2, -5,
					-- layer=2 filter=211 channel=42
					32, 13, -58, -47, -8, -40, -38, -31, 2,
					-- layer=2 filter=211 channel=43
					-8, 3, -34, 0, -9, 0, -6, -20, -4,
					-- layer=2 filter=211 channel=44
					8, -8, 0, -5, -3, -6, 10, 0, 7,
					-- layer=2 filter=211 channel=45
					-12, -14, -83, 7, 30, 15, 0, -14, -7,
					-- layer=2 filter=211 channel=46
					-27, -16, 18, -39, 9, -1, -7, 0, -18,
					-- layer=2 filter=211 channel=47
					-31, -16, -37, 55, 63, 60, 23, 81, 71,
					-- layer=2 filter=211 channel=48
					0, 0, -6, -1, -8, 4, -11, 2, 0,
					-- layer=2 filter=211 channel=49
					-5, 0, -24, -24, -3, -20, 21, 3, -24,
					-- layer=2 filter=211 channel=50
					-12, 13, 11, 16, -14, 8, 14, 14, 12,
					-- layer=2 filter=211 channel=51
					-4, -15, 2, 12, 5, 5, 0, 11, -11,
					-- layer=2 filter=211 channel=52
					-9, -33, 26, -14, -54, 12, 21, 3, 19,
					-- layer=2 filter=211 channel=53
					-8, -29, 15, -34, 0, 30, 6, 8, -30,
					-- layer=2 filter=211 channel=54
					9, 2, -19, -3, 17, -12, -5, -17, -12,
					-- layer=2 filter=211 channel=55
					-12, -2, 3, 0, -8, -1, -5, -2, 7,
					-- layer=2 filter=211 channel=56
					-29, -50, -25, 14, -8, -6, 6, 5, 15,
					-- layer=2 filter=211 channel=57
					13, -8, 2, -3, 7, 4, -8, -7, -5,
					-- layer=2 filter=211 channel=58
					-4, -27, -65, 29, 41, -8, -3, 53, 59,
					-- layer=2 filter=211 channel=59
					-23, -49, -17, -9, -15, 4, 22, 41, 14,
					-- layer=2 filter=211 channel=60
					-9, -98, -41, -32, -15, -25, 35, 14, 43,
					-- layer=2 filter=211 channel=61
					-26, -76, -21, -1, -46, -6, 42, 7, -20,
					-- layer=2 filter=211 channel=62
					2, -7, -9, 18, -20, -11, 17, -21, -10,
					-- layer=2 filter=211 channel=63
					-9, -51, 12, -32, -63, 16, -10, -3, 18,
					-- layer=2 filter=211 channel=64
					27, 64, 35, -22, -4, 1, -43, -79, -47,
					-- layer=2 filter=211 channel=65
					9, -57, 19, -6, -34, -20, 20, -56, -8,
					-- layer=2 filter=211 channel=66
					-39, -7, -9, 49, 6, 26, -34, -25, -10,
					-- layer=2 filter=211 channel=67
					-32, 10, 51, -24, 4, 3, -73, -47, -36,
					-- layer=2 filter=211 channel=68
					1, -8, 1, 8, 0, 9, -11, 9, 0,
					-- layer=2 filter=211 channel=69
					5, 29, -2, -46, -34, -22, -58, -55, -15,
					-- layer=2 filter=211 channel=70
					-48, -71, -61, 8, 16, 3, 19, 26, 9,
					-- layer=2 filter=211 channel=71
					-79, -60, -39, -2, 20, -10, 38, 30, 21,
					-- layer=2 filter=211 channel=72
					-34, -46, -47, -39, -18, 17, 1, 11, 17,
					-- layer=2 filter=211 channel=73
					6, 19, 4, -8, 10, 1, -2, 7, -5,
					-- layer=2 filter=211 channel=74
					-14, 0, 47, -90, -20, -9, -2, 20, 9,
					-- layer=2 filter=211 channel=75
					-69, -32, -14, -16, -9, -61, 0, -33, -6,
					-- layer=2 filter=211 channel=76
					42, 5, 84, -13, 18, 7, 21, 7, -31,
					-- layer=2 filter=211 channel=77
					4, 7, 2, 6, 3, 6, -1, 7, 6,
					-- layer=2 filter=211 channel=78
					28, 26, 8, 22, -11, -3, -11, -32, -22,
					-- layer=2 filter=211 channel=79
					-8, -10, -3, 1, 8, -5, -11, -8, -5,
					-- layer=2 filter=211 channel=80
					-9, 11, 1, -50, -20, -8, -1, 8, 10,
					-- layer=2 filter=211 channel=81
					0, -13, -7, 0, 10, 11, -6, 1, -8,
					-- layer=2 filter=211 channel=82
					-3, -8, -4, 11, 3, 2, -8, 5, 6,
					-- layer=2 filter=211 channel=83
					-23, -20, -51, -35, 0, 5, -5, -43, -24,
					-- layer=2 filter=211 channel=84
					3, -3, -3, 8, 6, 4, 0, 5, 6,
					-- layer=2 filter=211 channel=85
					6, -14, -9, -1, -4, -10, -11, 0, -1,
					-- layer=2 filter=211 channel=86
					4, 0, -1, -6, -7, 4, -3, -11, 0,
					-- layer=2 filter=211 channel=87
					-3, 34, 13, 0, -8, -32, 25, -51, 19,
					-- layer=2 filter=211 channel=88
					19, -18, 21, -9, -45, -18, -31, -8, 16,
					-- layer=2 filter=211 channel=89
					-37, -25, -32, -65, -21, -25, 20, 19, 24,
					-- layer=2 filter=211 channel=90
					-4, -8, 0, 8, 0, 7, 3, -6, 0,
					-- layer=2 filter=211 channel=91
					-21, -22, -28, -53, -6, -4, -16, 32, 32,
					-- layer=2 filter=211 channel=92
					0, -57, -48, -21, 8, -20, 8, 47, 45,
					-- layer=2 filter=211 channel=93
					52, 4, 95, 9, -9, 19, 17, -26, -28,
					-- layer=2 filter=211 channel=94
					-6, -61, -18, -1, -56, 38, 25, -21, 10,
					-- layer=2 filter=211 channel=95
					-1, 0, 11, 4, 6, 5, -13, 11, 15,
					-- layer=2 filter=211 channel=96
					13, -5, 4, 41, -35, 0, 17, -14, -32,
					-- layer=2 filter=211 channel=97
					20, 35, 10, -14, 50, 19, -57, -31, -21,
					-- layer=2 filter=211 channel=98
					-43, -30, -57, 11, 21, 20, 31, 40, 45,
					-- layer=2 filter=211 channel=99
					-21, -11, -3, -9, -45, 12, 23, 4, 33,
					-- layer=2 filter=211 channel=100
					-16, -11, -21, 10, 62, 47, 17, 43, -5,
					-- layer=2 filter=211 channel=101
					-18, -28, -30, 10, 23, -36, 26, 15, -1,
					-- layer=2 filter=211 channel=102
					17, 0, -18, 17, 27, -29, 28, -19, -17,
					-- layer=2 filter=211 channel=103
					-72, -58, -21, 13, -3, -15, -14, 23, -22,
					-- layer=2 filter=211 channel=104
					-25, -17, -45, -18, -8, 2, 36, 4, -9,
					-- layer=2 filter=211 channel=105
					65, 58, 41, -65, -11, -28, 22, -89, 28,
					-- layer=2 filter=211 channel=106
					-18, 4, -8, 22, 23, 2, -12, 13, 9,
					-- layer=2 filter=211 channel=107
					6, 28, -5, -28, -1, 44, 18, -1, -7,
					-- layer=2 filter=211 channel=108
					-46, -78, -92, 7, 16, 5, 35, 19, 8,
					-- layer=2 filter=211 channel=109
					19, 6, 6, 21, 0, 0, 14, 0, -3,
					-- layer=2 filter=211 channel=110
					11, 23, 23, -43, -2, 3, -63, -87, -57,
					-- layer=2 filter=211 channel=111
					0, -3, 3, 10, -5, -3, -10, -10, 7,
					-- layer=2 filter=211 channel=112
					-3, 6, 4, -6, 14, 14, 23, 35, 0,
					-- layer=2 filter=211 channel=113
					-24, -24, -14, -61, -41, 0, -17, -22, -43,
					-- layer=2 filter=211 channel=114
					3, 11, 0, 8, -6, 5, 8, 7, 0,
					-- layer=2 filter=211 channel=115
					1, -3, 2, 1, -6, -8, -3, -3, -8,
					-- layer=2 filter=211 channel=116
					11, 1, 9, 27, -10, -24, -16, -34, 7,
					-- layer=2 filter=211 channel=117
					-34, 1, -38, -3, 1, 25, -2, 9, 34,
					-- layer=2 filter=211 channel=118
					40, 34, 29, 1, 3, 9, -4, -15, 0,
					-- layer=2 filter=211 channel=119
					-30, 18, -54, -13, 12, -38, -6, 9, 2,
					-- layer=2 filter=211 channel=120
					0, 2, 9, 0, -4, -9, 0, 3, 7,
					-- layer=2 filter=211 channel=121
					-2, -5, -11, 0, -11, 0, 3, -8, 4,
					-- layer=2 filter=211 channel=122
					11, 13, 7, 9, -8, 5, -5, -6, -9,
					-- layer=2 filter=211 channel=123
					0, -20, -9, 5, 23, 17, -1, -26, 14,
					-- layer=2 filter=211 channel=124
					20, 44, 81, -11, 23, -21, 22, -21, -88,
					-- layer=2 filter=211 channel=125
					-8, 0, -9, 8, -4, -3, -4, 0, -1,
					-- layer=2 filter=211 channel=126
					50, -39, 32, -24, 25, 59, -24, 7, -7,
					-- layer=2 filter=211 channel=127
					2, 19, -23, 0, -25, -34, -40, -28, -25,
					-- layer=2 filter=212 channel=0
					-13, 15, 17, 13, 19, 14, -4, -12, -6,
					-- layer=2 filter=212 channel=1
					21, -23, 11, 11, -19, 1, 7, -14, -37,
					-- layer=2 filter=212 channel=2
					5, 9, 2, 3, -1, 0, 11, 1, 10,
					-- layer=2 filter=212 channel=3
					-73, -37, -21, -2, 13, 3, -43, -42, -43,
					-- layer=2 filter=212 channel=4
					-16, -13, 8, 6, 6, -14, -13, -24, 3,
					-- layer=2 filter=212 channel=5
					3, 19, -5, -1, -10, 4, -8, -15, 1,
					-- layer=2 filter=212 channel=6
					29, -20, -24, -9, 2, 37, -18, -22, 17,
					-- layer=2 filter=212 channel=7
					0, 0, 0, 37, 0, -15, 8, -41, 3,
					-- layer=2 filter=212 channel=8
					0, 0, -5, -2, -9, -2, 8, -4, -8,
					-- layer=2 filter=212 channel=9
					-62, -67, -26, -14, -39, 12, -47, -54, -26,
					-- layer=2 filter=212 channel=10
					-49, -32, -12, -6, -11, 3, -16, 5, 2,
					-- layer=2 filter=212 channel=11
					6, 30, 20, 3, 12, -5, -6, -21, 12,
					-- layer=2 filter=212 channel=12
					13, -4, 10, 11, 17, 15, 13, 0, 0,
					-- layer=2 filter=212 channel=13
					-4, 1, -3, 10, 10, 1, 6, -1, -2,
					-- layer=2 filter=212 channel=14
					27, -38, 4, 18, -9, -5, 24, 11, 9,
					-- layer=2 filter=212 channel=15
					-36, 8, 42, 13, 5, 4, -6, 28, 28,
					-- layer=2 filter=212 channel=16
					0, 47, 16, 0, -21, -4, 9, -7, -4,
					-- layer=2 filter=212 channel=17
					-6, -2, 5, 11, 6, 7, -5, 2, -1,
					-- layer=2 filter=212 channel=18
					-6, 29, 4, -6, 1, -30, -26, 4, -17,
					-- layer=2 filter=212 channel=19
					33, 14, 37, -19, -27, 0, -1, 19, 0,
					-- layer=2 filter=212 channel=20
					1, 8, -1, 7, 10, 6, 4, -6, -1,
					-- layer=2 filter=212 channel=21
					-9, 0, -1, 4, -1, 3, 0, -11, 19,
					-- layer=2 filter=212 channel=22
					1, 7, -2, 0, 8, 0, 2, 1, 4,
					-- layer=2 filter=212 channel=23
					-43, -18, -20, 18, 2, -3, -49, 11, -18,
					-- layer=2 filter=212 channel=24
					-59, 2, -16, 0, 7, 23, -36, -8, 24,
					-- layer=2 filter=212 channel=25
					-20, 23, 25, 25, 37, 34, 7, 23, 45,
					-- layer=2 filter=212 channel=26
					8, 0, 5, 4, 5, -1, -4, 5, 0,
					-- layer=2 filter=212 channel=27
					-24, -8, 0, 1, -22, -31, 1, -11, -12,
					-- layer=2 filter=212 channel=28
					12, -19, -21, 57, -4, -5, -21, 3, -33,
					-- layer=2 filter=212 channel=29
					0, 6, 9, -3, -7, -5, -10, -4, -6,
					-- layer=2 filter=212 channel=30
					0, -68, -49, -16, -47, 6, 11, -3, 14,
					-- layer=2 filter=212 channel=31
					-10, 67, 18, 14, 31, -8, 4, 45, 21,
					-- layer=2 filter=212 channel=32
					0, -8, 9, 10, 7, -6, 0, 9, 11,
					-- layer=2 filter=212 channel=33
					-20, -46, -32, -3, -46, -20, 36, -5, 19,
					-- layer=2 filter=212 channel=34
					-3, 27, 13, -31, -31, -14, 0, 12, -5,
					-- layer=2 filter=212 channel=35
					-33, -38, 3, 7, 14, -7, -25, -72, -46,
					-- layer=2 filter=212 channel=36
					8, 3, 3, 4, 6, -8, 8, 4, -10,
					-- layer=2 filter=212 channel=37
					6, 9, 20, -27, -3, -8, 0, -10, -5,
					-- layer=2 filter=212 channel=38
					-30, -28, -12, 0, -22, -14, 40, -6, -13,
					-- layer=2 filter=212 channel=39
					-20, -40, -9, 39, -10, -18, -32, -66, -44,
					-- layer=2 filter=212 channel=40
					-22, 21, 53, 36, 13, -8, -8, 5, 56,
					-- layer=2 filter=212 channel=41
					-8, -9, -6, 6, -3, -11, 1, 12, -9,
					-- layer=2 filter=212 channel=42
					-5, 13, 18, 22, -6, 14, 41, -13, -9,
					-- layer=2 filter=212 channel=43
					-47, 0, -11, -54, -24, -10, 11, 16, -37,
					-- layer=2 filter=212 channel=44
					5, -8, 6, -5, -1, -2, -4, -9, 4,
					-- layer=2 filter=212 channel=45
					39, 77, 28, -14, -3, 1, 46, 44, 43,
					-- layer=2 filter=212 channel=46
					-31, 13, 2, -23, 0, -1, -25, -19, -24,
					-- layer=2 filter=212 channel=47
					-31, -59, -61, -10, -39, -40, 17, -11, -12,
					-- layer=2 filter=212 channel=48
					1, 7, -8, -7, -9, 8, -2, 7, -4,
					-- layer=2 filter=212 channel=49
					-9, 20, 34, -23, -2, -8, -37, 14, 32,
					-- layer=2 filter=212 channel=50
					0, -11, 4, -22, 0, 1, -7, -18, 5,
					-- layer=2 filter=212 channel=51
					10, 18, 33, -8, 14, 12, -7, 10, 12,
					-- layer=2 filter=212 channel=52
					63, 36, 13, 14, 6, 20, 13, -29, -1,
					-- layer=2 filter=212 channel=53
					-18, 46, 77, 3, -9, 51, 14, -17, 21,
					-- layer=2 filter=212 channel=54
					44, 48, 25, 14, 34, 9, 24, 1, -9,
					-- layer=2 filter=212 channel=55
					-15, 3, 5, 1, 4, 7, -9, 2, -5,
					-- layer=2 filter=212 channel=56
					7, 29, 20, -3, -2, -1, -13, -37, -24,
					-- layer=2 filter=212 channel=57
					1, 1, 0, 4, 0, -12, 1, -6, -1,
					-- layer=2 filter=212 channel=58
					35, -4, 14, 25, 19, 22, 13, -4, -10,
					-- layer=2 filter=212 channel=59
					-10, 7, -17, -9, -55, -24, -17, -48, -19,
					-- layer=2 filter=212 channel=60
					18, -23, -21, -12, -60, -11, 16, 4, -24,
					-- layer=2 filter=212 channel=61
					3, 47, -43, 1, -42, -36, 19, -44, 6,
					-- layer=2 filter=212 channel=62
					16, 9, 28, -10, -12, 12, 6, 20, 30,
					-- layer=2 filter=212 channel=63
					-12, -14, -10, 22, 0, -15, -18, -8, -8,
					-- layer=2 filter=212 channel=64
					-29, -30, -6, 6, 2, 20, -16, -18, -2,
					-- layer=2 filter=212 channel=65
					13, 24, -13, -49, -26, -3, -17, -56, -12,
					-- layer=2 filter=212 channel=66
					25, 14, 43, 5, -19, 5, 49, -23, -25,
					-- layer=2 filter=212 channel=67
					-36, -21, -22, -2, 22, 28, -70, -38, -40,
					-- layer=2 filter=212 channel=68
					9, 5, 7, -8, -6, 4, 10, -9, -6,
					-- layer=2 filter=212 channel=69
					-34, -43, -7, -2, -26, 25, -22, -13, -3,
					-- layer=2 filter=212 channel=70
					42, -18, -4, 25, 13, -14, 0, -16, -22,
					-- layer=2 filter=212 channel=71
					-8, 36, 32, 13, -9, -6, -7, -29, -3,
					-- layer=2 filter=212 channel=72
					3, -33, -11, 69, 2, -53, 19, -8, 12,
					-- layer=2 filter=212 channel=73
					41, 75, 36, 50, 28, -3, 39, 25, 8,
					-- layer=2 filter=212 channel=74
					-27, -31, -67, 75, 52, 23, 15, 18, -31,
					-- layer=2 filter=212 channel=75
					59, 17, -3, 63, 61, -12, -4, -3, 34,
					-- layer=2 filter=212 channel=76
					50, -17, 29, 15, -4, 32, 35, -34, 3,
					-- layer=2 filter=212 channel=77
					-6, 9, -6, 4, 5, 10, -10, -1, -8,
					-- layer=2 filter=212 channel=78
					-16, 36, 31, -12, 3, -12, 5, 5, 35,
					-- layer=2 filter=212 channel=79
					8, -3, 2, 7, 10, 3, 3, -4, 11,
					-- layer=2 filter=212 channel=80
					-63, -12, -46, -35, 2, -11, -36, -44, -2,
					-- layer=2 filter=212 channel=81
					-3, 12, -10, 12, 14, 3, -5, -1, 7,
					-- layer=2 filter=212 channel=82
					-4, -3, 2, -4, -7, 3, 0, -1, -6,
					-- layer=2 filter=212 channel=83
					-74, -12, -5, 7, -27, -15, -32, -26, 16,
					-- layer=2 filter=212 channel=84
					-8, -9, 7, -10, 1, -1, 8, 3, 8,
					-- layer=2 filter=212 channel=85
					-8, 0, 0, 8, -9, 7, 0, -5, -10,
					-- layer=2 filter=212 channel=86
					-2, 4, 29, -12, 2, 2, -1, -10, 15,
					-- layer=2 filter=212 channel=87
					-56, -28, 5, -26, -9, -52, -40, -51, -11,
					-- layer=2 filter=212 channel=88
					-8, -100, -71, -38, -39, -50, 33, 13, -8,
					-- layer=2 filter=212 channel=89
					18, -23, -14, 30, -10, -8, 17, 12, 13,
					-- layer=2 filter=212 channel=90
					1, -5, 8, 10, -6, 8, -9, 2, 0,
					-- layer=2 filter=212 channel=91
					19, -21, 18, 35, -6, -10, 16, -16, -20,
					-- layer=2 filter=212 channel=92
					21, -17, 5, -2, -14, -7, 14, -13, -56,
					-- layer=2 filter=212 channel=93
					53, -21, 21, -6, 17, 21, -41, -15, -36,
					-- layer=2 filter=212 channel=94
					11, -4, -1, -2, -25, 16, -16, -20, 17,
					-- layer=2 filter=212 channel=95
					-3, 4, 3, -17, 1, 6, -14, -17, -5,
					-- layer=2 filter=212 channel=96
					18, 39, 22, -2, 37, 30, 42, 12, -1,
					-- layer=2 filter=212 channel=97
					-74, -37, -13, 25, -11, -7, 1, -15, 24,
					-- layer=2 filter=212 channel=98
					-12, -5, -26, 24, -20, -16, -23, -5, 8,
					-- layer=2 filter=212 channel=99
					30, 21, 32, 7, -12, 16, 23, 10, -15,
					-- layer=2 filter=212 channel=100
					-71, -76, -51, -18, -55, -33, 31, -23, -13,
					-- layer=2 filter=212 channel=101
					-9, 41, 63, 44, 14, 23, 7, -8, -2,
					-- layer=2 filter=212 channel=102
					-18, 2, 22, -13, 27, 10, -24, 7, -31,
					-- layer=2 filter=212 channel=103
					-26, 20, -15, 0, -11, -11, 11, 12, 3,
					-- layer=2 filter=212 channel=104
					-38, 31, 31, -2, -6, 7, -29, 20, 7,
					-- layer=2 filter=212 channel=105
					0, -23, -7, -31, -32, 21, 26, 6, -42,
					-- layer=2 filter=212 channel=106
					-1, -12, -11, 37, 21, 22, 5, 7, 17,
					-- layer=2 filter=212 channel=107
					0, 44, 11, -6, -5, -39, -3, -26, 0,
					-- layer=2 filter=212 channel=108
					-20, -27, -12, 0, -35, -16, 32, -2, -4,
					-- layer=2 filter=212 channel=109
					7, -18, -13, -3, -1, -1, -11, 2, 5,
					-- layer=2 filter=212 channel=110
					21, 23, 1, 9, -11, -10, 19, -18, 4,
					-- layer=2 filter=212 channel=111
					-4, 7, 12, 1, 8, 5, 1, -10, 3,
					-- layer=2 filter=212 channel=112
					-17, 44, -9, -30, 3, -40, -29, -32, 12,
					-- layer=2 filter=212 channel=113
					-4, -33, 24, -33, -47, -38, -31, -18, -8,
					-- layer=2 filter=212 channel=114
					1, -5, 1, -3, 12, -11, 10, 13, 6,
					-- layer=2 filter=212 channel=115
					7, 0, 8, -4, 4, 6, 5, -3, -5,
					-- layer=2 filter=212 channel=116
					-45, 2, 23, -37, 15, -36, -72, -41, -22,
					-- layer=2 filter=212 channel=117
					32, 35, -1, 80, -5, 8, 40, -23, -13,
					-- layer=2 filter=212 channel=118
					6, -15, 32, -33, -21, -10, 16, 0, -6,
					-- layer=2 filter=212 channel=119
					-4, 4, -26, -37, 9, -11, 49, -2, -17,
					-- layer=2 filter=212 channel=120
					6, -5, -6, -3, 7, 6, 0, 4, 6,
					-- layer=2 filter=212 channel=121
					9, 10, -4, 5, 5, -6, 2, -1, 10,
					-- layer=2 filter=212 channel=122
					-4, 3, -17, 2, 13, -10, 8, -2, 4,
					-- layer=2 filter=212 channel=123
					16, -13, -12, 43, 5, 8, 2, -23, 31,
					-- layer=2 filter=212 channel=124
					35, 41, 17, 68, 32, 14, 48, 19, 41,
					-- layer=2 filter=212 channel=125
					-6, -8, -1, 0, -2, 4, 1, -1, -4,
					-- layer=2 filter=212 channel=126
					17, 35, 11, 25, 32, 14, 92, 41, 33,
					-- layer=2 filter=212 channel=127
					-25, -35, -24, -19, -39, -34, 28, -3, -27,
					-- layer=2 filter=213 channel=0
					9, -17, -20, -17, -4, -13, -29, 12, 24,
					-- layer=2 filter=213 channel=1
					-3, 4, 6, -10, -9, 4, -10, -2, 0,
					-- layer=2 filter=213 channel=2
					-1, 3, 7, 2, -1, 3, 7, -10, 5,
					-- layer=2 filter=213 channel=3
					12, -8, 30, -18, -4, 19, -16, -29, 19,
					-- layer=2 filter=213 channel=4
					32, 8, 10, 2, 2, 8, -22, -41, -38,
					-- layer=2 filter=213 channel=5
					-22, -15, 0, 2, 6, -5, 21, 19, 17,
					-- layer=2 filter=213 channel=6
					21, 38, -35, 31, 65, 16, 56, 74, -6,
					-- layer=2 filter=213 channel=7
					-12, 3, 54, -15, -21, 77, -23, 0, 19,
					-- layer=2 filter=213 channel=8
					0, -5, 0, -7, 11, 6, 5, -9, 4,
					-- layer=2 filter=213 channel=9
					22, -30, -8, 9, -9, 23, 8, -14, 25,
					-- layer=2 filter=213 channel=10
					26, -30, -22, -13, -11, -7, -34, -14, 0,
					-- layer=2 filter=213 channel=11
					-2, -4, 0, -15, 0, 10, 5, 13, 10,
					-- layer=2 filter=213 channel=12
					-6, -5, 20, -10, 0, 30, -33, -30, 4,
					-- layer=2 filter=213 channel=13
					0, -4, 6, 10, 8, -5, -10, 7, -5,
					-- layer=2 filter=213 channel=14
					-8, -15, 5, -16, -28, 0, -12, -24, -3,
					-- layer=2 filter=213 channel=15
					-36, -41, -39, 0, -8, 0, 12, 6, 28,
					-- layer=2 filter=213 channel=16
					15, 33, 49, 77, 28, 8, 18, -40, -35,
					-- layer=2 filter=213 channel=17
					-5, 9, -8, -10, 2, 9, 4, -2, 8,
					-- layer=2 filter=213 channel=18
					-6, 32, 0, 10, 9, -34, -37, 9, -12,
					-- layer=2 filter=213 channel=19
					-5, 19, -36, 0, -18, -14, 16, 4, -21,
					-- layer=2 filter=213 channel=20
					10, 9, 4, 9, 2, 1, -2, 5, -5,
					-- layer=2 filter=213 channel=21
					-13, -5, -14, 5, -7, -6, 1, -20, -21,
					-- layer=2 filter=213 channel=22
					10, 7, -4, -4, -1, -1, 5, -5, -1,
					-- layer=2 filter=213 channel=23
					7, -7, 1, 18, 16, 13, -19, -29, -3,
					-- layer=2 filter=213 channel=24
					40, 1, 11, -15, -30, 4, -11, -7, 10,
					-- layer=2 filter=213 channel=25
					-5, -11, 27, -17, -27, 20, -14, -9, 20,
					-- layer=2 filter=213 channel=26
					-10, 1, -1, -6, -1, -6, 4, 8, 6,
					-- layer=2 filter=213 channel=27
					-5, -13, -21, -3, 9, 7, 11, 12, 24,
					-- layer=2 filter=213 channel=28
					13, -8, 33, 25, -23, 22, -40, -89, 0,
					-- layer=2 filter=213 channel=29
					0, -5, 3, 9, -6, 0, -1, 2, 7,
					-- layer=2 filter=213 channel=30
					15, 8, -3, -16, -14, 1, -39, -20, -38,
					-- layer=2 filter=213 channel=31
					-49, 38, 8, -4, 32, 8, -21, 9, 4,
					-- layer=2 filter=213 channel=32
					-2, -6, 0, 0, 0, 0, -6, 12, -4,
					-- layer=2 filter=213 channel=33
					6, -20, 46, -28, -41, 32, 49, -17, 32,
					-- layer=2 filter=213 channel=34
					2, 35, 12, -9, -45, 0, 6, -3, -6,
					-- layer=2 filter=213 channel=35
					6, 9, 31, 39, -7, 33, -61, -56, -84,
					-- layer=2 filter=213 channel=36
					-15, 9, -7, -2, 3, 9, -10, 1, -10,
					-- layer=2 filter=213 channel=37
					-6, -5, -5, 2, 0, 12, 23, 7, 30,
					-- layer=2 filter=213 channel=38
					-1, -12, -22, 7, -1, 8, 27, 14, 3,
					-- layer=2 filter=213 channel=39
					-8, 4, 9, 8, -2, 0, 7, -61, 7,
					-- layer=2 filter=213 channel=40
					6, 4, 14, -17, 3, 42, -27, 37, 4,
					-- layer=2 filter=213 channel=41
					-7, 0, -7, -3, 5, -5, 3, 3, -10,
					-- layer=2 filter=213 channel=42
					-3, -10, 7, 37, -4, 30, -5, -56, -32,
					-- layer=2 filter=213 channel=43
					-25, -15, 16, -17, -14, 32, -24, -15, 21,
					-- layer=2 filter=213 channel=44
					6, 4, 5, -5, -3, -4, -2, 6, 5,
					-- layer=2 filter=213 channel=45
					-15, 25, 43, 13, -7, 51, -21, -45, -39,
					-- layer=2 filter=213 channel=46
					44, 4, 16, 13, -49, -20, -29, -26, -31,
					-- layer=2 filter=213 channel=47
					55, 23, 53, 8, -4, 49, -3, -71, -26,
					-- layer=2 filter=213 channel=48
					11, -9, -2, 9, -8, -8, 0, 2, -4,
					-- layer=2 filter=213 channel=49
					-8, 22, 6, -6, 22, -22, -30, 25, -32,
					-- layer=2 filter=213 channel=50
					-27, -15, -17, 1, -18, -5, -6, -29, 0,
					-- layer=2 filter=213 channel=51
					-1, -14, 0, -2, -13, -3, -2, -1, 21,
					-- layer=2 filter=213 channel=52
					-17, -8, -30, 2, 27, 17, -20, -4, 16,
					-- layer=2 filter=213 channel=53
					5, 22, -75, 14, -9, -1, 10, 18, -61,
					-- layer=2 filter=213 channel=54
					-3, 8, 32, -2, -11, 18, -23, -7, -38,
					-- layer=2 filter=213 channel=55
					7, 19, 5, -6, -3, -6, 3, 9, 12,
					-- layer=2 filter=213 channel=56
					-10, 4, -2, -7, 7, 5, 15, 16, 31,
					-- layer=2 filter=213 channel=57
					0, 4, -3, -3, 8, 17, 7, -5, 2,
					-- layer=2 filter=213 channel=58
					-13, 0, 28, -1, -13, 25, -26, -61, 4,
					-- layer=2 filter=213 channel=59
					1, 26, -16, -11, 16, -6, -19, -9, -21,
					-- layer=2 filter=213 channel=60
					4, 16, 0, -13, -16, -16, -16, 9, -45,
					-- layer=2 filter=213 channel=61
					-5, 23, -40, -7, 13, -36, -33, 8, -23,
					-- layer=2 filter=213 channel=62
					7, 19, -21, -41, 21, -4, 10, 28, -51,
					-- layer=2 filter=213 channel=63
					6, 16, 27, -5, 15, -1, -29, -17, -9,
					-- layer=2 filter=213 channel=64
					8, 11, -3, 1, 24, -1, -15, -7, -38,
					-- layer=2 filter=213 channel=65
					34, 51, -27, 37, 18, -2, -1, 44, -38,
					-- layer=2 filter=213 channel=66
					-16, 4, 39, 2, 37, -46, -5, -38, 19,
					-- layer=2 filter=213 channel=67
					16, 0, -39, 53, 12, -28, 10, 8, -15,
					-- layer=2 filter=213 channel=68
					1, -9, -1, 0, 1, -7, 0, 4, -7,
					-- layer=2 filter=213 channel=69
					11, 21, 7, 7, -8, 4, 15, 0, -22,
					-- layer=2 filter=213 channel=70
					-5, 6, 0, 29, 4, 50, -51, -55, -34,
					-- layer=2 filter=213 channel=71
					-20, -10, -11, -5, 0, -8, 14, 3, 18,
					-- layer=2 filter=213 channel=72
					11, -41, 16, 1, -51, 2, 10, -27, -8,
					-- layer=2 filter=213 channel=73
					-2, 21, 6, 9, 30, 33, 4, 35, 0,
					-- layer=2 filter=213 channel=74
					9, -12, -18, 48, 11, -11, -14, -12, -44,
					-- layer=2 filter=213 channel=75
					35, 27, 98, 53, -14, 41, -43, -6, -30,
					-- layer=2 filter=213 channel=76
					31, 4, -38, -48, -7, 20, -26, -13, -90,
					-- layer=2 filter=213 channel=77
					-1, 6, -7, -9, -5, 1, 0, 3, 2,
					-- layer=2 filter=213 channel=78
					-17, -4, -2, -9, -4, 5, -5, 24, -3,
					-- layer=2 filter=213 channel=79
					0, -9, -7, 0, 8, -9, 0, 6, -4,
					-- layer=2 filter=213 channel=80
					-7, 2, -6, 0, -15, -35, -28, -53, -24,
					-- layer=2 filter=213 channel=81
					2, -10, -10, 0, 2, -2, -13, -2, -4,
					-- layer=2 filter=213 channel=82
					-8, 4, 9, 5, -12, 5, 12, 7, -5,
					-- layer=2 filter=213 channel=83
					17, 22, 9, 32, 47, 10, -29, -33, -45,
					-- layer=2 filter=213 channel=84
					0, 3, 3, -3, -3, 6, -4, -9, -6,
					-- layer=2 filter=213 channel=85
					5, -15, -10, 6, 2, -9, 2, 9, 0,
					-- layer=2 filter=213 channel=86
					10, 3, -2, 0, 15, -9, -4, -13, -3,
					-- layer=2 filter=213 channel=87
					28, 42, -44, 7, -18, -50, -26, -4, -82,
					-- layer=2 filter=213 channel=88
					-5, 9, -2, 5, -8, 18, -8, -11, -39,
					-- layer=2 filter=213 channel=89
					9, -7, -9, -10, -8, -14, -25, -42, -26,
					-- layer=2 filter=213 channel=90
					0, 9, 0, -4, 0, -10, -9, 8, -1,
					-- layer=2 filter=213 channel=91
					12, -19, 21, 17, -23, 23, -17, -29, 2,
					-- layer=2 filter=213 channel=92
					0, -21, -4, -15, -19, 2, -8, -17, 5,
					-- layer=2 filter=213 channel=93
					3, 33, 41, -1, -2, 35, 19, 43, -22,
					-- layer=2 filter=213 channel=94
					42, 24, -27, 11, 23, 12, 15, 9, -11,
					-- layer=2 filter=213 channel=95
					-1, -12, 0, -10, -4, -20, -8, -1, -21,
					-- layer=2 filter=213 channel=96
					50, 32, 41, 27, 65, 48, 45, 66, 16,
					-- layer=2 filter=213 channel=97
					21, -2, 40, -15, -15, 17, 14, -1, 5,
					-- layer=2 filter=213 channel=98
					23, 19, 18, 3, -35, 24, -31, -79, -44,
					-- layer=2 filter=213 channel=99
					22, -16, -27, 30, 23, 3, 16, 37, 20,
					-- layer=2 filter=213 channel=100
					-28, -2, -3, 47, 5, 19, -33, -11, -54,
					-- layer=2 filter=213 channel=101
					7, -19, 25, -28, -24, 26, -13, -16, 42,
					-- layer=2 filter=213 channel=102
					0, 29, 36, 26, 18, -14, 19, 17, -9,
					-- layer=2 filter=213 channel=103
					1, 8, -45, 11, 2, 3, -13, 2, 0,
					-- layer=2 filter=213 channel=104
					56, 29, -10, -6, 31, -27, 28, 19, -50,
					-- layer=2 filter=213 channel=105
					12, -39, -11, 1, -29, 26, -46, -48, -91,
					-- layer=2 filter=213 channel=106
					8, -6, 43, 3, -49, 28, 3, -34, 39,
					-- layer=2 filter=213 channel=107
					53, 72, 31, 9, -12, -7, 4, 16, -17,
					-- layer=2 filter=213 channel=108
					-22, -20, -2, 1, 7, 4, 2, 22, 30,
					-- layer=2 filter=213 channel=109
					1, 9, -7, -3, 3, -9, 11, 3, 3,
					-- layer=2 filter=213 channel=110
					14, 0, 29, 10, 30, 19, -36, -35, -19,
					-- layer=2 filter=213 channel=111
					0, 8, -5, 5, 6, -1, 3, -4, 0,
					-- layer=2 filter=213 channel=112
					21, -11, -22, 17, -25, -19, -7, 11, 20,
					-- layer=2 filter=213 channel=113
					0, 20, 2, -7, 17, -20, -45, -71, -57,
					-- layer=2 filter=213 channel=114
					7, 10, 13, -3, 11, 7, 7, -2, 7,
					-- layer=2 filter=213 channel=115
					6, -6, -8, -3, 4, -8, 0, 7, 9,
					-- layer=2 filter=213 channel=116
					13, 39, -31, 19, 0, -33, -29, -2, -14,
					-- layer=2 filter=213 channel=117
					-4, -16, -21, -7, -37, 27, -1, -48, -39,
					-- layer=2 filter=213 channel=118
					-20, -26, 3, -21, 5, 9, -19, -9, -11,
					-- layer=2 filter=213 channel=119
					13, 17, 12, 0, 0, -7, -37, -16, -32,
					-- layer=2 filter=213 channel=120
					-7, -9, 0, -5, 4, -1, -5, -5, 9,
					-- layer=2 filter=213 channel=121
					-3, -7, 6, -3, 9, 6, 6, 3, 11,
					-- layer=2 filter=213 channel=122
					6, 1, 1, -2, 9, -6, 12, 3, 7,
					-- layer=2 filter=213 channel=123
					1, 18, 39, -12, -17, 66, -3, -28, -15,
					-- layer=2 filter=213 channel=124
					0, -5, -16, 20, -6, 35, 9, 31, -32,
					-- layer=2 filter=213 channel=125
					1, -2, 0, 12, 6, -8, -4, -6, 3,
					-- layer=2 filter=213 channel=126
					43, -21, -19, 11, 20, 57, -2, 49, 44,
					-- layer=2 filter=213 channel=127
					23, 13, 17, -5, -16, 16, 0, -36, -20,
					-- layer=2 filter=214 channel=0
					16, -8, -10, 22, -4, -24, 35, -9, -3,
					-- layer=2 filter=214 channel=1
					-36, -13, 36, -5, 11, 52, -22, -2, 38,
					-- layer=2 filter=214 channel=2
					-1, 0, -9, 9, -6, -3, -8, -1, 0,
					-- layer=2 filter=214 channel=3
					31, 11, -33, 69, 27, -54, 22, -5, -30,
					-- layer=2 filter=214 channel=4
					-14, 6, -14, -24, -32, -13, -10, 9, 4,
					-- layer=2 filter=214 channel=5
					12, 25, 33, 0, 15, -28, 13, -10, -5,
					-- layer=2 filter=214 channel=6
					5, -68, -8, -38, -22, 5, -64, -3, -13,
					-- layer=2 filter=214 channel=7
					-36, 34, 27, -9, -41, 11, -25, -15, -18,
					-- layer=2 filter=214 channel=8
					0, -2, -8, -8, 5, 5, 3, -10, 8,
					-- layer=2 filter=214 channel=9
					12, 15, -14, 8, 0, -37, 0, -9, 20,
					-- layer=2 filter=214 channel=10
					21, -4, 5, 47, 4, -40, 19, -5, -14,
					-- layer=2 filter=214 channel=11
					24, 23, -10, 11, 15, -26, 12, 4, -33,
					-- layer=2 filter=214 channel=12
					-38, 21, 20, -14, 21, 67, -35, -3, 25,
					-- layer=2 filter=214 channel=13
					3, -4, 4, -9, -7, 0, 0, 4, -1,
					-- layer=2 filter=214 channel=14
					-10, -3, 17, -29, 9, 20, -19, -10, 0,
					-- layer=2 filter=214 channel=15
					24, 30, 4, 50, 12, 42, -16, -26, 52,
					-- layer=2 filter=214 channel=16
					-25, -22, 16, -21, -27, 2, -45, -25, 59,
					-- layer=2 filter=214 channel=17
					-2, -1, 7, -2, 2, -8, -2, 3, 6,
					-- layer=2 filter=214 channel=18
					-6, 47, 0, 12, 34, 30, -7, 27, 20,
					-- layer=2 filter=214 channel=19
					-29, -35, 30, -36, -10, 46, -42, 11, 27,
					-- layer=2 filter=214 channel=20
					-11, 7, 11, 8, 0, 6, -2, 6, 5,
					-- layer=2 filter=214 channel=21
					-8, 3, 12, 14, -17, -10, 2, 2, 12,
					-- layer=2 filter=214 channel=22
					7, 9, -2, 2, 0, -4, 9, 11, 3,
					-- layer=2 filter=214 channel=23
					-62, -38, -25, -17, -44, -22, -41, 10, 3,
					-- layer=2 filter=214 channel=24
					32, 2, -47, 43, 3, -71, 30, -25, -46,
					-- layer=2 filter=214 channel=25
					35, 15, -57, 31, 5, -75, 10, -16, -87,
					-- layer=2 filter=214 channel=26
					-3, 6, -2, -1, 6, -4, 10, -10, 5,
					-- layer=2 filter=214 channel=27
					-26, 4, 18, -48, 16, 19, -21, 26, 27,
					-- layer=2 filter=214 channel=28
					26, 24, -3, -28, 4, 20, 50, 37, 15,
					-- layer=2 filter=214 channel=29
					9, -7, -3, 3, 0, -7, -8, -7, -6,
					-- layer=2 filter=214 channel=30
					-45, 7, 1, -34, -6, 0, -33, -28, 28,
					-- layer=2 filter=214 channel=31
					45, 11, 53, 27, 36, 51, 0, 16, -13,
					-- layer=2 filter=214 channel=32
					3, 0, 1, -8, -1, -4, -7, 5, 11,
					-- layer=2 filter=214 channel=33
					6, 28, 1, 3, 5, 54, -19, -38, 13,
					-- layer=2 filter=214 channel=34
					-30, 7, 5, -32, 22, 50, 9, 0, 55,
					-- layer=2 filter=214 channel=35
					25, 9, 17, -29, -12, 40, 14, 11, 24,
					-- layer=2 filter=214 channel=36
					-9, -10, 5, 0, -12, -7, -12, -5, -6,
					-- layer=2 filter=214 channel=37
					23, -3, -15, 9, 15, -17, -3, 16, -2,
					-- layer=2 filter=214 channel=38
					-25, 0, 41, -24, 26, 36, -11, 27, 39,
					-- layer=2 filter=214 channel=39
					-33, 34, 37, 2, -18, -11, 12, 14, 28,
					-- layer=2 filter=214 channel=40
					16, 11, -5, -7, 36, -12, -4, 5, 41,
					-- layer=2 filter=214 channel=41
					0, -1, -7, -10, 12, 6, 0, 1, -3,
					-- layer=2 filter=214 channel=42
					11, -30, -39, -35, -27, 30, -11, 31, 76,
					-- layer=2 filter=214 channel=43
					35, 18, -14, 15, 20, -6, 16, -15, -14,
					-- layer=2 filter=214 channel=44
					-2, -9, 3, -6, -5, 2, -4, -10, 4,
					-- layer=2 filter=214 channel=45
					-48, 29, 63, -65, -11, 23, -13, -10, 22,
					-- layer=2 filter=214 channel=46
					-23, 2, 18, 5, 0, -1, -6, -19, 12,
					-- layer=2 filter=214 channel=47
					-26, -5, 0, -34, -7, 29, 12, -12, 12,
					-- layer=2 filter=214 channel=48
					8, 3, -3, -7, 6, 0, -4, 0, 9,
					-- layer=2 filter=214 channel=49
					-18, 36, -34, 14, 14, -1, -37, 5, -17,
					-- layer=2 filter=214 channel=50
					-6, -13, 8, -12, -19, 2, 4, -1, -17,
					-- layer=2 filter=214 channel=51
					23, 12, -10, 19, 16, -21, 19, -13, -26,
					-- layer=2 filter=214 channel=52
					-17, -15, -26, -2, -15, 9, 0, -4, 33,
					-- layer=2 filter=214 channel=53
					-28, -24, 7, 0, -47, 0, -85, 0, -11,
					-- layer=2 filter=214 channel=54
					0, 3, 19, 0, -2, 39, 0, 5, 18,
					-- layer=2 filter=214 channel=55
					4, -10, 14, 9, 4, 9, 8, 4, -10,
					-- layer=2 filter=214 channel=56
					36, 50, -2, 4, 7, -17, 38, 10, -23,
					-- layer=2 filter=214 channel=57
					2, 16, -16, -9, 21, 0, -3, 10, -3,
					-- layer=2 filter=214 channel=58
					8, 19, 80, -59, 11, 27, -13, 35, 37,
					-- layer=2 filter=214 channel=59
					3, -39, 14, -43, 45, 76, -3, 28, 66,
					-- layer=2 filter=214 channel=60
					-2, 20, 60, -34, 25, 36, -5, 33, 43,
					-- layer=2 filter=214 channel=61
					-26, -4, 28, -41, -10, 17, -11, -31, -7,
					-- layer=2 filter=214 channel=62
					-9, -18, 4, -51, -12, 9, -35, 12, -25,
					-- layer=2 filter=214 channel=63
					-57, -19, -12, -36, -27, -5, -3, -46, 10,
					-- layer=2 filter=214 channel=64
					-4, -11, -8, -4, -5, 6, -25, 0, 20,
					-- layer=2 filter=214 channel=65
					-44, -5, -36, -19, -30, 13, -34, -5, 23,
					-- layer=2 filter=214 channel=66
					-32, -7, -17, 3, -9, 21, 12, -26, 7,
					-- layer=2 filter=214 channel=67
					15, -12, -19, 16, -12, -50, 48, 6, 4,
					-- layer=2 filter=214 channel=68
					-1, 8, -7, 4, -3, 7, 4, -6, 11,
					-- layer=2 filter=214 channel=69
					-10, -36, -7, 0, -11, 5, -59, -7, 7,
					-- layer=2 filter=214 channel=70
					3, 33, 55, -30, -3, 30, 1, 15, 10,
					-- layer=2 filter=214 channel=71
					3, 6, -19, -38, -8, -23, -20, 6, -30,
					-- layer=2 filter=214 channel=72
					46, 29, 5, -25, -18, 12, -16, -5, -12,
					-- layer=2 filter=214 channel=73
					-60, -29, 1, -15, -4, 7, -61, -8, -28,
					-- layer=2 filter=214 channel=74
					-37, -23, -12, -1, -19, -33, -2, 2, 15,
					-- layer=2 filter=214 channel=75
					-55, -32, -14, -11, -27, 3, 10, -7, -29,
					-- layer=2 filter=214 channel=76
					20, 10, 7, 20, 35, 16, -25, 11, 39,
					-- layer=2 filter=214 channel=77
					1, -2, -10, -8, 9, 8, 1, -8, 5,
					-- layer=2 filter=214 channel=78
					13, 7, -38, 38, 10, -24, 4, 1, -37,
					-- layer=2 filter=214 channel=79
					-7, -6, -1, 0, 9, 8, 7, -7, -3,
					-- layer=2 filter=214 channel=80
					18, 6, 4, 4, -42, -27, -23, -16, 14,
					-- layer=2 filter=214 channel=81
					8, -5, -6, 10, -6, 9, -1, -9, 12,
					-- layer=2 filter=214 channel=82
					4, -7, -4, -7, 2, -8, 1, -1, -12,
					-- layer=2 filter=214 channel=83
					-32, -12, 1, -26, -46, 31, -47, -6, 28,
					-- layer=2 filter=214 channel=84
					-2, 9, 0, 6, 9, 10, -6, 6, 6,
					-- layer=2 filter=214 channel=85
					-1, 6, 4, 7, -12, -12, -8, -6, -7,
					-- layer=2 filter=214 channel=86
					-7, 3, -8, -8, 5, 2, -8, 4, -7,
					-- layer=2 filter=214 channel=87
					30, 19, 11, 17, -2, 20, -9, 55, 5,
					-- layer=2 filter=214 channel=88
					-78, -54, -6, -17, -2, 28, -18, -30, 8,
					-- layer=2 filter=214 channel=89
					-20, 8, 23, -30, -8, 19, -24, -1, 6,
					-- layer=2 filter=214 channel=90
					5, 0, 7, 0, -1, 4, 0, 4, -4,
					-- layer=2 filter=214 channel=91
					-12, -13, 41, -48, -2, 27, 20, 26, -4,
					-- layer=2 filter=214 channel=92
					-23, 15, 40, -16, 14, 49, -39, -32, 12,
					-- layer=2 filter=214 channel=93
					-2, -98, -22, -32, -48, -40, -13, -55, -42,
					-- layer=2 filter=214 channel=94
					-57, -29, -7, -77, -29, 26, -20, -62, -3,
					-- layer=2 filter=214 channel=95
					-4, 2, -7, 0, 0, -2, -8, 10, 13,
					-- layer=2 filter=214 channel=96
					-6, -43, -11, -57, -53, -9, -29, -28, 0,
					-- layer=2 filter=214 channel=97
					17, 0, -25, 35, 30, -45, -16, 16, -22,
					-- layer=2 filter=214 channel=98
					6, 33, -5, -33, 0, 18, 17, 20, 8,
					-- layer=2 filter=214 channel=99
					13, -30, 32, -40, 14, 13, -21, 11, 9,
					-- layer=2 filter=214 channel=100
					-45, 22, 15, -23, -6, 8, -60, 59, 56,
					-- layer=2 filter=214 channel=101
					56, 25, -16, 24, -38, -64, 22, -42, -33,
					-- layer=2 filter=214 channel=102
					-36, -10, 4, -36, -18, -6, -17, -5, -16,
					-- layer=2 filter=214 channel=103
					2, -56, 0, 23, -20, 5, 36, -57, 34,
					-- layer=2 filter=214 channel=104
					-8, 50, -21, -10, 16, -8, -24, -19, -9,
					-- layer=2 filter=214 channel=105
					10, 12, 21, -21, 15, 0, 61, 31, 64,
					-- layer=2 filter=214 channel=106
					36, -2, -8, 21, 0, -58, 42, 23, -45,
					-- layer=2 filter=214 channel=107
					0, -15, 10, 13, -6, -12, -7, -9, 24,
					-- layer=2 filter=214 channel=108
					-40, -24, 1, -85, -2, -7, -27, -5, 12,
					-- layer=2 filter=214 channel=109
					6, 10, 0, 0, 10, 9, 8, -1, -3,
					-- layer=2 filter=214 channel=110
					-8, -17, -15, -18, -26, 17, -24, -7, 78,
					-- layer=2 filter=214 channel=111
					5, -3, 6, -6, -6, 2, -5, -2, 2,
					-- layer=2 filter=214 channel=112
					3, 15, -25, 10, -27, -38, 42, -30, -23,
					-- layer=2 filter=214 channel=113
					-39, 21, -9, -21, -14, 36, -15, -36, 19,
					-- layer=2 filter=214 channel=114
					-3, -25, -5, 0, 1, -24, -12, -16, -7,
					-- layer=2 filter=214 channel=115
					-8, 8, 4, -5, 0, -6, 1, 3, 0,
					-- layer=2 filter=214 channel=116
					-8, 14, -11, -6, -23, 15, 6, 32, 25,
					-- layer=2 filter=214 channel=117
					-15, 19, 36, -8, -53, 26, -27, -35, -4,
					-- layer=2 filter=214 channel=118
					4, 11, -15, 42, 26, -31, 0, 9, -2,
					-- layer=2 filter=214 channel=119
					2, -26, 14, -33, 17, 35, -40, 0, 43,
					-- layer=2 filter=214 channel=120
					-5, 0, -6, -4, -6, 0, -5, -3, 9,
					-- layer=2 filter=214 channel=121
					-1, 6, 0, -7, -7, -8, 2, -2, 5,
					-- layer=2 filter=214 channel=122
					-4, 0, 2, 3, 0, 6, 1, 12, 13,
					-- layer=2 filter=214 channel=123
					7, 32, 24, -6, 2, 11, -32, 23, 16,
					-- layer=2 filter=214 channel=124
					20, -26, 16, 63, -3, 36, -12, -23, 61,
					-- layer=2 filter=214 channel=125
					-4, -12, 4, 6, 2, 6, 0, 7, -2,
					-- layer=2 filter=214 channel=126
					42, -16, 43, -18, -54, 36, -18, -9, -27,
					-- layer=2 filter=214 channel=127
					-89, -8, 8, -24, 0, 28, -30, -2, 21,
					-- layer=2 filter=215 channel=0
					2, 0, 23, 16, 17, 24, 3, -23, -7,
					-- layer=2 filter=215 channel=1
					28, 17, 51, 24, -27, 5, -29, -8, -4,
					-- layer=2 filter=215 channel=2
					-3, 5, -1, 10, 7, 7, 6, 4, -5,
					-- layer=2 filter=215 channel=3
					-5, -1, -8, 9, 15, 23, 40, 29, -1,
					-- layer=2 filter=215 channel=4
					-9, -6, -1, -20, 0, 48, 10, 5, 13,
					-- layer=2 filter=215 channel=5
					-20, -3, -14, 25, -10, 1, 16, 0, 2,
					-- layer=2 filter=215 channel=6
					8, 5, -4, -47, -109, -49, -82, -23, -53,
					-- layer=2 filter=215 channel=7
					11, 16, 25, 18, 31, 15, 9, 1, 26,
					-- layer=2 filter=215 channel=8
					-6, 8, -2, -5, -6, -6, 4, 5, 0,
					-- layer=2 filter=215 channel=9
					-23, 9, -7, 13, 11, 29, 25, 16, 11,
					-- layer=2 filter=215 channel=10
					-1, 8, 29, 20, 21, 14, 22, 3, 5,
					-- layer=2 filter=215 channel=11
					-2, -37, -17, -6, -6, 7, 30, 3, 6,
					-- layer=2 filter=215 channel=12
					6, -2, 20, 16, -21, -27, -35, -17, -20,
					-- layer=2 filter=215 channel=13
					-7, -9, -4, -5, -2, -8, 6, 6, 7,
					-- layer=2 filter=215 channel=14
					-4, -9, 13, 25, -23, -30, -34, -38, -40,
					-- layer=2 filter=215 channel=15
					1, 51, 19, -3, 17, -40, 8, -48, -55,
					-- layer=2 filter=215 channel=16
					-44, -8, -55, -37, 3, 6, 20, 43, 19,
					-- layer=2 filter=215 channel=17
					4, -7, 6, -3, 0, 6, 5, -7, 6,
					-- layer=2 filter=215 channel=18
					-20, 39, 25, -4, 16, -26, 9, -10, 10,
					-- layer=2 filter=215 channel=19
					2, 52, 26, 4, -19, -41, -41, 15, -16,
					-- layer=2 filter=215 channel=20
					0, 2, -4, 2, 1, 0, 2, -7, -5,
					-- layer=2 filter=215 channel=21
					-5, -5, 11, 2, -14, -5, -2, 8, 22,
					-- layer=2 filter=215 channel=22
					7, 1, -7, 0, -5, 0, -1, -4, 0,
					-- layer=2 filter=215 channel=23
					-12, 9, 23, -18, -1, 8, -14, 16, -11,
					-- layer=2 filter=215 channel=24
					-18, -42, -15, -8, -15, 12, 10, 26, 19,
					-- layer=2 filter=215 channel=25
					-26, -58, -44, -13, -12, -26, 29, 21, 16,
					-- layer=2 filter=215 channel=26
					10, -2, 2, -7, -10, 1, 6, -8, 4,
					-- layer=2 filter=215 channel=27
					-13, -62, -45, 24, -8, 7, 46, 20, 33,
					-- layer=2 filter=215 channel=28
					0, 22, 9, 24, 20, 29, 28, -4, -34,
					-- layer=2 filter=215 channel=29
					12, 5, -8, -4, 13, -3, -3, 8, -4,
					-- layer=2 filter=215 channel=30
					-7, 4, -8, -25, -8, -17, -19, -7, -7,
					-- layer=2 filter=215 channel=31
					-67, 7, -8, -71, -51, -9, -29, -24, 3,
					-- layer=2 filter=215 channel=32
					5, 4, 10, 4, 9, 3, 4, 0, 4,
					-- layer=2 filter=215 channel=33
					0, -11, 28, 2, 33, 17, 25, 9, -6,
					-- layer=2 filter=215 channel=34
					10, 31, 17, -10, 24, -3, 15, 22, 39,
					-- layer=2 filter=215 channel=35
					11, 14, -20, 1, 23, -6, 49, -11, -42,
					-- layer=2 filter=215 channel=36
					9, 2, -2, 3, 0, 8, -11, -8, 6,
					-- layer=2 filter=215 channel=37
					-17, -23, -15, 10, -24, 13, 26, -3, 2,
					-- layer=2 filter=215 channel=38
					-6, -16, -9, 37, -9, -10, 44, 16, 6,
					-- layer=2 filter=215 channel=39
					-19, -4, -24, -21, 14, -2, 14, 31, 35,
					-- layer=2 filter=215 channel=40
					14, 28, -1, -11, 16, -11, 2, 61, 31,
					-- layer=2 filter=215 channel=41
					-3, 5, 6, 8, 7, 2, -4, -1, 9,
					-- layer=2 filter=215 channel=42
					-28, -15, -30, 2, 3, 15, 21, 40, 10,
					-- layer=2 filter=215 channel=43
					-17, 25, 2, 19, -19, 17, 36, 33, 11,
					-- layer=2 filter=215 channel=44
					6, 7, 0, -9, 5, -10, -2, -4, 8,
					-- layer=2 filter=215 channel=45
					0, -35, -39, -6, -7, 10, 16, 30, 52,
					-- layer=2 filter=215 channel=46
					13, 0, 31, 13, -1, 31, 13, 11, -9,
					-- layer=2 filter=215 channel=47
					-4, -8, -15, 18, 11, 26, 47, -2, -7,
					-- layer=2 filter=215 channel=48
					7, -5, 2, -6, -9, 0, 2, 12, 5,
					-- layer=2 filter=215 channel=49
					-38, 39, -16, -10, -16, -55, -46, -12, -17,
					-- layer=2 filter=215 channel=50
					20, 11, 10, 15, 24, 25, -10, -7, 9,
					-- layer=2 filter=215 channel=51
					-27, -27, -31, 7, -14, -15, 29, -1, -6,
					-- layer=2 filter=215 channel=52
					-41, -23, 9, 10, 9, -16, -29, -12, -30,
					-- layer=2 filter=215 channel=53
					-24, 76, 23, -14, 13, -52, -4, -46, -37,
					-- layer=2 filter=215 channel=54
					13, -1, -4, 0, -9, 3, 6, 16, 17,
					-- layer=2 filter=215 channel=55
					1, 7, -2, 4, 0, 4, -10, 7, -4,
					-- layer=2 filter=215 channel=56
					-21, -4, -23, 11, 9, 4, 33, 8, 20,
					-- layer=2 filter=215 channel=57
					-7, -13, 1, 5, -3, 0, -7, -6, 6,
					-- layer=2 filter=215 channel=58
					8, -7, 23, 17, -24, -33, -27, -2, -3,
					-- layer=2 filter=215 channel=59
					16, 11, -16, 8, 2, 0, -7, 3, -11,
					-- layer=2 filter=215 channel=60
					38, 21, -31, -4, -9, -63, -44, -35, -69,
					-- layer=2 filter=215 channel=61
					-28, -57, -42, -30, -56, -47, -97, -56, -58,
					-- layer=2 filter=215 channel=62
					13, 32, 1, 5, 25, -23, 3, -48, 10,
					-- layer=2 filter=215 channel=63
					-7, -4, -16, -3, 13, 7, -40, 2, -7,
					-- layer=2 filter=215 channel=64
					-39, 4, -9, -38, -1, 15, -35, 5, 20,
					-- layer=2 filter=215 channel=65
					-26, -21, -49, -49, -90, -58, -103, -71, -29,
					-- layer=2 filter=215 channel=66
					22, 32, 18, 32, -59, 7, 15, -8, -3,
					-- layer=2 filter=215 channel=67
					29, 27, 64, -4, 22, 58, 20, 20, 18,
					-- layer=2 filter=215 channel=68
					-8, 7, 2, 0, -4, 8, 7, 6, 11,
					-- layer=2 filter=215 channel=69
					-2, 2, -9, 3, -9, 7, -25, 11, 17,
					-- layer=2 filter=215 channel=70
					-3, 1, -26, 7, 15, -13, 33, 7, 3,
					-- layer=2 filter=215 channel=71
					-21, -60, -41, -20, -5, 23, 27, 47, 58,
					-- layer=2 filter=215 channel=72
					-5, 15, 17, -15, 19, -3, -16, -52, -53,
					-- layer=2 filter=215 channel=73
					-53, 6, -23, -49, -61, -18, 20, -25, -16,
					-- layer=2 filter=215 channel=74
					17, 16, 25, 19, 11, 22, -22, 7, -27,
					-- layer=2 filter=215 channel=75
					-24, -4, 3, 33, 9, -6, -34, -30, -8,
					-- layer=2 filter=215 channel=76
					-39, 0, -5, 7, -9, -11, -2, -30, -20,
					-- layer=2 filter=215 channel=77
					5, -2, 4, -3, -4, 3, 11, 4, 8,
					-- layer=2 filter=215 channel=78
					0, -3, -45, -10, -6, -3, 10, -23, -16,
					-- layer=2 filter=215 channel=79
					-9, 3, -5, 0, 4, 1, 6, 6, -4,
					-- layer=2 filter=215 channel=80
					-19, 3, 22, -23, -17, 45, 13, 20, 10,
					-- layer=2 filter=215 channel=81
					7, 4, -2, -1, 3, 0, -1, -10, 9,
					-- layer=2 filter=215 channel=82
					0, 6, 0, -6, -8, -5, 3, -8, -2,
					-- layer=2 filter=215 channel=83
					-9, 2, 4, -18, -11, 5, -21, 4, 28,
					-- layer=2 filter=215 channel=84
					-4, -6, 2, 7, -10, 3, -2, 7, 6,
					-- layer=2 filter=215 channel=85
					0, -1, -8, 7, 19, 9, -2, 6, 10,
					-- layer=2 filter=215 channel=86
					6, 7, -16, -4, 12, -7, -14, -9, -10,
					-- layer=2 filter=215 channel=87
					42, 38, 31, -4, 53, 36, 45, -24, 11,
					-- layer=2 filter=215 channel=88
					6, 15, 29, 1, 9, 4, -45, -18, -10,
					-- layer=2 filter=215 channel=89
					6, 18, 21, 27, 4, -5, -3, -45, -72,
					-- layer=2 filter=215 channel=90
					-9, -7, 0, -9, -6, -9, 1, 7, 8,
					-- layer=2 filter=215 channel=91
					28, 25, -3, 41, 34, 17, 12, -11, -53,
					-- layer=2 filter=215 channel=92
					26, -11, 15, 28, -19, -27, 6, -22, -33,
					-- layer=2 filter=215 channel=93
					7, 34, -33, -33, 48, -41, -44, -69, 10,
					-- layer=2 filter=215 channel=94
					3, 26, 6, -3, -23, -36, -112, -41, -96,
					-- layer=2 filter=215 channel=95
					3, 6, 11, 10, 0, 0, 12, 14, 18,
					-- layer=2 filter=215 channel=96
					-15, 13, 1, -55, -16, -25, -131, -55, -59,
					-- layer=2 filter=215 channel=97
					4, 6, -2, 4, 10, 37, 13, 19, 7,
					-- layer=2 filter=215 channel=98
					4, -14, -25, 7, 4, 25, 22, -22, -27,
					-- layer=2 filter=215 channel=99
					-6, 21, -42, 5, -27, -77, -61, -84, -43,
					-- layer=2 filter=215 channel=100
					3, -12, 27, -12, -6, -6, 18, 12, -22,
					-- layer=2 filter=215 channel=101
					-27, -98, -65, 4, -4, -1, 30, 32, 33,
					-- layer=2 filter=215 channel=102
					-32, 19, -57, -68, 13, -84, -89, -77, -32,
					-- layer=2 filter=215 channel=103
					14, 6, 34, 19, 35, 29, -21, -24, -32,
					-- layer=2 filter=215 channel=104
					-17, 18, 42, -23, -25, -37, -53, -56, -67,
					-- layer=2 filter=215 channel=105
					7, -9, 22, 38, 15, 29, 43, -5, 15,
					-- layer=2 filter=215 channel=106
					-25, -34, -30, 3, 0, -1, 37, 26, 3,
					-- layer=2 filter=215 channel=107
					21, -23, -34, 17, -9, -12, -22, -33, -23,
					-- layer=2 filter=215 channel=108
					-26, 1, -34, -4, 4, 4, 0, 14, 35,
					-- layer=2 filter=215 channel=109
					-3, 0, 1, 15, -9, -4, 8, -8, 6,
					-- layer=2 filter=215 channel=110
					-50, -31, -22, -37, 14, 7, -35, -6, -23,
					-- layer=2 filter=215 channel=111
					-3, -5, -7, 4, 3, -13, -11, -4, 3,
					-- layer=2 filter=215 channel=112
					-16, -28, -33, 38, 1, -3, 44, 19, 17,
					-- layer=2 filter=215 channel=113
					-4, -36, 5, -14, 12, -21, -30, -33, -28,
					-- layer=2 filter=215 channel=114
					-3, -1, 5, -1, 6, 5, 2, 16, 6,
					-- layer=2 filter=215 channel=115
					9, 7, 8, 3, 0, 5, 8, -8, 0,
					-- layer=2 filter=215 channel=116
					10, 53, 32, -3, 55, 20, 27, -14, 2,
					-- layer=2 filter=215 channel=117
					38, 42, 13, 29, 25, -11, -42, -41, -49,
					-- layer=2 filter=215 channel=118
					-18, 2, 29, -23, 5, 41, 21, 6, -21,
					-- layer=2 filter=215 channel=119
					35, 4, 0, 47, -9, 6, 61, 18, 21,
					-- layer=2 filter=215 channel=120
					-8, 9, 1, 0, -6, 9, 0, 8, 1,
					-- layer=2 filter=215 channel=121
					-9, 7, -2, -8, 6, 8, -5, 6, 2,
					-- layer=2 filter=215 channel=122
					6, 12, -2, 0, -5, -7, 0, 4, -14,
					-- layer=2 filter=215 channel=123
					37, 25, 17, 21, 38, 14, -15, -8, 1,
					-- layer=2 filter=215 channel=124
					12, 63, 46, 38, 56, 0, 40, 0, 11,
					-- layer=2 filter=215 channel=125
					-3, -9, 0, -6, -3, -3, 10, 0, -3,
					-- layer=2 filter=215 channel=126
					60, 28, 51, -10, -38, 11, -43, 39, -84,
					-- layer=2 filter=215 channel=127
					-15, -7, 0, -12, -17, 11, -18, 2, 18,
					-- layer=2 filter=216 channel=0
					20, 4, 10, 6, 14, -8, 23, -1, 2,
					-- layer=2 filter=216 channel=1
					-29, 11, -1, 19, -6, 18, 18, 13, 7,
					-- layer=2 filter=216 channel=2
					-7, 11, -3, 5, -6, -9, -8, -3, 3,
					-- layer=2 filter=216 channel=3
					38, 18, 0, 24, -25, -10, -8, -11, 1,
					-- layer=2 filter=216 channel=4
					-12, -26, -37, 1, -18, -1, -2, 6, 21,
					-- layer=2 filter=216 channel=5
					4, -8, 9, 10, 1, -25, 10, -9, 5,
					-- layer=2 filter=216 channel=6
					10, -12, -16, 10, 30, 24, 48, 5, 16,
					-- layer=2 filter=216 channel=7
					43, 41, 12, 22, 38, -18, 0, -1, 1,
					-- layer=2 filter=216 channel=8
					2, -6, 4, 8, 1, 8, 2, -6, 2,
					-- layer=2 filter=216 channel=9
					38, 24, -8, 20, 17, 23, -17, -24, -14,
					-- layer=2 filter=216 channel=10
					49, 0, 15, 42, 4, -5, -10, -15, -2,
					-- layer=2 filter=216 channel=11
					22, 4, -6, 15, 7, -16, 19, 20, -3,
					-- layer=2 filter=216 channel=12
					5, -6, 10, 53, 38, 26, 17, 11, -2,
					-- layer=2 filter=216 channel=13
					7, 8, -6, 3, 4, -8, 9, 0, 6,
					-- layer=2 filter=216 channel=14
					15, 1, -11, 1, -7, 25, 34, 13, 6,
					-- layer=2 filter=216 channel=15
					-27, -2, -6, 8, -11, -18, 65, 59, 2,
					-- layer=2 filter=216 channel=16
					-2, -4, 34, -17, -46, -19, -48, -53, -69,
					-- layer=2 filter=216 channel=17
					-5, 5, 4, -9, -4, 10, -10, 1, -5,
					-- layer=2 filter=216 channel=18
					-94, -29, -8, -45, -61, -1, -61, -9, -5,
					-- layer=2 filter=216 channel=19
					4, 0, -10, 19, -6, -1, -10, -20, 19,
					-- layer=2 filter=216 channel=20
					9, -8, -2, -3, -4, -2, 3, 5, 8,
					-- layer=2 filter=216 channel=21
					4, 21, 6, 12, -8, 14, -2, 5, 8,
					-- layer=2 filter=216 channel=22
					8, 0, 4, 9, 0, -1, -9, -3, -4,
					-- layer=2 filter=216 channel=23
					-12, 24, -7, -64, 3, -37, -53, -26, -26,
					-- layer=2 filter=216 channel=24
					37, 9, 32, 29, 12, 8, -31, -13, 10,
					-- layer=2 filter=216 channel=25
					25, 19, 15, -6, -8, 4, 1, -5, 20,
					-- layer=2 filter=216 channel=26
					0, -9, -3, 2, 4, -10, -2, 5, 7,
					-- layer=2 filter=216 channel=27
					26, -4, 0, 29, 9, 28, 24, 0, 40,
					-- layer=2 filter=216 channel=28
					-12, 8, -20, -8, -2, -3, 5, -4, 5,
					-- layer=2 filter=216 channel=29
					2, 5, 11, -1, -5, -2, -8, -1, -6,
					-- layer=2 filter=216 channel=30
					-33, 10, -4, -22, 16, -10, -50, -30, -7,
					-- layer=2 filter=216 channel=31
					-45, -8, 43, 11, 70, -25, 52, 38, 18,
					-- layer=2 filter=216 channel=32
					-3, -1, -3, -7, 1, -8, -3, -4, -2,
					-- layer=2 filter=216 channel=33
					13, -23, -23, 15, -4, -1, 31, -2, -2,
					-- layer=2 filter=216 channel=34
					-69, -28, -17, -36, -20, 50, -55, -14, 0,
					-- layer=2 filter=216 channel=35
					-1, 0, 10, 9, 7, 0, -25, -27, -10,
					-- layer=2 filter=216 channel=36
					1, -3, 3, -1, 0, 6, -2, -1, -18,
					-- layer=2 filter=216 channel=37
					-13, -1, -5, -6, 6, -2, -4, 5, 0,
					-- layer=2 filter=216 channel=38
					24, 0, -6, 16, 4, 8, 30, -7, 10,
					-- layer=2 filter=216 channel=39
					-9, 29, 46, -15, -27, -82, -21, -35, 1,
					-- layer=2 filter=216 channel=40
					-40, -28, 15, -15, -2, 34, 17, -11, 34,
					-- layer=2 filter=216 channel=41
					7, 2, -6, 3, -7, -3, 0, 0, 5,
					-- layer=2 filter=216 channel=42
					19, -15, -11, -18, -27, -41, -18, -33, -36,
					-- layer=2 filter=216 channel=43
					-13, -5, 4, 2, -57, -5, -19, -29, 3,
					-- layer=2 filter=216 channel=44
					-2, 2, 9, -6, 0, -6, 4, -3, -2,
					-- layer=2 filter=216 channel=45
					17, 0, 48, -69, -34, 32, -38, -44, 2,
					-- layer=2 filter=216 channel=46
					4, -8, 14, 8, -26, -2, 8, 18, 10,
					-- layer=2 filter=216 channel=47
					14, -5, -8, -9, -8, -8, 9, -8, -32,
					-- layer=2 filter=216 channel=48
					-2, 9, 0, 8, -2, 0, -4, 11, -4,
					-- layer=2 filter=216 channel=49
					-37, 10, 2, 2, -16, -31, -19, 13, 15,
					-- layer=2 filter=216 channel=50
					2, 7, 3, 8, 11, 3, 20, 2, -8,
					-- layer=2 filter=216 channel=51
					10, 5, -4, -2, -8, -5, 6, 17, 8,
					-- layer=2 filter=216 channel=52
					-5, 30, 8, 6, -16, 12, 33, 4, -5,
					-- layer=2 filter=216 channel=53
					12, -14, -16, 19, 23, -40, 55, -16, 12,
					-- layer=2 filter=216 channel=54
					-2, 3, 22, 10, 0, 12, 20, 35, -19,
					-- layer=2 filter=216 channel=55
					-8, -2, 0, 4, 0, -4, 10, 3, -12,
					-- layer=2 filter=216 channel=56
					18, -8, -2, 16, -2, -9, 0, 9, -1,
					-- layer=2 filter=216 channel=57
					9, 0, 8, 11, 4, 5, 14, 3, 3,
					-- layer=2 filter=216 channel=58
					-13, -10, 9, 62, 52, 29, 29, 16, 15,
					-- layer=2 filter=216 channel=59
					-26, -25, -17, 0, -5, -7, -8, -3, -8,
					-- layer=2 filter=216 channel=60
					-33, 2, 2, -1, -31, -20, 11, -20, 2,
					-- layer=2 filter=216 channel=61
					-13, 36, 29, -23, -19, -1, -32, -24, -49,
					-- layer=2 filter=216 channel=62
					-44, -12, -34, -30, -24, -4, -4, 9, 19,
					-- layer=2 filter=216 channel=63
					24, 12, 25, -7, -22, -12, 12, -9, -39,
					-- layer=2 filter=216 channel=64
					22, 24, 0, 10, -8, -59, -46, -20, -24,
					-- layer=2 filter=216 channel=65
					-15, 44, 9, 8, 6, 22, 3, 20, -13,
					-- layer=2 filter=216 channel=66
					74, 15, -1, -52, 5, -36, -46, -5, -22,
					-- layer=2 filter=216 channel=67
					14, -37, -7, 21, -7, -3, -16, -59, -9,
					-- layer=2 filter=216 channel=68
					-6, 6, 8, -6, 2, -8, -5, -3, -3,
					-- layer=2 filter=216 channel=69
					8, -5, -16, -46, -53, -38, -19, -51, -22,
					-- layer=2 filter=216 channel=70
					15, 9, 32, 21, 20, 48, 4, 32, 20,
					-- layer=2 filter=216 channel=71
					7, -19, -12, 13, -31, 12, -10, -17, 12,
					-- layer=2 filter=216 channel=72
					71, 31, -32, 19, 7, -16, 31, 15, 1,
					-- layer=2 filter=216 channel=73
					26, 42, 75, -14, -10, -10, 1, -13, -17,
					-- layer=2 filter=216 channel=74
					35, 3, 24, 38, 10, -17, 10, -8, -61,
					-- layer=2 filter=216 channel=75
					-2, 13, -42, 39, 14, 21, 23, -9, -27,
					-- layer=2 filter=216 channel=76
					-17, -19, 16, 18, 42, 28, 14, 27, -30,
					-- layer=2 filter=216 channel=77
					3, -2, -7, -8, 9, -4, 3, 5, 4,
					-- layer=2 filter=216 channel=78
					-14, 0, -19, 16, 2, -17, -12, 24, -3,
					-- layer=2 filter=216 channel=79
					-4, 9, -5, -7, 10, -4, 9, -5, -8,
					-- layer=2 filter=216 channel=80
					0, 10, 8, -18, -4, -46, -62, -49, -39,
					-- layer=2 filter=216 channel=81
					4, 1, -7, 0, 1, 5, -3, -8, 1,
					-- layer=2 filter=216 channel=82
					8, 0, -12, 0, 2, 6, 0, 0, 0,
					-- layer=2 filter=216 channel=83
					-28, 30, -5, -49, -6, 44, -41, -7, 35,
					-- layer=2 filter=216 channel=84
					7, 0, 0, -8, -7, 10, -3, -4, 7,
					-- layer=2 filter=216 channel=85
					0, 9, 5, 15, 1, 11, 8, 2, 8,
					-- layer=2 filter=216 channel=86
					-7, -14, -5, -10, -13, -13, -7, -7, 4,
					-- layer=2 filter=216 channel=87
					-34, -50, -14, -38, -13, -23, -8, -17, -19,
					-- layer=2 filter=216 channel=88
					-17, -30, 12, -44, -12, 10, -20, -12, -44,
					-- layer=2 filter=216 channel=89
					15, -12, -27, 7, 23, -2, 23, 23, -12,
					-- layer=2 filter=216 channel=90
					0, 0, -4, 2, 0, -9, -3, 0, -1,
					-- layer=2 filter=216 channel=91
					4, -36, -38, 40, -17, -55, 49, 0, -4,
					-- layer=2 filter=216 channel=92
					2, -15, -12, 16, 3, -10, 38, 10, -8,
					-- layer=2 filter=216 channel=93
					-8, -33, -37, 2, -34, -15, 29, -61, -21,
					-- layer=2 filter=216 channel=94
					9, 15, 9, -3, 24, -5, 11, -4, 0,
					-- layer=2 filter=216 channel=95
					-20, -6, -17, -4, -4, -4, -18, -5, -4,
					-- layer=2 filter=216 channel=96
					-34, -1, 16, -30, 39, 38, 1, 24, 34,
					-- layer=2 filter=216 channel=97
					53, -12, 3, 47, 9, -3, 17, -18, -17,
					-- layer=2 filter=216 channel=98
					26, 26, 21, -1, -3, 4, 6, 5, 10,
					-- layer=2 filter=216 channel=99
					11, 13, -20, 20, 18, 16, 7, 14, -27,
					-- layer=2 filter=216 channel=100
					-7, -5, -14, 7, 1, 8, -16, -31, 0,
					-- layer=2 filter=216 channel=101
					-1, -2, 13, -3, -13, -12, 8, -2, -4,
					-- layer=2 filter=216 channel=102
					-38, 0, -6, 23, 6, -2, -6, -12, -29,
					-- layer=2 filter=216 channel=103
					-18, -12, 22, 19, 20, 14, 14, 34, 68,
					-- layer=2 filter=216 channel=104
					-82, -17, -19, -15, -13, -14, 3, 30, 5,
					-- layer=2 filter=216 channel=105
					-35, 1, -5, -32, 37, -12, -72, 38, -13,
					-- layer=2 filter=216 channel=106
					32, 7, -16, 20, 21, -42, 7, -10, -3,
					-- layer=2 filter=216 channel=107
					31, 34, 30, -50, -3, -2, -13, 12, 55,
					-- layer=2 filter=216 channel=108
					5, 7, 5, 3, 7, 40, 13, 6, 24,
					-- layer=2 filter=216 channel=109
					-3, 11, 3, -9, 0, 1, -1, -4, -3,
					-- layer=2 filter=216 channel=110
					7, 33, 19, -1, -2, -40, -54, -1, 0,
					-- layer=2 filter=216 channel=111
					4, 6, -6, 4, 7, -4, 10, -2, 5,
					-- layer=2 filter=216 channel=112
					15, 0, 26, 15, 12, -21, -20, -9, 24,
					-- layer=2 filter=216 channel=113
					-15, 23, 14, 14, -18, -18, -8, 7, -7,
					-- layer=2 filter=216 channel=114
					10, -2, 13, 12, 12, 13, 16, 19, 25,
					-- layer=2 filter=216 channel=115
					8, 2, 5, 9, -7, 1, 6, -4, 8,
					-- layer=2 filter=216 channel=116
					-71, 12, 21, -32, -30, 17, -16, 1, 5,
					-- layer=2 filter=216 channel=117
					33, 36, 2, -14, 41, 46, 12, -4, -17,
					-- layer=2 filter=216 channel=118
					-13, -19, 8, -4, -14, -2, -28, -8, 0,
					-- layer=2 filter=216 channel=119
					-38, -38, -20, -35, -82, -11, -50, -56, -42,
					-- layer=2 filter=216 channel=120
					5, 4, -3, -10, 0, 0, 3, 4, 4,
					-- layer=2 filter=216 channel=121
					-3, -7, -3, 5, -9, -4, 8, -6, -4,
					-- layer=2 filter=216 channel=122
					5, 9, 5, -2, 14, -10, 10, 5, 12,
					-- layer=2 filter=216 channel=123
					38, -1, -7, 13, 0, -7, 14, -9, -22,
					-- layer=2 filter=216 channel=124
					7, -61, -45, -34, 28, -25, 35, 31, -27,
					-- layer=2 filter=216 channel=125
					-8, 3, -11, 9, 6, 5, 0, 2, -7,
					-- layer=2 filter=216 channel=126
					-28, -77, -43, -11, -46, 9, -36, -60, -51,
					-- layer=2 filter=216 channel=127
					-18, 3, 14, -28, 10, 65, -5, 6, -3,
					-- layer=2 filter=217 channel=0
					-7, -15, -8, -17, -21, 3, -4, 7, 1,
					-- layer=2 filter=217 channel=1
					-9, -29, 3, -12, -26, -16, -44, 1, -23,
					-- layer=2 filter=217 channel=2
					1, 2, -2, -8, -7, -1, 8, 4, -6,
					-- layer=2 filter=217 channel=3
					-7, 2, 8, 18, -4, -25, -6, 1, -19,
					-- layer=2 filter=217 channel=4
					3, -12, 1, -48, -25, 19, -63, -35, -14,
					-- layer=2 filter=217 channel=5
					-12, 8, -13, 8, -8, 4, -13, 15, -11,
					-- layer=2 filter=217 channel=6
					26, 0, 4, 22, -14, -23, 37, 35, 7,
					-- layer=2 filter=217 channel=7
					-26, -10, 13, -36, -5, 38, -11, -47, 0,
					-- layer=2 filter=217 channel=8
					5, -5, 9, 4, -5, -6, -10, 1, 4,
					-- layer=2 filter=217 channel=9
					6, 30, 12, -15, -10, 14, -35, -23, 16,
					-- layer=2 filter=217 channel=10
					-14, 3, 26, 21, -10, 9, -26, 5, -2,
					-- layer=2 filter=217 channel=11
					-7, -9, -6, 23, 19, -7, 33, 21, 7,
					-- layer=2 filter=217 channel=12
					7, -5, 7, -3, -30, -14, -8, -3, -16,
					-- layer=2 filter=217 channel=13
					1, 1, 10, -3, 4, -4, -10, 7, -7,
					-- layer=2 filter=217 channel=14
					-1, -4, 4, 0, 15, 16, 13, 23, 4,
					-- layer=2 filter=217 channel=15
					24, 8, -58, 21, 28, -26, 31, -5, -48,
					-- layer=2 filter=217 channel=16
					-9, -19, 0, -70, 3, 63, -81, -17, 55,
					-- layer=2 filter=217 channel=17
					0, 4, -4, -4, -6, 4, -1, 9, 8,
					-- layer=2 filter=217 channel=18
					-5, 27, 2, -5, 22, -17, -3, -25, -50,
					-- layer=2 filter=217 channel=19
					-27, -26, -22, -15, -34, -14, -37, -10, -44,
					-- layer=2 filter=217 channel=20
					-6, 5, 5, -3, 8, -1, -6, -6, 2,
					-- layer=2 filter=217 channel=21
					5, -7, -13, -6, 7, -9, 2, 7, -2,
					-- layer=2 filter=217 channel=22
					-2, 1, 0, -2, 4, 5, 0, 0, 4,
					-- layer=2 filter=217 channel=23
					-9, -9, 18, -17, -30, 62, -62, -30, 9,
					-- layer=2 filter=217 channel=24
					-4, -7, 17, -32, 0, 15, -8, -15, 5,
					-- layer=2 filter=217 channel=25
					-18, -8, 1, 2, 4, 13, 32, 29, 13,
					-- layer=2 filter=217 channel=26
					-2, 8, 0, -3, 1, -4, -7, 0, -12,
					-- layer=2 filter=217 channel=27
					11, 12, 26, 30, 32, 14, 6, 9, -1,
					-- layer=2 filter=217 channel=28
					-27, 10, 17, 0, -20, 5, -19, 1, 17,
					-- layer=2 filter=217 channel=29
					0, 11, -8, -9, 2, 9, -6, -9, -4,
					-- layer=2 filter=217 channel=30
					-18, 8, 13, -12, -9, 16, -27, -35, -30,
					-- layer=2 filter=217 channel=31
					38, 2, 7, -1, 20, 15, 44, 55, 5,
					-- layer=2 filter=217 channel=32
					-8, 7, -4, 0, -8, 8, 1, -9, 6,
					-- layer=2 filter=217 channel=33
					53, 29, 16, 17, 19, 18, -21, 0, -41,
					-- layer=2 filter=217 channel=34
					-2, 48, 52, 21, 39, 38, -22, 17, 35,
					-- layer=2 filter=217 channel=35
					-37, 17, 14, 5, 24, 26, -21, 0, 8,
					-- layer=2 filter=217 channel=36
					-1, 10, 13, 11, 2, 11, -6, -7, 5,
					-- layer=2 filter=217 channel=37
					-7, 0, -18, 24, 12, 0, 5, 15, -3,
					-- layer=2 filter=217 channel=38
					-20, 2, -14, 3, 3, 15, -28, -12, -11,
					-- layer=2 filter=217 channel=39
					14, -7, 41, -25, 21, 72, -4, -6, 9,
					-- layer=2 filter=217 channel=40
					3, 29, 9, -22, 57, -2, -24, 12, -73,
					-- layer=2 filter=217 channel=41
					2, 0, 8, 3, 4, -7, -8, 6, -6,
					-- layer=2 filter=217 channel=42
					-3, -14, 34, -23, -10, 51, -37, -10, 51,
					-- layer=2 filter=217 channel=43
					-8, 25, 36, 3, 63, -21, -30, -26, -71,
					-- layer=2 filter=217 channel=44
					5, 9, 8, -8, 2, -9, -6, 11, -6,
					-- layer=2 filter=217 channel=45
					25, -8, 20, 17, -13, 10, 23, -30, -53,
					-- layer=2 filter=217 channel=46
					-19, -19, 2, -2, 7, 32, -30, -7, 19,
					-- layer=2 filter=217 channel=47
					-11, 14, 3, 6, -12, 30, -32, 15, 10,
					-- layer=2 filter=217 channel=48
					5, 6, -3, -12, -5, -3, -1, 1, -5,
					-- layer=2 filter=217 channel=49
					-47, -30, -18, -52, 4, 19, 27, 0, -26,
					-- layer=2 filter=217 channel=50
					-13, 17, -10, 0, -13, 12, 3, -2, 4,
					-- layer=2 filter=217 channel=51
					-23, -21, -16, 0, -8, -15, 16, 21, -9,
					-- layer=2 filter=217 channel=52
					-7, 0, -33, -16, -8, -15, 21, 1, 17,
					-- layer=2 filter=217 channel=53
					2, 49, -40, 18, -10, -18, -37, -21, -30,
					-- layer=2 filter=217 channel=54
					-18, -21, -33, -1, -14, 20, 13, 22, 24,
					-- layer=2 filter=217 channel=55
					12, -5, 3, 14, -8, 2, 5, -4, 10,
					-- layer=2 filter=217 channel=56
					-28, -12, -4, 11, 20, -1, 7, 21, 3,
					-- layer=2 filter=217 channel=57
					0, -6, 4, 5, 10, -2, 4, -3, 3,
					-- layer=2 filter=217 channel=58
					23, -3, 24, -5, -8, -2, -9, 13, -20,
					-- layer=2 filter=217 channel=59
					66, 48, 16, 9, 11, 23, -21, 5, -48,
					-- layer=2 filter=217 channel=60
					2, 14, -45, 3, -7, -14, 4, 31, -33,
					-- layer=2 filter=217 channel=61
					55, 0, -21, -13, 0, -5, 0, -10, -31,
					-- layer=2 filter=217 channel=62
					-41, -7, 15, 0, -7, -17, 11, 22, 17,
					-- layer=2 filter=217 channel=63
					30, -5, 15, -19, -8, 37, 15, -13, 12,
					-- layer=2 filter=217 channel=64
					-14, -11, -5, -53, -12, 37, -30, -9, 57,
					-- layer=2 filter=217 channel=65
					27, 0, -7, 44, -11, -11, 9, -12, 4,
					-- layer=2 filter=217 channel=66
					-39, 8, 29, 9, 11, 3, -20, -48, 20,
					-- layer=2 filter=217 channel=67
					-1, 6, 2, -24, -19, -26, -54, -63, -30,
					-- layer=2 filter=217 channel=68
					1, -8, 0, -6, 0, 9, 1, 6, 8,
					-- layer=2 filter=217 channel=69
					-18, -10, 16, -35, 8, 52, -12, 9, 56,
					-- layer=2 filter=217 channel=70
					-24, 6, -16, 16, 20, 30, 2, 13, -4,
					-- layer=2 filter=217 channel=71
					-9, -18, -12, 1, -6, -28, 8, -15, -23,
					-- layer=2 filter=217 channel=72
					-32, -17, 8, 12, 26, -5, -29, -15, 9,
					-- layer=2 filter=217 channel=73
					25, 5, 103, 0, 19, 11, 2, 1, 19,
					-- layer=2 filter=217 channel=74
					25, -2, 17, -31, -29, 3, -48, -72, -19,
					-- layer=2 filter=217 channel=75
					-30, -37, -17, -27, -30, -15, -38, -30, -27,
					-- layer=2 filter=217 channel=76
					25, 0, -23, 41, 56, -21, 9, -27, -43,
					-- layer=2 filter=217 channel=77
					-2, 3, 2, -4, 1, -6, -7, 8, 0,
					-- layer=2 filter=217 channel=78
					-39, -11, 10, 9, -3, 3, 25, 21, 1,
					-- layer=2 filter=217 channel=79
					4, 4, 5, 5, -8, -3, 3, -1, 5,
					-- layer=2 filter=217 channel=80
					11, -10, 0, -20, -10, 28, -37, -23, 12,
					-- layer=2 filter=217 channel=81
					2, -2, 9, 5, 5, 5, 2, 6, 12,
					-- layer=2 filter=217 channel=82
					-4, -5, 1, 3, -6, 7, -4, 2, 7,
					-- layer=2 filter=217 channel=83
					8, -20, -22, -13, -35, 17, -36, -31, -37,
					-- layer=2 filter=217 channel=84
					9, 8, -6, -8, 5, -1, 5, 0, -2,
					-- layer=2 filter=217 channel=85
					2, -1, 7, -2, 13, 12, 7, -5, -3,
					-- layer=2 filter=217 channel=86
					-6, -5, -7, -8, -11, -16, -10, -10, 6,
					-- layer=2 filter=217 channel=87
					35, 44, -11, 15, 58, -35, -1, 5, 13,
					-- layer=2 filter=217 channel=88
					35, 20, -1, 10, 6, -1, 6, -18, 9,
					-- layer=2 filter=217 channel=89
					17, 4, 16, -6, 34, -4, -19, 0, -6,
					-- layer=2 filter=217 channel=90
					6, 0, 5, -1, -7, -11, 0, -2, -8,
					-- layer=2 filter=217 channel=91
					20, -8, 17, 1, -11, -1, -17, -22, -3,
					-- layer=2 filter=217 channel=92
					-10, -15, 9, 14, -3, -11, -31, 4, -23,
					-- layer=2 filter=217 channel=93
					-17, -33, 52, 19, -6, 15, -40, 31, 1,
					-- layer=2 filter=217 channel=94
					24, 37, -12, -20, -36, 5, -26, -15, -3,
					-- layer=2 filter=217 channel=95
					1, 4, -14, 7, 4, -14, -4, 9, 4,
					-- layer=2 filter=217 channel=96
					43, -58, -36, 67, -4, -40, 27, 47, 26,
					-- layer=2 filter=217 channel=97
					0, 6, 0, -34, 51, 23, -24, -7, 12,
					-- layer=2 filter=217 channel=98
					-19, 21, -5, 0, -4, 22, 5, 21, 36,
					-- layer=2 filter=217 channel=99
					5, -1, -40, 28, -44, -13, -4, 25, -5,
					-- layer=2 filter=217 channel=100
					29, 0, 2, -2, 31, 51, -25, -4, -19,
					-- layer=2 filter=217 channel=101
					-23, 1, -4, 44, 9, -15, 11, 11, -17,
					-- layer=2 filter=217 channel=102
					-1, -28, -36, 26, -46, -17, 22, 17, 31,
					-- layer=2 filter=217 channel=103
					-38, -48, -52, 8, -23, -17, 5, 8, -39,
					-- layer=2 filter=217 channel=104
					14, 4, -19, -6, -10, -1, 2, -28, 0,
					-- layer=2 filter=217 channel=105
					16, 101, 22, -6, 45, 10, 12, 52, 20,
					-- layer=2 filter=217 channel=106
					7, -11, 27, 45, -19, 17, 0, -1, 12,
					-- layer=2 filter=217 channel=107
					0, -68, -20, -33, 7, -6, -10, -14, -2,
					-- layer=2 filter=217 channel=108
					-5, -17, -23, 23, -11, 4, 3, -13, -41,
					-- layer=2 filter=217 channel=109
					-4, 4, 1, 2, -6, -4, 1, -13, -8,
					-- layer=2 filter=217 channel=110
					-89, -42, 7, -41, -42, 51, -37, -36, 48,
					-- layer=2 filter=217 channel=111
					-7, 0, -2, -4, 1, 0, -6, 7, 5,
					-- layer=2 filter=217 channel=112
					36, -12, -41, -15, -10, 10, -4, 12, -25,
					-- layer=2 filter=217 channel=113
					-2, -31, 4, -6, -12, 12, -31, -7, -19,
					-- layer=2 filter=217 channel=114
					-8, -3, -3, -7, -14, 1, -10, -11, 0,
					-- layer=2 filter=217 channel=115
					-1, 7, 1, 12, -7, 6, 3, -3, -9,
					-- layer=2 filter=217 channel=116
					17, 45, -25, 43, 36, -76, 25, 18, 2,
					-- layer=2 filter=217 channel=117
					-27, -20, -24, -28, 7, 9, -29, -66, 0,
					-- layer=2 filter=217 channel=118
					-32, -15, 24, 0, 26, 7, -11, -1, -14,
					-- layer=2 filter=217 channel=119
					-12, -1, 14, -39, -2, 42, -40, -11, 5,
					-- layer=2 filter=217 channel=120
					2, 9, 3, -1, -10, -10, 8, -2, 0,
					-- layer=2 filter=217 channel=121
					-3, 2, -4, -7, 10, -5, -6, 7, -4,
					-- layer=2 filter=217 channel=122
					5, -4, 7, 0, -1, 3, -1, -6, 0,
					-- layer=2 filter=217 channel=123
					-40, -1, 18, -13, -18, -7, -17, -38, 7,
					-- layer=2 filter=217 channel=124
					-8, -39, -57, -31, -13, -2, -58, 0, -76,
					-- layer=2 filter=217 channel=125
					1, 9, -7, -4, 6, 9, 2, -3, 0,
					-- layer=2 filter=217 channel=126
					19, -17, 9, 6, 13, 8, 24, -39, -12,
					-- layer=2 filter=217 channel=127
					3, -4, -8, -8, 14, -4, -30, 11, -17,
					-- layer=2 filter=218 channel=0
					-14, -15, -16, -14, 5, -4, 5, -2, 1,
					-- layer=2 filter=218 channel=1
					2, 18, -3, 45, 13, -20, -24, -11, -2,
					-- layer=2 filter=218 channel=2
					7, -3, 8, -2, -4, -9, -7, -7, -11,
					-- layer=2 filter=218 channel=3
					-24, -11, 10, -58, -10, 3, -87, -37, -49,
					-- layer=2 filter=218 channel=4
					-65, -8, 16, -53, -6, -41, -11, 11, 2,
					-- layer=2 filter=218 channel=5
					3, 1, 8, 9, 8, 1, 9, 8, 1,
					-- layer=2 filter=218 channel=6
					9, 6, 9, -1, -34, 0, -1, 14, -3,
					-- layer=2 filter=218 channel=7
					5, 6, -8, -10, 0, -45, 12, 38, -29,
					-- layer=2 filter=218 channel=8
					3, 4, 4, 9, 1, -1, 8, 7, -5,
					-- layer=2 filter=218 channel=9
					-12, -33, -18, 4, -43, 10, -35, -31, -36,
					-- layer=2 filter=218 channel=10
					-8, -15, -10, -11, 16, -22, -18, -40, -40,
					-- layer=2 filter=218 channel=11
					5, 26, -5, 26, 24, 0, 15, 23, 20,
					-- layer=2 filter=218 channel=12
					9, -8, -8, 4, 13, -34, -46, 3, -30,
					-- layer=2 filter=218 channel=13
					4, 4, -5, -3, 9, 1, -1, 6, -6,
					-- layer=2 filter=218 channel=14
					9, -15, -31, 26, 0, -5, 19, -3, 8,
					-- layer=2 filter=218 channel=15
					-18, 9, 9, -31, 5, 0, 3, 4, 51,
					-- layer=2 filter=218 channel=16
					7, 35, 27, 36, 19, -9, 20, 22, 0,
					-- layer=2 filter=218 channel=17
					10, 1, -10, 0, -6, 9, 4, 0, 9,
					-- layer=2 filter=218 channel=18
					-38, -9, 19, -1, -19, 2, -12, 21, 8,
					-- layer=2 filter=218 channel=19
					15, 31, 17, 42, 8, -21, -23, -7, -3,
					-- layer=2 filter=218 channel=20
					-6, -10, -8, -6, 5, -10, -3, -3, 0,
					-- layer=2 filter=218 channel=21
					12, 7, 3, 2, 2, 14, 8, 5, -10,
					-- layer=2 filter=218 channel=22
					-7, -3, 5, 3, -10, 4, 2, 4, 0,
					-- layer=2 filter=218 channel=23
					-8, 21, 35, -61, -13, -53, 4, -51, -53,
					-- layer=2 filter=218 channel=24
					-2, -42, 9, -66, -35, 16, -70, 3, 6,
					-- layer=2 filter=218 channel=25
					14, 2, -5, -57, -17, -10, -25, 16, 16,
					-- layer=2 filter=218 channel=26
					3, -2, 5, -6, -8, 3, -14, -10, 5,
					-- layer=2 filter=218 channel=27
					2, -25, -22, 50, 19, 29, 14, 12, 42,
					-- layer=2 filter=218 channel=28
					-67, 0, -28, 48, 15, -6, 24, 15, -24,
					-- layer=2 filter=218 channel=29
					-9, 3, -8, -4, -7, 4, 6, -16, -2,
					-- layer=2 filter=218 channel=30
					20, -39, -22, -2, -47, -23, 25, -3, 18,
					-- layer=2 filter=218 channel=31
					-33, 4, -11, -19, 4, -49, 24, 36, 4,
					-- layer=2 filter=218 channel=32
					-9, 4, -2, -2, 1, 2, 1, 2, -6,
					-- layer=2 filter=218 channel=33
					-42, -24, 19, -9, 4, -35, -59, 24, -28,
					-- layer=2 filter=218 channel=34
					32, 33, 43, 10, -54, 33, 46, 0, -16,
					-- layer=2 filter=218 channel=35
					-44, -36, -39, 0, 0, -8, 23, 23, 36,
					-- layer=2 filter=218 channel=36
					6, 17, 6, 0, 8, -5, 0, -9, -22,
					-- layer=2 filter=218 channel=37
					5, 7, -13, 10, 9, 3, 7, 17, 28,
					-- layer=2 filter=218 channel=38
					-4, -47, -36, -8, 11, 6, 25, 4, 31,
					-- layer=2 filter=218 channel=39
					-7, -20, 29, 18, -10, -48, -20, -8, -61,
					-- layer=2 filter=218 channel=40
					2, -24, 71, -15, 15, 4, -3, -4, 7,
					-- layer=2 filter=218 channel=41
					5, -7, 0, 9, 1, 3, -3, 0, 6,
					-- layer=2 filter=218 channel=42
					15, 11, 38, -51, -16, -5, -36, -7, -20,
					-- layer=2 filter=218 channel=43
					-32, -26, 13, -11, -25, 12, -52, -27, 3,
					-- layer=2 filter=218 channel=44
					7, -4, 0, -12, 0, 5, 7, 2, -1,
					-- layer=2 filter=218 channel=45
					-20, -15, -9, 3, 30, 23, -27, -36, 6,
					-- layer=2 filter=218 channel=46
					-31, -38, -2, 45, -19, -16, 11, -38, -19,
					-- layer=2 filter=218 channel=47
					-20, 0, -13, 48, 65, 16, 23, 20, 4,
					-- layer=2 filter=218 channel=48
					0, -1, 2, -1, -7, 6, -8, 6, 3,
					-- layer=2 filter=218 channel=49
					-11, 0, 37, 63, 5, -13, 13, 43, 19,
					-- layer=2 filter=218 channel=50
					-8, -5, 5, -4, -2, 22, -18, -17, 12,
					-- layer=2 filter=218 channel=51
					29, 11, -20, -1, 12, -9, 15, 13, 34,
					-- layer=2 filter=218 channel=52
					38, -6, 9, 33, 3, 4, 17, -8, 31,
					-- layer=2 filter=218 channel=53
					0, -29, 0, 32, -28, -17, 4, -67, -52,
					-- layer=2 filter=218 channel=54
					-12, 38, 1, -7, 21, 8, -12, -1, -19,
					-- layer=2 filter=218 channel=55
					-8, 2, 8, -7, -1, -2, -3, 4, -2,
					-- layer=2 filter=218 channel=56
					16, 2, -17, 23, 10, 8, -7, 14, 0,
					-- layer=2 filter=218 channel=57
					-8, 6, -6, -3, -7, 10, 17, 4, 10,
					-- layer=2 filter=218 channel=58
					9, 17, 1, 8, 19, -4, -17, -10, -13,
					-- layer=2 filter=218 channel=59
					-10, 21, 1, 30, 9, 21, -18, -20, 20,
					-- layer=2 filter=218 channel=60
					6, 7, -16, 19, -20, 42, 40, 54, 9,
					-- layer=2 filter=218 channel=61
					-14, 4, -39, -2, -45, 26, 29, 43, 35,
					-- layer=2 filter=218 channel=62
					24, 0, 32, 1, -33, -1, -9, 6, -4,
					-- layer=2 filter=218 channel=63
					3, 1, -14, -4, -7, 5, -10, -28, -19,
					-- layer=2 filter=218 channel=64
					3, 17, 44, -93, -59, -23, -49, -48, 9,
					-- layer=2 filter=218 channel=65
					18, 12, -10, 10, -22, 28, 26, -10, 11,
					-- layer=2 filter=218 channel=66
					-49, -51, -33, -1, -6, 1, 12, 20, 8,
					-- layer=2 filter=218 channel=67
					18, -65, -44, -5, 4, -53, -19, -65, -48,
					-- layer=2 filter=218 channel=68
					-10, -9, -8, -1, 5, 7, -8, 6, -10,
					-- layer=2 filter=218 channel=69
					-1, -21, 33, -63, -44, 7, -6, -65, -17,
					-- layer=2 filter=218 channel=70
					-18, -13, -32, 12, 18, 0, 28, 20, -9,
					-- layer=2 filter=218 channel=71
					-1, -37, -31, 26, 10, 14, -18, 7, 23,
					-- layer=2 filter=218 channel=72
					4, 16, -8, 58, 1, -15, -21, -6, -10,
					-- layer=2 filter=218 channel=73
					18, 30, 14, -4, 6, -16, 56, 11, -4,
					-- layer=2 filter=218 channel=74
					-15, -30, -30, -1, 23, -48, -2, 0, -61,
					-- layer=2 filter=218 channel=75
					14, 4, -65, 21, -8, -46, 1, -77, -78,
					-- layer=2 filter=218 channel=76
					-3, -2, 10, -47, -27, -40, -4, -34, -21,
					-- layer=2 filter=218 channel=77
					-5, 7, -8, -4, 4, -5, -3, 8, -3,
					-- layer=2 filter=218 channel=78
					-2, -7, -19, -21, -5, 5, -1, -11, 9,
					-- layer=2 filter=218 channel=79
					-7, 9, 7, -9, -4, 9, -10, -7, 8,
					-- layer=2 filter=218 channel=80
					-15, -52, -17, 8, 14, -37, 38, 9, 2,
					-- layer=2 filter=218 channel=81
					5, -16, -1, 4, 4, -5, -11, -13, -12,
					-- layer=2 filter=218 channel=82
					7, -3, 7, 2, -10, -7, 3, 3, 0,
					-- layer=2 filter=218 channel=83
					-43, -10, 14, -35, 13, -21, -47, 7, 15,
					-- layer=2 filter=218 channel=84
					-6, -10, -3, -9, -3, 1, -4, 4, 10,
					-- layer=2 filter=218 channel=85
					6, 3, 0, 8, -5, 1, -4, 14, 16,
					-- layer=2 filter=218 channel=86
					-17, 0, 6, -3, -11, 16, 5, -14, 1,
					-- layer=2 filter=218 channel=87
					-8, -17, 27, -22, -5, 29, -40, 20, 14,
					-- layer=2 filter=218 channel=88
					-28, -54, 12, -83, -56, -26, 11, -26, 34,
					-- layer=2 filter=218 channel=89
					8, 26, -24, 38, -17, -64, -4, -4, -2,
					-- layer=2 filter=218 channel=90
					9, -3, 1, 6, 10, -1, 9, 4, 0,
					-- layer=2 filter=218 channel=91
					47, -15, -43, 17, -24, -57, -16, 7, -18,
					-- layer=2 filter=218 channel=92
					2, 2, -1, 21, 4, -41, -20, 2, 7,
					-- layer=2 filter=218 channel=93
					28, -28, 27, 22, -2, -4, -17, -46, -11,
					-- layer=2 filter=218 channel=94
					-28, 39, -1, -8, -53, 12, 18, -26, -15,
					-- layer=2 filter=218 channel=95
					8, 12, 8, -12, -15, -25, 23, 16, 11,
					-- layer=2 filter=218 channel=96
					-21, 12, -9, 16, -16, -28, 62, 27, -4,
					-- layer=2 filter=218 channel=97
					-2, -32, 16, -66, -10, -22, -48, 21, -21,
					-- layer=2 filter=218 channel=98
					-26, 17, -11, 22, 26, 8, 36, 13, 9,
					-- layer=2 filter=218 channel=99
					9, 45, -12, 13, 2, -24, 41, -9, -5,
					-- layer=2 filter=218 channel=100
					-28, -26, 12, -4, 11, 11, 40, 3, -18,
					-- layer=2 filter=218 channel=101
					19, -29, -28, 17, 8, -7, -2, 17, 5,
					-- layer=2 filter=218 channel=102
					14, 30, 7, 47, -33, -26, 16, 6, -7,
					-- layer=2 filter=218 channel=103
					5, -7, -71, -32, -4, 65, -12, -8, -5,
					-- layer=2 filter=218 channel=104
					-29, 13, 23, 13, 16, 13, -17, 16, -2,
					-- layer=2 filter=218 channel=105
					-40, 54, -36, -8, -28, -4, 2, -4, -14,
					-- layer=2 filter=218 channel=106
					16, -14, -5, -44, -15, -36, -31, -18, -24,
					-- layer=2 filter=218 channel=107
					-49, -30, -87, 3, 8, 26, -1, -31, 21,
					-- layer=2 filter=218 channel=108
					-8, -31, -34, 27, -19, 15, 24, 6, 14,
					-- layer=2 filter=218 channel=109
					19, -3, 0, 3, -8, -6, -1, -5, 10,
					-- layer=2 filter=218 channel=110
					8, 7, -14, -75, -78, -35, -33, 30, 34,
					-- layer=2 filter=218 channel=111
					8, 9, -5, 0, 2, 0, 0, 1, -8,
					-- layer=2 filter=218 channel=112
					33, -4, -33, 8, -22, -22, 21, -2, 22,
					-- layer=2 filter=218 channel=113
					24, -25, -9, 28, -41, -8, 13, -10, 31,
					-- layer=2 filter=218 channel=114
					9, 10, 10, 9, 12, 4, 17, 6, 5,
					-- layer=2 filter=218 channel=115
					2, 10, -10, 5, 5, -2, -3, -7, 2,
					-- layer=2 filter=218 channel=116
					-2, 7, -2, 2, 21, 30, -6, -1, 23,
					-- layer=2 filter=218 channel=117
					18, 25, -23, -4, 42, -43, 40, 16, -18,
					-- layer=2 filter=218 channel=118
					2, -41, -3, -38, 6, -2, -34, 19, 1,
					-- layer=2 filter=218 channel=119
					-56, -19, 7, -34, -32, 23, -2, 1, -36,
					-- layer=2 filter=218 channel=120
					-2, 0, 5, -7, 0, -6, -10, -1, 0,
					-- layer=2 filter=218 channel=121
					-7, -5, -4, 1, -5, 6, -8, -1, -1,
					-- layer=2 filter=218 channel=122
					4, -10, 0, -1, 4, 9, 12, -4, 5,
					-- layer=2 filter=218 channel=123
					23, 0, 32, 26, 0, -12, 18, -6, -20,
					-- layer=2 filter=218 channel=124
					-7, 13, 67, -45, 20, -24, -5, -11, -26,
					-- layer=2 filter=218 channel=125
					3, 8, -5, 3, -5, 10, -3, 7, -8,
					-- layer=2 filter=218 channel=126
					3, -55, -33, 27, -70, -16, -3, -17, -38,
					-- layer=2 filter=218 channel=127
					-12, 0, 8, -3, -4, 21, -14, -24, 9,
					-- layer=2 filter=219 channel=0
					-6, 8, 7, -2, -12, 2, -4, -4, 0,
					-- layer=2 filter=219 channel=1
					2, -10, -17, 4, -1, -4, 2, 0, -13,
					-- layer=2 filter=219 channel=2
					-8, -11, 0, -11, 7, -10, 1, 0, 4,
					-- layer=2 filter=219 channel=3
					-6, -7, -5, -7, -8, -1, -5, 2, 7,
					-- layer=2 filter=219 channel=4
					-6, 2, -3, 2, -5, -15, 1, 0, 0,
					-- layer=2 filter=219 channel=5
					-8, -2, 3, -9, 0, -1, -1, 4, -4,
					-- layer=2 filter=219 channel=6
					-6, -7, -1, -1, -6, -9, 0, 0, 2,
					-- layer=2 filter=219 channel=7
					-7, -5, 2, -9, 7, 7, 0, -11, -6,
					-- layer=2 filter=219 channel=8
					7, 2, 1, -7, 3, 1, -2, 4, -1,
					-- layer=2 filter=219 channel=9
					-11, 7, 3, 2, 1, -8, -9, -12, 3,
					-- layer=2 filter=219 channel=10
					-8, 4, -2, -1, -13, -2, 3, 6, 0,
					-- layer=2 filter=219 channel=11
					-11, 0, -17, -1, -3, -10, 5, -8, -7,
					-- layer=2 filter=219 channel=12
					-10, -7, -7, -11, -11, 0, -12, 0, -11,
					-- layer=2 filter=219 channel=13
					-4, -10, 0, -5, 9, 9, 5, 0, 4,
					-- layer=2 filter=219 channel=14
					-4, 0, 7, -1, 2, 8, -11, 0, -10,
					-- layer=2 filter=219 channel=15
					-1, -11, -10, -11, 7, 7, 6, 0, 0,
					-- layer=2 filter=219 channel=16
					4, -5, 2, -6, 6, -11, 4, -6, -11,
					-- layer=2 filter=219 channel=17
					5, 5, -4, 2, -10, 7, 4, -6, 9,
					-- layer=2 filter=219 channel=18
					-13, -5, -6, -8, 1, 2, -8, -6, 9,
					-- layer=2 filter=219 channel=19
					3, -4, -6, -7, -2, 6, 1, 1, 8,
					-- layer=2 filter=219 channel=20
					-6, -7, 4, 5, -9, -2, -6, -2, 9,
					-- layer=2 filter=219 channel=21
					-2, 0, 6, -3, -7, 6, -6, -2, 7,
					-- layer=2 filter=219 channel=22
					5, 3, 6, 1, 6, -9, -1, -6, 2,
					-- layer=2 filter=219 channel=23
					-11, -9, -3, -2, -5, -9, -13, 0, 5,
					-- layer=2 filter=219 channel=24
					-4, -1, -3, -10, 6, -7, -8, 0, -10,
					-- layer=2 filter=219 channel=25
					-3, -5, 8, 6, -10, 5, 5, 6, 6,
					-- layer=2 filter=219 channel=26
					-6, 6, 8, 1, 0, 10, -7, -5, -8,
					-- layer=2 filter=219 channel=27
					-9, 6, 1, 1, -9, -1, -7, -8, -11,
					-- layer=2 filter=219 channel=28
					-8, -10, -2, 0, 2, -15, 1, 4, -3,
					-- layer=2 filter=219 channel=29
					6, -5, 0, -9, -3, -6, -3, -5, -3,
					-- layer=2 filter=219 channel=30
					-7, -7, -10, -8, -11, -5, -1, 5, -5,
					-- layer=2 filter=219 channel=31
					7, 2, 8, -6, -4, -6, -5, -6, -4,
					-- layer=2 filter=219 channel=32
					-3, -6, 3, -3, 0, -7, -1, -5, 1,
					-- layer=2 filter=219 channel=33
					0, -7, -3, -5, -6, -8, 3, -7, 3,
					-- layer=2 filter=219 channel=34
					-4, -8, -8, 1, -9, -3, 7, -5, -10,
					-- layer=2 filter=219 channel=35
					0, 0, -7, -6, -10, 0, 0, -9, -11,
					-- layer=2 filter=219 channel=36
					6, 1, 0, -6, -6, -7, 2, -2, 6,
					-- layer=2 filter=219 channel=37
					-13, 0, -15, 2, -12, -4, -6, 1, 2,
					-- layer=2 filter=219 channel=38
					5, -10, -4, -6, -12, -4, -6, 8, 5,
					-- layer=2 filter=219 channel=39
					-4, -10, 2, -1, -2, -8, 1, -6, -8,
					-- layer=2 filter=219 channel=40
					0, -6, 1, 3, 7, 8, 0, 0, 1,
					-- layer=2 filter=219 channel=41
					5, -5, -7, 6, -7, -5, -1, -2, -5,
					-- layer=2 filter=219 channel=42
					7, 1, 2, 10, -6, 5, -7, -4, -6,
					-- layer=2 filter=219 channel=43
					0, -6, 4, 1, -10, -8, 6, 0, -8,
					-- layer=2 filter=219 channel=44
					-5, -2, 2, -5, -6, -3, -6, -2, 7,
					-- layer=2 filter=219 channel=45
					-11, 7, 3, -4, -5, 6, 0, 1, -6,
					-- layer=2 filter=219 channel=46
					3, -11, -11, -7, -3, -5, 7, 0, -2,
					-- layer=2 filter=219 channel=47
					-1, -6, 8, -18, -8, -1, 6, -11, -8,
					-- layer=2 filter=219 channel=48
					-2, -9, 2, -3, -4, -8, 2, -5, -8,
					-- layer=2 filter=219 channel=49
					3, 1, -5, -11, -8, 3, 6, -3, -5,
					-- layer=2 filter=219 channel=50
					-8, -4, 0, -5, 9, 0, -3, 0, -7,
					-- layer=2 filter=219 channel=51
					-9, 0, -3, 5, -4, -2, -10, -10, 0,
					-- layer=2 filter=219 channel=52
					-5, 0, -19, -12, -5, 5, -4, 5, 4,
					-- layer=2 filter=219 channel=53
					-10, 0, -11, 0, 0, -9, 6, 6, 7,
					-- layer=2 filter=219 channel=54
					-15, 2, 0, 0, -1, -8, -13, -10, -11,
					-- layer=2 filter=219 channel=55
					3, 1, 0, -5, -4, -3, -5, 7, 2,
					-- layer=2 filter=219 channel=56
					-5, -8, 0, -13, -11, 5, 2, 3, -7,
					-- layer=2 filter=219 channel=57
					-6, -9, 4, -6, 0, -1, 3, 5, -12,
					-- layer=2 filter=219 channel=58
					-4, 3, -4, -5, 9, 0, 0, 0, -1,
					-- layer=2 filter=219 channel=59
					-10, -11, -15, -2, -1, -8, -7, -2, -12,
					-- layer=2 filter=219 channel=60
					-10, 4, 1, -9, 3, -9, -8, -6, -2,
					-- layer=2 filter=219 channel=61
					-2, 0, 0, -6, -4, 4, -9, 9, 3,
					-- layer=2 filter=219 channel=62
					-11, 2, 2, -4, -4, -9, 1, 1, 1,
					-- layer=2 filter=219 channel=63
					-13, -7, -11, 4, 4, 2, -14, -16, -14,
					-- layer=2 filter=219 channel=64
					-6, 3, -6, -2, 4, 8, 6, 8, 6,
					-- layer=2 filter=219 channel=65
					-9, 0, 0, -1, 5, 1, -4, -11, -4,
					-- layer=2 filter=219 channel=66
					-10, 4, 3, -9, -11, -8, 6, -9, -4,
					-- layer=2 filter=219 channel=67
					5, 5, -8, -4, 0, 7, 3, 2, -1,
					-- layer=2 filter=219 channel=68
					-4, 6, -1, 3, 0, 8, 5, -6, -2,
					-- layer=2 filter=219 channel=69
					7, -6, -7, -4, 0, -3, -12, 0, -2,
					-- layer=2 filter=219 channel=70
					-7, -8, -14, -13, -7, 0, -14, -6, -5,
					-- layer=2 filter=219 channel=71
					-5, 6, 7, -8, -1, 0, 9, 0, 3,
					-- layer=2 filter=219 channel=72
					0, -8, -4, 8, -14, -4, -3, -6, 0,
					-- layer=2 filter=219 channel=73
					-8, -4, -6, -4, 1, 1, 8, 0, -4,
					-- layer=2 filter=219 channel=74
					2, 4, -5, -11, 0, 5, -10, 4, 5,
					-- layer=2 filter=219 channel=75
					-11, -2, -6, -11, 3, 0, -11, 5, 4,
					-- layer=2 filter=219 channel=76
					1, -7, 0, -7, -9, 6, -6, -6, -10,
					-- layer=2 filter=219 channel=77
					-10, -11, 6, 8, 4, 4, -6, -4, -7,
					-- layer=2 filter=219 channel=78
					-8, 4, -1, -4, -3, -3, 3, -8, 8,
					-- layer=2 filter=219 channel=79
					-12, -3, -6, -3, 3, 0, -6, 0, -2,
					-- layer=2 filter=219 channel=80
					-10, -8, -2, 0, -3, 4, 4, -3, 1,
					-- layer=2 filter=219 channel=81
					-9, 4, -12, -9, -3, 2, 0, -5, -7,
					-- layer=2 filter=219 channel=82
					4, -1, -10, 2, -4, 0, -6, 10, 5,
					-- layer=2 filter=219 channel=83
					4, -4, -13, -7, -6, -4, 5, -5, 6,
					-- layer=2 filter=219 channel=84
					1, -1, 4, 1, -9, -10, 4, -3, 2,
					-- layer=2 filter=219 channel=85
					-2, -4, -6, -11, -4, 1, 8, 4, -1,
					-- layer=2 filter=219 channel=86
					11, 11, -11, 9, 2, -2, 11, -12, -4,
					-- layer=2 filter=219 channel=87
					2, 0, -4, -6, 8, -3, -9, 7, -7,
					-- layer=2 filter=219 channel=88
					5, -5, 3, 3, -9, -1, 2, -13, 4,
					-- layer=2 filter=219 channel=89
					-12, -13, 3, 2, 1, 0, 0, -3, -4,
					-- layer=2 filter=219 channel=90
					-4, -9, 10, -8, 4, 10, 1, 0, -7,
					-- layer=2 filter=219 channel=91
					5, -11, -9, -3, -1, 3, 1, 0, -7,
					-- layer=2 filter=219 channel=92
					-15, -1, 0, 4, -7, 5, -11, -14, -7,
					-- layer=2 filter=219 channel=93
					-9, -11, 0, 4, -4, -4, -2, 8, 0,
					-- layer=2 filter=219 channel=94
					-2, -7, 2, -1, -7, -8, -3, -7, -1,
					-- layer=2 filter=219 channel=95
					7, 3, -8, 8, 1, -5, 3, 4, -4,
					-- layer=2 filter=219 channel=96
					-3, 2, -9, -11, 2, 6, -10, -10, 7,
					-- layer=2 filter=219 channel=97
					5, 5, -11, -11, 2, 7, 4, 2, -5,
					-- layer=2 filter=219 channel=98
					1, -12, -11, -13, -6, -7, -4, -5, -4,
					-- layer=2 filter=219 channel=99
					-8, -7, 3, 3, -4, 4, 6, -6, 5,
					-- layer=2 filter=219 channel=100
					-11, -4, -2, -1, -1, 6, -12, 2, 4,
					-- layer=2 filter=219 channel=101
					-5, -1, -5, -4, 7, -1, 1, 0, -3,
					-- layer=2 filter=219 channel=102
					-14, -15, -6, 2, -3, -8, -8, -10, -3,
					-- layer=2 filter=219 channel=103
					-12, -6, 3, -7, -9, -1, 3, 0, -5,
					-- layer=2 filter=219 channel=104
					-11, -1, 0, -7, 0, 2, 0, -9, -6,
					-- layer=2 filter=219 channel=105
					0, 2, -6, -2, -7, -10, -8, -7, -8,
					-- layer=2 filter=219 channel=106
					-9, 3, -1, -1, 4, 4, -11, 4, 1,
					-- layer=2 filter=219 channel=107
					0, 7, 1, -6, 2, -8, 6, -10, 1,
					-- layer=2 filter=219 channel=108
					-11, -10, 5, 5, -8, -11, -10, -7, -1,
					-- layer=2 filter=219 channel=109
					-1, 0, -9, -9, -7, 9, -10, -3, -9,
					-- layer=2 filter=219 channel=110
					3, -10, -10, -5, -5, -8, -13, 0, -5,
					-- layer=2 filter=219 channel=111
					7, 7, 8, -4, -8, 7, 3, 2, 0,
					-- layer=2 filter=219 channel=112
					1, -5, 4, 3, -8, 2, -11, -10, -2,
					-- layer=2 filter=219 channel=113
					6, -8, 1, -12, -3, -11, -11, -13, -7,
					-- layer=2 filter=219 channel=114
					-9, -6, 9, -8, -11, -7, -7, 0, 8,
					-- layer=2 filter=219 channel=115
					5, -3, 6, -9, 1, 6, -7, -3, -10,
					-- layer=2 filter=219 channel=116
					0, -6, -4, -1, -10, 0, -7, 8, -8,
					-- layer=2 filter=219 channel=117
					-2, -1, -17, 6, 8, -4, 5, -1, -1,
					-- layer=2 filter=219 channel=118
					-8, -7, 6, 1, -8, 5, 3, -2, 8,
					-- layer=2 filter=219 channel=119
					0, -4, 7, 0, -8, -5, 6, 8, -7,
					-- layer=2 filter=219 channel=120
					4, 10, -3, 4, 1, 6, -2, 1, 4,
					-- layer=2 filter=219 channel=121
					-5, -12, -3, -8, 6, -6, -11, 3, 2,
					-- layer=2 filter=219 channel=122
					-1, -8, 2, 0, 4, 6, -9, 3, -6,
					-- layer=2 filter=219 channel=123
					-11, 2, -1, -11, -3, -9, 4, 7, -4,
					-- layer=2 filter=219 channel=124
					-3, 4, 3, -6, -7, -1, 0, -4, 6,
					-- layer=2 filter=219 channel=125
					-4, 5, 4, 2, -9, -3, -9, -9, -2,
					-- layer=2 filter=219 channel=126
					-5, 0, 5, 8, -9, 0, -4, -5, 6,
					-- layer=2 filter=219 channel=127
					-9, 5, 2, 2, -13, -3, -3, -12, 2,
					-- layer=2 filter=220 channel=0
					-10, 4, 0, -59, -14, 3, -27, 26, 30,
					-- layer=2 filter=220 channel=1
					20, -9, -36, 49, -19, 1, 24, -6, -53,
					-- layer=2 filter=220 channel=2
					0, -5, -1, 1, 5, -5, -6, 0, 0,
					-- layer=2 filter=220 channel=3
					21, 21, -18, -6, 4, 1, -8, 20, -12,
					-- layer=2 filter=220 channel=4
					10, -15, 34, 11, -3, 42, 12, -23, 17,
					-- layer=2 filter=220 channel=5
					-25, -7, 38, -52, -12, 7, -16, -6, 51,
					-- layer=2 filter=220 channel=6
					-53, -9, 33, -4, -5, 12, -33, -45, 56,
					-- layer=2 filter=220 channel=7
					50, -21, -8, 10, -15, -47, 20, -9, 2,
					-- layer=2 filter=220 channel=8
					0, -7, 7, -5, -8, -9, -4, -6, 2,
					-- layer=2 filter=220 channel=9
					5, 25, -29, -40, -26, -33, -20, 1, -11,
					-- layer=2 filter=220 channel=10
					-18, -10, -3, -16, 17, 3, -18, 13, 9,
					-- layer=2 filter=220 channel=11
					-12, 8, 19, -29, 0, 42, -7, 13, 31,
					-- layer=2 filter=220 channel=12
					3, -25, 0, 12, -10, -9, 13, 0, -25,
					-- layer=2 filter=220 channel=13
					-1, 0, -2, -9, 3, -10, -9, 2, 6,
					-- layer=2 filter=220 channel=14
					34, -10, 11, 62, -3, 2, 52, -8, -23,
					-- layer=2 filter=220 channel=15
					-27, 42, 14, 22, -6, -12, 17, -26, -9,
					-- layer=2 filter=220 channel=16
					52, 12, -43, 12, -22, -52, 23, -5, -61,
					-- layer=2 filter=220 channel=17
					3, -5, -8, -3, 8, 8, 8, -3, 9,
					-- layer=2 filter=220 channel=18
					29, 12, 36, 18, 18, 6, 32, 28, 10,
					-- layer=2 filter=220 channel=19
					19, -4, -27, 26, -14, -9, 22, -3, -33,
					-- layer=2 filter=220 channel=20
					7, -10, -7, -5, -8, 7, 5, -7, 0,
					-- layer=2 filter=220 channel=21
					-12, 17, 8, 19, 8, 30, -5, 12, 29,
					-- layer=2 filter=220 channel=22
					0, 0, -4, 1, 0, -2, -2, 9, -1,
					-- layer=2 filter=220 channel=23
					-2, -10, -6, 30, 20, 14, 35, -16, -23,
					-- layer=2 filter=220 channel=24
					7, 3, -40, -13, -2, -43, -35, 12, -10,
					-- layer=2 filter=220 channel=25
					-31, -1, -29, -35, -6, -19, -25, 19, 1,
					-- layer=2 filter=220 channel=26
					0, 2, 1, -6, 4, 2, 3, -10, 2,
					-- layer=2 filter=220 channel=27
					-1, -14, 25, -2, -9, 19, -4, -2, 2,
					-- layer=2 filter=220 channel=28
					-3, -25, -14, 42, 10, -9, 9, -1, -19,
					-- layer=2 filter=220 channel=29
					3, -5, -2, -5, 10, -6, -7, -6, -4,
					-- layer=2 filter=220 channel=30
					-4, 6, 22, 4, -2, 12, -6, 14, 19,
					-- layer=2 filter=220 channel=31
					-91, -24, 0, 15, -24, -61, 44, 5, -14,
					-- layer=2 filter=220 channel=32
					-7, 2, -5, 3, -5, 1, -6, -11, 5,
					-- layer=2 filter=220 channel=33
					52, 17, 26, 45, -3, 37, 44, -18, -6,
					-- layer=2 filter=220 channel=34
					7, -11, 69, 17, -8, 8, -19, -26, 6,
					-- layer=2 filter=220 channel=35
					28, 0, 2, 76, 25, 11, 26, -8, 17,
					-- layer=2 filter=220 channel=36
					5, -4, -9, -17, 6, 5, -6, 12, -3,
					-- layer=2 filter=220 channel=37
					-14, -8, 24, -12, 4, 26, -6, -11, 36,
					-- layer=2 filter=220 channel=38
					-28, -5, 34, -9, -2, 37, -10, -6, 28,
					-- layer=2 filter=220 channel=39
					22, 3, -8, -6, -12, -28, -21, -32, -59,
					-- layer=2 filter=220 channel=40
					-39, -16, -39, -32, -6, 28, 26, -4, 2,
					-- layer=2 filter=220 channel=41
					-11, -1, -1, 5, 6, -10, 2, -5, 7,
					-- layer=2 filter=220 channel=42
					43, 8, -10, 57, -7, -31, 59, -11, -41,
					-- layer=2 filter=220 channel=43
					16, 12, 29, -17, 6, 37, -13, 27, 2,
					-- layer=2 filter=220 channel=44
					6, -3, 7, 6, -2, -5, 0, -4, -6,
					-- layer=2 filter=220 channel=45
					7, -23, -10, 48, -14, -18, 65, -14, -32,
					-- layer=2 filter=220 channel=46
					31, 8, -18, -5, 12, 3, 12, 10, -2,
					-- layer=2 filter=220 channel=47
					19, -4, 6, 10, 16, -21, 25, -3, -37,
					-- layer=2 filter=220 channel=48
					6, -4, 0, 0, -8, 0, -4, 1, 8,
					-- layer=2 filter=220 channel=49
					10, 3, 28, 11, 10, -8, 1, -22, -31,
					-- layer=2 filter=220 channel=50
					19, 16, 11, 12, -10, 11, -4, -6, -13,
					-- layer=2 filter=220 channel=51
					-27, -1, 24, -46, -4, 41, -20, 1, 44,
					-- layer=2 filter=220 channel=52
					-16, -21, 27, -5, 18, 30, 10, 1, 20,
					-- layer=2 filter=220 channel=53
					-3, 62, 11, -1, -7, 29, -30, 6, -7,
					-- layer=2 filter=220 channel=54
					17, -13, 19, 19, 14, 17, 19, 6, 8,
					-- layer=2 filter=220 channel=55
					-1, -6, 7, 11, 7, 10, 8, -7, 9,
					-- layer=2 filter=220 channel=56
					-34, -9, 43, -23, -8, 18, -18, 19, 29,
					-- layer=2 filter=220 channel=57
					8, -7, -8, -10, 0, 2, -6, -5, -3,
					-- layer=2 filter=220 channel=58
					-22, -34, 0, 7, -23, 15, -14, 20, -2,
					-- layer=2 filter=220 channel=59
					5, 1, 27, -26, -7, 40, -90, -37, -47,
					-- layer=2 filter=220 channel=60
					-77, -60, -33, -159, -30, -55, -65, -112, -18,
					-- layer=2 filter=220 channel=61
					2, 13, -35, -93, 8, -51, -69, -43, -22,
					-- layer=2 filter=220 channel=62
					6, -11, -12, 2, 37, 3, -5, -7, -7,
					-- layer=2 filter=220 channel=63
					-11, 11, 0, -25, -19, -7, -16, 0, -17,
					-- layer=2 filter=220 channel=64
					-3, 14, 2, 30, 21, -8, 20, 17, 16,
					-- layer=2 filter=220 channel=65
					-49, -23, -25, -54, 2, -19, -54, -46, 12,
					-- layer=2 filter=220 channel=66
					-60, -25, -86, -20, 11, 10, -24, -7, -36,
					-- layer=2 filter=220 channel=67
					-3, 45, 15, -31, 21, -16, -20, 15, 17,
					-- layer=2 filter=220 channel=68
					-5, -5, 8, -11, -5, 7, 9, 0, 10,
					-- layer=2 filter=220 channel=69
					26, 0, -9, 23, 10, -25, 26, 2, -32,
					-- layer=2 filter=220 channel=70
					12, -19, 3, 36, -3, 10, 31, -15, 8,
					-- layer=2 filter=220 channel=71
					2, 16, 37, -4, 0, 38, -14, -4, 7,
					-- layer=2 filter=220 channel=72
					25, -13, -11, -5, 33, 13, 18, 1, -14,
					-- layer=2 filter=220 channel=73
					-31, 26, -13, 25, -2, -49, 34, -35, -65,
					-- layer=2 filter=220 channel=74
					-21, 4, 31, -12, 17, -4, -1, 37, 11,
					-- layer=2 filter=220 channel=75
					49, 11, 14, 13, -30, -8, -16, -22, -19,
					-- layer=2 filter=220 channel=76
					-12, 9, 7, -29, -1, 6, -8, -14, 4,
					-- layer=2 filter=220 channel=77
					-3, -5, -2, -7, -1, 6, 8, -4, -3,
					-- layer=2 filter=220 channel=78
					-16, -2, 25, -11, -9, 17, -16, 17, 38,
					-- layer=2 filter=220 channel=79
					7, 8, 8, 0, 2, -3, -5, 5, -7,
					-- layer=2 filter=220 channel=80
					33, 29, 14, 35, -4, -2, 22, -2, -3,
					-- layer=2 filter=220 channel=81
					-5, 14, -1, 10, 0, 8, -2, 0, -1,
					-- layer=2 filter=220 channel=82
					-7, -11, -10, 7, -10, -4, -6, 11, 1,
					-- layer=2 filter=220 channel=83
					20, -9, 4, 31, 14, -7, 37, -10, -26,
					-- layer=2 filter=220 channel=84
					10, -2, -7, -1, -2, -4, 4, 11, 1,
					-- layer=2 filter=220 channel=85
					-3, 2, 4, 4, 0, 2, -5, 5, 2,
					-- layer=2 filter=220 channel=86
					14, 1, -16, 7, 2, -5, 10, -27, 0,
					-- layer=2 filter=220 channel=87
					-33, 0, 12, -50, 11, 52, -42, -28, 12,
					-- layer=2 filter=220 channel=88
					13, 33, 16, 8, 21, 4, 14, -11, 28,
					-- layer=2 filter=220 channel=89
					35, -21, -25, 42, 28, -15, 30, 14, -41,
					-- layer=2 filter=220 channel=90
					-1, 3, 10, 10, 0, -7, 5, 0, -9,
					-- layer=2 filter=220 channel=91
					23, -17, -31, 21, -14, -23, 3, 15, -14,
					-- layer=2 filter=220 channel=92
					42, -10, -17, 33, 1, -11, 35, -7, -54,
					-- layer=2 filter=220 channel=93
					-7, -36, -46, 61, -7, -40, -1, -4, -45,
					-- layer=2 filter=220 channel=94
					-8, -3, -31, -33, -33, -71, -37, -106, -89,
					-- layer=2 filter=220 channel=95
					0, 2, 13, 1, 10, 0, -3, -8, 6,
					-- layer=2 filter=220 channel=96
					-18, -4, 39, 4, -39, 59, -7, -9, 25,
					-- layer=2 filter=220 channel=97
					16, 32, 9, -12, -5, 27, 10, 7, 2,
					-- layer=2 filter=220 channel=98
					11, -12, -14, 40, 8, -24, 5, -6, -52,
					-- layer=2 filter=220 channel=99
					-3, 3, 26, 15, -1, -8, 5, -9, 12,
					-- layer=2 filter=220 channel=100
					-18, -20, 1, -51, -15, 6, 6, -35, -9,
					-- layer=2 filter=220 channel=101
					0, 31, 8, 10, 20, 21, 0, 13, -13,
					-- layer=2 filter=220 channel=102
					13, 0, 38, 12, -8, -9, 29, -17, -14,
					-- layer=2 filter=220 channel=103
					38, 12, 5, 40, -4, 25, 35, -6, 16,
					-- layer=2 filter=220 channel=104
					-2, 16, 23, -7, -8, -12, -28, -17, -8,
					-- layer=2 filter=220 channel=105
					-14, -23, 22, -43, 46, 25, 11, 10, 54,
					-- layer=2 filter=220 channel=106
					0, 6, -7, -22, 24, 5, -22, 29, -12,
					-- layer=2 filter=220 channel=107
					30, 34, -15, 12, 19, 21, 7, -44, -25,
					-- layer=2 filter=220 channel=108
					26, -25, -2, 8, -27, 0, -14, -53, -33,
					-- layer=2 filter=220 channel=109
					-10, 9, 2, -7, 1, 2, 0, 7, -5,
					-- layer=2 filter=220 channel=110
					33, 2, -40, 0, -2, -64, 1, -4, -27,
					-- layer=2 filter=220 channel=111
					8, 10, 0, -2, 3, 6, 1, -7, 4,
					-- layer=2 filter=220 channel=112
					-9, 25, 16, -66, 25, -14, -36, 3, 21,
					-- layer=2 filter=220 channel=113
					-20, 0, 0, 10, 2, 2, -31, 31, 1,
					-- layer=2 filter=220 channel=114
					-9, -11, 0, -26, -8, -4, -1, -17, 15,
					-- layer=2 filter=220 channel=115
					-9, -2, 8, 3, 9, 0, -13, 3, 3,
					-- layer=2 filter=220 channel=116
					3, 24, 22, -27, 4, 42, -35, -48, -6,
					-- layer=2 filter=220 channel=117
					23, -3, -2, 35, 11, -20, 31, -12, 10,
					-- layer=2 filter=220 channel=118
					-13, 19, 26, -7, 18, 35, 9, 32, 33,
					-- layer=2 filter=220 channel=119
					20, 19, 4, 33, 11, -19, 38, 17, -63,
					-- layer=2 filter=220 channel=120
					-10, 3, -2, 4, 0, 9, 5, 9, -8,
					-- layer=2 filter=220 channel=121
					0, 3, 4, -11, -2, 3, -12, -1, -8,
					-- layer=2 filter=220 channel=122
					-4, -5, -1, -1, -13, 6, 0, 4, 1,
					-- layer=2 filter=220 channel=123
					7, 8, 23, -20, 15, -20, -9, 0, -15,
					-- layer=2 filter=220 channel=124
					15, 33, 15, 30, 32, -5, 57, 24, 38,
					-- layer=2 filter=220 channel=125
					-7, -8, -4, -3, 5, 12, -2, 5, -2,
					-- layer=2 filter=220 channel=126
					8, -2, 11, -16, -6, -68, 27, -5, -45,
					-- layer=2 filter=220 channel=127
					6, -20, 19, 24, -17, 24, 3, -33, -18,
					-- layer=2 filter=221 channel=0
					-11, -3, 2, -9, -1, -15, -5, -12, -17,
					-- layer=2 filter=221 channel=1
					8, -11, -19, -5, -1, 4, -6, 9, -12,
					-- layer=2 filter=221 channel=2
					-4, 0, -5, 0, 5, 4, -1, 10, 9,
					-- layer=2 filter=221 channel=3
					-18, -8, 13, -3, -2, -9, -13, 4, 3,
					-- layer=2 filter=221 channel=4
					-15, -7, -18, -2, 4, -1, -9, -4, 13,
					-- layer=2 filter=221 channel=5
					0, 0, -5, -9, 6, 6, -18, 2, -13,
					-- layer=2 filter=221 channel=6
					-10, -28, -22, -3, -20, 1, 9, -20, 30,
					-- layer=2 filter=221 channel=7
					16, -7, -3, -17, -20, -11, 4, 6, -3,
					-- layer=2 filter=221 channel=8
					4, 0, -1, 7, -3, 8, -3, -2, -3,
					-- layer=2 filter=221 channel=9
					-6, 3, -11, 3, -10, -14, -3, -3, 3,
					-- layer=2 filter=221 channel=10
					-7, 0, -6, 1, 0, -16, -1, -10, 1,
					-- layer=2 filter=221 channel=11
					3, -6, -18, 1, -8, -9, -11, -17, -12,
					-- layer=2 filter=221 channel=12
					-2, 0, 2, -5, -10, -1, -5, -13, -10,
					-- layer=2 filter=221 channel=13
					2, -10, 3, -9, 5, 1, -5, -6, 4,
					-- layer=2 filter=221 channel=14
					-19, -13, -15, -1, -13, -8, -7, -11, -13,
					-- layer=2 filter=221 channel=15
					-9, -22, 3, -4, 0, 3, 3, -15, -15,
					-- layer=2 filter=221 channel=16
					-16, -6, -17, -11, 0, 6, 0, -1, -1,
					-- layer=2 filter=221 channel=17
					-2, -8, -8, -1, 6, -1, 0, 2, 9,
					-- layer=2 filter=221 channel=18
					9, -7, -17, -9, -7, -6, -5, -10, -16,
					-- layer=2 filter=221 channel=19
					3, -7, -22, -12, -11, -5, -1, 1, 6,
					-- layer=2 filter=221 channel=20
					4, 1, 1, 5, -3, -7, 0, 12, 3,
					-- layer=2 filter=221 channel=21
					-11, 8, 8, 0, 6, -1, 3, 5, -9,
					-- layer=2 filter=221 channel=22
					-7, 3, 2, 0, 5, 0, -7, 4, 8,
					-- layer=2 filter=221 channel=23
					3, -1, -5, -12, 2, 2, -8, 0, 6,
					-- layer=2 filter=221 channel=24
					-5, -8, 5, -13, 3, -9, 4, -6, -2,
					-- layer=2 filter=221 channel=25
					-20, -7, -10, -9, -7, -9, -19, -16, -3,
					-- layer=2 filter=221 channel=26
					-2, 8, -7, 5, -2, -3, 1, 9, 10,
					-- layer=2 filter=221 channel=27
					5, -5, -2, -13, -10, -6, -15, -4, -5,
					-- layer=2 filter=221 channel=28
					-16, -23, -7, -7, -12, -1, -4, -19, -7,
					-- layer=2 filter=221 channel=29
					0, -4, 0, 3, -2, 2, -2, 6, 1,
					-- layer=2 filter=221 channel=30
					-19, -15, 3, -16, -6, -10, -5, -17, -15,
					-- layer=2 filter=221 channel=31
					-5, -13, 0, -8, -9, -17, -13, 9, -14,
					-- layer=2 filter=221 channel=32
					-1, 8, -2, -4, 2, 11, 4, 8, -3,
					-- layer=2 filter=221 channel=33
					0, -12, -16, -11, -19, 0, 5, -7, 2,
					-- layer=2 filter=221 channel=34
					-5, -2, 1, -1, -4, -11, -7, -21, -18,
					-- layer=2 filter=221 channel=35
					-15, -14, -9, -2, 6, -6, -19, -8, -23,
					-- layer=2 filter=221 channel=36
					9, -12, 8, -8, 8, -5, 1, 1, -6,
					-- layer=2 filter=221 channel=37
					2, 4, -13, -14, -13, -5, -9, -9, -13,
					-- layer=2 filter=221 channel=38
					2, -10, -1, -14, -15, -1, -8, 2, -7,
					-- layer=2 filter=221 channel=39
					-5, 5, -14, -11, -2, -9, -6, -9, -8,
					-- layer=2 filter=221 channel=40
					-5, -5, 2, 8, -9, -17, -5, -9, -15,
					-- layer=2 filter=221 channel=41
					-6, 4, -2, -9, 9, 0, 7, -8, 5,
					-- layer=2 filter=221 channel=42
					3, -5, -6, -11, 9, 5, -17, 4, -1,
					-- layer=2 filter=221 channel=43
					-4, 4, -2, -3, -16, -3, -9, -10, -11,
					-- layer=2 filter=221 channel=44
					0, 0, -1, 4, 0, -1, 8, 0, 1,
					-- layer=2 filter=221 channel=45
					-4, -9, -13, 4, -9, -1, -12, -8, 0,
					-- layer=2 filter=221 channel=46
					-20, -14, -2, 0, 0, -8, 2, 4, -7,
					-- layer=2 filter=221 channel=47
					-2, -17, 3, -24, -5, -7, -8, -21, -12,
					-- layer=2 filter=221 channel=48
					-4, 0, 1, -6, 6, -5, -4, -3, 4,
					-- layer=2 filter=221 channel=49
					8, -10, -21, 9, -4, -9, 0, -16, -19,
					-- layer=2 filter=221 channel=50
					-4, -5, -2, 0, -13, 0, 4, -6, -3,
					-- layer=2 filter=221 channel=51
					-17, -13, -12, -6, -8, -6, -12, -7, -10,
					-- layer=2 filter=221 channel=52
					0, 0, -17, -2, -5, -13, -14, -4, -2,
					-- layer=2 filter=221 channel=53
					-3, -20, -6, -4, 1, -18, -1, -13, -6,
					-- layer=2 filter=221 channel=54
					3, -10, -11, -12, -11, -23, -17, 0, -16,
					-- layer=2 filter=221 channel=55
					-8, 2, -4, 8, 0, -8, 5, 4, 8,
					-- layer=2 filter=221 channel=56
					-9, 5, -7, -9, 0, -6, -2, -14, -17,
					-- layer=2 filter=221 channel=57
					1, -2, 1, 2, -8, 11, 11, 7, 2,
					-- layer=2 filter=221 channel=58
					-20, 3, -11, -13, -7, -5, -5, -3, -18,
					-- layer=2 filter=221 channel=59
					-8, -9, -23, 8, 0, 4, -18, 0, 6,
					-- layer=2 filter=221 channel=60
					-15, -9, 0, -16, -14, 18, -10, -13, -8,
					-- layer=2 filter=221 channel=61
					-3, -17, -9, 2, -23, -7, -5, -3, 12,
					-- layer=2 filter=221 channel=62
					-4, -8, -25, -4, -9, -15, 1, -5, 16,
					-- layer=2 filter=221 channel=63
					-4, -1, 9, -8, 0, 0, 5, 0, -11,
					-- layer=2 filter=221 channel=64
					-9, 3, 1, -11, 4, -5, -8, -6, 11,
					-- layer=2 filter=221 channel=65
					-14, -10, -12, 1, -18, -2, -16, 0, -2,
					-- layer=2 filter=221 channel=66
					0, 4, 3, 7, -3, 2, -3, 6, -2,
					-- layer=2 filter=221 channel=67
					-4, -10, -3, -7, -19, 4, -17, -13, 2,
					-- layer=2 filter=221 channel=68
					-8, 0, 9, 0, -5, -6, 10, -3, -2,
					-- layer=2 filter=221 channel=69
					-5, -10, -9, 0, -6, 3, 7, 6, -2,
					-- layer=2 filter=221 channel=70
					0, -16, 4, -3, -5, -7, -21, -9, -15,
					-- layer=2 filter=221 channel=71
					-4, 8, -4, -3, 5, 6, 2, -8, 7,
					-- layer=2 filter=221 channel=72
					-12, -22, -17, -28, -15, -18, -12, -6, 14,
					-- layer=2 filter=221 channel=73
					-2, -19, 4, -9, 0, -26, -9, -19, -15,
					-- layer=2 filter=221 channel=74
					3, -5, -17, -12, 4, 2, -10, -13, -16,
					-- layer=2 filter=221 channel=75
					-13, -15, 8, 0, 0, -1, 0, 2, -12,
					-- layer=2 filter=221 channel=76
					-12, -8, -16, -10, -23, -6, 5, -11, -20,
					-- layer=2 filter=221 channel=77
					5, 6, 4, 0, -2, 4, 8, -6, -10,
					-- layer=2 filter=221 channel=78
					-8, 0, -13, -10, -13, -6, -7, -15, -1,
					-- layer=2 filter=221 channel=79
					-5, -7, 3, 4, 6, -1, 8, 4, 8,
					-- layer=2 filter=221 channel=80
					-13, -2, -2, -4, -12, 2, -4, -5, 10,
					-- layer=2 filter=221 channel=81
					-2, -3, -6, 5, -11, 2, -5, -8, 5,
					-- layer=2 filter=221 channel=82
					-7, -6, -8, 0, 2, 2, 2, 2, 9,
					-- layer=2 filter=221 channel=83
					-11, -8, -5, -11, 0, -13, 0, 8, 5,
					-- layer=2 filter=221 channel=84
					1, 0, 2, 0, -8, 6, -3, 7, 9,
					-- layer=2 filter=221 channel=85
					-1, 9, 1, -9, 5, -5, -6, -2, 3,
					-- layer=2 filter=221 channel=86
					1, 1, 0, -7, -5, -1, -2, -9, -9,
					-- layer=2 filter=221 channel=87
					-1, -21, -8, -2, -9, -23, 5, -20, 1,
					-- layer=2 filter=221 channel=88
					-18, -13, -10, -17, 3, 0, -7, -17, -18,
					-- layer=2 filter=221 channel=89
					-16, -4, -10, 0, 1, -1, -6, -14, -3,
					-- layer=2 filter=221 channel=90
					-2, 3, 2, 0, -3, 9, -10, -9, 0,
					-- layer=2 filter=221 channel=91
					-5, -16, 1, -16, -14, -5, -8, -10, 1,
					-- layer=2 filter=221 channel=92
					-5, -1, -5, -14, -6, -8, -4, -4, 4,
					-- layer=2 filter=221 channel=93
					18, -17, 4, 10, -9, 1, 4, -2, 33,
					-- layer=2 filter=221 channel=94
					5, -3, -7, -11, -29, -14, 5, -5, 12,
					-- layer=2 filter=221 channel=95
					-5, -7, -3, 2, -7, 5, -9, 1, 0,
					-- layer=2 filter=221 channel=96
					4, -16, 10, 0, 2, 5, -3, -12, -14,
					-- layer=2 filter=221 channel=97
					-11, -10, 3, 5, -5, -14, 9, -6, 0,
					-- layer=2 filter=221 channel=98
					-26, -24, -5, -10, -1, -21, -16, -8, -10,
					-- layer=2 filter=221 channel=99
					7, -22, -31, 12, -20, -8, 8, -18, -17,
					-- layer=2 filter=221 channel=100
					-17, -6, -10, 6, 0, 4, -14, 8, -21,
					-- layer=2 filter=221 channel=101
					5, -3, -3, -7, 0, -2, 0, 0, -1,
					-- layer=2 filter=221 channel=102
					8, -8, -13, -6, -6, -17, 3, -2, 0,
					-- layer=2 filter=221 channel=103
					4, 6, 8, -9, -8, 1, -9, -9, 0,
					-- layer=2 filter=221 channel=104
					-3, -18, -18, -6, -19, -9, 2, -9, -17,
					-- layer=2 filter=221 channel=105
					-15, 0, 0, -2, 0, 3, -2, -11, 2,
					-- layer=2 filter=221 channel=106
					0, -3, -10, -19, 2, -7, -14, -14, -9,
					-- layer=2 filter=221 channel=107
					-1, 5, 4, -3, 7, -11, 6, -9, -7,
					-- layer=2 filter=221 channel=108
					-7, -5, 0, 4, -1, 6, -9, -12, -1,
					-- layer=2 filter=221 channel=109
					7, -2, 1, 7, 3, 9, 2, -1, 0,
					-- layer=2 filter=221 channel=110
					-4, -1, -2, -9, -14, -11, 2, -2, 4,
					-- layer=2 filter=221 channel=111
					1, 0, 3, 6, -1, -2, 0, -2, -1,
					-- layer=2 filter=221 channel=112
					-16, -10, 0, -19, -12, -8, -12, -7, -8,
					-- layer=2 filter=221 channel=113
					-17, -11, 8, 7, -11, -14, -5, -13, -11,
					-- layer=2 filter=221 channel=114
					6, -8, -4, 9, 6, -2, -8, 9, -4,
					-- layer=2 filter=221 channel=115
					6, -4, -8, -3, 3, -9, -10, 0, -7,
					-- layer=2 filter=221 channel=116
					-1, 0, -10, 1, 0, -12, -7, -23, 0,
					-- layer=2 filter=221 channel=117
					-3, -20, -8, -18, -28, -11, -4, -19, -22,
					-- layer=2 filter=221 channel=118
					-14, 1, -10, 4, -3, -3, -13, 2, 0,
					-- layer=2 filter=221 channel=119
					4, 0, -10, -7, -11, -9, 0, -9, -1,
					-- layer=2 filter=221 channel=120
					-4, 1, -3, -7, -4, 0, 7, 5, 8,
					-- layer=2 filter=221 channel=121
					10, 11, 11, -8, -3, 0, 5, -3, -2,
					-- layer=2 filter=221 channel=122
					-1, 6, -2, 8, 5, 4, 1, 0, 8,
					-- layer=2 filter=221 channel=123
					4, -24, -7, -7, -8, -8, -9, 1, 11,
					-- layer=2 filter=221 channel=124
					-10, -16, -4, -8, -12, -3, 12, 0, 14,
					-- layer=2 filter=221 channel=125
					-4, -6, 2, -9, -6, -2, -9, -9, 9,
					-- layer=2 filter=221 channel=126
					4, -1, 5, -6, -6, -18, -9, -12, -18,
					-- layer=2 filter=221 channel=127
					-8, -8, 5, 2, 7, 1, -16, -4, -14,
					-- layer=2 filter=222 channel=0
					-26, -17, -8, -13, -11, 2, 24, -5, -4,
					-- layer=2 filter=222 channel=1
					12, -1, -25, 22, 14, 8, -10, -2, -1,
					-- layer=2 filter=222 channel=2
					-3, -2, -2, 8, 1, -7, 6, 11, -4,
					-- layer=2 filter=222 channel=3
					-7, -41, -22, -13, -32, -19, -4, -5, 2,
					-- layer=2 filter=222 channel=4
					-30, -5, -27, -7, 16, -27, 34, -18, -30,
					-- layer=2 filter=222 channel=5
					0, -1, -19, 17, 0, -8, -2, -11, 0,
					-- layer=2 filter=222 channel=6
					13, 5, 14, 8, 39, 20, 7, 4, 25,
					-- layer=2 filter=222 channel=7
					-4, 11, 0, 5, 18, 42, -5, -40, -19,
					-- layer=2 filter=222 channel=8
					-7, -1, 9, -8, 0, 6, 4, -6, 0,
					-- layer=2 filter=222 channel=9
					5, -42, -10, -2, 0, 7, 1, 28, 32,
					-- layer=2 filter=222 channel=10
					-37, -13, -5, -4, 9, 4, 15, -17, -6,
					-- layer=2 filter=222 channel=11
					7, 21, -6, 13, 11, -1, -5, -3, -9,
					-- layer=2 filter=222 channel=12
					15, -3, -42, -7, -14, 10, -40, -13, -26,
					-- layer=2 filter=222 channel=13
					12, -1, 0, -3, 3, -6, 8, 6, 1,
					-- layer=2 filter=222 channel=14
					19, 10, -6, 13, -6, -6, -16, 0, 0,
					-- layer=2 filter=222 channel=15
					15, 4, 29, 55, -21, 6, -10, -64, 6,
					-- layer=2 filter=222 channel=16
					-5, -4, -24, 30, 19, 28, 23, 7, 7,
					-- layer=2 filter=222 channel=17
					-4, 0, -6, 10, -1, 0, 7, 6, -10,
					-- layer=2 filter=222 channel=18
					23, 12, 42, 9, 29, 12, 12, -25, 2,
					-- layer=2 filter=222 channel=19
					-18, 12, -22, 31, 22, 21, -22, 2, -26,
					-- layer=2 filter=222 channel=20
					7, 4, 2, 7, 3, -8, -2, -3, 8,
					-- layer=2 filter=222 channel=21
					14, 5, 19, 17, 16, 1, 15, 1, 1,
					-- layer=2 filter=222 channel=22
					-3, -8, 0, 7, -1, 10, 10, 5, 2,
					-- layer=2 filter=222 channel=23
					-19, -19, -26, 14, -5, -10, 0, 1, -3,
					-- layer=2 filter=222 channel=24
					13, -50, -4, -79, -71, -1, -20, -28, 35,
					-- layer=2 filter=222 channel=25
					-9, -37, -31, -33, -61, -3, -17, -19, 41,
					-- layer=2 filter=222 channel=26
					-2, -3, -1, -8, 2, -5, -9, 10, 0,
					-- layer=2 filter=222 channel=27
					-7, -8, -4, -3, -1, -6, 16, -2, -5,
					-- layer=2 filter=222 channel=28
					-28, 20, 34, 18, -30, -9, 40, 27, 11,
					-- layer=2 filter=222 channel=29
					-5, 4, -9, -7, 8, 1, 9, 3, -1,
					-- layer=2 filter=222 channel=30
					-16, -51, -2, -1, -12, 13, 8, 32, 19,
					-- layer=2 filter=222 channel=31
					-35, 20, -35, -5, -24, 49, -10, 10, 42,
					-- layer=2 filter=222 channel=32
					-1, -6, 0, 2, 3, -5, 0, 11, -5,
					-- layer=2 filter=222 channel=33
					6, 39, -22, 13, -10, -7, -3, -23, 5,
					-- layer=2 filter=222 channel=34
					-9, 65, 24, -13, 53, -2, -19, 21, 18,
					-- layer=2 filter=222 channel=35
					-6, -4, 7, 2, -9, -9, 30, -22, -3,
					-- layer=2 filter=222 channel=36
					-12, 0, 0, -14, -1, -6, -4, 9, 1,
					-- layer=2 filter=222 channel=37
					21, 21, -9, 3, 3, -1, 2, -2, -10,
					-- layer=2 filter=222 channel=38
					-3, 0, 26, 10, 5, 5, 28, 19, -6,
					-- layer=2 filter=222 channel=39
					-20, -25, -40, 28, 30, 40, -5, -24, 0,
					-- layer=2 filter=222 channel=40
					-5, -64, 34, -32, -4, 25, 10, 20, 40,
					-- layer=2 filter=222 channel=41
					5, -4, -1, 10, 6, -4, 6, 6, 9,
					-- layer=2 filter=222 channel=42
					-8, -14, -9, -10, -16, 42, -11, 14, 15,
					-- layer=2 filter=222 channel=43
					2, 16, -12, 24, 4, -33, 2, -6, -24,
					-- layer=2 filter=222 channel=44
					-4, -1, 0, -3, -1, 11, 2, -6, 1,
					-- layer=2 filter=222 channel=45
					-57, -51, -41, 9, -38, -8, 33, 35, 32,
					-- layer=2 filter=222 channel=46
					-26, -29, -21, 8, 14, -3, 26, 25, 2,
					-- layer=2 filter=222 channel=47
					-59, -30, -18, 18, -21, -2, 9, -3, 23,
					-- layer=2 filter=222 channel=48
					1, 1, -1, 10, -4, 6, 8, 7, 1,
					-- layer=2 filter=222 channel=49
					-4, -13, 15, -15, 38, 14, -17, -22, -37,
					-- layer=2 filter=222 channel=50
					12, 6, -14, -33, -5, 0, 13, 0, -14,
					-- layer=2 filter=222 channel=51
					0, 25, -5, 0, 18, -5, 8, -7, -5,
					-- layer=2 filter=222 channel=52
					19, 0, 6, -10, 8, -45, -8, -1, -38,
					-- layer=2 filter=222 channel=53
					-31, -22, -4, 9, 55, -14, 18, 35, 3,
					-- layer=2 filter=222 channel=54
					-5, 0, -57, -13, -3, -6, -11, -21, 2,
					-- layer=2 filter=222 channel=55
					7, -5, 6, -4, 10, -13, 0, -4, -2,
					-- layer=2 filter=222 channel=56
					20, 21, -15, 26, 8, 16, 11, -7, -1,
					-- layer=2 filter=222 channel=57
					-18, 0, -4, 6, 12, 0, -9, -2, -11,
					-- layer=2 filter=222 channel=58
					24, 3, -25, 21, -15, 4, -59, 8, -10,
					-- layer=2 filter=222 channel=59
					20, 53, 0, 34, 39, 19, -6, 25, -34,
					-- layer=2 filter=222 channel=60
					13, -8, 11, 18, 34, 19, 7, 8, -23,
					-- layer=2 filter=222 channel=61
					-1, -2, 0, 5, 8, 10, 41, 8, -7,
					-- layer=2 filter=222 channel=62
					-6, -13, -2, -5, 9, -17, -42, -17, -20,
					-- layer=2 filter=222 channel=63
					-18, -40, -19, 1, -14, 20, -2, 16, 26,
					-- layer=2 filter=222 channel=64
					-6, -41, -24, -19, 9, 30, -15, 13, 28,
					-- layer=2 filter=222 channel=65
					23, 1, 11, 30, 33, -1, 20, 14, 6,
					-- layer=2 filter=222 channel=66
					-3, 4, -8, 3, 27, 11, -20, -9, -27,
					-- layer=2 filter=222 channel=67
					5, 0, 2, 8, 10, 18, 36, 50, 29,
					-- layer=2 filter=222 channel=68
					7, 0, -3, -10, 7, 1, -6, -3, 3,
					-- layer=2 filter=222 channel=69
					2, -9, -8, 18, 31, 14, -23, 11, 0,
					-- layer=2 filter=222 channel=70
					-7, 0, -8, -6, -11, -38, 22, -2, 4,
					-- layer=2 filter=222 channel=71
					7, -6, 13, 13, 15, 27, 6, -1, 16,
					-- layer=2 filter=222 channel=72
					-2, 30, 22, 4, -8, 8, -23, -22, -41,
					-- layer=2 filter=222 channel=73
					-44, -4, 47, -21, 19, 14, -9, 25, 33,
					-- layer=2 filter=222 channel=74
					-24, -2, -6, -11, -4, 15, 36, 37, 0,
					-- layer=2 filter=222 channel=75
					2, -1, -26, -35, -22, -20, -6, -13, 59,
					-- layer=2 filter=222 channel=76
					-15, -15, 5, 15, 37, -26, -1, 10, 39,
					-- layer=2 filter=222 channel=77
					0, 5, 0, 0, 11, -8, 4, 4, 11,
					-- layer=2 filter=222 channel=78
					21, 25, -21, -2, -24, -17, 0, -1, 1,
					-- layer=2 filter=222 channel=79
					-7, 8, 4, 5, -8, 3, 9, -4, 9,
					-- layer=2 filter=222 channel=80
					-6, -12, -28, -8, 21, 23, 15, 24, 7,
					-- layer=2 filter=222 channel=81
					1, -9, 0, -2, 4, 0, 1, 2, 3,
					-- layer=2 filter=222 channel=82
					-8, 1, 0, 3, 8, -5, 7, 0, 3,
					-- layer=2 filter=222 channel=83
					12, -28, -17, -24, -37, -28, -4, 14, 6,
					-- layer=2 filter=222 channel=84
					6, 9, 4, -1, -2, 0, -6, -1, 10,
					-- layer=2 filter=222 channel=85
					-2, -1, 0, 7, -12, -12, -5, -2, -2,
					-- layer=2 filter=222 channel=86
					6, 7, -2, -16, 15, 23, -6, -8, -11,
					-- layer=2 filter=222 channel=87
					65, 47, 15, 71, 16, 6, 25, 18, -16,
					-- layer=2 filter=222 channel=88
					19, -8, -9, 8, -2, 12, 18, 29, 3,
					-- layer=2 filter=222 channel=89
					25, 24, -21, -4, 5, -6, -51, 6, -35,
					-- layer=2 filter=222 channel=90
					-9, -9, 1, 5, -1, 11, 1, 2, 12,
					-- layer=2 filter=222 channel=91
					40, -16, -21, -20, -24, 1, 15, -15, -40,
					-- layer=2 filter=222 channel=92
					14, 7, -29, 18, -10, -1, -28, -32, -31,
					-- layer=2 filter=222 channel=93
					40, 14, -47, -6, 9, -5, -31, -30, 31,
					-- layer=2 filter=222 channel=94
					-36, 19, 22, -5, -5, 17, 25, 24, 13,
					-- layer=2 filter=222 channel=95
					-1, -14, 0, -8, 0, -3, -6, 4, 8,
					-- layer=2 filter=222 channel=96
					-18, 29, -33, -18, 26, 18, 6, -7, -6,
					-- layer=2 filter=222 channel=97
					16, -3, -9, -6, -17, 4, -8, -9, 9,
					-- layer=2 filter=222 channel=98
					-9, -14, 5, 23, -36, 6, 18, 8, 16,
					-- layer=2 filter=222 channel=99
					-3, 8, 42, 8, 40, 22, 9, 8, 5,
					-- layer=2 filter=222 channel=100
					14, 17, 19, -13, -21, -10, 17, -6, 13,
					-- layer=2 filter=222 channel=101
					16, -7, -7, -15, 1, 34, -44, -24, 10,
					-- layer=2 filter=222 channel=102
					11, 36, -11, 24, 46, -32, -3, -19, -17,
					-- layer=2 filter=222 channel=103
					7, -10, 15, 60, -17, 31, 6, 12, 0,
					-- layer=2 filter=222 channel=104
					24, 38, 19, 16, 54, 7, 28, -13, 1,
					-- layer=2 filter=222 channel=105
					-3, -20, -1, 23, -34, 26, 51, 47, -11,
					-- layer=2 filter=222 channel=106
					13, 14, -15, -39, -65, -7, 8, -18, 38,
					-- layer=2 filter=222 channel=107
					-20, -35, 17, 37, 29, 32, -17, 13, -3,
					-- layer=2 filter=222 channel=108
					-13, -2, 5, -12, -5, -8, -16, -19, 5,
					-- layer=2 filter=222 channel=109
					-6, -9, 18, -14, -8, -12, -12, 0, 9,
					-- layer=2 filter=222 channel=110
					-17, -16, -17, -15, -9, 16, -27, -8, 38,
					-- layer=2 filter=222 channel=111
					3, -2, 0, 0, 12, -1, 0, 0, 2,
					-- layer=2 filter=222 channel=112
					6, -25, -1, -3, 15, 32, 22, -5, -17,
					-- layer=2 filter=222 channel=113
					-19, -41, 12, -15, -10, -8, 7, 13, 1,
					-- layer=2 filter=222 channel=114
					0, -5, 2, 2, 7, 10, 9, 16, 4,
					-- layer=2 filter=222 channel=115
					0, -1, -1, 1, 7, 10, 3, -3, 5,
					-- layer=2 filter=222 channel=116
					43, 30, 32, 53, 11, -27, 17, -21, -19,
					-- layer=2 filter=222 channel=117
					-15, 55, 13, 8, 1, 31, 13, 7, -11,
					-- layer=2 filter=222 channel=118
					-18, -2, -26, 1, 0, -12, 4, -1, -19,
					-- layer=2 filter=222 channel=119
					12, -26, 18, -3, 8, -9, 8, -12, 12,
					-- layer=2 filter=222 channel=120
					0, 5, 8, 2, -5, 2, 9, -5, -3,
					-- layer=2 filter=222 channel=121
					4, 3, 6, -4, 3, 5, 6, 11, 4,
					-- layer=2 filter=222 channel=122
					14, 0, 0, 0, 6, -2, -1, -2, 8,
					-- layer=2 filter=222 channel=123
					14, 6, 24, 29, 6, 35, -9, 4, 13,
					-- layer=2 filter=222 channel=124
					-7, 22, -41, 21, 7, 9, -52, -32, 15,
					-- layer=2 filter=222 channel=125
					-9, 0, 1, 0, -10, -4, 5, 4, -9,
					-- layer=2 filter=222 channel=126
					-47, -46, 21, 14, -28, 20, 6, -45, -12,
					-- layer=2 filter=222 channel=127
					-6, -13, -24, 5, 9, -25, -9, 8, -5,
					-- layer=2 filter=223 channel=0
					14, 25, -10, -19, -25, -34, -31, 1, -6,
					-- layer=2 filter=223 channel=1
					25, -9, 23, 18, -6, 12, -8, -16, -53,
					-- layer=2 filter=223 channel=2
					-3, -10, -2, 4, 4, -7, 3, -3, -10,
					-- layer=2 filter=223 channel=3
					51, -14, -51, 7, -55, -22, -3, 22, 13,
					-- layer=2 filter=223 channel=4
					8, 14, 1, -5, 12, -44, 17, 18, -10,
					-- layer=2 filter=223 channel=5
					-8, 31, 21, 4, 0, -15, -26, 5, 0,
					-- layer=2 filter=223 channel=6
					39, 24, -59, 45, 24, -33, 18, 15, 45,
					-- layer=2 filter=223 channel=7
					-18, 27, 9, -17, -9, 3, 51, 21, 19,
					-- layer=2 filter=223 channel=8
					-3, 4, -1, 0, 2, 1, 6, -4, -9,
					-- layer=2 filter=223 channel=9
					1, 0, 0, 53, 20, -33, -24, -10, -21,
					-- layer=2 filter=223 channel=10
					46, -15, -25, -12, -44, -71, 1, 5, -4,
					-- layer=2 filter=223 channel=11
					-4, -5, 15, 16, -22, -6, -2, -16, 5,
					-- layer=2 filter=223 channel=12
					16, 3, 21, 14, 1, 0, 13, -16, -20,
					-- layer=2 filter=223 channel=13
					-1, -8, 4, 0, 7, 8, -9, 7, 4,
					-- layer=2 filter=223 channel=14
					5, 9, 32, 11, 18, -12, -25, -29, -39,
					-- layer=2 filter=223 channel=15
					3, -29, -16, -10, 9, 25, -9, -22, -4,
					-- layer=2 filter=223 channel=16
					45, 30, -2, 8, 0, -35, -7, -11, 0,
					-- layer=2 filter=223 channel=17
					1, 0, -5, -8, 10, -4, 11, -8, 7,
					-- layer=2 filter=223 channel=18
					40, -47, -48, -13, -48, -17, -40, -16, 4,
					-- layer=2 filter=223 channel=19
					-24, 10, 9, 20, 11, 0, 30, -12, -8,
					-- layer=2 filter=223 channel=20
					-2, 10, -3, -6, 8, -10, -1, -11, 4,
					-- layer=2 filter=223 channel=21
					-3, 0, -5, 4, -13, -1, -6, -12, -1,
					-- layer=2 filter=223 channel=22
					4, 8, -1, -2, 10, 0, 9, -1, 8,
					-- layer=2 filter=223 channel=23
					27, 5, -26, 32, -34, -14, 20, 33, 23,
					-- layer=2 filter=223 channel=24
					57, 43, -27, 27, -25, -64, -3, -25, -31,
					-- layer=2 filter=223 channel=25
					41, 43, 14, 27, -1, -36, 23, -23, -2,
					-- layer=2 filter=223 channel=26
					-5, 0, -10, 0, 8, -7, 3, 0, 5,
					-- layer=2 filter=223 channel=27
					4, 11, 11, 8, -25, -3, -8, -51, -40,
					-- layer=2 filter=223 channel=28
					47, 36, 14, -62, -56, -71, 8, -7, 13,
					-- layer=2 filter=223 channel=29
					3, 3, 1, -8, 8, -9, 4, 1, -2,
					-- layer=2 filter=223 channel=30
					-2, -10, 0, -2, 2, -14, -6, -13, -77,
					-- layer=2 filter=223 channel=31
					34, -13, -36, -8, -41, 23, -14, -51, -25,
					-- layer=2 filter=223 channel=32
					4, 0, 6, 9, 0, 3, 0, -5, 8,
					-- layer=2 filter=223 channel=33
					-29, -21, 9, 6, 9, -20, 6, 15, 6,
					-- layer=2 filter=223 channel=34
					-39, 28, -25, 5, 18, -9, 31, 12, 14,
					-- layer=2 filter=223 channel=35
					20, 49, -16, -45, -28, -44, 12, 11, -2,
					-- layer=2 filter=223 channel=36
					-3, -4, -12, -2, 0, 6, -8, 0, -2,
					-- layer=2 filter=223 channel=37
					4, -13, -1, -4, 0, 35, -20, -21, 3,
					-- layer=2 filter=223 channel=38
					9, 31, 17, -1, -39, -8, -50, -53, -64,
					-- layer=2 filter=223 channel=39
					4, 15, -20, 20, -17, -44, 16, 4, 6,
					-- layer=2 filter=223 channel=40
					15, -31, -60, -57, -5, -37, -39, 31, 37,
					-- layer=2 filter=223 channel=41
					8, -1, 1, 6, 7, -3, 6, -4, -5,
					-- layer=2 filter=223 channel=42
					45, 25, -6, 23, -17, 13, 20, 34, 38,
					-- layer=2 filter=223 channel=43
					17, -20, -40, -89, -47, -17, -17, 41, 42,
					-- layer=2 filter=223 channel=44
					-1, -8, 0, -4, 2, 9, 4, 11, 7,
					-- layer=2 filter=223 channel=45
					3, 16, 18, 38, -24, -18, 14, -22, -25,
					-- layer=2 filter=223 channel=46
					-26, -6, -10, -22, -65, -73, 19, -1, -23,
					-- layer=2 filter=223 channel=47
					42, 21, -9, -15, -71, -58, -52, -65, -10,
					-- layer=2 filter=223 channel=48
					-1, 5, -10, 9, -4, 10, -2, 4, 3,
					-- layer=2 filter=223 channel=49
					15, -17, 20, 9, -58, -5, -56, -40, 8,
					-- layer=2 filter=223 channel=50
					-8, -13, 1, -3, -21, -7, 0, 10, 14,
					-- layer=2 filter=223 channel=51
					12, 10, 9, -7, -10, -7, -28, -13, 4,
					-- layer=2 filter=223 channel=52
					-31, -27, -17, -53, -28, 0, 42, 10, 25,
					-- layer=2 filter=223 channel=53
					-40, 43, -12, 0, -24, -2, 2, 11, -55,
					-- layer=2 filter=223 channel=54
					14, -26, -79, -4, -35, -21, 30, 9, 29,
					-- layer=2 filter=223 channel=55
					10, 6, -3, 12, 0, 5, 8, 8, 6,
					-- layer=2 filter=223 channel=56
					26, 0, 3, 16, -6, -8, -8, -14, 6,
					-- layer=2 filter=223 channel=57
					10, 0, -12, 5, -8, -3, -10, 0, 0,
					-- layer=2 filter=223 channel=58
					23, 0, 19, 17, 21, 23, 14, -1, -16,
					-- layer=2 filter=223 channel=59
					-2, 1, -2, 10, 3, 7, -11, 1, -10,
					-- layer=2 filter=223 channel=60
					7, 21, -7, 3, 15, 20, -42, -41, -25,
					-- layer=2 filter=223 channel=61
					5, 12, -16, -12, 9, -23, -39, -45, -4,
					-- layer=2 filter=223 channel=62
					-12, -29, -38, -5, -11, -26, 19, 3, 52,
					-- layer=2 filter=223 channel=63
					9, 0, -7, -3, -18, -24, -19, 1, 10,
					-- layer=2 filter=223 channel=64
					12, -3, -39, 31, 10, -25, -1, -2, -23,
					-- layer=2 filter=223 channel=65
					38, 2, -20, 0, 11, -15, 11, -8, 25,
					-- layer=2 filter=223 channel=66
					-11, -40, -19, 0, -41, -6, 9, -39, 15,
					-- layer=2 filter=223 channel=67
					-27, 27, 6, 22, 9, -12, -10, 13, -25,
					-- layer=2 filter=223 channel=68
					-5, -7, -5, -3, -8, 5, 4, 0, -11,
					-- layer=2 filter=223 channel=69
					-2, -5, -8, 10, -2, -31, -19, -5, -8,
					-- layer=2 filter=223 channel=70
					40, 34, -12, -51, -7, -31, 19, 24, 14,
					-- layer=2 filter=223 channel=71
					-24, 12, 16, 9, 0, -9, 33, -21, -34,
					-- layer=2 filter=223 channel=72
					37, 8, 7, -27, 48, 35, 19, 16, -15,
					-- layer=2 filter=223 channel=73
					-22, 16, 16, -36, -41, 57, -55, 2, -22,
					-- layer=2 filter=223 channel=74
					-14, -16, -5, -21, 24, 7, -72, -7, -45,
					-- layer=2 filter=223 channel=75
					15, 2, 0, -11, 6, -56, 47, 56, 24,
					-- layer=2 filter=223 channel=76
					-31, 25, 2, -19, -38, 15, -13, -3, 32,
					-- layer=2 filter=223 channel=77
					3, 0, -5, 5, 6, -6, 8, 0, -4,
					-- layer=2 filter=223 channel=78
					10, -2, -33, -28, -55, -18, 0, -16, 18,
					-- layer=2 filter=223 channel=79
					-8, -11, 5, -9, 3, 0, -8, 3, 5,
					-- layer=2 filter=223 channel=80
					-13, 14, -34, -33, -37, -58, -30, 15, 17,
					-- layer=2 filter=223 channel=81
					8, 2, -11, 6, -9, -8, -9, -7, -12,
					-- layer=2 filter=223 channel=82
					6, -8, -11, -1, -7, 3, 6, 10, -8,
					-- layer=2 filter=223 channel=83
					34, 13, -2, -24, -9, -34, -19, -3, -15,
					-- layer=2 filter=223 channel=84
					-3, 2, 0, 8, -10, 2, -7, 5, 11,
					-- layer=2 filter=223 channel=85
					-1, 0, -9, 13, -3, 7, 0, 3, -6,
					-- layer=2 filter=223 channel=86
					-3, 11, 2, 5, 22, 2, 12, 9, -1,
					-- layer=2 filter=223 channel=87
					7, 8, -20, 24, 10, -13, 2, 10, 37,
					-- layer=2 filter=223 channel=88
					-19, -9, 11, 5, -6, 31, -60, -4, -21,
					-- layer=2 filter=223 channel=89
					11, 0, 31, 17, 28, 34, 17, 1, -24,
					-- layer=2 filter=223 channel=90
					5, 9, -5, -11, -12, 2, 4, 11, 1,
					-- layer=2 filter=223 channel=91
					-8, 0, 7, 13, 33, 50, 31, 41, 5,
					-- layer=2 filter=223 channel=92
					3, -7, 38, 31, 27, 27, 1, -37, -22,
					-- layer=2 filter=223 channel=93
					-33, 5, -12, 8, 7, -26, 67, 32, 11,
					-- layer=2 filter=223 channel=94
					-14, 9, -24, 14, 23, 12, 5, 7, 19,
					-- layer=2 filter=223 channel=95
					7, 20, 8, 17, 6, 17, -1, 10, 2,
					-- layer=2 filter=223 channel=96
					2, -28, 13, 43, 47, 45, 19, 28, 13,
					-- layer=2 filter=223 channel=97
					30, 50, 5, 11, -22, -50, -20, -24, -27,
					-- layer=2 filter=223 channel=98
					24, 0, -17, -76, -42, -33, -27, -11, 16,
					-- layer=2 filter=223 channel=99
					-54, 17, 1, 0, 23, 30, 44, 8, 0,
					-- layer=2 filter=223 channel=100
					52, 32, -20, -7, -7, -17, 9, 1, 2,
					-- layer=2 filter=223 channel=101
					2, -2, -14, 26, 2, 16, 61, 16, -21,
					-- layer=2 filter=223 channel=102
					0, -21, -34, 33, 22, 19, 38, 5, 10,
					-- layer=2 filter=223 channel=103
					-34, -14, -17, 8, -4, 17, -4, 25, 32,
					-- layer=2 filter=223 channel=104
					18, -30, 31, -4, -28, 17, -2, 23, 54,
					-- layer=2 filter=223 channel=105
					19, -16, 27, -6, 21, 24, -10, -7, 60,
					-- layer=2 filter=223 channel=106
					29, 45, 0, 53, 19, 4, 29, 5, -41,
					-- layer=2 filter=223 channel=107
					-18, 15, 58, 9, -14, 9, 21, 39, 34,
					-- layer=2 filter=223 channel=108
					-21, -9, 11, 38, -10, 7, -10, -34, -46,
					-- layer=2 filter=223 channel=109
					-2, -6, 3, -9, 12, 7, -5, -3, 8,
					-- layer=2 filter=223 channel=110
					40, 20, -39, 26, 20, -4, 0, 7, -40,
					-- layer=2 filter=223 channel=111
					6, 0, 5, 1, 6, -10, 8, 4, 0,
					-- layer=2 filter=223 channel=112
					52, 37, 22, 2, -11, -9, -45, -55, -9,
					-- layer=2 filter=223 channel=113
					35, 5, 1, -29, -1, -3, -18, 11, -57,
					-- layer=2 filter=223 channel=114
					-13, -9, 2, -9, -8, -4, -17, -5, -7,
					-- layer=2 filter=223 channel=115
					0, -2, 6, -8, -8, 1, 1, 8, 2,
					-- layer=2 filter=223 channel=116
					8, -22, -39, 18, -10, -1, 4, 3, 37,
					-- layer=2 filter=223 channel=117
					-56, -13, 21, -20, -19, -27, 38, -2, -13,
					-- layer=2 filter=223 channel=118
					-16, -19, -38, -84, -78, -3, -39, 50, 52,
					-- layer=2 filter=223 channel=119
					22, 53, -12, 28, -10, -42, 18, -6, 0,
					-- layer=2 filter=223 channel=120
					3, -1, -7, -3, 2, -7, -7, 6, 8,
					-- layer=2 filter=223 channel=121
					5, -6, 4, 0, 3, -4, -8, -1, -2,
					-- layer=2 filter=223 channel=122
					5, 2, -11, -4, -13, 1, 5, 2, -1,
					-- layer=2 filter=223 channel=123
					-3, -6, -39, -41, 2, 2, -3, 39, 13,
					-- layer=2 filter=223 channel=124
					15, -34, -48, 18, -9, -6, 1, 23, 34,
					-- layer=2 filter=223 channel=125
					7, 6, -9, 3, 0, 5, 3, -5, 0,
					-- layer=2 filter=223 channel=126
					-15, 6, 18, 9, 30, 4, 0, -26, -3,
					-- layer=2 filter=223 channel=127
					16, -7, 13, -16, -10, -24, -31, 0, -8,
					-- layer=2 filter=224 channel=0
					2, -19, 2, 15, -3, 2, -1, 0, 0,
					-- layer=2 filter=224 channel=1
					-14, -19, -6, -4, -21, -4, 2, 4, 11,
					-- layer=2 filter=224 channel=2
					-3, 2, -6, -3, -2, 1, -4, 6, 3,
					-- layer=2 filter=224 channel=3
					2, 14, -6, 7, -22, -4, 5, 12, 3,
					-- layer=2 filter=224 channel=4
					-7, -17, -10, -6, -18, -1, -9, -3, -17,
					-- layer=2 filter=224 channel=5
					0, 2, -12, 2, -10, -18, -14, 2, -15,
					-- layer=2 filter=224 channel=6
					-2, -1, -13, -7, -7, -5, -22, 11, -16,
					-- layer=2 filter=224 channel=7
					10, 2, -17, -5, 1, 7, -5, -12, -7,
					-- layer=2 filter=224 channel=8
					-4, -1, 0, -2, -10, -4, -2, -6, -3,
					-- layer=2 filter=224 channel=9
					-7, -4, -16, -15, -5, -6, -4, 3, -1,
					-- layer=2 filter=224 channel=10
					-8, -2, 3, -3, -2, -6, 11, -11, -6,
					-- layer=2 filter=224 channel=11
					-10, -6, -7, 8, -10, -3, 1, 0, -12,
					-- layer=2 filter=224 channel=12
					-2, -12, -22, -8, 7, -14, -8, -4, 16,
					-- layer=2 filter=224 channel=13
					1, 5, -3, -11, -4, -11, -2, -8, -8,
					-- layer=2 filter=224 channel=14
					2, -14, -21, -3, 0, -4, -1, 3, 4,
					-- layer=2 filter=224 channel=15
					-4, 7, -9, -1, 6, -6, -17, 7, -16,
					-- layer=2 filter=224 channel=16
					-13, -2, -15, -11, -16, 0, -7, -23, -7,
					-- layer=2 filter=224 channel=17
					-6, -6, 7, -4, 1, 0, -2, 0, 6,
					-- layer=2 filter=224 channel=18
					-15, 7, -14, -12, 5, -5, -2, -16, -4,
					-- layer=2 filter=224 channel=19
					-13, -9, -7, -6, 2, -8, 4, -22, -23,
					-- layer=2 filter=224 channel=20
					-10, 1, -3, 2, -9, -7, 6, 0, -10,
					-- layer=2 filter=224 channel=21
					-5, -11, 5, -2, -7, -9, -3, 5, -1,
					-- layer=2 filter=224 channel=22
					-4, 6, -7, -2, 0, 3, -6, -10, 3,
					-- layer=2 filter=224 channel=23
					-9, -14, -14, -3, -14, -14, -14, -20, -7,
					-- layer=2 filter=224 channel=24
					0, -5, -4, 4, -7, 0, -6, -9, 2,
					-- layer=2 filter=224 channel=25
					-5, 8, 3, 0, -8, 0, 9, 5, 0,
					-- layer=2 filter=224 channel=26
					-7, 3, -7, -8, 0, -1, -3, -1, -5,
					-- layer=2 filter=224 channel=27
					-17, -7, -9, 1, -5, -25, 1, 18, -12,
					-- layer=2 filter=224 channel=28
					6, -7, 19, -8, -6, -17, -18, -8, -3,
					-- layer=2 filter=224 channel=29
					-12, -9, -8, 1, -7, 1, 8, -8, -7,
					-- layer=2 filter=224 channel=30
					-20, -18, 0, -7, -17, -5, -5, -8, -2,
					-- layer=2 filter=224 channel=31
					-1, -1, -2, -9, -3, 8, -19, 4, 6,
					-- layer=2 filter=224 channel=32
					-7, -10, 3, 2, 1, -10, -6, 10, -9,
					-- layer=2 filter=224 channel=33
					-8, -12, -13, -6, -5, 0, 1, 3, 1,
					-- layer=2 filter=224 channel=34
					-4, 6, 3, 0, -1, -8, -8, -5, -1,
					-- layer=2 filter=224 channel=35
					-5, -13, 6, -7, -10, -10, -14, -1, 10,
					-- layer=2 filter=224 channel=36
					-11, 6, -10, -4, -6, -2, -10, 1, -6,
					-- layer=2 filter=224 channel=37
					-6, 1, 4, 4, -7, 1, 0, 15, -12,
					-- layer=2 filter=224 channel=38
					-8, -20, -16, -1, 2, 1, 15, 11, -13,
					-- layer=2 filter=224 channel=39
					-2, -16, 1, -12, -7, -1, -17, -10, -17,
					-- layer=2 filter=224 channel=40
					0, 0, 4, 0, 4, 4, 6, 1, -4,
					-- layer=2 filter=224 channel=41
					-5, 2, 0, -7, -5, -10, -1, -1, -2,
					-- layer=2 filter=224 channel=42
					-11, 1, -3, -3, -19, -19, -15, -22, 2,
					-- layer=2 filter=224 channel=43
					-11, 14, -1, 0, -5, -13, -3, -3, -7,
					-- layer=2 filter=224 channel=44
					-8, 10, -7, -1, 7, 4, 3, 10, -9,
					-- layer=2 filter=224 channel=45
					-15, -3, -10, -3, -17, 3, -4, -10, -1,
					-- layer=2 filter=224 channel=46
					-14, -16, -17, -14, -19, -6, 9, -10, -11,
					-- layer=2 filter=224 channel=47
					1, 2, 0, 2, -7, -2, 0, 2, -1,
					-- layer=2 filter=224 channel=48
					-10, 8, 1, -6, 8, 8, -1, 4, 2,
					-- layer=2 filter=224 channel=49
					3, -3, -15, -12, 0, -10, -4, -16, -10,
					-- layer=2 filter=224 channel=50
					6, 8, -10, 3, -10, -1, 1, -3, 2,
					-- layer=2 filter=224 channel=51
					-12, -4, 3, 7, -11, -1, -12, -8, -18,
					-- layer=2 filter=224 channel=52
					0, -7, -7, -12, -5, 3, -13, -18, -9,
					-- layer=2 filter=224 channel=53
					2, -12, -22, 1, -5, -5, -21, -13, -7,
					-- layer=2 filter=224 channel=54
					0, -7, -7, -8, 4, -4, -18, -8, -10,
					-- layer=2 filter=224 channel=55
					8, 0, 2, 0, -1, -3, -5, 3, -9,
					-- layer=2 filter=224 channel=56
					-14, 7, 12, 4, -7, -13, 0, 12, -10,
					-- layer=2 filter=224 channel=57
					-6, -1, -7, -5, 0, -7, -7, 10, 10,
					-- layer=2 filter=224 channel=58
					-1, -5, -5, -3, -4, -3, -17, 0, -13,
					-- layer=2 filter=224 channel=59
					0, -18, -10, -1, 0, 6, -10, -2, -2,
					-- layer=2 filter=224 channel=60
					8, -1, -5, -15, -2, 2, -21, -3, -14,
					-- layer=2 filter=224 channel=61
					22, -1, -6, -7, -8, 0, -9, 7, -2,
					-- layer=2 filter=224 channel=62
					-4, 3, 0, -1, 4, -5, -5, 6, 0,
					-- layer=2 filter=224 channel=63
					-5, -13, -8, -4, -3, 4, -12, -19, -1,
					-- layer=2 filter=224 channel=64
					-7, 0, -14, -13, -1, -3, -14, -20, 0,
					-- layer=2 filter=224 channel=65
					5, -4, -4, -8, -1, 11, -3, -6, -15,
					-- layer=2 filter=224 channel=66
					-3, 2, -2, -4, -7, 0, -5, 5, 4,
					-- layer=2 filter=224 channel=67
					-13, -4, 4, -11, -20, 0, 8, -9, -12,
					-- layer=2 filter=224 channel=68
					-1, -7, -5, -7, -7, -11, -10, 5, 2,
					-- layer=2 filter=224 channel=69
					3, 2, -10, -19, -17, -9, -19, -11, -7,
					-- layer=2 filter=224 channel=70
					2, -12, 14, 10, 0, -4, -8, -3, 11,
					-- layer=2 filter=224 channel=71
					-2, -13, -16, 0, -16, -11, 12, -4, -8,
					-- layer=2 filter=224 channel=72
					-9, -18, -5, 0, 0, 4, -8, 6, -20,
					-- layer=2 filter=224 channel=73
					-16, -6, -3, -17, -1, -6, -11, 9, -7,
					-- layer=2 filter=224 channel=74
					-5, -11, -5, 5, -18, 5, 9, -4, -9,
					-- layer=2 filter=224 channel=75
					-17, 3, -3, 3, 17, 4, 0, -1, 0,
					-- layer=2 filter=224 channel=76
					2, 6, -17, -3, 11, -8, -9, 0, -7,
					-- layer=2 filter=224 channel=77
					-2, -1, -10, 3, 0, 5, 0, -10, -7,
					-- layer=2 filter=224 channel=78
					-15, -4, 0, -2, 2, 5, -2, -16, -1,
					-- layer=2 filter=224 channel=79
					-6, 6, -6, -10, -6, -5, 1, -3, -3,
					-- layer=2 filter=224 channel=80
					-14, -3, -4, -7, -2, -22, -4, -4, -4,
					-- layer=2 filter=224 channel=81
					4, 5, -10, -6, -2, 0, 2, 4, -2,
					-- layer=2 filter=224 channel=82
					-4, -6, 1, -12, 1, -7, -5, 0, 0,
					-- layer=2 filter=224 channel=83
					-5, -7, 1, -11, -4, -10, -21, 0, -1,
					-- layer=2 filter=224 channel=84
					-7, -9, 0, 6, 5, -8, 8, 1, -6,
					-- layer=2 filter=224 channel=85
					-6, 1, 8, 2, 10, -3, 1, 3, 4,
					-- layer=2 filter=224 channel=86
					-4, -10, -3, -5, 0, 6, -10, -6, 6,
					-- layer=2 filter=224 channel=87
					-5, 1, 1, 2, -18, -7, -5, -7, 2,
					-- layer=2 filter=224 channel=88
					-3, -2, -2, -9, -1, -11, -20, -17, 0,
					-- layer=2 filter=224 channel=89
					-10, 16, -8, -4, -14, -7, -4, 8, -10,
					-- layer=2 filter=224 channel=90
					8, 5, 6, 0, 1, -5, 0, 4, -10,
					-- layer=2 filter=224 channel=91
					-19, -11, -1, -13, -13, -7, -14, 9, 0,
					-- layer=2 filter=224 channel=92
					-10, 5, -9, -4, -3, 2, -6, -3, -9,
					-- layer=2 filter=224 channel=93
					-11, 0, -11, -1, -3, 4, -9, 2, 13,
					-- layer=2 filter=224 channel=94
					-12, -13, -12, -15, -3, -15, -4, 0, -5,
					-- layer=2 filter=224 channel=95
					7, 6, 0, 5, -11, 5, 0, 3, -8,
					-- layer=2 filter=224 channel=96
					-5, 11, -5, 1, -8, -18, -3, -19, -1,
					-- layer=2 filter=224 channel=97
					-7, -4, -5, 0, -6, -5, 0, -18, -6,
					-- layer=2 filter=224 channel=98
					0, 0, 0, 0, -4, -6, -5, -24, 12,
					-- layer=2 filter=224 channel=99
					-4, 2, -12, -10, 7, -8, 0, 2, 0,
					-- layer=2 filter=224 channel=100
					-3, -3, -16, -3, -18, -2, -12, -8, -13,
					-- layer=2 filter=224 channel=101
					-1, -13, -8, -4, -16, -14, -5, 4, 17,
					-- layer=2 filter=224 channel=102
					-7, 13, -8, 3, -10, -24, -9, -3, -15,
					-- layer=2 filter=224 channel=103
					-2, -11, 1, -1, 0, -8, -2, -4, 7,
					-- layer=2 filter=224 channel=104
					-13, 11, 1, -6, 4, -16, -15, -16, -7,
					-- layer=2 filter=224 channel=105
					4, -1, -17, -8, 10, -11, -3, -6, -14,
					-- layer=2 filter=224 channel=106
					4, -1, 2, -4, -20, -8, 0, 0, 5,
					-- layer=2 filter=224 channel=107
					4, -8, -9, 1, -10, 6, 5, 2, -11,
					-- layer=2 filter=224 channel=108
					-4, 16, -3, -11, -14, -3, -10, 2, -9,
					-- layer=2 filter=224 channel=109
					-5, 4, -2, -3, 2, -9, -5, -11, -11,
					-- layer=2 filter=224 channel=110
					-4, 0, -3, -12, -10, 0, -19, -4, 7,
					-- layer=2 filter=224 channel=111
					9, -8, 3, -4, 7, -10, -6, 3, -6,
					-- layer=2 filter=224 channel=112
					12, -9, 9, 5, -13, 0, -5, -5, 0,
					-- layer=2 filter=224 channel=113
					-7, -5, -12, -17, -9, 0, -8, -17, -1,
					-- layer=2 filter=224 channel=114
					-3, 0, 9, 8, 0, 1, 0, -6, 9,
					-- layer=2 filter=224 channel=115
					0, 9, -8, -2, 0, 5, -10, -5, 6,
					-- layer=2 filter=224 channel=116
					-4, 0, -5, -2, -7, -15, -3, -4, -3,
					-- layer=2 filter=224 channel=117
					-9, -13, -12, -18, 3, -1, -8, -16, 5,
					-- layer=2 filter=224 channel=118
					-3, 4, -5, -18, -28, -10, 6, -8, -20,
					-- layer=2 filter=224 channel=119
					1, 2, -1, -8, 0, -2, -9, 2, -18,
					-- layer=2 filter=224 channel=120
					0, 3, 0, 3, 7, -10, 0, 3, 5,
					-- layer=2 filter=224 channel=121
					-1, 8, -9, -10, -6, -3, 0, -7, 5,
					-- layer=2 filter=224 channel=122
					5, 3, 9, -3, 0, 2, -1, -3, -4,
					-- layer=2 filter=224 channel=123
					7, 2, -3, -3, -3, 0, -20, -8, -8,
					-- layer=2 filter=224 channel=124
					3, -19, -17, -9, -12, 2, -4, -3, -5,
					-- layer=2 filter=224 channel=125
					-6, 5, -10, 6, 1, -7, 0, -9, -4,
					-- layer=2 filter=224 channel=126
					-10, 8, -4, -13, -7, -12, -12, -12, -7,
					-- layer=2 filter=224 channel=127
					0, -2, -2, 0, -14, 1, -11, -10, 1,
					-- layer=2 filter=225 channel=0
					4, 18, -30, 3, -29, -56, 10, -20, -26,
					-- layer=2 filter=225 channel=1
					11, -7, 16, 13, -13, 23, -17, -8, -29,
					-- layer=2 filter=225 channel=2
					-6, -7, -4, 1, -6, 1, -8, -3, -11,
					-- layer=2 filter=225 channel=3
					-25, -5, -4, -45, -24, 13, 38, 26, 48,
					-- layer=2 filter=225 channel=4
					-2, -8, 11, -20, -34, -21, -28, -69, -62,
					-- layer=2 filter=225 channel=5
					12, 19, 7, -8, 13, 22, -8, -19, 0,
					-- layer=2 filter=225 channel=6
					-5, 18, 52, 21, 59, 32, -17, -8, -42,
					-- layer=2 filter=225 channel=7
					-24, -24, -36, 51, 22, -4, 21, 43, 15,
					-- layer=2 filter=225 channel=8
					-11, 4, -5, 11, 13, -8, -3, 7, -9,
					-- layer=2 filter=225 channel=9
					-23, -44, -17, -23, 18, 10, -24, 22, 29,
					-- layer=2 filter=225 channel=10
					-13, -21, 8, -20, -31, -49, 23, 9, 13,
					-- layer=2 filter=225 channel=11
					-1, 4, 7, -8, -21, 0, -22, -13, -2,
					-- layer=2 filter=225 channel=12
					-3, -13, 19, 17, -31, -6, 10, 6, -24,
					-- layer=2 filter=225 channel=13
					1, 8, 9, 2, -5, -7, -9, -9, -7,
					-- layer=2 filter=225 channel=14
					-6, 3, 8, 30, -13, -6, -9, -13, -25,
					-- layer=2 filter=225 channel=15
					5, 63, -35, -46, 23, 41, -3, -13, 43,
					-- layer=2 filter=225 channel=16
					35, 28, 11, -8, 14, -10, 10, -54, -29,
					-- layer=2 filter=225 channel=17
					5, 9, -7, 4, 2, -10, 6, -7, -9,
					-- layer=2 filter=225 channel=18
					-47, 1, -23, 0, -11, -13, -6, -39, -18,
					-- layer=2 filter=225 channel=19
					9, -5, -19, 15, 41, 18, 12, 9, 4,
					-- layer=2 filter=225 channel=20
					-4, -9, -3, -3, 0, -11, -7, 1, 9,
					-- layer=2 filter=225 channel=21
					-12, 4, -13, 2, 12, 22, 12, 12, 0,
					-- layer=2 filter=225 channel=22
					-9, -7, -7, 1, 2, 9, -8, -9, 0,
					-- layer=2 filter=225 channel=23
					14, 11, 30, -11, -35, -4, 36, 26, -31,
					-- layer=2 filter=225 channel=24
					-1, -23, 30, -18, -27, 1, -22, -1, 21,
					-- layer=2 filter=225 channel=25
					11, 34, 46, -12, -12, -2, -33, -13, -10,
					-- layer=2 filter=225 channel=26
					5, -8, 8, 8, 7, -3, -5, 3, -5,
					-- layer=2 filter=225 channel=27
					6, 30, -2, -21, -17, 11, -57, -33, 6,
					-- layer=2 filter=225 channel=28
					-40, -17, -85, -12, -8, -48, 56, 44, 27,
					-- layer=2 filter=225 channel=29
					3, 0, 3, -11, 7, 2, -6, -2, -4,
					-- layer=2 filter=225 channel=30
					37, -29, 9, -42, -9, -10, -9, -4, -15,
					-- layer=2 filter=225 channel=31
					-72, -18, -23, -20, -13, -79, 31, -37, -16,
					-- layer=2 filter=225 channel=32
					7, -1, 0, 4, -5, -10, -2, 3, 3,
					-- layer=2 filter=225 channel=33
					-14, -8, -6, -39, -37, -23, -26, -4, 9,
					-- layer=2 filter=225 channel=34
					-18, -38, -35, 15, 7, 25, -19, -19, -23,
					-- layer=2 filter=225 channel=35
					-43, -37, -17, 34, -20, -17, 46, 6, 16,
					-- layer=2 filter=225 channel=36
					5, 8, -9, -3, -7, -2, 5, 8, -1,
					-- layer=2 filter=225 channel=37
					29, 5, 11, -14, 15, 17, -31, 2, 3,
					-- layer=2 filter=225 channel=38
					17, -14, -2, -17, -27, 6, -39, -49, 6,
					-- layer=2 filter=225 channel=39
					-21, -7, -3, -24, -19, -65, 15, 9, -35,
					-- layer=2 filter=225 channel=40
					17, -34, 16, 14, -14, -34, -19, -6, 39,
					-- layer=2 filter=225 channel=41
					-4, -6, -8, -2, -3, 6, 5, -2, 7,
					-- layer=2 filter=225 channel=42
					33, 24, -3, -5, -31, -11, 73, 47, 11,
					-- layer=2 filter=225 channel=43
					-29, -5, -14, -91, 53, 40, -21, -2, 80,
					-- layer=2 filter=225 channel=44
					-3, 9, 0, -9, 6, -1, 2, -5, 0,
					-- layer=2 filter=225 channel=45
					21, 37, 2, -50, -3, 0, -46, -11, 20,
					-- layer=2 filter=225 channel=46
					16, -24, -5, -3, -14, -38, 21, -18, -44,
					-- layer=2 filter=225 channel=47
					42, 52, -8, -21, -48, -67, -12, 11, -16,
					-- layer=2 filter=225 channel=48
					3, 8, -7, -2, 7, 8, -4, 0, -8,
					-- layer=2 filter=225 channel=49
					-35, 10, 11, -8, 16, 19, -35, 0, -7,
					-- layer=2 filter=225 channel=50
					-1, 10, 14, 28, 14, 5, -1, -14, -1,
					-- layer=2 filter=225 channel=51
					17, -11, 10, 3, -28, -21, -1, -24, -22,
					-- layer=2 filter=225 channel=52
					-7, -14, 7, 0, 12, 10, 1, -6, 23,
					-- layer=2 filter=225 channel=53
					-12, 11, -12, -65, 46, -16, 16, 13, -21,
					-- layer=2 filter=225 channel=54
					15, -2, 36, 23, 3, -2, 17, -10, -16,
					-- layer=2 filter=225 channel=55
					-3, 2, 2, 0, -5, 13, 1, -3, 2,
					-- layer=2 filter=225 channel=56
					-34, -2, -29, -43, -30, -25, -35, -31, -6,
					-- layer=2 filter=225 channel=57
					1, -17, -7, -8, -3, -7, 5, -3, 3,
					-- layer=2 filter=225 channel=58
					7, 3, 15, 14, -10, -6, 22, 4, -4,
					-- layer=2 filter=225 channel=59
					20, -10, -17, 26, 29, 21, -4, -38, -23,
					-- layer=2 filter=225 channel=60
					33, -20, -28, 22, 21, -7, 23, 18, -46,
					-- layer=2 filter=225 channel=61
					14, -22, -28, 42, 35, -8, 21, 30, -1,
					-- layer=2 filter=225 channel=62
					-16, -3, 6, 33, 29, 44, 1, -45, 1,
					-- layer=2 filter=225 channel=63
					9, -4, -4, 23, 22, -45, 17, 6, -31,
					-- layer=2 filter=225 channel=64
					10, 7, 30, 8, -10, -27, 18, 4, -25,
					-- layer=2 filter=225 channel=65
					14, -32, 3, 13, 12, 20, 12, 22, -2,
					-- layer=2 filter=225 channel=66
					-40, -1, 25, 12, 35, 13, 9, 4, 14,
					-- layer=2 filter=225 channel=67
					10, -22, -10, -46, -35, 10, 1, -53, 18,
					-- layer=2 filter=225 channel=68
					2, 4, -4, -9, -7, -3, -2, -1, 0,
					-- layer=2 filter=225 channel=69
					0, 22, 38, -23, 5, -1, 11, 2, -11,
					-- layer=2 filter=225 channel=70
					-28, 16, -14, 0, -10, -33, 33, 11, 1,
					-- layer=2 filter=225 channel=71
					-26, 21, -5, -27, 33, 25, -78, -14, 46,
					-- layer=2 filter=225 channel=72
					11, 8, -59, 11, 16, 6, -1, 38, 18,
					-- layer=2 filter=225 channel=73
					19, -59, -106, -5, 18, -10, 34, 54, 1,
					-- layer=2 filter=225 channel=74
					14, -12, -28, -25, -20, -45, 23, -21, -17,
					-- layer=2 filter=225 channel=75
					-62, -22, 14, -15, 3, -8, 33, 11, -27,
					-- layer=2 filter=225 channel=76
					-13, -24, -45, -9, -9, -21, -37, -20, 46,
					-- layer=2 filter=225 channel=77
					10, 5, 5, 6, 9, -1, -10, 0, -13,
					-- layer=2 filter=225 channel=78
					-6, -19, 7, -2, -9, -12, 1, 1, -1,
					-- layer=2 filter=225 channel=79
					1, 2, -2, -5, -3, 9, 0, 7, 6,
					-- layer=2 filter=225 channel=80
					34, -12, -7, -17, -11, -31, -4, 13, -12,
					-- layer=2 filter=225 channel=81
					2, 15, 13, -4, -1, 1, -3, -4, 0,
					-- layer=2 filter=225 channel=82
					9, -7, -5, -4, -6, 7, 9, -4, -10,
					-- layer=2 filter=225 channel=83
					-3, 27, 23, -26, -4, -19, -10, 41, -37,
					-- layer=2 filter=225 channel=84
					0, 8, 3, 5, 2, -3, 2, 4, -8,
					-- layer=2 filter=225 channel=85
					-2, 3, 5, -7, 2, 0, -5, 2, -12,
					-- layer=2 filter=225 channel=86
					-14, 7, 5, 0, 8, 28, 20, -15, 11,
					-- layer=2 filter=225 channel=87
					-5, 11, -38, -21, -13, 17, -63, -74, 1,
					-- layer=2 filter=225 channel=88
					22, -9, -5, -36, 3, -24, -10, -1, 4,
					-- layer=2 filter=225 channel=89
					-13, -19, -20, 25, -7, 2, -12, -25, 8,
					-- layer=2 filter=225 channel=90
					4, 6, 8, 8, -3, 7, -6, 8, 9,
					-- layer=2 filter=225 channel=91
					0, 13, -12, 11, -20, 0, -9, -1, 11,
					-- layer=2 filter=225 channel=92
					12, 4, 3, 27, -27, 17, -34, -7, -23,
					-- layer=2 filter=225 channel=93
					-58, 12, 0, -4, -8, 25, -3, 18, 10,
					-- layer=2 filter=225 channel=94
					29, 2, 16, 41, 39, 61, 0, 24, -37,
					-- layer=2 filter=225 channel=95
					0, 8, 3, 8, 8, 2, -7, 7, 4,
					-- layer=2 filter=225 channel=96
					11, 15, 14, 33, 23, 28, -5, -5, -40,
					-- layer=2 filter=225 channel=97
					15, -28, 6, -27, -47, -21, 3, -43, -16,
					-- layer=2 filter=225 channel=98
					-16, -19, -72, 16, -23, -44, 32, 22, -4,
					-- layer=2 filter=225 channel=99
					0, -19, -13, 26, 46, 3, -4, 2, 24,
					-- layer=2 filter=225 channel=100
					13, -16, -32, -31, -38, 2, 57, -9, 35,
					-- layer=2 filter=225 channel=101
					-29, 6, 20, -8, -16, 27, -9, 14, 55,
					-- layer=2 filter=225 channel=102
					5, 17, 0, 0, 30, 26, -3, -20, -64,
					-- layer=2 filter=225 channel=103
					0, -27, 5, 32, -1, -51, 55, 53, -2,
					-- layer=2 filter=225 channel=104
					-26, 32, 3, -32, 31, 32, -39, -15, -23,
					-- layer=2 filter=225 channel=105
					-37, -60, -23, 6, 19, -13, 28, -45, 16,
					-- layer=2 filter=225 channel=106
					-23, 0, 17, -29, -37, -26, 3, -11, -37,
					-- layer=2 filter=225 channel=107
					-21, 4, -5, 0, -3, 40, 45, 19, 16,
					-- layer=2 filter=225 channel=108
					0, 0, 10, -15, 26, 6, -64, -5, -37,
					-- layer=2 filter=225 channel=109
					11, -7, -5, 4, 11, 12, -3, -3, 4,
					-- layer=2 filter=225 channel=110
					14, 1, 10, 5, 18, -10, 17, 29, -17,
					-- layer=2 filter=225 channel=111
					-11, -9, 3, -3, 1, -3, 5, -5, -2,
					-- layer=2 filter=225 channel=112
					26, -26, -37, 14, -32, -48, 9, -35, -13,
					-- layer=2 filter=225 channel=113
					24, 16, -9, -8, 9, -27, 23, 8, -28,
					-- layer=2 filter=225 channel=114
					6, -9, 2, 1, 2, -6, 4, 10, -2,
					-- layer=2 filter=225 channel=115
					-3, -2, 9, 8, -3, -4, -8, -3, -8,
					-- layer=2 filter=225 channel=116
					-6, 16, -32, -39, 10, 39, -26, -29, -19,
					-- layer=2 filter=225 channel=117
					-41, -54, -53, 22, 2, -23, 59, 20, 4,
					-- layer=2 filter=225 channel=118
					20, -20, -13, -71, 18, -2, -12, 3, 17,
					-- layer=2 filter=225 channel=119
					0, 35, 1, 9, -70, 18, 19, -47, -16,
					-- layer=2 filter=225 channel=120
					8, 0, -5, 0, -8, 6, 8, -7, -10,
					-- layer=2 filter=225 channel=121
					-6, 6, 10, 6, -8, -5, -1, -1, 12,
					-- layer=2 filter=225 channel=122
					0, -11, 7, 14, 6, 2, 5, -9, -1,
					-- layer=2 filter=225 channel=123
					8, -18, -71, 4, 26, -39, 17, 17, -9,
					-- layer=2 filter=225 channel=124
					-67, 14, -9, -8, -11, 15, 12, -18, 49,
					-- layer=2 filter=225 channel=125
					-2, -8, -7, 4, -7, 0, -1, 1, 2,
					-- layer=2 filter=225 channel=126
					83, -25, -3, 9, -16, 34, 13, 12, 21,
					-- layer=2 filter=225 channel=127
					15, 0, 13, -35, -12, 41, 7, 20, -26,
					-- layer=2 filter=226 channel=0
					0, -1, 0, 0, -6, 1, 16, 5, 22,
					-- layer=2 filter=226 channel=1
					-6, -26, 14, -10, -6, -34, -7, -18, -5,
					-- layer=2 filter=226 channel=2
					-2, 0, 8, -5, 6, -2, -6, -6, 3,
					-- layer=2 filter=226 channel=3
					22, -3, -1, -24, -27, 12, -5, 28, 0,
					-- layer=2 filter=226 channel=4
					18, 12, 14, -11, 14, -2, 10, 8, -17,
					-- layer=2 filter=226 channel=5
					4, 6, -5, -34, -11, -24, 0, -17, -34,
					-- layer=2 filter=226 channel=6
					19, 1, 13, 35, 24, 55, -25, 22, 25,
					-- layer=2 filter=226 channel=7
					42, 8, -14, 46, 29, 12, -10, 28, 1,
					-- layer=2 filter=226 channel=8
					-3, 9, 10, -3, 1, -5, -5, 6, -2,
					-- layer=2 filter=226 channel=9
					18, -27, 38, -46, -34, -22, 5, -5, -15,
					-- layer=2 filter=226 channel=10
					22, 13, 22, 5, 4, 25, -13, 12, 29,
					-- layer=2 filter=226 channel=11
					20, 16, -12, -32, -20, -41, -22, -7, -23,
					-- layer=2 filter=226 channel=12
					-4, 16, 43, 30, 5, -21, 2, -6, 5,
					-- layer=2 filter=226 channel=13
					5, 8, 0, 10, 8, -6, 4, -8, 12,
					-- layer=2 filter=226 channel=14
					-3, -4, 22, 19, -6, -35, 39, -10, -8,
					-- layer=2 filter=226 channel=15
					5, -6, -10, -26, -29, -31, -14, -40, -98,
					-- layer=2 filter=226 channel=16
					7, -31, -45, -20, -3, 21, -22, -14, -27,
					-- layer=2 filter=226 channel=17
					-9, 4, 1, 1, -3, -5, 6, -8, 5,
					-- layer=2 filter=226 channel=18
					-37, 18, 4, -74, 4, 4, -29, -32, -21,
					-- layer=2 filter=226 channel=19
					37, -19, -6, -13, -14, 15, -10, -36, 19,
					-- layer=2 filter=226 channel=20
					-3, 4, -4, -4, 5, -5, 5, 6, -4,
					-- layer=2 filter=226 channel=21
					3, 27, 22, 9, 9, 23, 10, 12, 1,
					-- layer=2 filter=226 channel=22
					-10, -8, -1, -2, -8, -3, -3, -6, -5,
					-- layer=2 filter=226 channel=23
					14, 24, -10, 16, 23, 2, 35, 2, 30,
					-- layer=2 filter=226 channel=24
					-19, 2, 0, 8, 8, 35, 32, 29, 30,
					-- layer=2 filter=226 channel=25
					-7, 0, 0, -13, -5, 7, 19, 33, 16,
					-- layer=2 filter=226 channel=26
					6, -3, 8, 0, 9, 0, -4, -1, -4,
					-- layer=2 filter=226 channel=27
					-21, -8, -13, -50, -40, -42, -9, -31, -54,
					-- layer=2 filter=226 channel=28
					23, 40, 43, 38, 23, 43, -5, 0, -11,
					-- layer=2 filter=226 channel=29
					-6, 6, 1, 0, -7, 0, 12, 5, 3,
					-- layer=2 filter=226 channel=30
					-20, 4, -15, 7, 6, -28, -8, -4, -32,
					-- layer=2 filter=226 channel=31
					-4, 33, 33, 27, 38, -20, 63, -11, -24,
					-- layer=2 filter=226 channel=32
					0, -6, 10, 7, 1, -3, -5, 0, 12,
					-- layer=2 filter=226 channel=33
					-3, -22, 1, 27, 15, -25, 3, 17, -31,
					-- layer=2 filter=226 channel=34
					-3, 51, -18, -4, 32, 6, -6, -6, 42,
					-- layer=2 filter=226 channel=35
					22, 17, 23, 11, 38, 19, -5, 11, -6,
					-- layer=2 filter=226 channel=36
					8, 14, 8, -3, -2, 1, -5, -12, -4,
					-- layer=2 filter=226 channel=37
					-2, -1, -30, -32, -35, -19, -23, 5, -20,
					-- layer=2 filter=226 channel=38
					-9, -5, -20, -34, -37, 5, -8, 0, -18,
					-- layer=2 filter=226 channel=39
					31, 6, -31, 6, 2, -7, -11, -15, 21,
					-- layer=2 filter=226 channel=40
					-11, -2, -56, -32, -57, -6, 0, -56, -90,
					-- layer=2 filter=226 channel=41
					8, 2, 6, -2, 11, 5, 6, 1, 5,
					-- layer=2 filter=226 channel=42
					20, -9, 12, -2, -24, -9, 20, 5, -5,
					-- layer=2 filter=226 channel=43
					-13, -15, -33, -29, -23, -7, -56, 13, -27,
					-- layer=2 filter=226 channel=44
					7, 5, -5, 2, 10, 7, -12, -3, 0,
					-- layer=2 filter=226 channel=45
					5, -24, -78, 48, 24, -12, 14, 48, -10,
					-- layer=2 filter=226 channel=46
					-12, -3, 10, -15, -6, 1, 7, -20, 7,
					-- layer=2 filter=226 channel=47
					-2, -37, -10, 26, 1, -3, -3, 4, 15,
					-- layer=2 filter=226 channel=48
					8, -4, 6, 6, -1, -2, 9, -3, -4,
					-- layer=2 filter=226 channel=49
					6, 16, 33, -71, -37, -17, 3, -37, 17,
					-- layer=2 filter=226 channel=50
					16, 4, 1, 15, -2, 0, -2, 15, 11,
					-- layer=2 filter=226 channel=51
					9, 18, 4, -1, -19, -15, -2, 11, -26,
					-- layer=2 filter=226 channel=52
					-14, -66, -62, -8, -20, -11, -13, -7, 2,
					-- layer=2 filter=226 channel=53
					5, 4, 21, -50, -1, -29, -78, -79, 19,
					-- layer=2 filter=226 channel=54
					54, 12, 8, 20, 30, -10, 7, 39, 25,
					-- layer=2 filter=226 channel=55
					-7, 0, 5, 10, -2, 3, 15, -7, 13,
					-- layer=2 filter=226 channel=56
					0, 0, -15, -37, -26, -55, -25, -36, -45,
					-- layer=2 filter=226 channel=57
					11, 1, -2, -4, 1, 10, -5, 9, 0,
					-- layer=2 filter=226 channel=58
					14, 26, 5, 28, -17, -6, -5, 0, 17,
					-- layer=2 filter=226 channel=59
					1, -17, -30, -18, -8, -16, -33, 26, -21,
					-- layer=2 filter=226 channel=60
					1, -3, 12, -40, -17, 51, -58, 16, 14,
					-- layer=2 filter=226 channel=61
					-30, -15, 4, -25, 4, 0, -35, 4, -19,
					-- layer=2 filter=226 channel=62
					18, 10, 22, 7, 36, 24, -9, -52, 43,
					-- layer=2 filter=226 channel=63
					8, 0, -23, 32, 3, 16, 2, 6, 17,
					-- layer=2 filter=226 channel=64
					-16, -1, -20, -11, 6, -1, 27, 23, 27,
					-- layer=2 filter=226 channel=65
					-15, 40, 24, 4, -22, 17, -3, 7, -11,
					-- layer=2 filter=226 channel=66
					-5, 24, 39, 18, 0, -27, -36, 44, -25,
					-- layer=2 filter=226 channel=67
					-13, -7, -6, -36, -42, -34, -12, -9, -42,
					-- layer=2 filter=226 channel=68
					-4, 10, 9, -6, -4, -9, 1, 0, -3,
					-- layer=2 filter=226 channel=69
					0, -9, -14, 11, 2, -5, 6, -11, 17,
					-- layer=2 filter=226 channel=70
					8, 17, 34, 27, 20, 21, 21, 15, -15,
					-- layer=2 filter=226 channel=71
					0, -30, -63, -29, -6, -80, -105, -94, -84,
					-- layer=2 filter=226 channel=72
					34, 16, 22, 18, 0, 13, 7, 8, -23,
					-- layer=2 filter=226 channel=73
					47, -24, -43, 89, 22, -2, 64, 14, -21,
					-- layer=2 filter=226 channel=74
					4, -3, -7, -1, -33, 9, 11, 7, 14,
					-- layer=2 filter=226 channel=75
					-28, -69, -16, -33, -15, -20, 6, 21, 40,
					-- layer=2 filter=226 channel=76
					-11, -38, -52, -20, 3, 31, 7, -59, 30,
					-- layer=2 filter=226 channel=77
					-3, -1, -10, 2, 5, 8, -3, 5, 5,
					-- layer=2 filter=226 channel=78
					28, 24, -17, -12, 3, -14, 19, 16, 4,
					-- layer=2 filter=226 channel=79
					11, 5, 5, 8, 4, 9, 11, -2, -1,
					-- layer=2 filter=226 channel=80
					13, -18, 14, 0, -20, 22, -6, 7, -3,
					-- layer=2 filter=226 channel=81
					2, -9, 2, 2, 9, -14, 6, -14, -5,
					-- layer=2 filter=226 channel=82
					-1, 11, 8, -2, 2, 0, -3, -3, -4,
					-- layer=2 filter=226 channel=83
					2, 9, 17, 27, 14, 16, 16, 14, -28,
					-- layer=2 filter=226 channel=84
					2, -2, -4, -11, -4, 0, 4, 1, 9,
					-- layer=2 filter=226 channel=85
					-2, 14, -7, -8, 0, 0, 1, 5, 1,
					-- layer=2 filter=226 channel=86
					10, -3, -11, 1, 5, -9, 12, -10, 4,
					-- layer=2 filter=226 channel=87
					8, -5, 3, -32, 14, 34, -8, 14, 19,
					-- layer=2 filter=226 channel=88
					14, 19, -10, 13, 8, -36, 9, -5, -19,
					-- layer=2 filter=226 channel=89
					0, -14, 8, -17, -5, -36, 11, -16, -28,
					-- layer=2 filter=226 channel=90
					9, 8, 0, 0, 1, -1, 4, -7, 4,
					-- layer=2 filter=226 channel=91
					-4, 0, 20, 10, -22, -3, -19, -19, 9,
					-- layer=2 filter=226 channel=92
					7, 5, 16, 22, 1, -24, -4, -10, -24,
					-- layer=2 filter=226 channel=93
					15, 27, -4, 15, 21, -3, 20, -8, 0,
					-- layer=2 filter=226 channel=94
					-13, 4, 5, -16, 27, 20, -113, -1, -8,
					-- layer=2 filter=226 channel=95
					-3, 11, -4, -1, 9, 0, -6, 1, 5,
					-- layer=2 filter=226 channel=96
					42, 17, 19, 15, -14, -31, 69, 11, 40,
					-- layer=2 filter=226 channel=97
					10, -32, 2, -12, -32, 12, 13, 1, 0,
					-- layer=2 filter=226 channel=98
					1, -15, 25, 34, 20, 27, 29, 9, 25,
					-- layer=2 filter=226 channel=99
					-18, -69, -68, -13, -5, -13, -17, -1, 29,
					-- layer=2 filter=226 channel=100
					20, -7, -5, -15, 5, 25, -7, -11, -30,
					-- layer=2 filter=226 channel=101
					12, -46, -54, -76, -65, -45, -72, -112, -92,
					-- layer=2 filter=226 channel=102
					24, 21, 22, -54, -32, -35, -15, -25, 36,
					-- layer=2 filter=226 channel=103
					10, -5, 12, 39, -25, -8, 9, 9, 2,
					-- layer=2 filter=226 channel=104
					0, 39, 27, -48, -11, -3, -66, -59, -8,
					-- layer=2 filter=226 channel=105
					12, -77, -7, -15, 25, 8, -5, -20, -25,
					-- layer=2 filter=226 channel=106
					16, 40, 14, -35, -39, -14, -35, -24, 5,
					-- layer=2 filter=226 channel=107
					11, 19, 19, 58, -9, 1, 3, 23, 19,
					-- layer=2 filter=226 channel=108
					2, -11, 12, -37, -53, -97, -5, -37, -4,
					-- layer=2 filter=226 channel=109
					-2, 7, -4, 7, 10, 2, 1, -5, 4,
					-- layer=2 filter=226 channel=110
					5, 0, 2, -28, 11, 5, 2, 8, -2,
					-- layer=2 filter=226 channel=111
					0, 7, 11, -1, -9, -2, -8, -8, 6,
					-- layer=2 filter=226 channel=112
					-52, -18, 40, -19, -24, -6, -23, -27, -3,
					-- layer=2 filter=226 channel=113
					-21, 40, -4, 17, -8, -2, -4, 13, 0,
					-- layer=2 filter=226 channel=114
					18, 3, 12, 0, 10, 11, -2, -3, 17,
					-- layer=2 filter=226 channel=115
					9, 3, 3, 3, -10, 7, -8, -1, -8,
					-- layer=2 filter=226 channel=116
					3, 10, -12, -36, 13, 27, -46, -31, 4,
					-- layer=2 filter=226 channel=117
					1, -27, -37, 4, -61, -82, -14, -7, -27,
					-- layer=2 filter=226 channel=118
					31, -3, 2, 5, -10, 35, -6, 16, 33,
					-- layer=2 filter=226 channel=119
					-14, 14, 10, -4, -4, -26, 6, 7, -7,
					-- layer=2 filter=226 channel=120
					0, -1, 7, -1, -5, -4, 4, 2, -1,
					-- layer=2 filter=226 channel=121
					9, 12, -9, 11, -5, -8, -5, -4, -3,
					-- layer=2 filter=226 channel=122
					1, 4, -2, -7, 7, -8, 10, 2, 5,
					-- layer=2 filter=226 channel=123
					9, -22, -15, 21, 25, 18, -2, 13, 32,
					-- layer=2 filter=226 channel=124
					-33, -51, -15, -2, 13, -25, 33, -13, -25,
					-- layer=2 filter=226 channel=125
					-9, 8, -3, 1, 4, 3, 6, 1, 10,
					-- layer=2 filter=226 channel=126
					-61, -15, 3, -14, -52, -27, -63, -2, -19,
					-- layer=2 filter=226 channel=127
					-24, -11, 12, 40, -10, -1, 5, 11, -18,
					-- layer=2 filter=227 channel=0
					-32, 3, 6, -26, 5, 19, 1, 11, 16,
					-- layer=2 filter=227 channel=1
					-8, 11, -4, -10, -71, -18, 25, -21, -34,
					-- layer=2 filter=227 channel=2
					1, 7, -6, 4, 6, -12, -2, 6, 0,
					-- layer=2 filter=227 channel=3
					-28, 2, 39, -22, 5, 81, -36, 12, 76,
					-- layer=2 filter=227 channel=4
					-73, -10, -33, -27, -21, -1, -57, 0, 2,
					-- layer=2 filter=227 channel=5
					-7, 1, -5, -11, 7, -15, -5, 10, 39,
					-- layer=2 filter=227 channel=6
					31, -18, -22, 48, -52, -24, 18, -52, -74,
					-- layer=2 filter=227 channel=7
					-54, 1, 18, 30, 27, 18, 7, -35, -7,
					-- layer=2 filter=227 channel=8
					-2, 4, -5, 1, -10, 0, 3, 7, -9,
					-- layer=2 filter=227 channel=9
					-53, -7, 15, -26, -45, 45, 3, 1, 66,
					-- layer=2 filter=227 channel=10
					-19, -14, 26, -7, -4, 50, 0, 16, 45,
					-- layer=2 filter=227 channel=11
					-8, 8, 11, -16, 9, 7, 19, 3, -24,
					-- layer=2 filter=227 channel=12
					-22, -13, -15, -7, -26, -53, 67, -22, 8,
					-- layer=2 filter=227 channel=13
					8, -1, -8, -1, -6, 9, 3, -7, 7,
					-- layer=2 filter=227 channel=14
					-10, -3, 16, -16, -38, -46, 11, -13, -33,
					-- layer=2 filter=227 channel=15
					-74, -13, -61, 12, 27, 18, 35, -4, -57,
					-- layer=2 filter=227 channel=16
					-21, 1, 18, -20, 41, 31, -44, 9, 31,
					-- layer=2 filter=227 channel=17
					0, -8, 5, -6, -9, 9, -1, -11, 2,
					-- layer=2 filter=227 channel=18
					-34, -31, -32, -18, 7, -20, 11, 27, -94,
					-- layer=2 filter=227 channel=19
					3, 21, 40, 1, -37, -29, 25, 2, -39,
					-- layer=2 filter=227 channel=20
					-2, -3, 1, -11, 10, -5, 0, -3, 4,
					-- layer=2 filter=227 channel=21
					-2, 8, -15, -15, -8, -3, -16, 12, -7,
					-- layer=2 filter=227 channel=22
					-8, 5, 1, 3, -11, -4, 6, 3, 9,
					-- layer=2 filter=227 channel=23
					14, 14, -23, 0, -23, 8, -30, -30, 8,
					-- layer=2 filter=227 channel=24
					-40, -23, -14, -32, 0, 25, -5, 4, 25,
					-- layer=2 filter=227 channel=25
					-31, -21, -16, -13, 27, 37, -20, -14, 8,
					-- layer=2 filter=227 channel=26
					4, -2, -3, 7, -5, 4, -7, 6, 8,
					-- layer=2 filter=227 channel=27
					1, 18, 26, -16, -1, 0, -4, 4, -11,
					-- layer=2 filter=227 channel=28
					-37, -65, 28, 16, 22, 29, -59, -7, 10,
					-- layer=2 filter=227 channel=29
					-11, 3, -2, 7, 5, 0, 0, -4, -11,
					-- layer=2 filter=227 channel=30
					10, -29, -22, -50, -45, -5, -9, 7, 26,
					-- layer=2 filter=227 channel=31
					-23, 60, 12, 1, 31, 24, 40, 46, 48,
					-- layer=2 filter=227 channel=32
					-7, 3, 9, 8, 9, -12, 2, -1, 0,
					-- layer=2 filter=227 channel=33
					13, -28, -6, -35, 18, 35, 21, -30, 28,
					-- layer=2 filter=227 channel=34
					55, 5, -5, 29, 42, -5, -22, 52, -56,
					-- layer=2 filter=227 channel=35
					-49, 2, 16, 21, 46, 46, -44, 9, -9,
					-- layer=2 filter=227 channel=36
					-9, -4, -16, -9, -16, 2, -6, -5, 6,
					-- layer=2 filter=227 channel=37
					10, 0, -5, 7, -2, -12, 4, 8, -14,
					-- layer=2 filter=227 channel=38
					12, 0, -18, 18, -41, -29, 5, 7, -14,
					-- layer=2 filter=227 channel=39
					-27, -12, 21, -45, 10, 7, 7, -30, 4,
					-- layer=2 filter=227 channel=40
					-16, -13, -27, -52, 27, 20, 12, 40, -62,
					-- layer=2 filter=227 channel=41
					4, -9, -3, 1, 9, -2, -10, -5, 5,
					-- layer=2 filter=227 channel=42
					-32, 12, -2, -41, 28, 14, -12, -31, 14,
					-- layer=2 filter=227 channel=43
					-65, -10, 23, -69, 28, 54, -70, -4, 47,
					-- layer=2 filter=227 channel=44
					5, 4, -5, -9, -2, 1, -8, -6, -7,
					-- layer=2 filter=227 channel=45
					3, 44, -12, -15, 23, -7, 12, 0, 0,
					-- layer=2 filter=227 channel=46
					-4, -18, -3, -68, 16, 30, -38, 9, 23,
					-- layer=2 filter=227 channel=47
					-23, -106, -52, 3, -1, 8, -29, -3, -18,
					-- layer=2 filter=227 channel=48
					0, -4, 1, 7, -1, 1, -5, 0, 5,
					-- layer=2 filter=227 channel=49
					-46, -38, -21, -51, -28, -16, 27, -24, -42,
					-- layer=2 filter=227 channel=50
					-4, -23, -10, -2, -18, -28, -7, -16, 7,
					-- layer=2 filter=227 channel=51
					-8, 7, -2, -3, 15, 0, -11, 9, -4,
					-- layer=2 filter=227 channel=52
					-25, 13, -15, -5, 7, -34, -8, 5, -53,
					-- layer=2 filter=227 channel=53
					12, 26, -19, 8, -6, -76, -12, 30, -4,
					-- layer=2 filter=227 channel=54
					15, 11, -8, 41, 28, -5, -9, 16, -43,
					-- layer=2 filter=227 channel=55
					10, -2, 2, 13, -9, 7, -7, 4, 10,
					-- layer=2 filter=227 channel=56
					-17, 6, 2, -32, 1, 6, -4, 2, -6,
					-- layer=2 filter=227 channel=57
					10, 0, -6, -1, -4, 0, 8, 8, -7,
					-- layer=2 filter=227 channel=58
					-8, 10, 2, -16, -22, -25, 53, -1, -5,
					-- layer=2 filter=227 channel=59
					32, 25, -2, 22, -1, -3, 48, -44, -56,
					-- layer=2 filter=227 channel=60
					31, -41, -63, 53, -33, -52, -7, -30, -46,
					-- layer=2 filter=227 channel=61
					5, -47, -35, 50, -38, -40, 31, -37, -46,
					-- layer=2 filter=227 channel=62
					15, -18, -21, 4, 11, -10, 34, 17, -104,
					-- layer=2 filter=227 channel=63
					-8, 6, 4, -22, -25, -21, -15, -20, 9,
					-- layer=2 filter=227 channel=64
					-9, 3, 2, 0, 3, 20, -16, -26, -4,
					-- layer=2 filter=227 channel=65
					0, -48, -76, 62, -69, -16, 18, -62, -29,
					-- layer=2 filter=227 channel=66
					-38, 15, 8, 10, 47, 22, 13, -18, 39,
					-- layer=2 filter=227 channel=67
					-4, -19, -4, -60, -27, 31, -19, 8, 66,
					-- layer=2 filter=227 channel=68
					5, -11, 3, 5, -1, -1, -9, 5, -11,
					-- layer=2 filter=227 channel=69
					-5, 20, 14, -37, -5, 14, -9, -17, 0,
					-- layer=2 filter=227 channel=70
					-73, -28, 0, 7, 25, 11, 2, 9, 6,
					-- layer=2 filter=227 channel=71
					13, 50, 20, -1, 17, 0, -12, -18, -4,
					-- layer=2 filter=227 channel=72
					-15, -17, 18, 29, 21, 22, -54, -45, -50,
					-- layer=2 filter=227 channel=73
					16, -8, 0, 14, -7, -11, -6, 2, 12,
					-- layer=2 filter=227 channel=74
					-21, -24, 22, -60, 18, 8, 21, 15, 45,
					-- layer=2 filter=227 channel=75
					-30, -23, 29, -41, -85, -63, 50, -26, 7,
					-- layer=2 filter=227 channel=76
					1, 36, -14, 34, 30, -23, 37, 87, -42,
					-- layer=2 filter=227 channel=77
					-6, 0, -10, 3, -12, -9, 5, 6, -4,
					-- layer=2 filter=227 channel=78
					-10, -27, -33, -1, 11, -5, 12, 0, -19,
					-- layer=2 filter=227 channel=79
					-6, 6, 7, 6, 3, -10, 8, -8, 2,
					-- layer=2 filter=227 channel=80
					-42, -6, 18, -22, -10, 11, -34, -7, 17,
					-- layer=2 filter=227 channel=81
					-1, 4, -1, -3, -13, -6, 5, 0, -7,
					-- layer=2 filter=227 channel=82
					1, -4, 3, 0, -11, -3, 9, -3, 7,
					-- layer=2 filter=227 channel=83
					11, -4, -12, -22, -21, -31, -1, -21, 32,
					-- layer=2 filter=227 channel=84
					-1, -10, 0, 0, 1, 4, -7, 8, -1,
					-- layer=2 filter=227 channel=85
					-3, 11, 0, -11, -4, 7, -11, -9, 4,
					-- layer=2 filter=227 channel=86
					3, 9, 1, 10, -15, 6, 1, 8, -15,
					-- layer=2 filter=227 channel=87
					-39, 28, -4, 18, 27, 12, 56, 59, -133,
					-- layer=2 filter=227 channel=88
					1, -3, -15, -29, -20, 4, 31, 17, 22,
					-- layer=2 filter=227 channel=89
					-13, 11, 10, 0, -1, -11, 59, -56, -23,
					-- layer=2 filter=227 channel=90
					-2, 0, 6, -1, 4, 1, -6, 5, 1,
					-- layer=2 filter=227 channel=91
					-17, -38, -2, 0, -22, -12, 1, -18, 17,
					-- layer=2 filter=227 channel=92
					-28, -16, 0, 12, -29, -14, 29, -14, -32,
					-- layer=2 filter=227 channel=93
					17, -14, -63, 18, -95, -17, -57, -16, -58,
					-- layer=2 filter=227 channel=94
					14, 8, 31, 19, -24, -73, 19, -31, -46,
					-- layer=2 filter=227 channel=95
					0, -12, -20, -7, 4, -24, -23, 0, -3,
					-- layer=2 filter=227 channel=96
					14, 62, -60, 26, 23, -55, 22, 32, -55,
					-- layer=2 filter=227 channel=97
					-69, -8, -9, -109, 0, 74, -11, 1, 36,
					-- layer=2 filter=227 channel=98
					-25, -49, -6, 13, 11, 25, -47, -20, -43,
					-- layer=2 filter=227 channel=99
					-22, 15, 1, -9, -26, 12, 24, -16, -77,
					-- layer=2 filter=227 channel=100
					-3, -25, -24, -26, -19, -27, 0, -12, 26,
					-- layer=2 filter=227 channel=101
					-40, 15, 21, -57, 49, 45, -42, -28, 26,
					-- layer=2 filter=227 channel=102
					16, 45, -22, 2, 24, -17, -5, 26, -59,
					-- layer=2 filter=227 channel=103
					-35, -30, 7, 46, -31, -8, 0, 32, -13,
					-- layer=2 filter=227 channel=104
					-28, 12, -40, -11, 0, -104, 10, -7, -108,
					-- layer=2 filter=227 channel=105
					8, 48, 37, 2, 19, -7, 72, 53, 32,
					-- layer=2 filter=227 channel=106
					-38, -11, -9, 0, -15, 33, -17, -4, 26,
					-- layer=2 filter=227 channel=107
					16, -50, -23, -4, -6, 76, -43, -31, 27,
					-- layer=2 filter=227 channel=108
					1, 13, -19, -16, -33, -51, 0, -27, -45,
					-- layer=2 filter=227 channel=109
					7, 0, -4, 15, -3, 2, -19, 8, 2,
					-- layer=2 filter=227 channel=110
					4, 8, 15, 15, 12, 23, -30, 4, -7,
					-- layer=2 filter=227 channel=111
					-8, 2, 3, 10, -5, 8, 1, 4, -7,
					-- layer=2 filter=227 channel=112
					-9, -59, -47, 4, -43, 21, 6, 22, 19,
					-- layer=2 filter=227 channel=113
					-22, -24, -22, -17, -34, 2, -17, 0, -3,
					-- layer=2 filter=227 channel=114
					16, 11, -2, -3, -3, -5, -3, -7, 8,
					-- layer=2 filter=227 channel=115
					3, -7, -9, -8, 4, -8, 6, -4, 6,
					-- layer=2 filter=227 channel=116
					-40, 22, -23, 30, 36, -26, 19, 88, -82,
					-- layer=2 filter=227 channel=117
					-4, 7, 30, 29, 7, 12, -36, -49, -32,
					-- layer=2 filter=227 channel=118
					-48, -18, -11, -31, -5, 42, -25, 32, 47,
					-- layer=2 filter=227 channel=119
					-43, -18, -11, -40, 23, 4, -24, 20, -12,
					-- layer=2 filter=227 channel=120
					6, -5, -3, -6, -8, 10, 5, -3, -4,
					-- layer=2 filter=227 channel=121
					1, 5, 4, -7, 7, -11, 7, -8, -2,
					-- layer=2 filter=227 channel=122
					9, 8, -7, -1, -17, 7, 10, 11, -9,
					-- layer=2 filter=227 channel=123
					-6, -13, -12, 8, 21, 9, -12, -32, -22,
					-- layer=2 filter=227 channel=124
					-21, 8, -21, 21, 1, 15, 55, -20, -17,
					-- layer=2 filter=227 channel=125
					-7, -9, 2, 7, -10, 10, 1, 3, -2,
					-- layer=2 filter=227 channel=126
					-9, 0, 24, 0, -9, -4, -11, 6, -31,
					-- layer=2 filter=227 channel=127
					-4, 2, -26, 28, 5, -15, 30, -22, -7,
					-- layer=2 filter=228 channel=0
					2, 4, 0, 2, 0, -8, -11, 4, -1,
					-- layer=2 filter=228 channel=1
					3, -9, 1, -13, -14, -21, -20, -2, 10,
					-- layer=2 filter=228 channel=2
					-1, -8, -10, -2, -7, -10, 6, -10, 8,
					-- layer=2 filter=228 channel=3
					-17, -12, -14, -6, -7, -14, -9, -7, -9,
					-- layer=2 filter=228 channel=4
					6, -7, -2, -2, -5, 0, -11, -2, 0,
					-- layer=2 filter=228 channel=5
					-8, -12, -15, 4, -10, -7, 4, 2, 1,
					-- layer=2 filter=228 channel=6
					0, -1, 0, -21, 1, -2, -12, -14, -10,
					-- layer=2 filter=228 channel=7
					7, 1, -3, -2, 12, 6, -6, -2, -3,
					-- layer=2 filter=228 channel=8
					1, 2, -4, -9, -8, -9, 0, -6, 9,
					-- layer=2 filter=228 channel=9
					-11, -2, -5, -5, -7, 0, -2, 0, -12,
					-- layer=2 filter=228 channel=10
					-11, -6, -18, -18, -9, -9, -2, -12, -7,
					-- layer=2 filter=228 channel=11
					-4, 7, -11, -8, -7, -10, -15, -8, -2,
					-- layer=2 filter=228 channel=12
					7, -4, 5, -11, -8, 1, -11, -10, -3,
					-- layer=2 filter=228 channel=13
					4, -10, 6, -7, -4, -5, -4, -1, 3,
					-- layer=2 filter=228 channel=14
					-7, -1, -6, -6, -17, -14, 0, -8, 0,
					-- layer=2 filter=228 channel=15
					7, -11, -11, -4, -8, -8, 7, 6, -2,
					-- layer=2 filter=228 channel=16
					-10, -7, 1, -13, -7, 0, -12, 0, 2,
					-- layer=2 filter=228 channel=17
					1, 6, -6, -4, -9, -1, 1, 4, -7,
					-- layer=2 filter=228 channel=18
					-14, -8, -3, 0, 0, 0, -5, -4, -11,
					-- layer=2 filter=228 channel=19
					0, 11, 11, -4, -7, 9, 3, -2, -2,
					-- layer=2 filter=228 channel=20
					-11, -5, -4, -7, 3, -9, 0, -5, -11,
					-- layer=2 filter=228 channel=21
					10, 1, 8, 2, -8, -6, 1, 4, -7,
					-- layer=2 filter=228 channel=22
					-6, 0, 8, 1, 8, -5, 10, -10, 8,
					-- layer=2 filter=228 channel=23
					-9, 0, -18, -5, -15, -14, 2, -7, -2,
					-- layer=2 filter=228 channel=24
					-6, -9, -14, -5, -1, -13, -15, -6, -10,
					-- layer=2 filter=228 channel=25
					13, 13, 5, -17, -6, -12, -19, -20, -18,
					-- layer=2 filter=228 channel=26
					0, 8, 2, 2, 9, 6, 8, 5, -4,
					-- layer=2 filter=228 channel=27
					-5, -1, 14, -3, 0, 15, -12, 4, 7,
					-- layer=2 filter=228 channel=28
					-14, -6, -19, 5, 0, -6, -15, -15, -1,
					-- layer=2 filter=228 channel=29
					1, 0, -7, 4, 1, 7, -4, 1, 4,
					-- layer=2 filter=228 channel=30
					1, -17, -7, -12, -12, 0, 4, -9, 6,
					-- layer=2 filter=228 channel=31
					-11, -5, 2, -11, 0, -6, -12, 3, -9,
					-- layer=2 filter=228 channel=32
					-7, -7, 8, 4, 2, -4, 0, 3, 0,
					-- layer=2 filter=228 channel=33
					3, -8, -5, -5, 0, 5, 6, 0, 0,
					-- layer=2 filter=228 channel=34
					-10, -9, 1, -4, -3, -3, 2, -3, 5,
					-- layer=2 filter=228 channel=35
					-10, -9, -2, -2, 8, 6, -11, -17, -22,
					-- layer=2 filter=228 channel=36
					-11, 6, -4, -2, 0, 1, -2, 8, -1,
					-- layer=2 filter=228 channel=37
					-13, -4, -1, -15, 2, -7, 3, 0, -9,
					-- layer=2 filter=228 channel=38
					-1, -7, -3, -13, 2, 12, 4, 8, 0,
					-- layer=2 filter=228 channel=39
					-13, -7, 1, -8, -14, -18, -5, -9, 2,
					-- layer=2 filter=228 channel=40
					-7, 8, 3, 13, 4, 1, -4, 2, -4,
					-- layer=2 filter=228 channel=41
					-4, 0, -2, 12, -7, -9, -4, -1, 8,
					-- layer=2 filter=228 channel=42
					-4, -1, -3, 0, -3, -2, -10, -8, 4,
					-- layer=2 filter=228 channel=43
					-4, -2, -4, 0, -11, -1, -10, -3, -5,
					-- layer=2 filter=228 channel=44
					9, 0, 1, 10, -10, 5, -5, -4, 8,
					-- layer=2 filter=228 channel=45
					-9, -2, -3, 0, -2, 1, -8, -3, -11,
					-- layer=2 filter=228 channel=46
					-1, -1, 2, -8, 6, -9, -9, 6, -11,
					-- layer=2 filter=228 channel=47
					-7, -4, -16, 8, 5, 11, -12, -14, -12,
					-- layer=2 filter=228 channel=48
					5, 7, 1, -9, 1, -2, -8, 0, 6,
					-- layer=2 filter=228 channel=49
					-15, -1, -18, -19, -9, -6, 5, -2, 0,
					-- layer=2 filter=228 channel=50
					1, 4, 0, -5, -3, -1, -7, 0, -10,
					-- layer=2 filter=228 channel=51
					-8, -1, -5, -11, -7, -13, -10, -5, 0,
					-- layer=2 filter=228 channel=52
					-4, -6, -1, 3, -10, 2, 5, 6, 2,
					-- layer=2 filter=228 channel=53
					-10, 0, 7, -7, -6, 5, 8, -7, -7,
					-- layer=2 filter=228 channel=54
					-4, 2, 2, 2, -15, 0, -16, 2, -11,
					-- layer=2 filter=228 channel=55
					9, 0, 2, 1, 5, -2, -4, -8, -2,
					-- layer=2 filter=228 channel=56
					-10, -7, -4, 6, 0, -9, 7, 4, 3,
					-- layer=2 filter=228 channel=57
					1, -8, -9, -7, -10, 4, 2, -4, 6,
					-- layer=2 filter=228 channel=58
					6, 0, -4, 3, -9, -13, -17, -11, 3,
					-- layer=2 filter=228 channel=59
					0, -4, 10, -3, 5, -4, -6, -5, 17,
					-- layer=2 filter=228 channel=60
					-8, -10, 5, -7, 2, -5, -11, -4, -6,
					-- layer=2 filter=228 channel=61
					-1, -1, 11, -6, 6, 1, -4, -12, -1,
					-- layer=2 filter=228 channel=62
					-15, -6, -11, 0, 10, -3, -15, -9, 0,
					-- layer=2 filter=228 channel=63
					-18, -8, -1, -8, -15, -10, 0, -11, 1,
					-- layer=2 filter=228 channel=64
					-6, -2, -9, -5, -17, -5, 0, -11, -2,
					-- layer=2 filter=228 channel=65
					1, 4, -6, -9, 1, -7, -1, -13, -7,
					-- layer=2 filter=228 channel=66
					-5, 8, 1, 7, -1, 10, -5, 6, -11,
					-- layer=2 filter=228 channel=67
					0, 1, 6, -2, 0, 1, -14, 4, 1,
					-- layer=2 filter=228 channel=68
					2, 7, 7, -5, -4, -12, 8, -4, 7,
					-- layer=2 filter=228 channel=69
					-11, -14, -3, -16, -3, -23, -11, 0, -6,
					-- layer=2 filter=228 channel=70
					-2, -11, -13, 10, 5, 17, -6, 0, -9,
					-- layer=2 filter=228 channel=71
					0, 0, 0, -7, 2, 3, -7, -16, -13,
					-- layer=2 filter=228 channel=72
					3, -9, 0, -6, -1, -4, -2, -4, -15,
					-- layer=2 filter=228 channel=73
					3, 11, 12, -11, -8, -8, 0, 0, 9,
					-- layer=2 filter=228 channel=74
					-14, -5, -8, -17, -14, -15, -2, -13, -13,
					-- layer=2 filter=228 channel=75
					13, 13, -1, 1, -7, 10, -14, 5, 13,
					-- layer=2 filter=228 channel=76
					-5, 7, 0, -6, -11, 0, 6, 5, -8,
					-- layer=2 filter=228 channel=77
					-8, -5, 4, -7, 5, 6, -2, 8, -4,
					-- layer=2 filter=228 channel=78
					6, -12, -13, -5, -2, 5, 7, -7, -5,
					-- layer=2 filter=228 channel=79
					2, -8, -9, -8, 2, -6, 7, -2, -10,
					-- layer=2 filter=228 channel=80
					-2, -2, -8, -15, -1, -14, -4, -10, -15,
					-- layer=2 filter=228 channel=81
					-5, 6, -1, 0, 1, -7, -6, 0, -4,
					-- layer=2 filter=228 channel=82
					3, 8, -10, -3, 0, 3, -4, 8, -7,
					-- layer=2 filter=228 channel=83
					-7, 0, 5, 1, -5, -4, 0, -5, -8,
					-- layer=2 filter=228 channel=84
					4, -8, -5, 7, -2, 4, 0, -1, 8,
					-- layer=2 filter=228 channel=85
					5, 7, -3, 7, 5, -4, 0, 10, -2,
					-- layer=2 filter=228 channel=86
					0, -3, 0, 3, 5, 1, -6, -3, 9,
					-- layer=2 filter=228 channel=87
					0, 8, -10, 7, 9, 8, -7, 3, -7,
					-- layer=2 filter=228 channel=88
					-18, -3, -14, -12, -15, -14, 0, -15, 2,
					-- layer=2 filter=228 channel=89
					-9, -5, -1, -14, -12, -16, -6, -1, -9,
					-- layer=2 filter=228 channel=90
					10, -3, -9, 1, -2, -6, 0, 9, 3,
					-- layer=2 filter=228 channel=91
					2, -7, -2, -8, 0, -12, -7, 4, 9,
					-- layer=2 filter=228 channel=92
					-2, -13, -9, -13, 5, -2, -17, 3, 3,
					-- layer=2 filter=228 channel=93
					0, 0, 0, -3, 0, 2, -3, 0, -10,
					-- layer=2 filter=228 channel=94
					0, -8, -1, 0, -3, -6, -5, -1, 3,
					-- layer=2 filter=228 channel=95
					-3, -10, -7, 6, -5, 7, 1, 6, 2,
					-- layer=2 filter=228 channel=96
					-3, -13, 7, 3, 0, -19, -6, 1, 9,
					-- layer=2 filter=228 channel=97
					0, -4, 3, -5, -13, 0, 0, -10, -1,
					-- layer=2 filter=228 channel=98
					-13, -2, -8, 0, 3, -9, -7, -5, -4,
					-- layer=2 filter=228 channel=99
					1, 1, 2, -2, -3, -2, -2, -12, 6,
					-- layer=2 filter=228 channel=100
					-3, -1, -6, -4, 0, 7, -1, 9, -9,
					-- layer=2 filter=228 channel=101
					5, 9, 2, -8, 6, 2, -11, 0, 0,
					-- layer=2 filter=228 channel=102
					-10, -5, 3, -1, -8, -1, 3, -15, -8,
					-- layer=2 filter=228 channel=103
					8, 1, -9, 5, 0, -4, -11, 2, -5,
					-- layer=2 filter=228 channel=104
					-8, -14, -10, -2, 3, -11, -1, 8, 4,
					-- layer=2 filter=228 channel=105
					0, -2, 0, -12, 3, 9, 5, -2, 4,
					-- layer=2 filter=228 channel=106
					18, -3, -2, -8, -12, -2, -10, -17, -15,
					-- layer=2 filter=228 channel=107
					7, -2, 9, 0, 5, -10, -9, 9, 3,
					-- layer=2 filter=228 channel=108
					-1, -1, -1, -13, 1, 0, -5, -4, -2,
					-- layer=2 filter=228 channel=109
					-1, 7, 2, 7, 0, -9, 3, -4, 8,
					-- layer=2 filter=228 channel=110
					-12, 1, -13, -12, 0, -5, -7, 0, -14,
					-- layer=2 filter=228 channel=111
					-3, -4, -7, 0, 6, -9, -6, 5, 4,
					-- layer=2 filter=228 channel=112
					-1, 7, -7, -6, -3, -11, -2, -4, -10,
					-- layer=2 filter=228 channel=113
					-9, -9, 3, 10, 5, 7, -10, -4, 5,
					-- layer=2 filter=228 channel=114
					-4, -4, 0, -9, -6, 1, 3, 0, 3,
					-- layer=2 filter=228 channel=115
					0, 2, -8, -3, 1, 6, 1, -9, -9,
					-- layer=2 filter=228 channel=116
					-7, -4, -3, 3, -6, 2, -1, 1, 8,
					-- layer=2 filter=228 channel=117
					-14, -3, 10, 2, 1, 3, -10, -9, -4,
					-- layer=2 filter=228 channel=118
					3, -15, 5, 4, -10, 6, -12, 0, 0,
					-- layer=2 filter=228 channel=119
					-3, 0, -6, 9, 2, -3, -10, -6, -5,
					-- layer=2 filter=228 channel=120
					-7, -1, -5, -4, 0, 10, -1, 10, 3,
					-- layer=2 filter=228 channel=121
					10, 7, -7, 4, 4, 3, -10, 8, -2,
					-- layer=2 filter=228 channel=122
					7, 6, 3, 5, 6, -7, -1, 0, 8,
					-- layer=2 filter=228 channel=123
					12, 5, 7, -8, -1, 5, -10, 0, -12,
					-- layer=2 filter=228 channel=124
					8, 7, -7, 1, -9, -6, -14, -9, -8,
					-- layer=2 filter=228 channel=125
					-7, -5, 10, -10, 11, 5, 3, 8, 0,
					-- layer=2 filter=228 channel=126
					3, -2, -3, 4, -7, 6, 0, -2, 3,
					-- layer=2 filter=228 channel=127
					-2, -12, -9, -9, -2, -18, -7, 1, 5,
					-- layer=2 filter=229 channel=0
					18, 11, 5, 19, -11, -3, -2, 0, -21,
					-- layer=2 filter=229 channel=1
					-12, -1, 42, -1, -1, 29, -31, 0, 23,
					-- layer=2 filter=229 channel=2
					0, -6, -12, -3, -2, -4, -10, -2, 7,
					-- layer=2 filter=229 channel=3
					27, -17, -4, 26, 0, -27, 26, 13, 19,
					-- layer=2 filter=229 channel=4
					4, 5, -8, -2, -10, 15, -97, -78, -65,
					-- layer=2 filter=229 channel=5
					34, 9, -10, -5, -15, -25, 22, -1, -29,
					-- layer=2 filter=229 channel=6
					-2, 24, 20, 6, -19, 33, 22, -38, 34,
					-- layer=2 filter=229 channel=7
					48, -7, -13, 6, -26, 19, -28, 12, -30,
					-- layer=2 filter=229 channel=8
					-2, 7, -9, -5, -3, -4, -9, -4, -4,
					-- layer=2 filter=229 channel=9
					1, -29, -18, 30, 49, 0, -8, 27, 30,
					-- layer=2 filter=229 channel=10
					24, -1, 18, -15, -27, -5, -26, -8, -24,
					-- layer=2 filter=229 channel=11
					9, 0, -20, 19, -20, -7, 14, 15, 2,
					-- layer=2 filter=229 channel=12
					7, 3, 14, 30, 28, 22, -21, 2, 6,
					-- layer=2 filter=229 channel=13
					0, -7, -2, 7, 6, -1, 0, 0, 3,
					-- layer=2 filter=229 channel=14
					11, -7, -1, 23, 22, 24, -12, 14, 25,
					-- layer=2 filter=229 channel=15
					-13, 0, -64, 38, 10, 26, -10, 2, -8,
					-- layer=2 filter=229 channel=16
					0, 19, 7, -28, 0, 20, -55, -39, -6,
					-- layer=2 filter=229 channel=17
					9, 7, -4, 3, -9, 3, 1, 8, 0,
					-- layer=2 filter=229 channel=18
					-9, 14, -28, 0, -9, 4, -35, -70, -21,
					-- layer=2 filter=229 channel=19
					2, 4, 66, -22, 49, 40, -5, -34, 36,
					-- layer=2 filter=229 channel=20
					-4, -5, 5, -1, 0, 6, -2, -6, 7,
					-- layer=2 filter=229 channel=21
					5, -1, -2, 21, 15, 15, -10, 4, 21,
					-- layer=2 filter=229 channel=22
					4, 4, -2, -7, -7, -1, 7, 0, -1,
					-- layer=2 filter=229 channel=23
					1, 20, 19, -7, 46, 34, -66, -42, -42,
					-- layer=2 filter=229 channel=24
					30, 11, 9, 24, 5, -24, 9, 15, 11,
					-- layer=2 filter=229 channel=25
					55, 3, -16, 18, -12, -29, 30, 20, 28,
					-- layer=2 filter=229 channel=26
					9, -2, 2, -2, -5, -7, 0, 9, -1,
					-- layer=2 filter=229 channel=27
					3, 13, 33, 2, 4, 30, -9, -18, -1,
					-- layer=2 filter=229 channel=28
					-1, -21, -34, -10, -20, -25, -13, 1, 0,
					-- layer=2 filter=229 channel=29
					5, -6, -9, -7, -2, 0, 4, -10, -8,
					-- layer=2 filter=229 channel=30
					-14, 3, 25, -46, 31, 48, -75, -52, -41,
					-- layer=2 filter=229 channel=31
					39, 13, -8, 36, -1, 21, -17, -31, -1,
					-- layer=2 filter=229 channel=32
					9, -1, -6, 5, 8, 10, 5, -2, 10,
					-- layer=2 filter=229 channel=33
					20, -3, -36, 23, -37, -11, 33, -4, 14,
					-- layer=2 filter=229 channel=34
					23, 34, -16, -28, 44, -20, 24, -7, -45,
					-- layer=2 filter=229 channel=35
					13, 13, 24, 15, 2, -12, -42, -28, -25,
					-- layer=2 filter=229 channel=36
					5, -1, -11, -4, 2, 2, -4, -9, 5,
					-- layer=2 filter=229 channel=37
					-1, 2, 12, 10, -15, -24, 26, 6, 9,
					-- layer=2 filter=229 channel=38
					-21, 23, 17, 3, 1, 26, 16, -42, -17,
					-- layer=2 filter=229 channel=39
					10, 21, 24, -44, 14, 23, -52, -51, -17,
					-- layer=2 filter=229 channel=40
					-2, 26, -12, 27, 71, -25, -7, -50, 2,
					-- layer=2 filter=229 channel=41
					7, -2, -6, 6, 7, -7, -3, 3, 3,
					-- layer=2 filter=229 channel=42
					-12, 13, 29, 24, 27, 7, -66, -1, -13,
					-- layer=2 filter=229 channel=43
					5, -5, -6, 3, 33, -3, 3, -4, -19,
					-- layer=2 filter=229 channel=44
					0, -7, 10, -5, -9, -8, -6, -4, -8,
					-- layer=2 filter=229 channel=45
					18, -4, -23, -5, 5, 58, -74, -68, 32,
					-- layer=2 filter=229 channel=46
					11, 40, 33, -45, -1, 3, -8, -34, -46,
					-- layer=2 filter=229 channel=47
					-3, -11, -25, -54, -25, 8, -3, 1, -17,
					-- layer=2 filter=229 channel=48
					6, -9, 5, 1, 4, -8, 7, 4, 2,
					-- layer=2 filter=229 channel=49
					15, -4, 14, 4, 3, 20, -24, 1, 5,
					-- layer=2 filter=229 channel=50
					-6, -7, -11, 5, 2, -14, 12, 0, -8,
					-- layer=2 filter=229 channel=51
					17, -15, -20, 27, 0, -25, 28, 7, -2,
					-- layer=2 filter=229 channel=52
					-36, -44, -23, 24, -8, 10, -14, -5, 28,
					-- layer=2 filter=229 channel=53
					-78, -18, 20, -3, -28, 28, 16, -32, 54,
					-- layer=2 filter=229 channel=54
					6, -7, -7, 0, 4, 16, 18, -6, -13,
					-- layer=2 filter=229 channel=55
					-10, -1, 7, 3, 2, 0, -2, 3, 5,
					-- layer=2 filter=229 channel=56
					7, 0, 3, 24, -15, -9, 26, -9, 8,
					-- layer=2 filter=229 channel=57
					-4, 1, 6, -3, -7, 6, 15, 0, -7,
					-- layer=2 filter=229 channel=58
					12, 10, 40, 14, 27, 16, -11, -35, 0,
					-- layer=2 filter=229 channel=59
					-74, -28, 4, -29, 46, 7, 12, -21, 34,
					-- layer=2 filter=229 channel=60
					22, 7, 23, -6, 17, 9, 0, -29, -13,
					-- layer=2 filter=229 channel=61
					-29, -14, -13, -18, -3, -12, -56, -22, -24,
					-- layer=2 filter=229 channel=62
					7, -1, 51, 5, -12, 4, 46, -42, -20,
					-- layer=2 filter=229 channel=63
					-45, 11, 0, -56, -9, 26, -54, -31, -35,
					-- layer=2 filter=229 channel=64
					-18, 21, 28, -20, 23, 41, -55, -23, -18,
					-- layer=2 filter=229 channel=65
					-18, 32, 13, -7, 3, 4, -18, 6, -10,
					-- layer=2 filter=229 channel=66
					38, -66, 1, -16, -8, -45, -31, -5, -10,
					-- layer=2 filter=229 channel=67
					-22, -11, -6, 8, 18, 11, -23, -68, -31,
					-- layer=2 filter=229 channel=68
					4, 6, -4, 10, 7, 0, 5, -4, 0,
					-- layer=2 filter=229 channel=69
					1, 10, 11, 6, 55, 24, -37, 16, 20,
					-- layer=2 filter=229 channel=70
					8, 0, 17, 7, -25, -15, -16, -4, -4,
					-- layer=2 filter=229 channel=71
					16, 6, 3, 6, 1, 22, 13, 9, 39,
					-- layer=2 filter=229 channel=72
					22, 8, -33, 3, -4, -8, 9, 44, 42,
					-- layer=2 filter=229 channel=73
					42, -27, -18, 0, 1, 10, -17, -25, 5,
					-- layer=2 filter=229 channel=74
					-27, 0, -4, -40, 6, 6, -66, -90, -60,
					-- layer=2 filter=229 channel=75
					16, -8, 0, 6, -1, 4, -80, -11, 32,
					-- layer=2 filter=229 channel=76
					22, 27, -10, 62, -105, 49, -45, -69, -10,
					-- layer=2 filter=229 channel=77
					9, 2, -6, -7, 8, 6, 7, 3, -1,
					-- layer=2 filter=229 channel=78
					12, -14, -8, 25, -24, -41, 12, 7, 1,
					-- layer=2 filter=229 channel=79
					-3, -7, -4, 2, 11, -4, 2, 11, 9,
					-- layer=2 filter=229 channel=80
					-19, 0, 35, -52, -8, -6, -80, -59, -61,
					-- layer=2 filter=229 channel=81
					9, 9, -7, 0, -1, 4, -5, 4, -6,
					-- layer=2 filter=229 channel=82
					10, -6, 0, 3, -6, -3, 2, 7, 5,
					-- layer=2 filter=229 channel=83
					-27, 11, 14, -25, 40, 17, -65, -46, -37,
					-- layer=2 filter=229 channel=84
					1, -2, 5, 7, 4, 9, 7, 4, -6,
					-- layer=2 filter=229 channel=85
					-16, -4, -10, 2, 5, -3, -1, 0, -15,
					-- layer=2 filter=229 channel=86
					-3, -6, -19, -5, -11, -8, -9, 9, -5,
					-- layer=2 filter=229 channel=87
					6, 14, 18, 31, 5, 32, -21, -37, -48,
					-- layer=2 filter=229 channel=88
					-74, 2, 7, -20, 41, 21, -92, -29, -3,
					-- layer=2 filter=229 channel=89
					-1, 22, 2, -1, 7, -2, -25, 6, 12,
					-- layer=2 filter=229 channel=90
					1, -8, 10, -3, 4, 0, 5, -5, -6,
					-- layer=2 filter=229 channel=91
					29, -5, 17, 19, -13, -11, -26, -6, 33,
					-- layer=2 filter=229 channel=92
					25, 6, 1, 12, 17, 26, -12, -1, 23,
					-- layer=2 filter=229 channel=93
					3, 9, 66, -39, -19, 72, 9, 23, 2,
					-- layer=2 filter=229 channel=94
					-10, -21, -1, -35, 23, 26, 8, 10, 27,
					-- layer=2 filter=229 channel=95
					-10, -19, -21, 0, -16, -21, -16, -5, -13,
					-- layer=2 filter=229 channel=96
					-1, 11, 41, -27, -9, 11, 2, 38, -4,
					-- layer=2 filter=229 channel=97
					22, -5, 18, 18, 0, -29, -19, 29, 0,
					-- layer=2 filter=229 channel=98
					11, -24, -6, -4, -26, 1, -19, 34, 11,
					-- layer=2 filter=229 channel=99
					-68, -21, 10, 1, 0, -2, -21, 19, 37,
					-- layer=2 filter=229 channel=100
					-42, 11, 42, -11, 16, 12, -14, -71, -65,
					-- layer=2 filter=229 channel=101
					35, -15, 3, 42, -11, -8, 3, 17, 25,
					-- layer=2 filter=229 channel=102
					6, 21, 0, -18, -26, -6, -19, 0, -27,
					-- layer=2 filter=229 channel=103
					-18, -3, 2, -9, -4, -4, -53, -21, 0,
					-- layer=2 filter=229 channel=104
					15, -15, -3, -3, -35, 31, 9, -26, -27,
					-- layer=2 filter=229 channel=105
					22, -11, -21, 18, 55, 34, -37, -53, 16,
					-- layer=2 filter=229 channel=106
					46, 12, -19, 29, -11, -13, 17, 15, 10,
					-- layer=2 filter=229 channel=107
					24, 11, 19, 33, 34, -5, 44, 14, -5,
					-- layer=2 filter=229 channel=108
					-11, -12, 1, -12, 8, 18, -12, -22, -12,
					-- layer=2 filter=229 channel=109
					0, 1, 11, 4, 9, -2, -2, -7, -2,
					-- layer=2 filter=229 channel=110
					4, 35, 42, -8, 9, 39, -49, 5, 2,
					-- layer=2 filter=229 channel=111
					4, 5, 5, -1, -10, 2, 7, 0, 1,
					-- layer=2 filter=229 channel=112
					14, 8, -16, 15, -11, -43, 32, 22, -3,
					-- layer=2 filter=229 channel=113
					-18, -1, 12, -37, 29, 33, -49, -2, 3,
					-- layer=2 filter=229 channel=114
					-1, -5, 3, -4, -18, 9, -8, 12, 6,
					-- layer=2 filter=229 channel=115
					-7, 9, 7, 7, -5, 2, 2, -1, 8,
					-- layer=2 filter=229 channel=116
					0, 15, 13, 11, -2, 27, -30, -15, -43,
					-- layer=2 filter=229 channel=117
					57, -55, -35, -36, -5, 37, -26, 47, -14,
					-- layer=2 filter=229 channel=118
					24, 0, 33, 29, 1, 8, 9, -18, 0,
					-- layer=2 filter=229 channel=119
					3, 0, 5, 13, 12, 3, -30, -83, -40,
					-- layer=2 filter=229 channel=120
					-6, -6, -4, 5, -8, 10, -6, -2, -1,
					-- layer=2 filter=229 channel=121
					3, 0, 6, -2, 8, -8, 3, 0, 4,
					-- layer=2 filter=229 channel=122
					-4, -1, 5, 5, 7, -8, 8, 3, 3,
					-- layer=2 filter=229 channel=123
					-29, -16, -34, -12, -20, -9, -15, -5, -14,
					-- layer=2 filter=229 channel=124
					13, -9, -40, 54, -26, 2, -16, -9, -30,
					-- layer=2 filter=229 channel=125
					4, -8, 4, 10, 1, -15, 2, -6, 11,
					-- layer=2 filter=229 channel=126
					-24, 52, 46, 1, 23, -7, -22, -14, -1,
					-- layer=2 filter=229 channel=127
					-18, 12, 12, 6, 56, -7, -8, -28, 58,
					-- layer=2 filter=230 channel=0
					-3, -12, -2, -10, -8, 5, -8, 5, -4,
					-- layer=2 filter=230 channel=1
					-12, -5, -2, 3, -1, 3, 2, 0, -1,
					-- layer=2 filter=230 channel=2
					-8, 4, 11, 5, 4, 6, 7, 0, -8,
					-- layer=2 filter=230 channel=3
					-4, -10, -4, 1, 8, -10, -2, 0, 1,
					-- layer=2 filter=230 channel=4
					2, 4, 7, 0, -3, 2, -11, 7, 0,
					-- layer=2 filter=230 channel=5
					-10, -6, -14, -7, 3, 5, -6, -6, 8,
					-- layer=2 filter=230 channel=6
					-9, 2, -10, -1, 5, 4, -2, 1, 1,
					-- layer=2 filter=230 channel=7
					-8, 8, -1, -7, -13, -10, -9, -8, -12,
					-- layer=2 filter=230 channel=8
					4, 2, 5, 3, 7, 7, 10, 1, 4,
					-- layer=2 filter=230 channel=9
					-7, 3, 3, 5, -8, 10, 7, -1, -10,
					-- layer=2 filter=230 channel=10
					-10, -9, -12, 0, -7, -5, -3, -6, -5,
					-- layer=2 filter=230 channel=11
					1, -2, -10, -17, -3, -17, -6, -15, -11,
					-- layer=2 filter=230 channel=12
					0, -4, -10, 4, 4, -6, 0, -8, 6,
					-- layer=2 filter=230 channel=13
					0, -1, 6, -5, 1, -6, 9, -9, 0,
					-- layer=2 filter=230 channel=14
					2, -7, 5, -1, 7, -6, 9, -10, -5,
					-- layer=2 filter=230 channel=15
					0, 6, 0, -8, 6, -3, 1, 5, 10,
					-- layer=2 filter=230 channel=16
					-3, -7, -7, -10, 0, -7, -8, -1, -9,
					-- layer=2 filter=230 channel=17
					7, 7, 8, -1, -2, -1, 7, 7, -10,
					-- layer=2 filter=230 channel=18
					-2, 0, -8, -8, 2, 4, -3, 3, -5,
					-- layer=2 filter=230 channel=19
					-11, 0, 11, -13, 0, -11, 5, -9, 0,
					-- layer=2 filter=230 channel=20
					0, 5, -2, 2, 10, 6, -2, -6, 8,
					-- layer=2 filter=230 channel=21
					-4, 1, 0, 2, -11, 0, -7, 10, -8,
					-- layer=2 filter=230 channel=22
					6, 0, -6, 0, 8, 4, 7, 1, -4,
					-- layer=2 filter=230 channel=23
					7, 8, -10, 5, 1, -7, 2, 7, 4,
					-- layer=2 filter=230 channel=24
					-5, -3, -2, -11, -7, 3, -4, -9, -9,
					-- layer=2 filter=230 channel=25
					1, -5, -3, 0, -14, -5, -11, -1, -14,
					-- layer=2 filter=230 channel=26
					-6, 9, 4, -3, -6, -4, 3, 5, 0,
					-- layer=2 filter=230 channel=27
					-8, 1, -6, -5, -13, -2, 0, -4, -8,
					-- layer=2 filter=230 channel=28
					-8, -1, -7, 1, -12, -6, -12, -9, 0,
					-- layer=2 filter=230 channel=29
					-8, 5, 1, 10, 0, 10, -7, 7, 4,
					-- layer=2 filter=230 channel=30
					-7, -9, -5, -7, -6, -7, -1, 5, -5,
					-- layer=2 filter=230 channel=31
					-1, -10, 1, -1, -8, 1, 8, 4, 5,
					-- layer=2 filter=230 channel=32
					0, 0, 5, 8, 0, -8, 0, 5, 8,
					-- layer=2 filter=230 channel=33
					-8, 5, -5, -3, 2, 2, -8, 7, 8,
					-- layer=2 filter=230 channel=34
					-16, 5, 9, -6, -5, 0, -2, -10, 1,
					-- layer=2 filter=230 channel=35
					-8, 0, 0, -7, 0, -12, -1, -7, -11,
					-- layer=2 filter=230 channel=36
					-8, 5, -9, 2, 2, -10, 4, 4, 3,
					-- layer=2 filter=230 channel=37
					0, -17, -8, 0, 0, 2, 1, -4, -11,
					-- layer=2 filter=230 channel=38
					-2, -2, -11, -9, -2, 5, 0, 1, 6,
					-- layer=2 filter=230 channel=39
					-2, 5, -3, -5, 0, -5, 10, -9, -4,
					-- layer=2 filter=230 channel=40
					-4, -3, 1, -5, 4, -3, -9, 1, -7,
					-- layer=2 filter=230 channel=41
					-7, -4, -3, 7, 2, -2, -8, 6, -2,
					-- layer=2 filter=230 channel=42
					-1, 2, -10, 0, -12, -5, 7, 4, -7,
					-- layer=2 filter=230 channel=43
					-6, -3, 5, -8, -10, 0, 6, -1, 5,
					-- layer=2 filter=230 channel=44
					-5, -4, 1, -1, 0, 4, 9, -8, 3,
					-- layer=2 filter=230 channel=45
					-7, 0, 6, 5, 6, -2, -6, 6, 10,
					-- layer=2 filter=230 channel=46
					0, -2, -9, -8, -7, -7, 7, 2, 2,
					-- layer=2 filter=230 channel=47
					4, 3, -3, -2, -2, 1, -5, -8, -7,
					-- layer=2 filter=230 channel=48
					7, -7, -4, -7, -6, 3, 5, -6, -6,
					-- layer=2 filter=230 channel=49
					3, 0, 7, 8, 5, 6, -9, -7, -7,
					-- layer=2 filter=230 channel=50
					-6, -8, 1, 5, 0, -10, -4, 7, 7,
					-- layer=2 filter=230 channel=51
					0, -14, 6, -4, 2, 2, -1, -4, -4,
					-- layer=2 filter=230 channel=52
					-2, -15, -2, -15, -2, 1, 3, -13, -8,
					-- layer=2 filter=230 channel=53
					3, 2, -11, -8, 0, -10, -5, -8, 2,
					-- layer=2 filter=230 channel=54
					-12, -6, 2, -3, -10, 4, -2, 4, -12,
					-- layer=2 filter=230 channel=55
					9, -4, 7, 8, -5, 0, -5, -10, 8,
					-- layer=2 filter=230 channel=56
					0, -15, 1, -1, -7, -6, -10, -10, -11,
					-- layer=2 filter=230 channel=57
					-3, 8, 7, 0, 3, -4, -4, 4, 6,
					-- layer=2 filter=230 channel=58
					0, 2, -8, -12, 1, 5, -14, 1, 4,
					-- layer=2 filter=230 channel=59
					3, -5, -7, -7, -12, 1, -2, 0, -12,
					-- layer=2 filter=230 channel=60
					-6, -6, -1, 3, -6, -2, -5, -9, 2,
					-- layer=2 filter=230 channel=61
					6, 3, -2, 0, -8, 11, 5, -7, -8,
					-- layer=2 filter=230 channel=62
					3, -13, 2, -1, -8, -9, 2, -8, 3,
					-- layer=2 filter=230 channel=63
					0, -6, 0, -4, -8, -2, 5, 9, 5,
					-- layer=2 filter=230 channel=64
					1, -10, -3, -5, -7, -4, -6, 3, 6,
					-- layer=2 filter=230 channel=65
					-1, -3, -5, -2, 2, -11, 8, 9, 4,
					-- layer=2 filter=230 channel=66
					-4, -2, -2, 4, -7, -5, 0, 1, -4,
					-- layer=2 filter=230 channel=67
					-5, -4, 1, -11, 2, -2, 0, -3, 8,
					-- layer=2 filter=230 channel=68
					8, 0, -9, 9, 6, 6, -5, -2, -6,
					-- layer=2 filter=230 channel=69
					-1, -11, 5, -7, 0, 7, -2, 8, 2,
					-- layer=2 filter=230 channel=70
					-7, 0, -6, -3, -13, -7, -6, -5, -6,
					-- layer=2 filter=230 channel=71
					-3, -9, 7, 3, 0, -4, 9, 0, -1,
					-- layer=2 filter=230 channel=72
					0, -1, -4, -1, 5, -13, 5, -6, -5,
					-- layer=2 filter=230 channel=73
					-1, 0, 7, 5, 3, -5, 9, -5, -2,
					-- layer=2 filter=230 channel=74
					-5, -4, 3, -2, 7, -4, -4, 6, 5,
					-- layer=2 filter=230 channel=75
					2, 4, -3, -11, -8, -8, -8, -4, 5,
					-- layer=2 filter=230 channel=76
					1, -11, -5, -8, -5, 10, -8, -8, -8,
					-- layer=2 filter=230 channel=77
					-2, -5, 3, 2, -2, -6, 0, 8, 11,
					-- layer=2 filter=230 channel=78
					-2, -11, -2, 0, 6, 4, -6, 4, -10,
					-- layer=2 filter=230 channel=79
					10, -7, -8, 3, -4, -3, -3, -2, 6,
					-- layer=2 filter=230 channel=80
					4, -10, 3, 2, -4, -5, 4, 1, 2,
					-- layer=2 filter=230 channel=81
					1, 6, -9, 12, 0, -2, 10, -9, 9,
					-- layer=2 filter=230 channel=82
					7, -3, 1, -1, -9, -7, 7, -7, 4,
					-- layer=2 filter=230 channel=83
					4, -2, 3, 1, -8, 8, -3, -7, -7,
					-- layer=2 filter=230 channel=84
					-3, -6, 4, 8, 5, 0, -6, -3, 0,
					-- layer=2 filter=230 channel=85
					2, -9, 1, -2, 0, -4, -11, 8, -5,
					-- layer=2 filter=230 channel=86
					1, 5, -7, 1, -8, -10, -10, -1, -11,
					-- layer=2 filter=230 channel=87
					-6, -7, 5, 8, -6, 9, -1, 1, -10,
					-- layer=2 filter=230 channel=88
					6, -5, -9, -1, -5, -5, -4, -8, 7,
					-- layer=2 filter=230 channel=89
					-5, 2, -4, -3, -3, -3, 6, 4, -7,
					-- layer=2 filter=230 channel=90
					0, -1, 4, 8, 1, 0, -1, 9, 10,
					-- layer=2 filter=230 channel=91
					-2, -4, -5, -8, -10, 5, -7, 0, -14,
					-- layer=2 filter=230 channel=92
					-11, -9, -7, 1, -5, -1, -10, -1, -1,
					-- layer=2 filter=230 channel=93
					7, -5, -6, 9, -2, -5, -6, -4, 3,
					-- layer=2 filter=230 channel=94
					0, -10, -6, 0, -6, 1, -8, -12, 2,
					-- layer=2 filter=230 channel=95
					-5, -2, -6, 0, -1, -7, -5, 9, 1,
					-- layer=2 filter=230 channel=96
					-6, 6, -4, -8, 0, -5, -3, -3, -10,
					-- layer=2 filter=230 channel=97
					2, -11, 1, -1, -2, 0, 0, -5, -5,
					-- layer=2 filter=230 channel=98
					2, -10, -12, -9, -7, -8, -16, -2, 3,
					-- layer=2 filter=230 channel=99
					0, 2, -4, -10, -10, 2, -14, -6, 5,
					-- layer=2 filter=230 channel=100
					-10, 1, -8, 4, -1, 7, -2, -15, -8,
					-- layer=2 filter=230 channel=101
					-12, -7, -2, 4, 0, -1, 7, -1, -8,
					-- layer=2 filter=230 channel=102
					0, -6, -14, -2, -13, -3, -8, -4, 4,
					-- layer=2 filter=230 channel=103
					-9, 9, -3, 6, -9, -4, 0, 1, 10,
					-- layer=2 filter=230 channel=104
					-8, -8, -10, -5, -2, -4, 0, -5, 5,
					-- layer=2 filter=230 channel=105
					-7, 1, 6, -8, 0, -9, 1, -2, -11,
					-- layer=2 filter=230 channel=106
					-3, 4, -11, -10, -11, -6, -2, 4, -3,
					-- layer=2 filter=230 channel=107
					10, 3, 0, 3, 3, -3, -2, -6, -3,
					-- layer=2 filter=230 channel=108
					-7, -3, -6, -7, 0, -5, 6, -1, 2,
					-- layer=2 filter=230 channel=109
					6, -9, -2, 1, 11, 2, -8, 5, 2,
					-- layer=2 filter=230 channel=110
					-2, 3, 4, 1, -5, 0, -4, -3, 7,
					-- layer=2 filter=230 channel=111
					-5, -4, -6, -5, 4, -3, -5, 1, -5,
					-- layer=2 filter=230 channel=112
					8, -9, -1, -12, 0, -3, 8, 11, 0,
					-- layer=2 filter=230 channel=113
					-2, -10, -3, -8, 8, -4, -4, 0, -3,
					-- layer=2 filter=230 channel=114
					1, 0, -9, 6, -5, 7, 9, -5, 1,
					-- layer=2 filter=230 channel=115
					4, -6, -4, 10, 5, 2, -3, 10, 0,
					-- layer=2 filter=230 channel=116
					-6, -5, -8, -4, -11, 0, 4, -4, 2,
					-- layer=2 filter=230 channel=117
					-2, -7, 7, 3, -7, -5, 8, 0, -4,
					-- layer=2 filter=230 channel=118
					-1, -9, 7, -1, 2, -9, 4, -4, 8,
					-- layer=2 filter=230 channel=119
					3, 1, -6, 4, -11, -6, 9, -3, 9,
					-- layer=2 filter=230 channel=120
					-1, 8, 7, 0, -6, -9, -5, 9, 1,
					-- layer=2 filter=230 channel=121
					9, -6, -7, 3, -5, -2, -6, 2, 1,
					-- layer=2 filter=230 channel=122
					7, 0, 1, 9, -2, -7, -2, 7, 9,
					-- layer=2 filter=230 channel=123
					3, -1, -14, -3, 4, -7, -5, 0, 6,
					-- layer=2 filter=230 channel=124
					-6, -8, 8, -7, 5, -1, 7, 4, 2,
					-- layer=2 filter=230 channel=125
					-4, 2, 4, -8, -1, -5, 7, -8, -7,
					-- layer=2 filter=230 channel=126
					3, 3, -10, 10, -7, -7, -4, 1, -6,
					-- layer=2 filter=230 channel=127
					-1, 3, 7, -1, -7, -3, 0, 0, -6,
					-- layer=2 filter=231 channel=0
					-7, 3, 4, -10, 0, 5, 4, 0, 7,
					-- layer=2 filter=231 channel=1
					0, 6, -3, 4, 3, -1, -8, -9, 0,
					-- layer=2 filter=231 channel=2
					7, 6, 6, 3, -1, 0, -7, 1, 0,
					-- layer=2 filter=231 channel=3
					4, -5, -5, 0, 2, 0, -3, 5, 1,
					-- layer=2 filter=231 channel=4
					-1, 3, 2, 3, 8, -1, 8, 0, -9,
					-- layer=2 filter=231 channel=5
					3, -9, -2, 5, -13, 4, -6, -2, 0,
					-- layer=2 filter=231 channel=6
					-1, -8, 3, -9, 1, -2, 8, -6, 3,
					-- layer=2 filter=231 channel=7
					8, -1, -6, -10, 6, -1, 1, -8, 0,
					-- layer=2 filter=231 channel=8
					1, 2, 7, 1, -4, 8, -2, 2, 8,
					-- layer=2 filter=231 channel=9
					-7, -9, -2, -6, 1, -7, 8, -9, -10,
					-- layer=2 filter=231 channel=10
					-1, -10, 2, 11, 3, 3, -11, 0, -10,
					-- layer=2 filter=231 channel=11
					-9, -7, -2, 0, -9, -1, -1, 2, -6,
					-- layer=2 filter=231 channel=12
					-5, 0, -1, -6, 9, -4, -6, 0, 2,
					-- layer=2 filter=231 channel=13
					1, -3, 3, 5, -1, 4, -3, -7, -11,
					-- layer=2 filter=231 channel=14
					6, 1, -12, -3, -7, 1, 4, 5, -2,
					-- layer=2 filter=231 channel=15
					-9, -3, 7, -2, -11, -6, -1, 4, 1,
					-- layer=2 filter=231 channel=16
					3, 8, 8, -6, 6, -8, -2, 8, 7,
					-- layer=2 filter=231 channel=17
					-5, -4, -2, -5, -5, -4, 8, 2, 7,
					-- layer=2 filter=231 channel=18
					6, -2, -2, 4, 0, -7, 5, 0, -9,
					-- layer=2 filter=231 channel=19
					0, -7, 5, -3, 1, 0, -4, 0, -11,
					-- layer=2 filter=231 channel=20
					1, 6, -1, -2, -1, 2, -8, 0, 3,
					-- layer=2 filter=231 channel=21
					-5, 8, -10, -1, 2, 3, -3, -2, -5,
					-- layer=2 filter=231 channel=22
					-7, 5, -4, -1, 0, -2, 7, 7, 2,
					-- layer=2 filter=231 channel=23
					-9, -1, 7, -11, -8, 5, -3, -9, 0,
					-- layer=2 filter=231 channel=24
					7, -4, 6, -8, -10, 0, -2, 5, 2,
					-- layer=2 filter=231 channel=25
					-8, -2, -8, -8, -1, -6, 5, -12, -10,
					-- layer=2 filter=231 channel=26
					-6, 6, 5, 4, 2, 4, -7, -6, -8,
					-- layer=2 filter=231 channel=27
					-4, -6, 0, 1, -11, 4, 3, 4, 0,
					-- layer=2 filter=231 channel=28
					-3, 6, -1, -10, 0, -6, 3, -10, -11,
					-- layer=2 filter=231 channel=29
					9, -9, -4, 5, 7, 1, 1, 2, 4,
					-- layer=2 filter=231 channel=30
					-13, 7, 2, 5, 0, -4, -10, 2, -8,
					-- layer=2 filter=231 channel=31
					0, -9, 3, 3, 1, 5, 2, 0, -6,
					-- layer=2 filter=231 channel=32
					5, -3, -7, -8, -3, 8, 0, 5, 3,
					-- layer=2 filter=231 channel=33
					-4, 7, -5, -9, -6, 2, 4, 7, 7,
					-- layer=2 filter=231 channel=34
					2, -7, 1, -9, 2, -5, 0, -11, -4,
					-- layer=2 filter=231 channel=35
					-11, -3, 0, -9, -5, -1, -5, 0, -2,
					-- layer=2 filter=231 channel=36
					-7, 8, 0, -5, -2, -1, 1, 0, 7,
					-- layer=2 filter=231 channel=37
					4, -1, 0, -4, -4, -9, -6, -5, -7,
					-- layer=2 filter=231 channel=38
					0, 0, -12, -10, -6, -13, 0, -2, -7,
					-- layer=2 filter=231 channel=39
					-5, 3, 1, -3, -11, -7, -7, 2, 5,
					-- layer=2 filter=231 channel=40
					-8, 3, 7, -11, 6, 8, -2, 4, -3,
					-- layer=2 filter=231 channel=41
					6, -2, -3, 10, -10, 5, -2, -6, -8,
					-- layer=2 filter=231 channel=42
					-7, -11, 2, 0, 3, -3, 6, -8, 1,
					-- layer=2 filter=231 channel=43
					-3, -8, 5, -6, 3, -12, -5, -6, -2,
					-- layer=2 filter=231 channel=44
					0, -10, -1, 2, -10, -7, 8, 8, 7,
					-- layer=2 filter=231 channel=45
					7, -4, -7, 7, -8, -10, 0, -1, 8,
					-- layer=2 filter=231 channel=46
					2, 2, 0, 0, -12, 7, -5, 8, 6,
					-- layer=2 filter=231 channel=47
					0, 0, -3, -13, 5, 0, -11, 1, -1,
					-- layer=2 filter=231 channel=48
					9, -2, -7, 7, -6, -5, 10, 4, 4,
					-- layer=2 filter=231 channel=49
					-12, 5, -2, 8, -4, -5, 6, 1, 2,
					-- layer=2 filter=231 channel=50
					-4, 8, 0, 11, 9, -6, -9, -3, 3,
					-- layer=2 filter=231 channel=51
					-5, -9, -8, 0, 6, -10, -6, 1, 0,
					-- layer=2 filter=231 channel=52
					-10, -11, -7, -1, -12, -1, -5, -1, 0,
					-- layer=2 filter=231 channel=53
					1, 7, -11, 1, 5, -3, 5, 0, 7,
					-- layer=2 filter=231 channel=54
					-6, -12, 2, 2, 6, -1, -5, 7, 5,
					-- layer=2 filter=231 channel=55
					7, 5, 7, 11, -8, 8, -1, 5, 0,
					-- layer=2 filter=231 channel=56
					-11, -10, -2, -3, -6, -11, -9, -8, 5,
					-- layer=2 filter=231 channel=57
					2, -5, -8, -5, 2, -7, -1, -10, -6,
					-- layer=2 filter=231 channel=58
					-1, -12, -11, -2, -3, -4, 7, -4, -11,
					-- layer=2 filter=231 channel=59
					5, 0, 0, 0, -8, -1, 7, 6, 4,
					-- layer=2 filter=231 channel=60
					7, -1, 1, -12, 5, 4, -11, -1, -9,
					-- layer=2 filter=231 channel=61
					-10, 6, -9, -7, 6, -9, -1, 2, 3,
					-- layer=2 filter=231 channel=62
					-9, -8, 4, -5, 0, 8, -8, -3, -3,
					-- layer=2 filter=231 channel=63
					-9, -10, 1, -11, -9, 6, 5, -9, 0,
					-- layer=2 filter=231 channel=64
					-5, -5, -7, 3, 7, 1, 0, -7, 2,
					-- layer=2 filter=231 channel=65
					-12, 3, 2, 1, 0, -11, -6, -7, -8,
					-- layer=2 filter=231 channel=66
					-9, 0, -4, 2, 9, -5, 2, -11, 1,
					-- layer=2 filter=231 channel=67
					1, 0, -6, -6, 4, -2, -4, -1, -9,
					-- layer=2 filter=231 channel=68
					-1, -5, 1, 0, 1, -1, -7, -7, -7,
					-- layer=2 filter=231 channel=69
					-7, -3, -9, -2, 4, -10, -11, -7, 8,
					-- layer=2 filter=231 channel=70
					-4, 5, 5, -1, -7, 0, 3, -2, -8,
					-- layer=2 filter=231 channel=71
					-7, -11, 3, -5, -1, -13, 7, -2, -6,
					-- layer=2 filter=231 channel=72
					-2, -8, 5, 6, -10, 2, -9, -8, 0,
					-- layer=2 filter=231 channel=73
					3, -2, -6, 6, -10, 8, -9, -8, 8,
					-- layer=2 filter=231 channel=74
					-10, 8, 1, -6, -9, 3, -1, 4, -6,
					-- layer=2 filter=231 channel=75
					-6, 3, -1, -4, 5, 0, 1, -6, 0,
					-- layer=2 filter=231 channel=76
					0, -1, 3, -13, -10, -6, -1, -11, 3,
					-- layer=2 filter=231 channel=77
					2, -7, -9, -5, 7, 0, -1, 7, -10,
					-- layer=2 filter=231 channel=78
					-8, -8, -6, 5, -2, -9, -3, -9, -6,
					-- layer=2 filter=231 channel=79
					-3, 1, -6, -9, 0, -6, -10, -1, 9,
					-- layer=2 filter=231 channel=80
					-11, 0, 4, -10, -2, 8, -4, 0, 4,
					-- layer=2 filter=231 channel=81
					-10, 7, 1, 3, 4, 2, -2, 3, 5,
					-- layer=2 filter=231 channel=82
					5, 8, 2, 7, -5, 1, 6, -9, 1,
					-- layer=2 filter=231 channel=83
					8, -2, 3, -2, 7, 2, 1, 5, -9,
					-- layer=2 filter=231 channel=84
					-10, 6, -3, -9, -7, 2, 0, -4, 0,
					-- layer=2 filter=231 channel=85
					8, 0, -2, 4, -9, -6, -9, -1, -10,
					-- layer=2 filter=231 channel=86
					-7, -4, 0, 0, -4, 2, -9, 10, -10,
					-- layer=2 filter=231 channel=87
					6, 8, -9, 0, -9, 4, 1, -3, -3,
					-- layer=2 filter=231 channel=88
					-12, 3, 7, 2, -5, 4, 5, -12, -3,
					-- layer=2 filter=231 channel=89
					-1, -7, -7, 0, -8, -6, -2, -10, 5,
					-- layer=2 filter=231 channel=90
					6, 6, -3, -6, -5, -4, 9, 5, 0,
					-- layer=2 filter=231 channel=91
					-4, -4, 1, 2, 4, 3, 6, -9, -3,
					-- layer=2 filter=231 channel=92
					-9, 1, -2, -4, 4, 8, 5, 7, -7,
					-- layer=2 filter=231 channel=93
					-2, 8, 8, 1, -3, 5, 5, -11, -9,
					-- layer=2 filter=231 channel=94
					4, -4, -9, -11, -9, -8, 0, 0, -8,
					-- layer=2 filter=231 channel=95
					3, 1, 2, 4, -8, -4, -8, -4, -8,
					-- layer=2 filter=231 channel=96
					-5, -2, -2, -9, 7, 9, -11, -6, -10,
					-- layer=2 filter=231 channel=97
					7, -8, -1, -4, -1, -3, -1, -1, -4,
					-- layer=2 filter=231 channel=98
					0, -9, -12, -9, -12, 1, -1, -5, -2,
					-- layer=2 filter=231 channel=99
					-9, 5, -9, -5, 0, -13, -11, -5, 0,
					-- layer=2 filter=231 channel=100
					0, -1, -11, -13, -14, -6, -9, -2, -7,
					-- layer=2 filter=231 channel=101
					6, -4, -14, 9, 3, -3, 1, 3, -3,
					-- layer=2 filter=231 channel=102
					-10, -4, -10, -2, -3, -11, 3, -5, -5,
					-- layer=2 filter=231 channel=103
					-5, 0, -6, -7, 8, -11, -8, -10, 0,
					-- layer=2 filter=231 channel=104
					5, -8, 0, -2, -5, -1, 6, -4, 6,
					-- layer=2 filter=231 channel=105
					-1, 9, 9, -7, -3, 5, -2, -8, -1,
					-- layer=2 filter=231 channel=106
					5, -14, 5, -10, -3, 1, -13, 1, 3,
					-- layer=2 filter=231 channel=107
					-3, 6, 5, -2, 0, -6, -8, 3, 4,
					-- layer=2 filter=231 channel=108
					4, 0, -5, 5, 4, 0, 3, -7, 2,
					-- layer=2 filter=231 channel=109
					6, -10, -1, -3, -5, -2, -6, 3, -4,
					-- layer=2 filter=231 channel=110
					-9, 3, 3, -6, 8, -7, 1, -3, 6,
					-- layer=2 filter=231 channel=111
					3, -7, 2, 7, 0, -4, -7, 0, 7,
					-- layer=2 filter=231 channel=112
					1, -7, -9, -8, -2, -6, 2, -7, -8,
					-- layer=2 filter=231 channel=113
					0, -10, -3, -9, 2, -5, -7, 0, 4,
					-- layer=2 filter=231 channel=114
					-11, -7, 10, -7, 0, -6, 3, -9, 0,
					-- layer=2 filter=231 channel=115
					8, -7, 2, -8, -7, 8, 10, -10, -7,
					-- layer=2 filter=231 channel=116
					-6, 0, -11, 8, -8, 6, 0, -12, 5,
					-- layer=2 filter=231 channel=117
					-7, -11, -11, -9, 5, -11, -5, 0, -9,
					-- layer=2 filter=231 channel=118
					-4, -11, 4, 1, -3, 2, -4, 7, -1,
					-- layer=2 filter=231 channel=119
					5, 6, -11, -13, -10, -7, -10, 5, -11,
					-- layer=2 filter=231 channel=120
					1, 4, -6, 0, 0, -2, -3, -7, -9,
					-- layer=2 filter=231 channel=121
					-6, -5, 5, -6, 2, -1, 3, 3, -5,
					-- layer=2 filter=231 channel=122
					-8, -4, 0, 4, 8, 9, 9, 7, -10,
					-- layer=2 filter=231 channel=123
					-11, -5, -12, -1, 2, -14, 5, 5, 1,
					-- layer=2 filter=231 channel=124
					2, -11, 0, -1, -8, -11, -7, -6, 4,
					-- layer=2 filter=231 channel=125
					-3, -1, -7, 7, 2, 5, -5, -4, 2,
					-- layer=2 filter=231 channel=126
					0, -6, -2, -10, 0, -10, -1, 1, 3,
					-- layer=2 filter=231 channel=127
					3, -5, -3, -1, -11, -1, -12, -3, 3,
					-- layer=2 filter=232 channel=0
					31, 3, 41, 19, -11, 8, -15, -20, 20,
					-- layer=2 filter=232 channel=1
					-9, 0, -11, 12, -11, -18, 47, -50, -20,
					-- layer=2 filter=232 channel=2
					-8, -6, 0, 9, 7, 7, 0, 12, -11,
					-- layer=2 filter=232 channel=3
					-24, -20, 4, 2, 10, 26, 54, 34, 52,
					-- layer=2 filter=232 channel=4
					-6, -30, -33, -33, -3, -9, -9, -5, -25,
					-- layer=2 filter=232 channel=5
					50, 8, 13, 14, -1, 15, -33, -8, -13,
					-- layer=2 filter=232 channel=6
					-18, -7, 3, 19, -19, 23, -13, -69, 19,
					-- layer=2 filter=232 channel=7
					-57, -35, 0, -4, 5, -4, -31, -37, -48,
					-- layer=2 filter=232 channel=8
					7, -4, 6, 3, -11, 6, -9, 5, -9,
					-- layer=2 filter=232 channel=9
					-32, -21, -24, 10, -2, -17, -7, 12, 31,
					-- layer=2 filter=232 channel=10
					22, 6, 5, -3, -15, -1, 25, 8, 38,
					-- layer=2 filter=232 channel=11
					-38, -17, -5, -20, 25, 23, -15, 5, -2,
					-- layer=2 filter=232 channel=12
					1, 14, -27, 8, -19, -50, 22, -53, -27,
					-- layer=2 filter=232 channel=13
					0, -9, -3, 6, -3, -3, -11, 3, 2,
					-- layer=2 filter=232 channel=14
					-38, -21, -30, -2, 1, -19, 18, -25, -54,
					-- layer=2 filter=232 channel=15
					36, 16, 62, -9, -15, 13, -26, 19, -1,
					-- layer=2 filter=232 channel=16
					-20, -43, -19, 73, 34, -5, 34, 4, 8,
					-- layer=2 filter=232 channel=17
					0, 1, 0, 7, -7, -1, -1, 6, -10,
					-- layer=2 filter=232 channel=18
					-41, -68, 9, -53, 0, 20, 27, 25, 17,
					-- layer=2 filter=232 channel=19
					-17, -18, 4, 6, 17, 4, -5, -9, 0,
					-- layer=2 filter=232 channel=20
					-9, -10, 1, 7, -4, -3, 8, 2, -6,
					-- layer=2 filter=232 channel=21
					-2, 11, 2, 13, 0, 5, -17, -14, 0,
					-- layer=2 filter=232 channel=22
					10, -3, -7, -9, -12, 9, -3, 2, 9,
					-- layer=2 filter=232 channel=23
					30, -77, -12, 50, 36, -30, 24, 18, 26,
					-- layer=2 filter=232 channel=24
					-23, -47, -42, -47, -25, 6, 35, 42, 68,
					-- layer=2 filter=232 channel=25
					-31, -29, -37, -42, -21, 34, 13, 32, 65,
					-- layer=2 filter=232 channel=26
					-6, -10, 1, 0, 5, -6, -8, 10, 2,
					-- layer=2 filter=232 channel=27
					13, 26, 33, 47, 36, 12, -12, -21, -23,
					-- layer=2 filter=232 channel=28
					-20, -52, -11, 3, 28, 0, 28, 1, -7,
					-- layer=2 filter=232 channel=29
					-10, 4, -9, -12, -4, -11, 2, 7, 8,
					-- layer=2 filter=232 channel=30
					25, 2, 5, 22, -56, -49, -13, 49, 11,
					-- layer=2 filter=232 channel=31
					-7, -38, -42, 37, -27, -50, 12, 4, -34,
					-- layer=2 filter=232 channel=32
					-3, -5, 0, -7, -9, 9, -8, 6, -3,
					-- layer=2 filter=232 channel=33
					-14, 12, 50, -3, 35, -5, 19, 41, 4,
					-- layer=2 filter=232 channel=34
					-21, -45, 39, -45, 31, 44, -15, 33, -15,
					-- layer=2 filter=232 channel=35
					-34, -28, -25, -9, 43, 6, 18, 35, 31,
					-- layer=2 filter=232 channel=36
					-6, 4, -5, -5, 6, 13, -7, -15, -6,
					-- layer=2 filter=232 channel=37
					6, 5, 14, -3, 27, 22, -24, -2, -7,
					-- layer=2 filter=232 channel=38
					49, 34, 1, 14, -20, 3, -52, -30, -29,
					-- layer=2 filter=232 channel=39
					16, -36, -34, 39, 24, -18, 18, 22, -9,
					-- layer=2 filter=232 channel=40
					-16, -25, 36, -3, -14, -36, 13, 36, -6,
					-- layer=2 filter=232 channel=41
					-4, -2, 2, 8, 7, 1, 4, 4, 6,
					-- layer=2 filter=232 channel=42
					-30, -26, -20, 37, 3, -62, 33, -2, -47,
					-- layer=2 filter=232 channel=43
					-19, 0, 0, -9, 50, 24, 31, 27, 13,
					-- layer=2 filter=232 channel=44
					-8, 9, -6, 8, -4, 3, 9, -4, -8,
					-- layer=2 filter=232 channel=45
					-20, 18, 24, -5, -5, -38, 60, 41, 1,
					-- layer=2 filter=232 channel=46
					19, 0, 7, 7, -22, 0, -52, -15, -3,
					-- layer=2 filter=232 channel=47
					-40, 31, 38, 19, 30, -18, 6, -47, -17,
					-- layer=2 filter=232 channel=48
					8, 10, -6, -1, -3, 5, -3, -4, 7,
					-- layer=2 filter=232 channel=49
					-21, -46, 24, -38, 1, 23, 48, 32, 20,
					-- layer=2 filter=232 channel=50
					-20, 4, 0, -3, 5, -17, 1, 8, -9,
					-- layer=2 filter=232 channel=51
					6, 6, -4, -31, -6, 27, -20, -21, -2,
					-- layer=2 filter=232 channel=52
					-7, 0, 7, -42, 12, 0, -34, 10, 0,
					-- layer=2 filter=232 channel=53
					-13, -24, 5, -16, -22, 67, 0, 20, 24,
					-- layer=2 filter=232 channel=54
					-39, -31, -22, -7, -14, 29, 7, 8, 6,
					-- layer=2 filter=232 channel=55
					11, -7, -3, -4, 6, 0, -1, -6, 3,
					-- layer=2 filter=232 channel=56
					-16, -7, 11, -33, 15, 28, -5, -2, -5,
					-- layer=2 filter=232 channel=57
					5, 1, 5, 3, 4, -2, 2, 1, 1,
					-- layer=2 filter=232 channel=58
					12, 25, -26, 19, -24, -56, -3, -37, -40,
					-- layer=2 filter=232 channel=59
					13, 19, 7, 49, 17, 1, 26, 1, -11,
					-- layer=2 filter=232 channel=60
					1, 20, -12, 14, -30, 18, -52, -21, -64,
					-- layer=2 filter=232 channel=61
					-13, -12, 20, -7, -16, 15, -15, -58, -1,
					-- layer=2 filter=232 channel=62
					-46, -38, -17, -34, 2, 9, 7, 39, -1,
					-- layer=2 filter=232 channel=63
					32, -40, -25, 43, 19, 4, -32, -2, 26,
					-- layer=2 filter=232 channel=64
					-22, -42, -6, -7, 0, -35, 32, 42, 0,
					-- layer=2 filter=232 channel=65
					18, -33, -31, 0, -45, -3, -3, -33, -10,
					-- layer=2 filter=232 channel=66
					6, -19, -39, -4, -36, -13, -24, -38, -11,
					-- layer=2 filter=232 channel=67
					28, 2, -24, 7, -31, -21, -32, 0, 28,
					-- layer=2 filter=232 channel=68
					0, -11, 9, 7, -7, -9, 0, 8, 0,
					-- layer=2 filter=232 channel=69
					-39, -40, 6, 8, -40, -45, 53, 6, -28,
					-- layer=2 filter=232 channel=70
					-4, 4, 11, 13, 34, 0, -1, -1, -5,
					-- layer=2 filter=232 channel=71
					-32, 4, 18, -11, 46, 16, 7, 21, -10,
					-- layer=2 filter=232 channel=72
					-36, -67, 17, -24, -14, -7, -21, -12, -53,
					-- layer=2 filter=232 channel=73
					21, 42, 58, -16, 4, 43, 25, 5, -1,
					-- layer=2 filter=232 channel=74
					6, 6, -20, -3, -25, -40, -29, -10, 14,
					-- layer=2 filter=232 channel=75
					-59, -87, -60, 29, -14, -49, 61, -10, -73,
					-- layer=2 filter=232 channel=76
					9, -8, 12, -9, -38, 10, -25, -35, 17,
					-- layer=2 filter=232 channel=77
					0, 0, -8, -1, -11, -6, 0, -5, 3,
					-- layer=2 filter=232 channel=78
					-30, -24, -5, -51, -3, 19, -9, 17, 26,
					-- layer=2 filter=232 channel=79
					6, -7, -11, -1, 8, 5, 7, -6, 3,
					-- layer=2 filter=232 channel=80
					-14, -26, -9, 23, 11, -16, 30, 32, -27,
					-- layer=2 filter=232 channel=81
					0, -8, -4, 9, 15, 5, 4, 18, 7,
					-- layer=2 filter=232 channel=82
					-2, 2, 0, -7, -6, -5, 1, -13, 0,
					-- layer=2 filter=232 channel=83
					4, -11, -10, 28, 14, -46, 24, 26, -21,
					-- layer=2 filter=232 channel=84
					-7, -10, 0, -3, -5, -7, -1, -3, 7,
					-- layer=2 filter=232 channel=85
					18, 8, 9, -1, 2, -3, -17, 11, 2,
					-- layer=2 filter=232 channel=86
					2, 8, 1, 1, 9, -11, 11, 0, 3,
					-- layer=2 filter=232 channel=87
					10, 4, 6, -16, 48, 8, 27, 27, 50,
					-- layer=2 filter=232 channel=88
					13, 9, -34, 39, -14, -45, 20, 39, 17,
					-- layer=2 filter=232 channel=89
					-17, 5, -2, 21, 11, -33, 44, -21, -16,
					-- layer=2 filter=232 channel=90
					11, -6, -10, 5, -10, -8, -7, -1, 10,
					-- layer=2 filter=232 channel=91
					5, 29, 0, 31, 23, -51, 36, -1, -52,
					-- layer=2 filter=232 channel=92
					5, 26, -22, 11, -15, -50, 33, -34, -55,
					-- layer=2 filter=232 channel=93
					15, -22, -10, 2, 5, 23, -53, -32, 10,
					-- layer=2 filter=232 channel=94
					-20, -22, 0, 48, -34, 20, -13, -29, -21,
					-- layer=2 filter=232 channel=95
					11, -4, 12, 0, 2, 17, 11, -1, 2,
					-- layer=2 filter=232 channel=96
					18, 6, 8, -21, -16, 15, -14, -18, -2,
					-- layer=2 filter=232 channel=97
					-30, -19, -13, -5, 9, 1, 35, 38, 44,
					-- layer=2 filter=232 channel=98
					-54, 1, 49, 9, 45, 14, 21, -8, -7,
					-- layer=2 filter=232 channel=99
					-12, 14, 22, -7, 22, 1, 24, 5, 28,
					-- layer=2 filter=232 channel=100
					86, 45, -9, 11, -25, -37, -22, 16, -44,
					-- layer=2 filter=232 channel=101
					-56, -48, -34, -55, 10, 6, 0, 19, 50,
					-- layer=2 filter=232 channel=102
					-8, -27, 15, -29, 5, 16, 0, 17, -1,
					-- layer=2 filter=232 channel=103
					7, 32, 18, 66, -20, -69, 33, -20, -46,
					-- layer=2 filter=232 channel=104
					-3, 2, 0, -7, 13, 1, 9, 5, 39,
					-- layer=2 filter=232 channel=105
					-30, 4, -36, 28, -15, -13, 0, -34, 54,
					-- layer=2 filter=232 channel=106
					-32, -15, -18, -32, 0, 27, 9, 9, 72,
					-- layer=2 filter=232 channel=107
					-28, 25, 29, -4, -13, -8, 15, 0, -19,
					-- layer=2 filter=232 channel=108
					0, 17, 12, -10, 12, -9, 7, -13, -26,
					-- layer=2 filter=232 channel=109
					1, 0, 2, 9, -5, -1, -21, 4, -3,
					-- layer=2 filter=232 channel=110
					-40, -40, -41, -16, -15, -34, 7, -30, -22,
					-- layer=2 filter=232 channel=111
					-8, -12, 7, -9, 6, -6, -4, 4, -7,
					-- layer=2 filter=232 channel=112
					-19, -1, 19, -20, -16, 55, 0, 14, 19,
					-- layer=2 filter=232 channel=113
					27, -18, -6, 1, -21, -33, -22, 36, 19,
					-- layer=2 filter=232 channel=114
					10, 5, 18, 8, 15, 5, 4, 4, 10,
					-- layer=2 filter=232 channel=115
					-2, 3, 3, 0, -1, -1, 0, 0, -2,
					-- layer=2 filter=232 channel=116
					61, 18, 26, 4, 48, 8, 35, 35, 25,
					-- layer=2 filter=232 channel=117
					-48, 20, 37, -47, -14, 13, -15, -11, -65,
					-- layer=2 filter=232 channel=118
					-25, -1, 0, -22, 22, 19, 21, 19, 14,
					-- layer=2 filter=232 channel=119
					-29, -66, 5, -8, -49, -41, 60, 31, -11,
					-- layer=2 filter=232 channel=120
					0, 9, 5, -8, -9, 0, -9, 5, 8,
					-- layer=2 filter=232 channel=121
					-9, -6, -3, -4, -6, 4, 10, -2, -1,
					-- layer=2 filter=232 channel=122
					0, 1, -11, -14, 6, 0, 6, 9, -9,
					-- layer=2 filter=232 channel=123
					-27, -32, 13, 12, 15, 0, -46, -6, -25,
					-- layer=2 filter=232 channel=124
					23, 3, -6, -10, -5, -19, -27, -42, -9,
					-- layer=2 filter=232 channel=125
					10, -7, 3, -4, -1, -1, 1, 3, 10,
					-- layer=2 filter=232 channel=126
					-12, 11, 44, -61, -18, -13, -7, 5, 0,
					-- layer=2 filter=232 channel=127
					-3, -27, -18, -4, -3, -26, 37, 19, 25,
					-- layer=2 filter=233 channel=0
					-22, 1, -9, -9, 16, 5, -13, 0, -23,
					-- layer=2 filter=233 channel=1
					0, -4, 39, 3, -15, 6, -18, 13, 20,
					-- layer=2 filter=233 channel=2
					9, -6, 3, 3, -3, -10, 8, 4, -8,
					-- layer=2 filter=233 channel=3
					-2, -30, -36, 11, 8, -18, 0, -23, -12,
					-- layer=2 filter=233 channel=4
					3, -8, 19, 7, -9, 12, -15, -44, -15,
					-- layer=2 filter=233 channel=5
					-29, -30, 9, -5, 20, 18, 0, 27, 21,
					-- layer=2 filter=233 channel=6
					43, 52, 6, 53, 13, 66, 60, 33, 11,
					-- layer=2 filter=233 channel=7
					11, 37, 24, 57, 52, 26, -89, -68, 35,
					-- layer=2 filter=233 channel=8
					3, 10, -6, -9, 9, 0, -1, 3, -5,
					-- layer=2 filter=233 channel=9
					22, -14, 15, 4, 5, 20, 29, 10, -1,
					-- layer=2 filter=233 channel=10
					0, -8, -4, -1, 17, -20, -13, -11, -17,
					-- layer=2 filter=233 channel=11
					-20, -16, -4, -5, -16, -1, 15, -5, 4,
					-- layer=2 filter=233 channel=12
					46, 18, 43, -2, -9, 35, 3, 6, 47,
					-- layer=2 filter=233 channel=13
					9, -1, 0, 10, 3, 11, 0, 6, -6,
					-- layer=2 filter=233 channel=14
					43, 1, 12, 5, -24, -2, 0, -5, 3,
					-- layer=2 filter=233 channel=15
					-15, -26, -12, -6, -6, -25, 24, 23, -31,
					-- layer=2 filter=233 channel=16
					-25, -6, 10, 1, -53, -32, -12, -49, -14,
					-- layer=2 filter=233 channel=17
					0, -6, 8, -6, 3, -8, -9, -9, -3,
					-- layer=2 filter=233 channel=18
					-17, 18, 52, 9, -19, -1, -15, -12, -18,
					-- layer=2 filter=233 channel=19
					-24, 31, 10, 5, -23, -31, -2, -4, -10,
					-- layer=2 filter=233 channel=20
					-5, 0, -7, 2, -2, 3, 5, -8, -3,
					-- layer=2 filter=233 channel=21
					3, 12, 10, 1, 1, -3, 8, -16, -22,
					-- layer=2 filter=233 channel=22
					-8, -9, 8, -5, 2, 2, 4, 1, 3,
					-- layer=2 filter=233 channel=23
					-4, -13, -17, -9, -32, 33, -29, -47, -3,
					-- layer=2 filter=233 channel=24
					11, -4, -18, -4, -6, -19, 3, 7, -2,
					-- layer=2 filter=233 channel=25
					-29, -20, -38, -22, -5, -34, 21, 33, 2,
					-- layer=2 filter=233 channel=26
					-4, 9, 7, -10, 4, 6, -2, 2, -4,
					-- layer=2 filter=233 channel=27
					-14, -27, -8, -20, -9, -23, 33, 30, 27,
					-- layer=2 filter=233 channel=28
					50, 27, 16, 25, 5, -11, -56, -56, -49,
					-- layer=2 filter=233 channel=29
					5, 11, 0, -1, -4, 10, -6, -7, 4,
					-- layer=2 filter=233 channel=30
					-2, 2, 4, -2, 13, 3, -6, 18, -22,
					-- layer=2 filter=233 channel=31
					-27, 4, -64, -4, -37, -30, 18, 4, 43,
					-- layer=2 filter=233 channel=32
					-3, -4, 3, -9, 7, 1, -4, 0, 3,
					-- layer=2 filter=233 channel=33
					11, -31, 25, 25, 25, -15, -11, -33, 29,
					-- layer=2 filter=233 channel=34
					13, 41, 41, 25, 12, -3, -31, -14, -52,
					-- layer=2 filter=233 channel=35
					32, 29, -9, 20, 4, 22, -73, -83, -73,
					-- layer=2 filter=233 channel=36
					4, -3, 11, -6, 9, -2, 0, -4, -6,
					-- layer=2 filter=233 channel=37
					-15, -17, -5, 2, -4, 5, 33, 9, 20,
					-- layer=2 filter=233 channel=38
					-13, -4, -5, 10, 10, -15, 44, 45, 26,
					-- layer=2 filter=233 channel=39
					6, -15, 19, 37, 2, 22, -18, -30, 30,
					-- layer=2 filter=233 channel=40
					-19, -75, -29, 1, -25, 56, 5, -37, -13,
					-- layer=2 filter=233 channel=41
					-5, -1, 8, -1, 0, 4, -6, 6, 7,
					-- layer=2 filter=233 channel=42
					0, -25, 12, -15, 10, 25, -17, -14, 23,
					-- layer=2 filter=233 channel=43
					-53, -1, -19, -8, -7, 4, 10, 4, -18,
					-- layer=2 filter=233 channel=44
					0, 2, -6, -6, 8, 1, -10, 9, -8,
					-- layer=2 filter=233 channel=45
					-43, -67, -58, 4, 18, -26, 31, 55, 82,
					-- layer=2 filter=233 channel=46
					-1, 9, 19, 9, 6, -6, -10, -3, -46,
					-- layer=2 filter=233 channel=47
					1, -14, 17, 45, 6, 3, -50, -24, 24,
					-- layer=2 filter=233 channel=48
					-4, -2, -10, 2, 8, 3, -5, 3, 1,
					-- layer=2 filter=233 channel=49
					-23, -6, 2, 5, -15, -11, -13, -3, -37,
					-- layer=2 filter=233 channel=50
					2, -2, -8, -15, -6, -16, -9, -4, -19,
					-- layer=2 filter=233 channel=51
					-8, -17, 0, -6, -22, 3, -6, -5, -6,
					-- layer=2 filter=233 channel=52
					-71, -22, 39, 22, -8, 30, 1, 9, 1,
					-- layer=2 filter=233 channel=53
					-1, 20, -20, 35, 30, -24, 7, 47, 11,
					-- layer=2 filter=233 channel=54
					-32, -2, -18, -12, 5, 0, -55, -51, 13,
					-- layer=2 filter=233 channel=55
					16, -1, 9, -7, 3, -1, 6, 12, 1,
					-- layer=2 filter=233 channel=56
					-2, 0, 8, 19, -2, -11, 14, 14, 10,
					-- layer=2 filter=233 channel=57
					-11, -7, 7, -4, -9, -2, -3, 13, -2,
					-- layer=2 filter=233 channel=58
					39, 19, 18, -7, 3, 27, 4, 9, 32,
					-- layer=2 filter=233 channel=59
					13, 12, 35, -54, 21, 17, 10, 2, 6,
					-- layer=2 filter=233 channel=60
					-1, 20, 14, -25, -3, -2, -14, -7, -4,
					-- layer=2 filter=233 channel=61
					-10, -21, -37, -69, -4, 0, -53, -11, -6,
					-- layer=2 filter=233 channel=62
					0, 45, 18, -6, 18, -9, -17, 10, -33,
					-- layer=2 filter=233 channel=63
					-18, -5, 10, -12, -1, 5, -30, -22, 18,
					-- layer=2 filter=233 channel=64
					15, -1, 9, 7, 35, 31, -27, -25, 0,
					-- layer=2 filter=233 channel=65
					32, -5, -23, -15, -9, 14, 6, 9, -10,
					-- layer=2 filter=233 channel=66
					5, -7, 20, 7, 16, -13, 2, -35, -55,
					-- layer=2 filter=233 channel=67
					10, 21, 24, -2, -14, 2, 22, 12, 0,
					-- layer=2 filter=233 channel=68
					-5, 2, 2, 7, 12, 0, 6, -7, 9,
					-- layer=2 filter=233 channel=69
					6, -24, -4, 16, -4, 7, -16, -8, -10,
					-- layer=2 filter=233 channel=70
					12, -9, -26, 9, 9, 3, -61, -74, -34,
					-- layer=2 filter=233 channel=71
					17, 6, -36, -33, -32, -20, 24, 34, 26,
					-- layer=2 filter=233 channel=72
					42, 7, 36, 56, 23, -8, -34, -55, -22,
					-- layer=2 filter=233 channel=73
					6, -40, -11, -20, -43, -44, -27, -8, 25,
					-- layer=2 filter=233 channel=74
					8, 11, 24, -5, -6, 22, 4, -12, -1,
					-- layer=2 filter=233 channel=75
					20, 32, -2, 7, -14, 20, -5, -53, -17,
					-- layer=2 filter=233 channel=76
					-38, -44, 3, -27, -1, 0, -34, -30, 38,
					-- layer=2 filter=233 channel=77
					1, -3, -6, 3, 5, -5, -5, -5, 3,
					-- layer=2 filter=233 channel=78
					-15, 4, 16, -12, -17, 20, -23, -22, -12,
					-- layer=2 filter=233 channel=79
					-4, 5, -8, -10, 2, 8, 5, 4, -2,
					-- layer=2 filter=233 channel=80
					10, 1, -3, 18, -30, -25, -8, -55, -18,
					-- layer=2 filter=233 channel=81
					-3, 13, 0, -4, 2, 9, 13, 4, -3,
					-- layer=2 filter=233 channel=82
					-1, -7, 6, -11, -3, 10, -3, 2, 3,
					-- layer=2 filter=233 channel=83
					10, 20, 5, -28, -19, -1, -33, -32, -32,
					-- layer=2 filter=233 channel=84
					11, -8, 0, 7, -8, 0, 4, 8, -5,
					-- layer=2 filter=233 channel=85
					-4, 7, -1, 1, -24, -3, 11, 7, 7,
					-- layer=2 filter=233 channel=86
					-9, -8, 1, -5, -9, 12, 7, -3, -8,
					-- layer=2 filter=233 channel=87
					43, 50, 12, 7, 9, 6, 16, -39, -13,
					-- layer=2 filter=233 channel=88
					1, -5, 18, -7, -10, 28, 1, 11, -10,
					-- layer=2 filter=233 channel=89
					46, 12, 18, 0, -7, 20, -5, -14, -5,
					-- layer=2 filter=233 channel=90
					6, -7, -6, 5, -4, 3, -5, 7, 11,
					-- layer=2 filter=233 channel=91
					40, 26, 36, 13, 24, 2, 9, 4, 22,
					-- layer=2 filter=233 channel=92
					24, 9, 40, -2, 1, 12, 0, 0, 14,
					-- layer=2 filter=233 channel=93
					-29, 7, 18, 3, 18, 32, 21, -2, -22,
					-- layer=2 filter=233 channel=94
					-22, 35, 5, -21, 6, 21, -26, 7, 2,
					-- layer=2 filter=233 channel=95
					2, 5, 11, 4, 5, 1, 18, 7, 18,
					-- layer=2 filter=233 channel=96
					13, 47, 23, -22, 43, 53, -17, 0, 34,
					-- layer=2 filter=233 channel=97
					15, 0, 32, 25, 14, -14, 9, -11, 0,
					-- layer=2 filter=233 channel=98
					26, 6, -22, 28, -14, -6, -107, -128, -60,
					-- layer=2 filter=233 channel=99
					-29, -15, -3, 8, 2, -15, -10, -8, -1,
					-- layer=2 filter=233 channel=100
					14, 26, 21, -41, -9, 7, 2, -2, 0,
					-- layer=2 filter=233 channel=101
					-7, -21, -23, -47, -40, -32, -13, -23, 19,
					-- layer=2 filter=233 channel=102
					5, 29, 9, 7, 19, -1, -35, -8, -17,
					-- layer=2 filter=233 channel=103
					15, 47, 41, 21, 39, 49, 34, -16, 48,
					-- layer=2 filter=233 channel=104
					10, 17, -13, 7, 2, -16, -3, -28, -19,
					-- layer=2 filter=233 channel=105
					-33, -26, 0, -32, 5, 17, 23, -10, 16,
					-- layer=2 filter=233 channel=106
					-17, -3, -11, 3, -17, -58, -11, -21, 7,
					-- layer=2 filter=233 channel=107
					5, -3, 9, 33, 29, 19, 10, 20, 47,
					-- layer=2 filter=233 channel=108
					-12, -7, -23, -16, 6, 16, -1, 33, 24,
					-- layer=2 filter=233 channel=109
					6, 4, 3, -17, -2, 2, 8, 10, 17,
					-- layer=2 filter=233 channel=110
					12, -8, 11, -43, -29, 7, -44, -23, -1,
					-- layer=2 filter=233 channel=111
					6, 4, 1, -2, 3, 0, 4, 7, 3,
					-- layer=2 filter=233 channel=112
					2, -46, -41, -6, -4, 0, 11, 11, 3,
					-- layer=2 filter=233 channel=113
					7, -30, 0, -8, -3, -8, -25, -24, -36,
					-- layer=2 filter=233 channel=114
					-4, -2, 6, -9, 12, 5, 2, 16, 9,
					-- layer=2 filter=233 channel=115
					-1, 4, 5, -12, -11, 8, -12, 5, 2,
					-- layer=2 filter=233 channel=116
					22, 20, -2, 30, -1, -16, 2, -5, -7,
					-- layer=2 filter=233 channel=117
					-16, 33, -7, 38, 31, -22, -59, -71, 13,
					-- layer=2 filter=233 channel=118
					-13, 0, -4, 1, 1, -22, 1, -25, -31,
					-- layer=2 filter=233 channel=119
					-13, -6, 0, -22, -1, 3, -30, 10, -43,
					-- layer=2 filter=233 channel=120
					-8, 2, 6, 7, 2, -5, -8, -2, -4,
					-- layer=2 filter=233 channel=121
					-9, 0, -4, 6, -6, 3, 10, -1, 3,
					-- layer=2 filter=233 channel=122
					5, -1, 6, -4, -3, 7, 3, -12, -1,
					-- layer=2 filter=233 channel=123
					21, 6, 56, 50, 31, 47, -77, -51, 15,
					-- layer=2 filter=233 channel=124
					9, -8, 19, -3, 19, 6, 21, -23, 27,
					-- layer=2 filter=233 channel=125
					-6, 10, -4, 1, 10, 3, 0, 8, 10,
					-- layer=2 filter=233 channel=126
					-13, 31, 56, -37, 29, 9, -3, 6, 22,
					-- layer=2 filter=233 channel=127
					-22, 0, 17, -5, -25, 24, -12, -6, 10,
					-- layer=2 filter=234 channel=0
					-10, 22, -3, 29, 11, -8, 25, 9, 0,
					-- layer=2 filter=234 channel=1
					6, -30, -14, 10, -11, -9, -16, -23, -6,
					-- layer=2 filter=234 channel=2
					-8, -2, -6, 0, 5, 11, -11, 5, -4,
					-- layer=2 filter=234 channel=3
					19, 2, 14, 1, -26, -4, 32, 6, 17,
					-- layer=2 filter=234 channel=4
					-20, -15, -5, -4, -25, -17, -14, -11, -7,
					-- layer=2 filter=234 channel=5
					14, 32, -2, -14, -12, -4, 0, 19, -6,
					-- layer=2 filter=234 channel=6
					-5, 6, -29, 25, 57, 15, 8, 24, -6,
					-- layer=2 filter=234 channel=7
					11, -22, -18, 22, -38, 1, 0, -36, -18,
					-- layer=2 filter=234 channel=8
					-9, 0, -1, 7, 0, 8, -9, 7, 5,
					-- layer=2 filter=234 channel=9
					-20, -10, 30, 13, -13, 23, -11, 0, -13,
					-- layer=2 filter=234 channel=10
					17, 24, 19, 22, 2, -12, 24, -2, 18,
					-- layer=2 filter=234 channel=11
					2, 2, -15, 4, 15, -6, 3, 10, -12,
					-- layer=2 filter=234 channel=12
					10, -14, -18, 14, -38, -22, -5, -24, -35,
					-- layer=2 filter=234 channel=13
					6, 0, -6, 2, 4, 9, 1, 11, -7,
					-- layer=2 filter=234 channel=14
					13, -34, -7, 22, -8, -15, 3, -18, -19,
					-- layer=2 filter=234 channel=15
					1, 34, -14, 40, 19, -10, -13, -10, -51,
					-- layer=2 filter=234 channel=16
					-13, -8, 23, -12, -69, -23, -38, -38, 14,
					-- layer=2 filter=234 channel=17
					-1, -2, 10, -9, 9, 9, -8, 7, -4,
					-- layer=2 filter=234 channel=18
					-5, 41, -34, 1, 36, -51, 0, 29, -2,
					-- layer=2 filter=234 channel=19
					41, 17, 18, 23, 7, 7, 16, 21, 32,
					-- layer=2 filter=234 channel=20
					1, -6, 4, -2, 1, 3, -4, 1, 4,
					-- layer=2 filter=234 channel=21
					8, 15, 1, 8, 2, -4, 7, 3, 13,
					-- layer=2 filter=234 channel=22
					6, -2, 5, -8, -1, -8, -11, -11, 10,
					-- layer=2 filter=234 channel=23
					-44, -16, -4, -15, -2, -21, -20, -5, 4,
					-- layer=2 filter=234 channel=24
					-1, 9, 1, 1, -12, -18, 13, 20, 36,
					-- layer=2 filter=234 channel=25
					-12, -9, -2, -3, -22, -30, 23, -9, 13,
					-- layer=2 filter=234 channel=26
					-3, 9, 5, -6, 4, 0, 1, -6, -11,
					-- layer=2 filter=234 channel=27
					17, -11, 20, 8, 6, 33, 0, 3, 0,
					-- layer=2 filter=234 channel=28
					22, -9, -18, 45, -11, -20, 30, -4, 8,
					-- layer=2 filter=234 channel=29
					0, -3, 11, 11, 7, -2, 0, 8, 11,
					-- layer=2 filter=234 channel=30
					4, -4, 12, -6, -17, -5, -25, -15, -2,
					-- layer=2 filter=234 channel=31
					2, -11, -16, 35, -10, -6, 10, 100, -28,
					-- layer=2 filter=234 channel=32
					5, 5, -8, 11, 13, 0, 9, -6, 6,
					-- layer=2 filter=234 channel=33
					29, -57, -28, 26, -17, 5, 16, -15, -4,
					-- layer=2 filter=234 channel=34
					-24, 17, 14, -15, 24, 36, -45, 18, 19,
					-- layer=2 filter=234 channel=35
					22, -3, -32, 19, -7, 0, 26, -11, 30,
					-- layer=2 filter=234 channel=36
					-7, 6, 1, -6, -4, -10, 9, -4, 9,
					-- layer=2 filter=234 channel=37
					-5, -7, 8, -1, 16, -4, -9, 8, -2,
					-- layer=2 filter=234 channel=38
					7, -13, -3, 9, -4, 1, 8, -8, -9,
					-- layer=2 filter=234 channel=39
					21, -1, 7, -10, 9, 14, -25, -4, -2,
					-- layer=2 filter=234 channel=40
					-16, 8, 2, -3, 5, 13, -22, 1, 62,
					-- layer=2 filter=234 channel=41
					-7, 5, -6, -7, 2, 2, 2, -5, 4,
					-- layer=2 filter=234 channel=42
					4, 9, -3, 13, -18, 28, -1, -17, 12,
					-- layer=2 filter=234 channel=43
					29, 30, -5, -23, 21, -2, 25, 25, 39,
					-- layer=2 filter=234 channel=44
					8, -8, 9, 7, 0, 6, -6, 0, 1,
					-- layer=2 filter=234 channel=45
					24, -36, -2, -3, -48, -4, 39, -15, -11,
					-- layer=2 filter=234 channel=46
					-11, 18, 2, -19, -13, -12, -8, -16, -10,
					-- layer=2 filter=234 channel=47
					20, -60, -38, 27, -23, -21, 15, -18, -15,
					-- layer=2 filter=234 channel=48
					2, -6, -7, -3, 0, 7, -6, -3, -3,
					-- layer=2 filter=234 channel=49
					-13, 34, -10, 24, 19, -43, -43, -12, -25,
					-- layer=2 filter=234 channel=50
					-3, -4, 11, 5, -3, 25, -13, -24, -13,
					-- layer=2 filter=234 channel=51
					-10, -6, -10, 14, 2, 6, 17, 5, 14,
					-- layer=2 filter=234 channel=52
					-1, -18, -32, -6, 13, 8, 3, 14, 19,
					-- layer=2 filter=234 channel=53
					-15, 16, 7, 51, -2, -42, 5, 32, -1,
					-- layer=2 filter=234 channel=54
					-9, -22, -56, 2, -8, 0, 27, 20, 25,
					-- layer=2 filter=234 channel=55
					-10, -2, -4, 9, 4, 3, -5, -2, -12,
					-- layer=2 filter=234 channel=56
					-3, 3, 5, 11, 2, 2, 13, 7, -14,
					-- layer=2 filter=234 channel=57
					-13, 1, -7, 5, 12, 15, -8, -5, 1,
					-- layer=2 filter=234 channel=58
					21, -18, -24, -18, -34, -21, -13, -34, -36,
					-- layer=2 filter=234 channel=59
					12, -22, 0, -24, 21, 37, -3, 16, 30,
					-- layer=2 filter=234 channel=60
					-14, -12, -8, -26, 15, 46, -1, -10, -28,
					-- layer=2 filter=234 channel=61
					-5, 16, 12, 2, 34, 15, 12, -2, 25,
					-- layer=2 filter=234 channel=62
					-43, 7, -54, -31, 30, -3, -55, 27, 0,
					-- layer=2 filter=234 channel=63
					-28, -4, 8, -14, 33, 5, 2, 14, 14,
					-- layer=2 filter=234 channel=64
					-12, -5, 0, 8, 0, 10, -18, -7, 37,
					-- layer=2 filter=234 channel=65
					-16, -28, 13, 2, 34, 42, 5, 32, 7,
					-- layer=2 filter=234 channel=66
					-30, 7, 11, -19, -18, -13, -9, -32, 48,
					-- layer=2 filter=234 channel=67
					-26, 3, 4, -7, 13, 3, -16, -16, -17,
					-- layer=2 filter=234 channel=68
					3, -6, 8, 0, 11, -8, -6, 0, 10,
					-- layer=2 filter=234 channel=69
					-2, -1, -2, 19, 18, 11, -24, -30, 19,
					-- layer=2 filter=234 channel=70
					16, 10, -13, 9, -31, 16, 16, -30, -3,
					-- layer=2 filter=234 channel=71
					0, -5, 6, 6, -25, 23, 2, -11, 1,
					-- layer=2 filter=234 channel=72
					19, -60, -47, 35, -17, 9, 41, -12, -14,
					-- layer=2 filter=234 channel=73
					-43, 3, 15, -3, -14, -21, 3, -34, -24,
					-- layer=2 filter=234 channel=74
					0, 1, -9, 16, 17, -16, 15, -6, 0,
					-- layer=2 filter=234 channel=75
					0, -42, 5, -11, -39, -58, -21, -6, -2,
					-- layer=2 filter=234 channel=76
					-18, -43, 17, 0, 45, 25, 11, 42, 7,
					-- layer=2 filter=234 channel=77
					-3, 7, 0, 4, 3, 12, 11, 5, 7,
					-- layer=2 filter=234 channel=78
					-18, 7, -37, -8, 10, 0, 1, 5, -4,
					-- layer=2 filter=234 channel=79
					9, -8, 1, -4, -6, 5, -3, 9, -5,
					-- layer=2 filter=234 channel=80
					5, 14, 17, 4, -13, 4, -6, -22, 16,
					-- layer=2 filter=234 channel=81
					-11, -2, 2, -3, 3, -2, 0, -7, 8,
					-- layer=2 filter=234 channel=82
					-9, 1, 2, -11, 0, -9, -7, 5, 2,
					-- layer=2 filter=234 channel=83
					-4, -16, -2, 12, -46, 8, -11, -33, 1,
					-- layer=2 filter=234 channel=84
					6, -5, 5, 5, 2, -3, 0, -6, -3,
					-- layer=2 filter=234 channel=85
					3, -12, -2, -16, -5, -5, -2, -6, -3,
					-- layer=2 filter=234 channel=86
					3, 17, 0, -2, 1, -10, 0, -8, -12,
					-- layer=2 filter=234 channel=87
					-23, -10, -45, -16, 74, 24, -29, 33, 4,
					-- layer=2 filter=234 channel=88
					-28, -1, 30, 15, -3, 0, -3, 15, 28,
					-- layer=2 filter=234 channel=89
					4, -25, -31, 6, -2, -7, -2, -7, 5,
					-- layer=2 filter=234 channel=90
					4, -7, 1, 2, -9, 0, 7, 4, 9,
					-- layer=2 filter=234 channel=91
					13, -26, -3, -7, -72, 2, 27, -27, -19,
					-- layer=2 filter=234 channel=92
					1, -38, -29, 6, -30, -11, -21, -28, -26,
					-- layer=2 filter=234 channel=93
					0, -17, -16, 7, 15, -40, -16, 17, -46,
					-- layer=2 filter=234 channel=94
					-34, -41, -3, 8, 29, 0, 8, 7, -9,
					-- layer=2 filter=234 channel=95
					-7, 6, 5, -1, 4, 7, -6, 11, 1,
					-- layer=2 filter=234 channel=96
					-24, -5, 20, 13, 74, 43, -14, 24, 37,
					-- layer=2 filter=234 channel=97
					25, 16, 0, 7, 0, -1, 36, -14, 27,
					-- layer=2 filter=234 channel=98
					11, -37, -27, 28, -18, -2, 15, -17, -8,
					-- layer=2 filter=234 channel=99
					-23, -26, -1, 15, 3, 36, 25, -5, 23,
					-- layer=2 filter=234 channel=100
					1, 2, -10, -26, -28, 43, 14, -17, 0,
					-- layer=2 filter=234 channel=101
					11, 18, 2, -9, -30, -3, -13, -23, -14,
					-- layer=2 filter=234 channel=102
					-46, -10, 13, 9, 31, -5, -32, 40, 1,
					-- layer=2 filter=234 channel=103
					61, 1, -29, -40, -53, -11, 23, -8, -3,
					-- layer=2 filter=234 channel=104
					-20, 16, -25, 58, 24, -15, 9, 25, -46,
					-- layer=2 filter=234 channel=105
					-37, -6, 28, 8, 11, 65, -21, 7, 18,
					-- layer=2 filter=234 channel=106
					19, 0, 9, -4, -28, -10, 29, 9, -13,
					-- layer=2 filter=234 channel=107
					22, 35, 4, 28, -19, 6, -7, -5, -14,
					-- layer=2 filter=234 channel=108
					1, -35, 38, 27, 0, 15, -10, -20, -4,
					-- layer=2 filter=234 channel=109
					-5, -7, 27, -5, -7, 9, -23, 0, 0,
					-- layer=2 filter=234 channel=110
					-41, -33, -9, 11, 3, 28, 1, 11, 61,
					-- layer=2 filter=234 channel=111
					8, -12, 2, -5, 5, 7, -8, 0, 9,
					-- layer=2 filter=234 channel=112
					21, 22, 0, 13, 0, 2, 17, 16, 5,
					-- layer=2 filter=234 channel=113
					6, 11, 31, 27, -15, -1, -16, -2, -3,
					-- layer=2 filter=234 channel=114
					-4, 1, 7, 1, 12, 17, 3, -6, 14,
					-- layer=2 filter=234 channel=115
					2, -7, -2, 5, 1, -1, 12, -11, 7,
					-- layer=2 filter=234 channel=116
					-32, 3, -10, -19, 46, 15, -37, 1, -13,
					-- layer=2 filter=234 channel=117
					4, -22, -49, 7, -28, -14, 29, -32, -5,
					-- layer=2 filter=234 channel=118
					-1, 11, 13, 2, 9, 3, 9, 16, 23,
					-- layer=2 filter=234 channel=119
					13, 9, -30, -5, 10, -8, -11, -1, 47,
					-- layer=2 filter=234 channel=120
					-9, 3, 0, -10, 0, 0, -3, 7, -5,
					-- layer=2 filter=234 channel=121
					-2, 9, -4, -9, -5, -6, 2, 1, -7,
					-- layer=2 filter=234 channel=122
					-9, 9, 1, 7, 8, 12, 6, 13, 14,
					-- layer=2 filter=234 channel=123
					-4, -28, -32, 28, 5, 3, -6, -5, 9,
					-- layer=2 filter=234 channel=124
					9, -20, -63, 34, -20, -6, -2, -3, -26,
					-- layer=2 filter=234 channel=125
					9, -7, -8, -4, 7, 6, 9, 4, 4,
					-- layer=2 filter=234 channel=126
					-6, -25, -22, 16, 34, -25, 0, 24, 9,
					-- layer=2 filter=234 channel=127
					-10, -28, 10, -13, -25, -22, -38, 4, -3,
					-- layer=2 filter=235 channel=0
					-8, 4, 11, -1, 3, -3, 23, -7, -22,
					-- layer=2 filter=235 channel=1
					10, -6, -25, -9, -11, -5, -16, -25, 12,
					-- layer=2 filter=235 channel=2
					-2, 5, 0, -5, 8, 8, -8, -4, 0,
					-- layer=2 filter=235 channel=3
					-33, 11, 20, 14, -6, 3, 20, 2, 0,
					-- layer=2 filter=235 channel=4
					-1, -5, -17, 14, 16, 18, 24, 43, 10,
					-- layer=2 filter=235 channel=5
					32, 17, 13, 20, 9, -4, 0, 2, -34,
					-- layer=2 filter=235 channel=6
					18, 6, -3, 8, 18, 39, 7, 4, 9,
					-- layer=2 filter=235 channel=7
					22, 39, 30, 22, -5, 0, -25, -46, -26,
					-- layer=2 filter=235 channel=8
					10, 7, 6, -7, 0, 1, 4, -3, 5,
					-- layer=2 filter=235 channel=9
					-10, 17, 9, -34, 5, 0, 2, -6, 4,
					-- layer=2 filter=235 channel=10
					-18, -5, 9, 1, 18, -8, 38, -8, -1,
					-- layer=2 filter=235 channel=11
					45, 1, -11, 6, 13, -8, -7, 0, -12,
					-- layer=2 filter=235 channel=12
					37, 2, -42, -50, -12, 5, -42, -14, 3,
					-- layer=2 filter=235 channel=13
					0, -6, 5, 8, 3, 0, -6, -9, 4,
					-- layer=2 filter=235 channel=14
					15, -10, -17, -52, -19, 5, -48, -33, 2,
					-- layer=2 filter=235 channel=15
					-24, 18, -26, 14, -13, -10, -66, -26, -16,
					-- layer=2 filter=235 channel=16
					-12, -21, 3, 21, 3, 6, -12, 3, 2,
					-- layer=2 filter=235 channel=17
					-6, -2, 3, 0, -8, 1, 6, -8, 4,
					-- layer=2 filter=235 channel=18
					-5, 41, -9, 20, 27, -13, -32, 17, 14,
					-- layer=2 filter=235 channel=19
					10, 2, -49, 31, 28, 17, -14, -25, 43,
					-- layer=2 filter=235 channel=20
					-2, -1, 6, -4, 8, -3, -6, 0, 10,
					-- layer=2 filter=235 channel=21
					21, 19, 12, 16, 0, 3, 9, 8, 0,
					-- layer=2 filter=235 channel=22
					3, 5, -5, -7, 3, -3, 1, -2, -4,
					-- layer=2 filter=235 channel=23
					-13, -30, -9, 4, 5, 18, -33, 2, 13,
					-- layer=2 filter=235 channel=24
					-35, 6, 30, -31, -6, 14, 0, 9, 33,
					-- layer=2 filter=235 channel=25
					-5, -1, 0, -42, -39, 21, 6, 13, 57,
					-- layer=2 filter=235 channel=26
					3, -2, -10, -9, -2, 0, -2, 1, -3,
					-- layer=2 filter=235 channel=27
					-10, 30, 21, 15, 5, 5, 22, -32, -16,
					-- layer=2 filter=235 channel=28
					-8, -18, -26, -18, -6, -13, 2, -22, 1,
					-- layer=2 filter=235 channel=29
					1, 4, -6, 2, -8, 9, 1, -4, -5,
					-- layer=2 filter=235 channel=30
					-34, -6, -25, 5, -7, 25, 7, 9, 17,
					-- layer=2 filter=235 channel=31
					-34, -43, 40, -2, -10, 61, -65, 92, -7,
					-- layer=2 filter=235 channel=32
					6, -5, 0, 3, 0, 1, -5, 7, 0,
					-- layer=2 filter=235 channel=33
					-19, -20, 2, -27, -24, 13, -16, -27, 0,
					-- layer=2 filter=235 channel=34
					36, 28, 31, 33, 10, 27, 4, -4, 10,
					-- layer=2 filter=235 channel=35
					27, 5, 7, 33, 16, 21, 25, 10, 14,
					-- layer=2 filter=235 channel=36
					0, 4, 4, -8, -11, -10, -6, -5, 5,
					-- layer=2 filter=235 channel=37
					26, 4, -2, 6, 0, 5, -15, -17, -15,
					-- layer=2 filter=235 channel=38
					2, 4, -5, 5, -18, -1, 8, -19, -4,
					-- layer=2 filter=235 channel=39
					-59, -41, -13, -10, 6, 36, 0, -1, 4,
					-- layer=2 filter=235 channel=40
					4, -49, -52, -14, 6, 19, -22, 35, 81,
					-- layer=2 filter=235 channel=41
					9, 0, 8, -4, -7, 8, -11, -2, 2,
					-- layer=2 filter=235 channel=42
					-19, -48, -4, -9, -6, 16, -34, 27, 26,
					-- layer=2 filter=235 channel=43
					29, 44, -14, 25, 21, -36, -5, -6, -22,
					-- layer=2 filter=235 channel=44
					1, 3, -2, -1, 5, 10, 7, -4, -9,
					-- layer=2 filter=235 channel=45
					-75, -16, 3, -7, -48, 11, 39, 2, -4,
					-- layer=2 filter=235 channel=46
					-4, 5, -11, -2, -3, -7, 17, 3, -4,
					-- layer=2 filter=235 channel=47
					-30, -73, -62, -39, -55, 9, -28, -21, -32,
					-- layer=2 filter=235 channel=48
					0, -8, 0, 1, 0, 4, -6, -4, 6,
					-- layer=2 filter=235 channel=49
					-2, 32, -20, 3, 41, -7, -50, -2, 13,
					-- layer=2 filter=235 channel=50
					1, 14, -15, -2, -7, -10, -14, -17, 3,
					-- layer=2 filter=235 channel=51
					22, 13, 0, -15, -24, 10, -30, -18, -23,
					-- layer=2 filter=235 channel=52
					29, 20, -18, 19, -3, 10, 1, -31, 6,
					-- layer=2 filter=235 channel=53
					10, 12, -35, 0, -1, 0, -50, 24, 68,
					-- layer=2 filter=235 channel=54
					16, -8, -29, 0, 13, 5, 9, 16, 1,
					-- layer=2 filter=235 channel=55
					2, -10, 4, -7, -15, 0, 11, 0, 0,
					-- layer=2 filter=235 channel=56
					38, 7, -3, 9, 9, -15, -20, -34, -8,
					-- layer=2 filter=235 channel=57
					-5, 14, 3, 2, 14, 3, 5, 1, 0,
					-- layer=2 filter=235 channel=58
					56, -4, -6, -27, 4, 0, -16, -3, -17,
					-- layer=2 filter=235 channel=59
					34, 34, 1, -2, 35, 1, 16, 6, 31,
					-- layer=2 filter=235 channel=60
					45, 12, -26, 25, -1, 12, -16, -3, -20,
					-- layer=2 filter=235 channel=61
					3, 16, 0, 10, -8, 6, 16, -1, -31,
					-- layer=2 filter=235 channel=62
					-6, -3, -30, -17, 26, 8, -14, -12, 18,
					-- layer=2 filter=235 channel=63
					-30, -63, -15, 9, 11, 7, 6, 38, 38,
					-- layer=2 filter=235 channel=64
					-55, -30, -25, -11, -15, 25, -8, 0, 31,
					-- layer=2 filter=235 channel=65
					2, -6, -19, -9, 8, 35, 23, 23, 0,
					-- layer=2 filter=235 channel=66
					21, -8, 72, 0, 19, -28, 16, -27, -33,
					-- layer=2 filter=235 channel=67
					-5, -8, 6, -32, -18, -22, 14, -21, -40,
					-- layer=2 filter=235 channel=68
					-10, -3, 1, 8, 0, 7, 6, 10, 8,
					-- layer=2 filter=235 channel=69
					-32, -31, -21, -21, -24, 18, -8, 3, 18,
					-- layer=2 filter=235 channel=70
					17, 7, -13, 24, 23, 14, 21, -9, 4,
					-- layer=2 filter=235 channel=71
					-22, 1, -16, 8, 3, 0, 3, -21, -13,
					-- layer=2 filter=235 channel=72
					-29, -1, -14, 27, -3, -16, -48, -17, -28,
					-- layer=2 filter=235 channel=73
					-31, 21, 56, -7, -46, -9, 7, 5, -27,
					-- layer=2 filter=235 channel=74
					-13, 3, -2, -16, 2, -5, 23, 0, 0,
					-- layer=2 filter=235 channel=75
					0, -43, -36, -90, -38, 0, -54, -46, -3,
					-- layer=2 filter=235 channel=76
					-23, -34, -11, -9, 13, 19, -34, 8, 49,
					-- layer=2 filter=235 channel=77
					6, 10, -6, 3, 4, 10, -4, -4, 9,
					-- layer=2 filter=235 channel=78
					34, 9, -11, 6, -4, -11, -24, -2, -2,
					-- layer=2 filter=235 channel=79
					0, 0, 3, 1, 11, 1, 6, 2, -3,
					-- layer=2 filter=235 channel=80
					6, -25, 19, 11, 9, 14, 20, 22, 4,
					-- layer=2 filter=235 channel=81
					-26, -11, -23, -20, -9, -13, -3, -5, -10,
					-- layer=2 filter=235 channel=82
					5, 5, 11, 1, -8, 2, 8, 4, -9,
					-- layer=2 filter=235 channel=83
					-10, -30, -14, -9, 20, 30, 5, 13, 37,
					-- layer=2 filter=235 channel=84
					10, 2, 0, 5, -10, -8, 7, -2, -6,
					-- layer=2 filter=235 channel=85
					1, 16, -13, -14, -6, 1, 1, -1, 0,
					-- layer=2 filter=235 channel=86
					-3, 9, 0, -18, -8, -8, -10, -14, 5,
					-- layer=2 filter=235 channel=87
					35, 34, -52, 1, 38, 9, -30, 25, 7,
					-- layer=2 filter=235 channel=88
					-17, -28, -38, -18, -43, 5, 9, 26, 46,
					-- layer=2 filter=235 channel=89
					23, -15, -36, -31, 11, -3, -49, -33, 16,
					-- layer=2 filter=235 channel=90
					6, 8, -2, 0, 0, 0, 2, -1, 8,
					-- layer=2 filter=235 channel=91
					17, -19, -15, -20, -5, -32, -20, -19, -18,
					-- layer=2 filter=235 channel=92
					20, -13, -33, -10, 0, -8, -38, -16, 0,
					-- layer=2 filter=235 channel=93
					58, -11, -66, -24, -37, -6, 10, -32, -31,
					-- layer=2 filter=235 channel=94
					-3, -4, -8, 34, 21, 24, -7, -5, 5,
					-- layer=2 filter=235 channel=95
					2, 3, -4, 5, -2, -3, -7, 7, -1,
					-- layer=2 filter=235 channel=96
					33, -17, -24, 9, 12, 30, -36, 19, 47,
					-- layer=2 filter=235 channel=97
					-14, -8, 9, 1, -9, 35, 6, -11, 0,
					-- layer=2 filter=235 channel=98
					11, -14, -30, 4, -28, 9, 9, -19, -17,
					-- layer=2 filter=235 channel=99
					18, -20, -38, -15, -6, -6, -16, -7, -2,
					-- layer=2 filter=235 channel=100
					-1, -11, 8, -1, 19, 27, 12, 21, 19,
					-- layer=2 filter=235 channel=101
					34, 28, -6, 1, -15, 17, -8, 5, 26,
					-- layer=2 filter=235 channel=102
					1, 25, -29, 26, 29, 25, -36, -10, 25,
					-- layer=2 filter=235 channel=103
					43, -5, 57, 13, 20, -12, -3, 7, -1,
					-- layer=2 filter=235 channel=104
					0, 23, -44, 19, 12, 29, -39, 7, 26,
					-- layer=2 filter=235 channel=105
					-5, -64, 34, -6, 43, 22, 6, 53, 47,
					-- layer=2 filter=235 channel=106
					26, 12, 24, -33, -5, 3, 18, -7, 18,
					-- layer=2 filter=235 channel=107
					30, -46, 55, -15, 45, 23, -19, 22, 50,
					-- layer=2 filter=235 channel=108
					-15, 8, -18, 5, 20, 13, -36, -36, 15,
					-- layer=2 filter=235 channel=109
					-5, 4, 13, -5, 4, 9, -13, 0, 3,
					-- layer=2 filter=235 channel=110
					-18, -45, -15, -23, -17, 24, -17, -22, 49,
					-- layer=2 filter=235 channel=111
					-6, 2, -1, -8, 9, -6, -6, 5, -4,
					-- layer=2 filter=235 channel=112
					24, 10, 15, 1, -8, 6, 0, -22, -39,
					-- layer=2 filter=235 channel=113
					-26, -34, 15, -11, -31, 14, 6, 23, 4,
					-- layer=2 filter=235 channel=114
					1, 20, 6, 6, 10, 8, 7, 9, 4,
					-- layer=2 filter=235 channel=115
					-3, 6, -11, 10, 5, 9, -5, 2, 8,
					-- layer=2 filter=235 channel=116
					5, 27, -19, 22, 23, -23, -20, -6, 10,
					-- layer=2 filter=235 channel=117
					15, 47, 0, -21, -45, -21, -38, -76, -78,
					-- layer=2 filter=235 channel=118
					-24, 22, 0, 19, 18, -15, 16, 4, -14,
					-- layer=2 filter=235 channel=119
					1, -10, -6, 7, 0, -6, 27, 20, 13,
					-- layer=2 filter=235 channel=120
					-2, -8, -7, 0, 2, -9, 5, 9, -7,
					-- layer=2 filter=235 channel=121
					6, 0, -1, 11, 8, 7, -2, 1, 4,
					-- layer=2 filter=235 channel=122
					12, -5, 4, 17, -2, 3, 2, -9, 0,
					-- layer=2 filter=235 channel=123
					9, -16, -24, -5, -11, -21, -16, -21, -33,
					-- layer=2 filter=235 channel=124
					4, 1, -25, -30, 25, 10, -85, -23, -24,
					-- layer=2 filter=235 channel=125
					-14, 5, -6, 2, -6, -7, -2, 0, 14,
					-- layer=2 filter=235 channel=126
					27, -30, 4, -5, -47, -18, -20, -22, 0,
					-- layer=2 filter=235 channel=127
					-14, -23, -21, -27, 5, 0, 8, 5, 47,
					-- layer=2 filter=236 channel=0
					15, 6, 3, 11, -7, 2, -1, 9, -6,
					-- layer=2 filter=236 channel=1
					-16, 6, -7, -23, -18, -23, 17, 0, 14,
					-- layer=2 filter=236 channel=2
					0, 3, 7, -10, -3, 9, -11, 8, 0,
					-- layer=2 filter=236 channel=3
					-11, 5, 16, 17, -18, -12, 8, -17, -6,
					-- layer=2 filter=236 channel=4
					-13, 26, 9, -10, -17, -12, 9, -21, 18,
					-- layer=2 filter=236 channel=5
					15, 11, -3, 0, -22, 8, 10, -3, -21,
					-- layer=2 filter=236 channel=6
					19, 6, 6, 45, 59, 36, 50, 41, 50,
					-- layer=2 filter=236 channel=7
					12, -12, 8, -13, 0, 20, -2, -9, 0,
					-- layer=2 filter=236 channel=8
					7, 9, -5, 8, -1, 0, -5, 0, 5,
					-- layer=2 filter=236 channel=9
					-4, 24, 0, 6, -32, -13, 7, -4, 6,
					-- layer=2 filter=236 channel=10
					26, 21, 16, 31, 3, -5, -4, -15, -13,
					-- layer=2 filter=236 channel=11
					-7, -3, -5, -15, -6, -17, 1, 6, 2,
					-- layer=2 filter=236 channel=12
					-16, 6, -6, -32, -21, -50, 7, -5, 0,
					-- layer=2 filter=236 channel=13
					10, -9, 10, -4, 0, 1, 5, -5, 6,
					-- layer=2 filter=236 channel=14
					-6, 0, -7, -23, -35, -33, 11, -6, 29,
					-- layer=2 filter=236 channel=15
					-15, -32, 14, -2, -56, -7, -22, 14, 6,
					-- layer=2 filter=236 channel=16
					30, 33, 71, -16, -44, 46, -35, -11, -18,
					-- layer=2 filter=236 channel=17
					-1, 0, 6, -10, 5, 1, 4, 0, -7,
					-- layer=2 filter=236 channel=18
					-6, 15, -45, -28, -5, -23, -36, -30, -2,
					-- layer=2 filter=236 channel=19
					3, 7, 2, 32, 34, 0, 28, -4, 1,
					-- layer=2 filter=236 channel=20
					0, 7, -9, 10, -7, 7, 9, 2, 7,
					-- layer=2 filter=236 channel=21
					9, 9, 4, 1, 12, 18, 0, -1, 29,
					-- layer=2 filter=236 channel=22
					-8, 6, 2, 11, 3, 8, -5, -7, -6,
					-- layer=2 filter=236 channel=23
					-23, 8, 15, -17, -16, 34, -33, -30, -14,
					-- layer=2 filter=236 channel=24
					-14, 11, 35, -7, -9, 23, -3, -4, 27,
					-- layer=2 filter=236 channel=25
					3, -2, 20, 1, -18, -5, 23, 13, 34,
					-- layer=2 filter=236 channel=26
					-4, -3, -7, 8, 0, -2, -7, -6, 0,
					-- layer=2 filter=236 channel=27
					12, 3, -10, 37, -1, 1, 13, -14, -12,
					-- layer=2 filter=236 channel=28
					27, 19, -7, 13, -2, 11, -14, -26, 3,
					-- layer=2 filter=236 channel=29
					-3, -1, 5, -2, -4, -5, -5, -6, 8,
					-- layer=2 filter=236 channel=30
					-28, 10, 1, -12, -42, -12, -2, -41, -18,
					-- layer=2 filter=236 channel=31
					-69, -26, 63, 9, 23, -26, 19, 34, 27,
					-- layer=2 filter=236 channel=32
					6, 0, 4, -10, 3, -2, 3, 8, 11,
					-- layer=2 filter=236 channel=33
					23, -37, -6, -6, -2, 27, 29, 5, 58,
					-- layer=2 filter=236 channel=34
					22, 1, -21, -9, 45, 8, -41, -15, 22,
					-- layer=2 filter=236 channel=35
					18, -2, -6, 20, 28, 10, -19, -26, -13,
					-- layer=2 filter=236 channel=36
					3, 9, 16, -14, -7, -1, 2, 1, 17,
					-- layer=2 filter=236 channel=37
					-5, -20, -9, 15, -13, -1, 5, -9, -3,
					-- layer=2 filter=236 channel=38
					12, 6, 16, 25, -14, -5, 23, -16, -17,
					-- layer=2 filter=236 channel=39
					5, -35, 13, -25, -39, 3, -43, -16, -26,
					-- layer=2 filter=236 channel=40
					25, -45, -27, -19, 41, 37, -47, 21, 26,
					-- layer=2 filter=236 channel=41
					-2, -4, -12, 3, -10, -8, -10, 10, 9,
					-- layer=2 filter=236 channel=42
					-10, 37, 22, -6, -46, 37, -13, 4, -13,
					-- layer=2 filter=236 channel=43
					0, 21, -9, 16, -18, 3, 0, -2, 13,
					-- layer=2 filter=236 channel=44
					11, -2, -8, 9, 6, -4, 0, 9, 8,
					-- layer=2 filter=236 channel=45
					-2, 3, 9, 8, -25, -6, -2, -15, -17,
					-- layer=2 filter=236 channel=46
					-24, -27, -18, 25, -18, -11, -25, -12, 5,
					-- layer=2 filter=236 channel=47
					16, -3, -21, -5, -10, -1, -17, -50, -4,
					-- layer=2 filter=236 channel=48
					0, -8, 4, 10, 6, -9, 7, 0, 7,
					-- layer=2 filter=236 channel=49
					-2, 29, 6, -31, 0, 28, -52, -13, -3,
					-- layer=2 filter=236 channel=50
					-3, 16, -6, 6, 3, 11, -5, 2, 0,
					-- layer=2 filter=236 channel=51
					0, -11, -11, -1, -9, 0, -2, 4, 0,
					-- layer=2 filter=236 channel=52
					-23, -12, -23, -13, 2, -42, -1, -1, 29,
					-- layer=2 filter=236 channel=53
					-48, 15, -19, 5, -44, -11, 27, -9, 48,
					-- layer=2 filter=236 channel=54
					-19, -24, -40, 1, 5, 20, -10, 12, -2,
					-- layer=2 filter=236 channel=55
					-3, -6, 5, -3, -10, -14, 5, 10, -8,
					-- layer=2 filter=236 channel=56
					-7, 18, 3, -20, -14, 0, -2, 7, 8,
					-- layer=2 filter=236 channel=57
					7, 2, 1, 8, -5, 4, -4, -7, 3,
					-- layer=2 filter=236 channel=58
					-14, 4, 13, -15, -17, -37, 5, -8, -2,
					-- layer=2 filter=236 channel=59
					-14, -14, -30, 43, -3, -35, 0, 23, 7,
					-- layer=2 filter=236 channel=60
					14, -30, -8, 6, -17, -15, -12, -14, -31,
					-- layer=2 filter=236 channel=61
					-19, -1, -6, 6, -15, -58, -15, -44, -47,
					-- layer=2 filter=236 channel=62
					8, 0, -2, 0, 62, 8, 5, 11, 0,
					-- layer=2 filter=236 channel=63
					-18, -32, 6, 2, 0, -1, 2, -18, -9,
					-- layer=2 filter=236 channel=64
					-39, -11, 32, -12, -30, 49, 0, -18, 3,
					-- layer=2 filter=236 channel=65
					-4, -28, 20, 9, 22, -28, 18, 27, -17,
					-- layer=2 filter=236 channel=66
					28, -16, 0, -17, -33, 17, -2, 26, 0,
					-- layer=2 filter=236 channel=67
					7, 16, -9, 28, -17, -9, 26, -26, -7,
					-- layer=2 filter=236 channel=68
					-4, -5, -4, 7, -8, 5, -8, 1, 4,
					-- layer=2 filter=236 channel=69
					-26, 24, 34, -16, -18, 25, -1, -16, 4,
					-- layer=2 filter=236 channel=70
					23, 12, 2, 14, 7, 11, 2, 4, -12,
					-- layer=2 filter=236 channel=71
					-3, 14, 0, 27, -4, 1, 3, -36, -5,
					-- layer=2 filter=236 channel=72
					15, -32, -40, 0, 7, 25, -8, -9, 8,
					-- layer=2 filter=236 channel=73
					10, 48, 74, 1, 19, 44, -7, -29, 30,
					-- layer=2 filter=236 channel=74
					-1, 1, -13, 20, -6, -20, 28, -3, -19,
					-- layer=2 filter=236 channel=75
					17, 14, 5, 4, -3, -11, 28, 14, 40,
					-- layer=2 filter=236 channel=76
					-4, -33, 19, 24, -4, -19, 36, -23, 10,
					-- layer=2 filter=236 channel=77
					10, 8, 0, -2, 0, 6, 0, -2, 4,
					-- layer=2 filter=236 channel=78
					-22, -4, -23, -4, -6, -24, -1, 19, 3,
					-- layer=2 filter=236 channel=79
					0, -7, -7, 11, 6, -8, 0, 4, 2,
					-- layer=2 filter=236 channel=80
					-4, -1, 9, -18, -27, -9, -10, -34, -12,
					-- layer=2 filter=236 channel=81
					1, -6, -1, 3, 10, -5, 2, -6, 5,
					-- layer=2 filter=236 channel=82
					9, 10, -3, -8, -10, 8, -7, -3, -5,
					-- layer=2 filter=236 channel=83
					-36, 16, -13, 12, -8, 23, 13, -26, 0,
					-- layer=2 filter=236 channel=84
					-9, 0, -7, 2, 5, -11, 2, -6, -5,
					-- layer=2 filter=236 channel=85
					-3, -2, 6, 8, 0, -5, -3, 12, 5,
					-- layer=2 filter=236 channel=86
					2, -3, -7, -12, 0, -2, -19, -21, -5,
					-- layer=2 filter=236 channel=87
					-10, -14, -47, -3, 0, -37, -8, -22, 1,
					-- layer=2 filter=236 channel=88
					-24, -25, 4, 8, -13, -9, 19, 1, 3,
					-- layer=2 filter=236 channel=89
					6, 0, -14, 1, 15, -22, 17, -9, 21,
					-- layer=2 filter=236 channel=90
					-4, -6, 9, 0, 5, -7, 2, 2, 0,
					-- layer=2 filter=236 channel=91
					21, -12, 1, 33, 14, -25, 39, 11, 0,
					-- layer=2 filter=236 channel=92
					12, 9, -2, -14, -12, -28, 24, -5, 6,
					-- layer=2 filter=236 channel=93
					8, -16, 29, -11, -2, 43, -34, -33, -4,
					-- layer=2 filter=236 channel=94
					-10, 22, -14, 27, -3, -11, -8, -23, -32,
					-- layer=2 filter=236 channel=95
					-8, 7, -4, 0, 3, -6, 3, -9, 6,
					-- layer=2 filter=236 channel=96
					41, 37, 33, 42, 90, 20, 52, 55, 51,
					-- layer=2 filter=236 channel=97
					-6, 23, 15, -7, -35, -5, 28, -14, 33,
					-- layer=2 filter=236 channel=98
					17, 1, 0, 4, 16, 22, -25, -24, 1,
					-- layer=2 filter=236 channel=99
					-17, 12, -4, 32, 13, -11, 25, -10, 10,
					-- layer=2 filter=236 channel=100
					12, 0, -3, 46, -15, -14, 4, -42, -58,
					-- layer=2 filter=236 channel=101
					-2, -17, 4, 6, -15, -12, -1, -13, 0,
					-- layer=2 filter=236 channel=102
					-12, 0, 4, -52, 24, -12, -11, -7, 17,
					-- layer=2 filter=236 channel=103
					26, 19, 0, -4, -21, -11, 23, 38, 36,
					-- layer=2 filter=236 channel=104
					-16, 9, -12, 9, 1, 28, -15, 1, 15,
					-- layer=2 filter=236 channel=105
					13, 7, -23, 29, -33, 22, -41, -34, -4,
					-- layer=2 filter=236 channel=106
					10, -9, 24, -12, -25, -23, 37, -7, 27,
					-- layer=2 filter=236 channel=107
					0, 26, -23, -10, -4, 12, 12, -7, -21,
					-- layer=2 filter=236 channel=108
					5, 13, 17, -3, -14, -18, 2, -24, 13,
					-- layer=2 filter=236 channel=109
					3, 6, 23, -12, 0, -1, -9, 3, 0,
					-- layer=2 filter=236 channel=110
					-5, -3, 28, -10, 6, 41, 5, -5, 8,
					-- layer=2 filter=236 channel=111
					9, 13, -4, -13, -5, -8, 1, -7, -8,
					-- layer=2 filter=236 channel=112
					-14, 8, 2, 8, -44, 1, -10, 19, -4,
					-- layer=2 filter=236 channel=113
					-25, -39, 26, -16, -27, -20, -47, -18, -36,
					-- layer=2 filter=236 channel=114
					-4, 20, 1, 2, 2, 2, 10, 11, 8,
					-- layer=2 filter=236 channel=115
					-4, 1, -9, 7, 7, 5, 4, -8, 6,
					-- layer=2 filter=236 channel=116
					-7, 1, -28, -30, -10, -44, -26, -31, 24,
					-- layer=2 filter=236 channel=117
					-8, -24, -17, -18, 10, -6, -14, -11, 36,
					-- layer=2 filter=236 channel=118
					13, 34, 15, 35, 28, 1, 8, 20, 25,
					-- layer=2 filter=236 channel=119
					15, 39, 21, -16, 2, 7, -1, -26, 22,
					-- layer=2 filter=236 channel=120
					-3, 6, -2, -5, -4, 8, 7, -2, -4,
					-- layer=2 filter=236 channel=121
					-2, 6, -6, 6, -6, -6, -5, 8, 3,
					-- layer=2 filter=236 channel=122
					-2, -5, -1, 0, 8, 11, 10, 0, -3,
					-- layer=2 filter=236 channel=123
					-4, -45, -26, 1, -18, 8, -6, -27, 37,
					-- layer=2 filter=236 channel=124
					-30, -37, -29, -5, -19, 1, 18, 18, -1,
					-- layer=2 filter=236 channel=125
					3, -6, -1, 8, -5, -2, -7, -7, -3,
					-- layer=2 filter=236 channel=126
					4, -4, 22, -5, -18, -75, -16, -87, -26,
					-- layer=2 filter=236 channel=127
					-25, -28, -4, -25, -15, -36, 17, 3, -3,
					-- layer=2 filter=237 channel=0
					7, -30, -22, -35, -6, -16, -14, 11, -10,
					-- layer=2 filter=237 channel=1
					-6, -11, -8, -9, -9, 13, 4, -49, -33,
					-- layer=2 filter=237 channel=2
					-5, 1, -10, -3, -7, -11, -2, -4, 6,
					-- layer=2 filter=237 channel=3
					-28, -27, -31, 16, -4, 9, -4, -20, -36,
					-- layer=2 filter=237 channel=4
					20, -20, -35, 1, 4, -20, 24, 20, 15,
					-- layer=2 filter=237 channel=5
					-3, 6, 26, -47, -10, -12, -7, -11, -22,
					-- layer=2 filter=237 channel=6
					2, 9, -8, -15, 2, -7, 10, 34, 44,
					-- layer=2 filter=237 channel=7
					14, 0, 9, -3, 9, 6, -5, -6, 0,
					-- layer=2 filter=237 channel=8
					8, -6, -8, 6, -1, 0, 0, -5, 4,
					-- layer=2 filter=237 channel=9
					-5, -12, 11, -17, -28, -11, 5, 22, 39,
					-- layer=2 filter=237 channel=10
					-10, -39, -40, -3, 2, -3, 3, -2, -13,
					-- layer=2 filter=237 channel=11
					-9, 32, 10, -10, -16, 8, -11, -10, -25,
					-- layer=2 filter=237 channel=12
					17, 27, -21, -32, -14, -26, -28, -22, 2,
					-- layer=2 filter=237 channel=13
					6, -6, -3, -1, -8, -1, -2, 1, 3,
					-- layer=2 filter=237 channel=14
					-4, 33, 12, -42, -12, -24, -6, -57, -28,
					-- layer=2 filter=237 channel=15
					-4, 17, -9, 25, -27, 22, -52, -4, -12,
					-- layer=2 filter=237 channel=16
					24, -51, -22, 30, 20, -15, 28, 31, 9,
					-- layer=2 filter=237 channel=17
					-9, 1, -7, -7, -2, 5, -4, -5, -9,
					-- layer=2 filter=237 channel=18
					11, 38, 10, 8, 5, 25, 15, 5, 12,
					-- layer=2 filter=237 channel=19
					-31, 3, -27, 8, 22, 49, -26, -13, -8,
					-- layer=2 filter=237 channel=20
					6, 0, 2, 5, -5, -5, 2, -2, 3,
					-- layer=2 filter=237 channel=21
					0, -3, -6, 20, 0, -1, 1, -16, -1,
					-- layer=2 filter=237 channel=22
					4, -8, -9, -7, 16, 8, 0, -3, 3,
					-- layer=2 filter=237 channel=23
					35, -14, -27, 27, 27, 10, -5, 28, 24,
					-- layer=2 filter=237 channel=24
					30, -21, -13, 18, -45, -37, 12, -4, -56,
					-- layer=2 filter=237 channel=25
					14, -2, 5, 18, -40, -20, 36, -23, -68,
					-- layer=2 filter=237 channel=26
					7, -1, -2, -2, -10, -4, 4, -7, 6,
					-- layer=2 filter=237 channel=27
					2, -13, -5, 24, 11, 23, 10, -20, 27,
					-- layer=2 filter=237 channel=28
					6, 49, -15, 10, 4, -7, -16, -27, -8,
					-- layer=2 filter=237 channel=29
					-4, -10, 0, 0, 7, 4, 8, -1, 0,
					-- layer=2 filter=237 channel=30
					29, -42, -30, 22, 6, 28, 46, 17, 9,
					-- layer=2 filter=237 channel=31
					28, 22, -21, 20, -32, -4, -33, 38, 38,
					-- layer=2 filter=237 channel=32
					7, 1, 7, -8, -3, 12, -2, 0, 3,
					-- layer=2 filter=237 channel=33
					6, -15, 26, 20, 6, -6, 9, -20, -23,
					-- layer=2 filter=237 channel=34
					-29, 56, -1, -4, 10, 20, 26, -14, 8,
					-- layer=2 filter=237 channel=35
					-36, 31, 11, 3, 22, -15, -28, -23, 12,
					-- layer=2 filter=237 channel=36
					13, 1, 2, -12, -11, 4, -7, 0, -12,
					-- layer=2 filter=237 channel=37
					-8, 10, 8, -12, -11, 4, 7, 0, -6,
					-- layer=2 filter=237 channel=38
					-4, 27, 47, 2, 9, 7, -12, -9, -1,
					-- layer=2 filter=237 channel=39
					44, -40, -25, -2, 25, -12, 28, 4, -1,
					-- layer=2 filter=237 channel=40
					-23, -1, -43, 16, -17, -31, 30, -12, 17,
					-- layer=2 filter=237 channel=41
					6, -4, 5, 10, -7, -8, -3, -3, -9,
					-- layer=2 filter=237 channel=42
					13, -24, -39, 13, 31, 15, -9, 31, -9,
					-- layer=2 filter=237 channel=43
					-33, -4, -57, -31, -10, -18, 19, -28, 0,
					-- layer=2 filter=237 channel=44
					1, -3, 0, -7, -9, 6, 3, 4, -3,
					-- layer=2 filter=237 channel=45
					-6, -12, -50, 64, -26, -24, 1, -12, -22,
					-- layer=2 filter=237 channel=46
					9, -34, -11, 14, 6, 0, 44, 4, 16,
					-- layer=2 filter=237 channel=47
					-1, 2, -35, -1, -25, -32, 12, -1, 1,
					-- layer=2 filter=237 channel=48
					0, 0, 6, -6, 2, 6, 0, -3, -8,
					-- layer=2 filter=237 channel=49
					4, 30, -18, -15, 11, 2, 16, 21, 53,
					-- layer=2 filter=237 channel=50
					-2, -8, -13, -10, 6, -11, 2, 13, -12,
					-- layer=2 filter=237 channel=51
					2, -7, 36, -27, 3, 1, -17, -12, -5,
					-- layer=2 filter=237 channel=52
					-3, 5, 23, -18, -26, -7, -29, -29, 18,
					-- layer=2 filter=237 channel=53
					65, -2, -36, 5, 4, 15, 22, -16, -29,
					-- layer=2 filter=237 channel=54
					-29, 0, -16, -34, -26, -20, -37, -6, -32,
					-- layer=2 filter=237 channel=55
					14, -4, 1, 10, 2, -4, 5, 7, 0,
					-- layer=2 filter=237 channel=56
					-2, 31, 0, -15, -23, -3, 0, -2, -12,
					-- layer=2 filter=237 channel=57
					-3, 1, -5, -12, 5, -1, -1, 5, 3,
					-- layer=2 filter=237 channel=58
					20, 54, 2, -32, -14, -21, -47, -24, 17,
					-- layer=2 filter=237 channel=59
					36, 54, 34, 10, -25, -5, -30, -13, 11,
					-- layer=2 filter=237 channel=60
					11, 43, 32, -18, 15, 32, -57, -20, -16,
					-- layer=2 filter=237 channel=61
					-4, 26, 21, 0, 10, 3, -26, 41, 42,
					-- layer=2 filter=237 channel=62
					-13, 19, 2, -37, -2, -12, -11, 3, 12,
					-- layer=2 filter=237 channel=63
					20, -31, -53, 12, -1, -4, 9, 30, 4,
					-- layer=2 filter=237 channel=64
					16, -30, -31, 29, 8, 6, 32, 21, 28,
					-- layer=2 filter=237 channel=65
					12, 31, 60, -4, -9, 2, 6, 57, 44,
					-- layer=2 filter=237 channel=66
					28, -7, 9, 10, -10, -49, -3, -7, -22,
					-- layer=2 filter=237 channel=67
					17, -31, 15, 14, -3, -34, 26, 31, 11,
					-- layer=2 filter=237 channel=68
					-7, -4, -9, 6, -7, -6, 9, -4, 6,
					-- layer=2 filter=237 channel=69
					-2, -28, -42, 13, 23, -14, 30, 23, 9,
					-- layer=2 filter=237 channel=70
					1, 31, -12, 19, 22, -33, -23, -20, 4,
					-- layer=2 filter=237 channel=71
					26, 34, 11, 1, -7, 17, 34, -15, -6,
					-- layer=2 filter=237 channel=72
					-19, 4, 0, 4, 68, 11, -45, -18, -62,
					-- layer=2 filter=237 channel=73
					-2, 30, -22, 32, 14, 36, 61, 31, 30,
					-- layer=2 filter=237 channel=74
					-4, -8, -12, 4, 19, -11, 25, 26, 7,
					-- layer=2 filter=237 channel=75
					-3, -1, -30, -38, -15, -14, -65, -87, -50,
					-- layer=2 filter=237 channel=76
					-29, 15, 0, 16, -30, 62, 11, 14, 32,
					-- layer=2 filter=237 channel=77
					1, 4, 8, -8, 7, 7, -5, 0, -2,
					-- layer=2 filter=237 channel=78
					-14, 14, -12, -30, -29, -3, -7, -13, 0,
					-- layer=2 filter=237 channel=79
					5, -1, 9, 1, -1, 3, 5, -9, 0,
					-- layer=2 filter=237 channel=80
					11, -41, -54, 1, 8, -5, 34, 37, 19,
					-- layer=2 filter=237 channel=81
					5, -6, -4, -2, -15, -2, 1, 1, -3,
					-- layer=2 filter=237 channel=82
					1, 1, 6, -1, 7, 0, -3, 10, -3,
					-- layer=2 filter=237 channel=83
					13, -7, -68, 66, 18, -16, 18, -9, 22,
					-- layer=2 filter=237 channel=84
					6, 6, 7, 6, -4, -8, -1, -7, -10,
					-- layer=2 filter=237 channel=85
					15, -13, -1, -1, -4, -11, -6, -7, 5,
					-- layer=2 filter=237 channel=86
					14, 15, 8, 13, -6, 1, 12, 12, 0,
					-- layer=2 filter=237 channel=87
					80, 45, -2, 36, 8, 53, -20, 5, 5,
					-- layer=2 filter=237 channel=88
					36, -34, -50, 52, -8, -6, 4, 4, 29,
					-- layer=2 filter=237 channel=89
					0, 34, 3, -25, -8, -16, -14, -31, -38,
					-- layer=2 filter=237 channel=90
					-4, -5, 5, 1, 0, 0, 1, -5, -1,
					-- layer=2 filter=237 channel=91
					-14, 16, -19, -72, -11, -31, -57, -16, -35,
					-- layer=2 filter=237 channel=92
					0, 4, -20, -38, 24, -11, -7, -9, -19,
					-- layer=2 filter=237 channel=93
					-35, -16, -23, -46, -40, -5, 2, -18, -1,
					-- layer=2 filter=237 channel=94
					11, -6, -10, 22, 30, 14, -6, 48, 13,
					-- layer=2 filter=237 channel=95
					9, 3, -4, 13, -4, 0, 10, 6, -5,
					-- layer=2 filter=237 channel=96
					29, 8, 0, 15, 5, 23, -6, 2, -5,
					-- layer=2 filter=237 channel=97
					12, -11, -3, 4, 22, -6, 15, 46, 14,
					-- layer=2 filter=237 channel=98
					-34, -18, -7, -3, 11, -23, -12, 8, 11,
					-- layer=2 filter=237 channel=99
					4, -1, 53, 2, -32, 41, -30, -22, -19,
					-- layer=2 filter=237 channel=100
					-8, 0, -31, 27, 1, -15, -9, -2, -21,
					-- layer=2 filter=237 channel=101
					9, 4, 33, -44, -12, 19, 42, -39, -61,
					-- layer=2 filter=237 channel=102
					4, 7, 16, 22, -16, 38, 4, -7, 58,
					-- layer=2 filter=237 channel=103
					-27, -38, -30, -33, -25, 2, 17, 19, -33,
					-- layer=2 filter=237 channel=104
					-1, 16, -57, 27, 27, 30, 7, 11, 6,
					-- layer=2 filter=237 channel=105
					20, -42, 35, -15, -15, 19, -2, -13, 30,
					-- layer=2 filter=237 channel=106
					58, 25, 24, 2, -53, -70, 3, -47, -79,
					-- layer=2 filter=237 channel=107
					1, -57, -18, 32, -20, -35, -18, -9, -51,
					-- layer=2 filter=237 channel=108
					19, -6, -4, 15, -23, 8, 4, -67, -29,
					-- layer=2 filter=237 channel=109
					18, -17, -3, 15, 7, 0, -3, 0, -8,
					-- layer=2 filter=237 channel=110
					43, -7, -24, 32, 16, -21, -12, -9, -15,
					-- layer=2 filter=237 channel=111
					0, 0, 0, 3, 6, 2, 8, -4, -9,
					-- layer=2 filter=237 channel=112
					-44, -8, 26, -26, 15, 3, -14, 30, 33,
					-- layer=2 filter=237 channel=113
					2, -26, -8, 8, 32, 24, 25, 3, 20,
					-- layer=2 filter=237 channel=114
					-21, -13, -2, -9, -14, -23, -4, -1, 5,
					-- layer=2 filter=237 channel=115
					2, 1, 8, -1, -10, 4, 9, -7, -4,
					-- layer=2 filter=237 channel=116
					43, 57, -16, 35, 43, 49, -14, -2, 34,
					-- layer=2 filter=237 channel=117
					-41, -43, -50, 15, -15, 26, -19, -1, -39,
					-- layer=2 filter=237 channel=118
					-6, 1, -18, -18, -30, 4, 6, 11, 13,
					-- layer=2 filter=237 channel=119
					6, 4, -36, 24, 3, -5, 31, 6, -12,
					-- layer=2 filter=237 channel=120
					-3, -1, 2, -6, 0, 0, 1, -8, -6,
					-- layer=2 filter=237 channel=121
					-5, -11, -2, 3, 8, 2, 0, -11, 8,
					-- layer=2 filter=237 channel=122
					-9, 6, -9, -14, 5, 5, 3, 1, -10,
					-- layer=2 filter=237 channel=123
					-7, -19, 3, -18, 10, -10, -21, 23, -16,
					-- layer=2 filter=237 channel=124
					20, -18, -10, 15, -56, -22, -24, 31, -49,
					-- layer=2 filter=237 channel=125
					-5, -9, 2, -5, 0, 8, 6, 0, -2,
					-- layer=2 filter=237 channel=126
					17, 1, 15, -13, 14, 19, 58, -12, -37,
					-- layer=2 filter=237 channel=127
					41, 5, -11, 45, -8, 18, 23, -14, 0,
					-- layer=2 filter=238 channel=0
					24, -14, -35, 14, 4, -24, 8, -5, -15,
					-- layer=2 filter=238 channel=1
					-19, -1, 14, 23, 11, -24, -14, -1, -26,
					-- layer=2 filter=238 channel=2
					1, 1, -11, 0, 4, 9, 0, -11, -12,
					-- layer=2 filter=238 channel=3
					7, -13, 16, 23, 18, -20, -12, -11, 1,
					-- layer=2 filter=238 channel=4
					16, -12, 16, -53, -6, -17, -54, -50, 17,
					-- layer=2 filter=238 channel=5
					24, -9, -6, 16, 18, -21, 24, 30, -27,
					-- layer=2 filter=238 channel=6
					-57, -30, -5, -36, -47, -39, 17, -53, -17,
					-- layer=2 filter=238 channel=7
					-23, -7, -10, -8, 11, -21, -21, -20, 35,
					-- layer=2 filter=238 channel=8
					-7, 7, 1, -11, 10, 4, -6, -4, 5,
					-- layer=2 filter=238 channel=9
					3, 11, -14, -17, -6, 8, -30, -28, 38,
					-- layer=2 filter=238 channel=10
					20, 11, -2, 22, 10, -16, 3, -16, 8,
					-- layer=2 filter=238 channel=11
					2, 2, -3, 29, 30, -7, 22, 1, -31,
					-- layer=2 filter=238 channel=12
					-23, 28, 35, -9, -41, -7, -25, 18, -32,
					-- layer=2 filter=238 channel=13
					9, -11, -5, 0, 1, 1, -1, 10, -9,
					-- layer=2 filter=238 channel=14
					7, 0, -6, 15, 10, -17, -9, 0, -17,
					-- layer=2 filter=238 channel=15
					-40, 26, 45, 19, 44, -5, 16, 2, 8,
					-- layer=2 filter=238 channel=16
					15, 1, 7, -4, -22, 22, -62, -1, 46,
					-- layer=2 filter=238 channel=17
					-6, 3, 6, -1, -5, -4, -8, 4, 7,
					-- layer=2 filter=238 channel=18
					0, 23, 37, -37, 40, 20, 6, 31, 21,
					-- layer=2 filter=238 channel=19
					4, -1, -7, -25, 9, -21, -69, -20, -27,
					-- layer=2 filter=238 channel=20
					-3, 2, 0, 10, 6, 6, -11, 0, 4,
					-- layer=2 filter=238 channel=21
					-5, 10, 0, 1, 3, 1, 6, 3, -5,
					-- layer=2 filter=238 channel=22
					-3, 0, 3, 0, -9, 11, -2, 5, -1,
					-- layer=2 filter=238 channel=23
					-5, 6, 12, -23, -19, 24, -28, -41, 31,
					-- layer=2 filter=238 channel=24
					8, 3, 6, 13, -13, -20, 13, -21, 4,
					-- layer=2 filter=238 channel=25
					5, 11, -12, 28, -2, -30, 23, -23, -31,
					-- layer=2 filter=238 channel=26
					4, -4, -4, 8, -9, 9, 7, 7, -6,
					-- layer=2 filter=238 channel=27
					-6, 6, -4, 11, 11, -56, -17, 7, -37,
					-- layer=2 filter=238 channel=28
					44, 5, 0, -15, 27, -11, 21, -20, 17,
					-- layer=2 filter=238 channel=29
					-8, -5, -10, -4, 0, 0, 7, 4, 4,
					-- layer=2 filter=238 channel=30
					-18, 1, -18, -3, -34, -13, -21, -29, 7,
					-- layer=2 filter=238 channel=31
					-19, -17, -21, -26, 13, 4, -50, -52, -105,
					-- layer=2 filter=238 channel=32
					2, 7, -6, -4, 2, -8, 0, 7, -6,
					-- layer=2 filter=238 channel=33
					-7, 11, 12, 50, 46, -35, 7, -36, -4,
					-- layer=2 filter=238 channel=34
					-61, -56, 17, -53, 66, -1, 62, 64, -42,
					-- layer=2 filter=238 channel=35
					-16, -18, 8, -12, 38, 29, 17, 11, -8,
					-- layer=2 filter=238 channel=36
					5, -3, 4, 3, -1, 4, -5, -10, -11,
					-- layer=2 filter=238 channel=37
					1, -9, 2, 15, 32, -5, 25, 14, -22,
					-- layer=2 filter=238 channel=38
					-5, -5, -27, 32, -13, -14, -24, -11, -68,
					-- layer=2 filter=238 channel=39
					11, -8, -1, 3, -3, 53, -34, -7, 66,
					-- layer=2 filter=238 channel=40
					-64, -28, 60, -32, 42, 0, -16, 36, -22,
					-- layer=2 filter=238 channel=41
					4, -9, 12, 4, -8, -6, -3, -6, -13,
					-- layer=2 filter=238 channel=42
					29, -5, 15, -3, -8, 30, -22, 0, 47,
					-- layer=2 filter=238 channel=43
					-16, 3, 30, -7, 66, 17, -25, 21, 0,
					-- layer=2 filter=238 channel=44
					7, -4, -7, -4, 6, 11, 1, -9, -9,
					-- layer=2 filter=238 channel=45
					-7, 10, -29, 6, 19, -4, -17, -19, -11,
					-- layer=2 filter=238 channel=46
					10, -11, -11, 29, -27, 20, -12, -25, 1,
					-- layer=2 filter=238 channel=47
					63, 9, -8, -4, 41, -15, 1, -28, -3,
					-- layer=2 filter=238 channel=48
					6, 3, 11, 4, -1, -2, -9, -4, -4,
					-- layer=2 filter=238 channel=49
					10, 0, 4, -25, 21, 21, -7, 10, 35,
					-- layer=2 filter=238 channel=50
					5, 1, 30, -22, 9, -6, -21, 0, -13,
					-- layer=2 filter=238 channel=51
					21, -23, -27, 30, 22, -26, 34, 7, -25,
					-- layer=2 filter=238 channel=52
					4, -10, -34, 15, 12, -27, 22, 10, -34,
					-- layer=2 filter=238 channel=53
					-3, -51, -6, 49, -28, -32, -13, -32, -18,
					-- layer=2 filter=238 channel=54
					2, -6, -15, 1, 16, -4, 16, -23, -38,
					-- layer=2 filter=238 channel=55
					-7, 5, 13, 7, -3, 2, 9, 1, 10,
					-- layer=2 filter=238 channel=56
					-3, -3, -3, 21, 32, 13, 21, 20, -2,
					-- layer=2 filter=238 channel=57
					-11, -10, -5, 3, 17, 3, 7, 15, 9,
					-- layer=2 filter=238 channel=58
					-16, 12, 28, 1, -19, -20, -18, 36, -24,
					-- layer=2 filter=238 channel=59
					0, 12, 27, 59, 70, -27, -20, 27, 15,
					-- layer=2 filter=238 channel=60
					22, 39, -3, 42, 60, 18, 18, 70, -8,
					-- layer=2 filter=238 channel=61
					8, -3, -51, 25, 27, -15, 21, 22, 39,
					-- layer=2 filter=238 channel=62
					-45, -19, 12, -16, -10, -8, 7, -15, -11,
					-- layer=2 filter=238 channel=63
					0, -8, 11, -20, -13, 0, -29, -41, 16,
					-- layer=2 filter=238 channel=64
					0, 9, 3, -26, -21, 19, -41, -30, 38,
					-- layer=2 filter=238 channel=65
					-38, -17, -21, -9, -35, -22, 3, 6, 14,
					-- layer=2 filter=238 channel=66
					68, -35, -7, 15, -5, 23, 46, 15, 77,
					-- layer=2 filter=238 channel=67
					3, 18, -26, 49, -27, -4, -2, -35, 6,
					-- layer=2 filter=238 channel=68
					0, -11, 8, 4, -2, -3, -8, -12, 0,
					-- layer=2 filter=238 channel=69
					-5, -16, 14, 1, 2, 28, -43, -17, 65,
					-- layer=2 filter=238 channel=70
					-9, -30, -3, -12, 26, 15, 19, 2, -4,
					-- layer=2 filter=238 channel=71
					5, 18, -2, 35, 13, -58, -10, 10, -28,
					-- layer=2 filter=238 channel=72
					-8, -29, -20, 0, 25, -23, -16, -33, 36,
					-- layer=2 filter=238 channel=73
					1, -30, -21, 18, 10, 18, 1, 5, 35,
					-- layer=2 filter=238 channel=74
					-22, 12, 0, 18, -19, -3, -48, -11, -13,
					-- layer=2 filter=238 channel=75
					-22, -22, -36, -68, -22, 25, -41, -34, 33,
					-- layer=2 filter=238 channel=76
					-49, -25, 17, -5, -19, -21, -15, -31, -19,
					-- layer=2 filter=238 channel=77
					1, -11, 3, 0, 3, -5, 10, -6, -5,
					-- layer=2 filter=238 channel=78
					-11, -3, -9, 5, 4, -16, 29, -3, -18,
					-- layer=2 filter=238 channel=79
					-2, -2, 5, 8, 3, 6, -1, 4, -6,
					-- layer=2 filter=238 channel=80
					14, -1, -4, -19, -17, 24, -64, -13, 49,
					-- layer=2 filter=238 channel=81
					4, 15, 2, -1, 0, 16, 10, 17, 1,
					-- layer=2 filter=238 channel=82
					11, 1, -3, -5, 3, -16, 0, 3, 2,
					-- layer=2 filter=238 channel=83
					0, -4, -19, -34, -39, -11, -74, -43, 8,
					-- layer=2 filter=238 channel=84
					4, -11, -8, -7, -4, -5, -10, -3, 8,
					-- layer=2 filter=238 channel=85
					-3, -5, 8, 1, -4, -8, 6, 15, -17,
					-- layer=2 filter=238 channel=86
					-8, 11, 13, 0, 23, -3, -5, 1, 0,
					-- layer=2 filter=238 channel=87
					-103, 51, 59, 33, 57, 19, 42, 4, 11,
					-- layer=2 filter=238 channel=88
					-23, 16, -3, 7, -27, 8, -14, -19, 5,
					-- layer=2 filter=238 channel=89
					-2, 3, 18, 24, 20, -37, -11, 24, -11,
					-- layer=2 filter=238 channel=90
					4, -8, -5, -1, 5, -8, -10, 1, 0,
					-- layer=2 filter=238 channel=91
					-14, 2, 33, -40, -19, 10, -1, 45, 7,
					-- layer=2 filter=238 channel=92
					-13, 2, 16, 15, 17, -5, 2, 30, -10,
					-- layer=2 filter=238 channel=93
					-58, -6, 7, -79, -68, -39, -36, -5, 4,
					-- layer=2 filter=238 channel=94
					-31, -51, -42, 8, 1, 17, -32, -37, 4,
					-- layer=2 filter=238 channel=95
					-15, 7, -5, -12, -23, -11, -12, -21, -8,
					-- layer=2 filter=238 channel=96
					-33, -64, -65, -26, -65, -64, -23, -36, -60,
					-- layer=2 filter=238 channel=97
					11, -2, 15, 11, -5, 15, -41, -41, 19,
					-- layer=2 filter=238 channel=98
					14, 1, 14, -3, 26, -1, 21, 0, 13,
					-- layer=2 filter=238 channel=99
					-2, 17, -10, 15, 7, -10, 25, 38, -12,
					-- layer=2 filter=238 channel=100
					-17, 18, -20, -12, -2, 14, -42, -10, -28,
					-- layer=2 filter=238 channel=101
					8, 14, 0, 25, 14, -24, 11, -5, -36,
					-- layer=2 filter=238 channel=102
					-14, -23, 8, -62, -21, 0, -30, 6, 10,
					-- layer=2 filter=238 channel=103
					-19, -18, 41, -55, -49, 3, -2, -18, -44,
					-- layer=2 filter=238 channel=104
					-20, 3, 6, 26, 1, 6, 1, -28, 3,
					-- layer=2 filter=238 channel=105
					-15, 23, 1, 17, 6, -4, 15, -27, 29,
					-- layer=2 filter=238 channel=106
					10, 17, 4, 30, -17, -38, 26, -8, -41,
					-- layer=2 filter=238 channel=107
					-45, -51, -20, 24, -17, 44, -30, -50, -19,
					-- layer=2 filter=238 channel=108
					-3, -1, -24, -59, -10, -67, -37, -15, -32,
					-- layer=2 filter=238 channel=109
					4, 0, -4, 1, 16, -14, -18, -4, -16,
					-- layer=2 filter=238 channel=110
					13, -4, 0, -30, -24, 7, -32, -20, 1,
					-- layer=2 filter=238 channel=111
					2, 2, -4, 4, -9, 0, -9, -3, -3,
					-- layer=2 filter=238 channel=112
					35, 19, -48, 37, 12, -15, 24, -6, -31,
					-- layer=2 filter=238 channel=113
					-3, -8, -14, -22, -55, 0, -28, -5, 26,
					-- layer=2 filter=238 channel=114
					0, 1, -1, 9, 4, -21, -22, -13, -10,
					-- layer=2 filter=238 channel=115
					6, 8, -5, -4, -5, 11, -2, 7, 2,
					-- layer=2 filter=238 channel=116
					-57, 16, 16, 7, 30, -17, 18, 28, -17,
					-- layer=2 filter=238 channel=117
					6, -15, 6, -5, 15, 17, -6, -46, 22,
					-- layer=2 filter=238 channel=118
					-5, -14, 33, -19, 17, 11, -13, 17, 23,
					-- layer=2 filter=238 channel=119
					-2, -4, 7, -34, 23, 40, -38, -15, 16,
					-- layer=2 filter=238 channel=120
					5, -4, -4, -3, 10, -8, 6, 4, 10,
					-- layer=2 filter=238 channel=121
					-8, -1, -3, -5, 8, -3, 7, 11, 1,
					-- layer=2 filter=238 channel=122
					-3, 4, 0, 12, -8, -8, 0, 1, -14,
					-- layer=2 filter=238 channel=123
					-27, -14, 3, 10, 10, -18, -8, -5, 28,
					-- layer=2 filter=238 channel=124
					-43, 18, 45, 34, 3, 12, 4, -37, 20,
					-- layer=2 filter=238 channel=125
					7, -11, -4, 5, -7, -7, 4, 0, 0,
					-- layer=2 filter=238 channel=126
					23, 2, 3, -1, 59, 59, -58, 30, 52,
					-- layer=2 filter=238 channel=127
					-20, -28, 6, -8, -7, 21, -34, -7, 24,
					-- layer=2 filter=239 channel=0
					-3, 1, -9, 23, -9, 23, 17, -2, 8,
					-- layer=2 filter=239 channel=1
					-29, -17, -18, -11, -30, -38, -37, 42, -20,
					-- layer=2 filter=239 channel=2
					3, 0, 5, -6, 5, -1, 9, -3, -3,
					-- layer=2 filter=239 channel=3
					-7, 19, -34, -20, -29, 7, -19, -44, -20,
					-- layer=2 filter=239 channel=4
					17, -19, 8, -8, 28, 3, 31, 14, 39,
					-- layer=2 filter=239 channel=5
					-13, -22, -3, 5, 6, 19, 15, 5, -2,
					-- layer=2 filter=239 channel=6
					-3, 36, 6, 21, 32, 15, 72, 67, 56,
					-- layer=2 filter=239 channel=7
					-14, 6, -7, -28, -42, -17, 21, -23, 13,
					-- layer=2 filter=239 channel=8
					0, -1, 0, 3, 0, -11, -5, 4, -3,
					-- layer=2 filter=239 channel=9
					-15, -15, -5, -19, 12, -20, -5, -2, 13,
					-- layer=2 filter=239 channel=10
					15, 10, -12, -4, 1, 4, 0, 1, 19,
					-- layer=2 filter=239 channel=11
					-17, -15, 0, 9, -4, 14, 13, 12, 24,
					-- layer=2 filter=239 channel=12
					-39, -30, -28, -20, -32, -56, -15, -22, -19,
					-- layer=2 filter=239 channel=13
					-6, -3, 3, -6, -2, -8, 4, -11, 5,
					-- layer=2 filter=239 channel=14
					-53, -48, -49, -3, -3, -49, -17, 14, -12,
					-- layer=2 filter=239 channel=15
					3, -39, -29, 48, 10, -17, -10, -86, -12,
					-- layer=2 filter=239 channel=16
					-7, 13, 7, 9, -2, 3, -7, -25, 5,
					-- layer=2 filter=239 channel=17
					-8, 8, 6, -9, 0, -1, 0, 8, 3,
					-- layer=2 filter=239 channel=18
					-5, -35, 7, 5, 4, 13, -14, -25, -8,
					-- layer=2 filter=239 channel=19
					-16, 19, -6, 31, 28, 16, -52, 18, -8,
					-- layer=2 filter=239 channel=20
					0, -8, -7, -4, 0, 5, -3, -11, 4,
					-- layer=2 filter=239 channel=21
					-2, 8, -1, 0, -9, -12, -18, -4, -25,
					-- layer=2 filter=239 channel=22
					1, -5, 0, -6, -6, 10, 0, 0, 1,
					-- layer=2 filter=239 channel=23
					15, 10, -2, -3, -7, 0, 27, 18, 44,
					-- layer=2 filter=239 channel=24
					4, 3, -28, -11, -41, 29, -37, -25, 1,
					-- layer=2 filter=239 channel=25
					-23, -9, -4, -23, -13, -6, -52, -52, -26,
					-- layer=2 filter=239 channel=26
					3, 5, -4, 8, 8, -2, -4, 3, 4,
					-- layer=2 filter=239 channel=27
					-29, -13, 10, 3, 0, 0, 10, 22, 7,
					-- layer=2 filter=239 channel=28
					-7, 40, -17, 21, 21, -8, 39, 9, 14,
					-- layer=2 filter=239 channel=29
					-2, 3, 0, 1, 4, -6, 1, 8, 8,
					-- layer=2 filter=239 channel=30
					-31, -3, -16, 5, 1, 5, 14, -1, 14,
					-- layer=2 filter=239 channel=31
					-32, 6, -30, -28, 48, -46, 47, -1, 46,
					-- layer=2 filter=239 channel=32
					-8, 11, -5, 1, -10, -2, -4, -9, -8,
					-- layer=2 filter=239 channel=33
					0, -19, -23, -47, -50, -20, 28, -42, 8,
					-- layer=2 filter=239 channel=34
					2, -13, 38, 6, 39, 30, 28, 14, 33,
					-- layer=2 filter=239 channel=35
					-4, 3, 23, 7, 24, -4, 5, 17, 5,
					-- layer=2 filter=239 channel=36
					-6, 4, -5, -10, 0, 7, 1, 2, 5,
					-- layer=2 filter=239 channel=37
					-30, -6, 3, 9, -8, 10, 21, 15, 7,
					-- layer=2 filter=239 channel=38
					-20, -50, -27, 14, 10, -16, 26, 27, 3,
					-- layer=2 filter=239 channel=39
					-8, -4, -4, -25, -7, -12, -13, -15, 6,
					-- layer=2 filter=239 channel=40
					25, 5, 13, 66, 53, 44, 20, -53, -2,
					-- layer=2 filter=239 channel=41
					1, -6, -2, 7, 6, -4, 7, 8, -9,
					-- layer=2 filter=239 channel=42
					-9, -35, -22, -36, -50, -34, -15, -29, 4,
					-- layer=2 filter=239 channel=43
					-30, -9, -43, -39, -15, -15, -2, -33, 18,
					-- layer=2 filter=239 channel=44
					3, -5, 9, 1, -7, 0, -10, 0, 3,
					-- layer=2 filter=239 channel=45
					-12, 2, -14, -11, 10, -5, -4, -10, 24,
					-- layer=2 filter=239 channel=46
					2, 6, -13, 7, 10, -10, 4, -2, -14,
					-- layer=2 filter=239 channel=47
					30, 43, 27, -16, 12, -17, 15, -31, 11,
					-- layer=2 filter=239 channel=48
					-8, -5, 8, -3, -3, 5, -5, -7, 4,
					-- layer=2 filter=239 channel=49
					0, -72, -1, -22, -1, -23, -59, -43, -13,
					-- layer=2 filter=239 channel=50
					5, 5, -5, -14, 5, -10, -4, -2, -20,
					-- layer=2 filter=239 channel=51
					-33, -26, -9, -2, -6, 13, 7, 15, 3,
					-- layer=2 filter=239 channel=52
					-37, 5, 7, 12, -1, -7, 0, 17, 15,
					-- layer=2 filter=239 channel=53
					6, 5, -36, -29, 7, -63, -20, -42, -15,
					-- layer=2 filter=239 channel=54
					15, -20, 12, 15, 19, 1, 28, 33, 41,
					-- layer=2 filter=239 channel=55
					-2, 0, -1, -10, 6, -5, -4, 5, -8,
					-- layer=2 filter=239 channel=56
					-40, -19, -27, 26, -14, 0, 1, 16, 11,
					-- layer=2 filter=239 channel=57
					-4, 2, 1, -2, -7, -6, 8, 4, 7,
					-- layer=2 filter=239 channel=58
					-27, -14, -68, -15, -12, -11, -38, -27, -14,
					-- layer=2 filter=239 channel=59
					-6, 15, 25, 27, -32, -17, -39, 21, 2,
					-- layer=2 filter=239 channel=60
					5, -14, 14, -22, 18, -10, -15, -19, -39,
					-- layer=2 filter=239 channel=61
					-11, 9, 25, 1, 21, 22, 14, -24, -1,
					-- layer=2 filter=239 channel=62
					20, -17, -2, 18, 15, 36, 9, 50, 26,
					-- layer=2 filter=239 channel=63
					20, 7, 7, 5, -6, 13, 21, 5, 24,
					-- layer=2 filter=239 channel=64
					-2, -1, -14, 3, -10, -29, -6, 2, -20,
					-- layer=2 filter=239 channel=65
					-1, 38, 48, 29, 31, 32, 42, 23, -1,
					-- layer=2 filter=239 channel=66
					2, 6, -24, 0, -7, 0, -18, 33, -16,
					-- layer=2 filter=239 channel=67
					11, 16, -21, 12, -3, -5, 7, 0, -12,
					-- layer=2 filter=239 channel=68
					4, 4, 8, 1, -8, -6, 7, 10, 3,
					-- layer=2 filter=239 channel=69
					16, -6, -12, -8, -6, -9, -25, 7, -3,
					-- layer=2 filter=239 channel=70
					0, 1, 16, 13, 17, 23, 4, 7, 17,
					-- layer=2 filter=239 channel=71
					-36, -2, 22, -44, -69, -42, 10, -43, -23,
					-- layer=2 filter=239 channel=72
					-34, -31, -33, 0, -22, -16, 21, -2, -24,
					-- layer=2 filter=239 channel=73
					6, 36, -8, -1, 23, 33, -44, -29, 32,
					-- layer=2 filter=239 channel=74
					-6, -13, -5, 28, 13, 6, 4, -11, 3,
					-- layer=2 filter=239 channel=75
					-46, -104, -68, -21, -56, -35, -13, -29, -7,
					-- layer=2 filter=239 channel=76
					29, 17, 22, 11, 38, -20, -36, 10, 41,
					-- layer=2 filter=239 channel=77
					-4, -6, -4, -1, -9, -4, -3, 0, -3,
					-- layer=2 filter=239 channel=78
					-21, -17, -28, -2, -14, -22, -15, -10, -13,
					-- layer=2 filter=239 channel=79
					1, 8, 1, -3, 3, 5, 0, -7, 0,
					-- layer=2 filter=239 channel=80
					14, 10, 5, 8, 2, 3, 14, 0, -13,
					-- layer=2 filter=239 channel=81
					-1, 0, -13, -16, -1, -18, -7, -7, 0,
					-- layer=2 filter=239 channel=82
					-1, -2, -3, -2, -6, 8, -7, 7, 3,
					-- layer=2 filter=239 channel=83
					-4, 14, -1, 29, -1, 8, 29, -12, 31,
					-- layer=2 filter=239 channel=84
					3, 0, 1, 0, -11, -11, 8, 9, 11,
					-- layer=2 filter=239 channel=85
					0, 11, -7, 9, -7, -6, -5, -3, -6,
					-- layer=2 filter=239 channel=86
					6, 21, -4, 14, 1, 7, -4, 0, -7,
					-- layer=2 filter=239 channel=87
					63, -2, -5, 30, 35, -7, -43, 14, 31,
					-- layer=2 filter=239 channel=88
					-2, 8, -8, 19, 25, 24, 31, -10, 5,
					-- layer=2 filter=239 channel=89
					-46, -30, -21, -14, -23, -50, -38, -6, -23,
					-- layer=2 filter=239 channel=90
					-2, -2, 4, 0, 13, 6, 4, -3, 4,
					-- layer=2 filter=239 channel=91
					-54, -50, -71, -88, -60, -74, -60, -76, -77,
					-- layer=2 filter=239 channel=92
					-55, -28, -42, -26, -20, -65, -40, -11, -35,
					-- layer=2 filter=239 channel=93
					-27, 4, -7, -30, -78, -14, -34, -44, -65,
					-- layer=2 filter=239 channel=94
					4, -21, 21, 22, -3, 0, 35, 51, 11,
					-- layer=2 filter=239 channel=95
					-3, -25, -10, -2, -12, -12, 15, -8, 3,
					-- layer=2 filter=239 channel=96
					5, 16, 6, 81, 19, 22, 29, 49, -3,
					-- layer=2 filter=239 channel=97
					22, -10, -27, -8, -7, -4, -31, -47, -9,
					-- layer=2 filter=239 channel=98
					7, 36, 27, 12, 27, -15, 30, 5, 23,
					-- layer=2 filter=239 channel=99
					39, 38, 56, 0, -7, -37, -9, 11, -18,
					-- layer=2 filter=239 channel=100
					10, -37, -13, 35, 13, 13, 18, 22, 12,
					-- layer=2 filter=239 channel=101
					36, 9, 64, -21, -11, 22, -14, -11, -31,
					-- layer=2 filter=239 channel=102
					8, -18, 21, 33, 19, -24, -2, 62, -32,
					-- layer=2 filter=239 channel=103
					-45, 11, 1, -15, 11, -22, 23, 16, 22,
					-- layer=2 filter=239 channel=104
					-4, -76, -10, 2, 6, -13, -7, 7, 15,
					-- layer=2 filter=239 channel=105
					25, -6, 46, 52, 23, 60, -33, -37, 20,
					-- layer=2 filter=239 channel=106
					-23, -24, -40, -39, -25, 16, -56, -72, -29,
					-- layer=2 filter=239 channel=107
					-12, 19, 3, 33, -1, -11, -5, -35, -50,
					-- layer=2 filter=239 channel=108
					-59, -17, 1, -6, 0, -13, 0, 9, -5,
					-- layer=2 filter=239 channel=109
					12, -11, -12, 5, -11, -6, 0, -8, 5,
					-- layer=2 filter=239 channel=110
					5, -16, -13, -49, -43, -50, -88, -64, -45,
					-- layer=2 filter=239 channel=111
					-2, -8, -7, 2, -6, -6, -3, -1, 3,
					-- layer=2 filter=239 channel=112
					-6, -42, 11, 6, 0, -3, -10, -30, 5,
					-- layer=2 filter=239 channel=113
					-5, -16, 16, -14, 13, 2, 1, -3, 15,
					-- layer=2 filter=239 channel=114
					1, 2, 9, 6, 0, -1, 14, -2, 1,
					-- layer=2 filter=239 channel=115
					3, 0, 1, -4, 2, -4, -4, 9, -8,
					-- layer=2 filter=239 channel=116
					21, 9, -25, 6, 23, 0, -23, 5, -13,
					-- layer=2 filter=239 channel=117
					-32, -4, -5, -34, -2, -31, 8, 0, -35,
					-- layer=2 filter=239 channel=118
					13, 10, -17, -27, -2, 14, -23, -6, 5,
					-- layer=2 filter=239 channel=119
					37, -14, 16, 25, 40, 30, 25, 13, 41,
					-- layer=2 filter=239 channel=120
					2, 0, 7, -2, -8, -2, 7, -1, -10,
					-- layer=2 filter=239 channel=121
					1, 5, -3, 0, -4, 0, 0, -5, -4,
					-- layer=2 filter=239 channel=122
					-15, -4, -4, -6, -3, 13, 3, 5, 0,
					-- layer=2 filter=239 channel=123
					1, -29, -8, 6, 5, -10, 21, 9, 5,
					-- layer=2 filter=239 channel=124
					16, -27, -47, -16, 13, -64, -15, -49, 19,
					-- layer=2 filter=239 channel=125
					-3, -5, -6, 5, 5, 8, 9, 12, 8,
					-- layer=2 filter=239 channel=126
					-38, -11, -63, -71, -26, 3, -51, -53, -69,
					-- layer=2 filter=239 channel=127
					8, 4, -5, 0, 13, 13, 8, 25, 11,
					-- layer=2 filter=240 channel=0
					-6, -7, 8, -21, -7, 30, 0, 12, 20,
					-- layer=2 filter=240 channel=1
					-44, -2, 7, -39, -54, -6, -1, -20, 21,
					-- layer=2 filter=240 channel=2
					3, -1, 1, 5, 9, 5, 4, -4, -7,
					-- layer=2 filter=240 channel=3
					22, 7, 1, 17, -24, -24, -38, -15, 5,
					-- layer=2 filter=240 channel=4
					-24, -41, -26, 18, 4, 11, 26, 0, 3,
					-- layer=2 filter=240 channel=5
					-12, 9, 12, -19, 14, 19, -26, -31, 16,
					-- layer=2 filter=240 channel=6
					23, -3, 4, 23, 58, 48, -11, 6, 67,
					-- layer=2 filter=240 channel=7
					-17, -34, -10, 26, 1, 6, 12, 27, 24,
					-- layer=2 filter=240 channel=8
					-3, -5, 11, -11, -4, 1, -5, 4, 1,
					-- layer=2 filter=240 channel=9
					26, 11, -2, 42, -26, -8, -19, -4, 23,
					-- layer=2 filter=240 channel=10
					32, 20, 33, 14, -9, 12, -11, 1, 22,
					-- layer=2 filter=240 channel=11
					5, 16, 19, -1, 16, 22, 8, 4, 20,
					-- layer=2 filter=240 channel=12
					-25, 4, 16, 8, 16, -7, 15, -6, 37,
					-- layer=2 filter=240 channel=13
					9, -1, -9, -5, 11, -3, -2, -7, 9,
					-- layer=2 filter=240 channel=14
					-32, 5, 6, 14, 7, -8, 13, 5, 15,
					-- layer=2 filter=240 channel=15
					-24, -43, -3, 0, -53, -15, 7, -70, 18,
					-- layer=2 filter=240 channel=16
					8, -22, -18, -12, -5, -47, 1, -55, -35,
					-- layer=2 filter=240 channel=17
					2, -2, -4, 4, -3, 4, 1, -7, 2,
					-- layer=2 filter=240 channel=18
					21, 7, -1, -32, -30, -22, -25, -66, -79,
					-- layer=2 filter=240 channel=19
					-17, -6, 22, -37, -70, -12, -24, -13, -41,
					-- layer=2 filter=240 channel=20
					0, -6, 5, 4, 0, -2, -6, -12, 5,
					-- layer=2 filter=240 channel=21
					1, -1, -5, 0, -14, -1, 4, -12, -12,
					-- layer=2 filter=240 channel=22
					4, 10, 1, -6, -8, -1, 2, -6, -4,
					-- layer=2 filter=240 channel=23
					-12, -33, -23, 14, -14, -22, 9, -5, -6,
					-- layer=2 filter=240 channel=24
					53, 21, 4, 19, -14, -10, -32, -14, -18,
					-- layer=2 filter=240 channel=25
					27, 31, -6, 31, 10, -3, -6, 13, 4,
					-- layer=2 filter=240 channel=26
					4, 4, -9, -5, 4, 6, 5, 2, 1,
					-- layer=2 filter=240 channel=27
					-37, -5, -36, -20, -32, -3, 4, 0, 4,
					-- layer=2 filter=240 channel=28
					6, -22, 7, 33, 10, 13, 10, 30, 39,
					-- layer=2 filter=240 channel=29
					0, 0, 1, 2, 6, 1, 4, -2, 1,
					-- layer=2 filter=240 channel=30
					30, 30, -19, -19, -20, -14, -11, -13, -16,
					-- layer=2 filter=240 channel=31
					29, 34, 75, -49, 66, 2, -61, -39, -3,
					-- layer=2 filter=240 channel=32
					0, -9, -5, -7, 7, 0, -5, 4, -9,
					-- layer=2 filter=240 channel=33
					-19, -21, 2, 32, -52, 5, 44, 8, 24,
					-- layer=2 filter=240 channel=34
					-24, 14, 44, -19, 9, 44, -21, 0, -30,
					-- layer=2 filter=240 channel=35
					14, 8, 4, 18, 32, -5, 11, 7, 9,
					-- layer=2 filter=240 channel=36
					5, -5, -1, -6, 4, -11, -13, 1, 0,
					-- layer=2 filter=240 channel=37
					-20, 10, 1, 0, 3, 14, 3, -24, 11,
					-- layer=2 filter=240 channel=38
					-62, -5, -18, -15, 15, -31, -16, -26, 5,
					-- layer=2 filter=240 channel=39
					0, 8, -33, -1, -59, -9, -52, -76, -32,
					-- layer=2 filter=240 channel=40
					29, 32, 6, -49, 12, -5, -58, -69, -49,
					-- layer=2 filter=240 channel=41
					-5, 1, -10, -2, 10, 7, 0, 4, -10,
					-- layer=2 filter=240 channel=42
					18, -24, -35, 3, 12, -13, -5, -45, -28,
					-- layer=2 filter=240 channel=43
					20, 33, 19, -26, -3, 15, -19, -16, -41,
					-- layer=2 filter=240 channel=44
					-9, -2, 6, 5, -6, -5, 1, -2, 4,
					-- layer=2 filter=240 channel=45
					48, -6, -32, -17, -49, -31, 24, -64, -19,
					-- layer=2 filter=240 channel=46
					4, 24, -18, -17, -8, 9, -10, -19, -12,
					-- layer=2 filter=240 channel=47
					-45, -49, -39, -17, -38, -23, -25, -5, -19,
					-- layer=2 filter=240 channel=48
					9, 5, -1, -8, 10, 0, 8, -3, 0,
					-- layer=2 filter=240 channel=49
					-15, 14, 3, -73, -39, -67, -10, -98, -42,
					-- layer=2 filter=240 channel=50
					-4, -24, -10, 8, -7, 1, -20, 0, 3,
					-- layer=2 filter=240 channel=51
					-21, 0, 18, 15, 22, 31, -8, 19, 10,
					-- layer=2 filter=240 channel=52
					20, 23, 28, 19, -8, 46, -10, -8, 13,
					-- layer=2 filter=240 channel=53
					31, 47, 32, -76, 1, 15, -65, -89, -33,
					-- layer=2 filter=240 channel=54
					0, 19, 21, -9, 27, 8, 8, 26, 31,
					-- layer=2 filter=240 channel=55
					-3, 4, 0, 0, -9, 9, -13, -4, -5,
					-- layer=2 filter=240 channel=56
					7, 2, 24, -17, -9, 9, -32, -17, -10,
					-- layer=2 filter=240 channel=57
					14, -6, -3, -5, -8, -10, 5, 0, -2,
					-- layer=2 filter=240 channel=58
					-6, 0, 11, 12, -9, 18, 20, -15, 30,
					-- layer=2 filter=240 channel=59
					-52, -15, 33, -25, -40, -47, -21, -31, -27,
					-- layer=2 filter=240 channel=60
					-18, -18, 5, -55, -29, -44, -18, -36, -4,
					-- layer=2 filter=240 channel=61
					49, 0, 0, 21, -33, -2, -42, -46, -26,
					-- layer=2 filter=240 channel=62
					11, 24, 24, -7, 31, 49, 29, -23, 7,
					-- layer=2 filter=240 channel=63
					19, -33, -11, -13, -55, -19, -17, -21, 0,
					-- layer=2 filter=240 channel=64
					29, 12, -11, 19, -9, -17, -10, -24, -31,
					-- layer=2 filter=240 channel=65
					42, 18, 21, 53, 13, 18, 5, -15, 0,
					-- layer=2 filter=240 channel=66
					17, 25, -50, 18, 34, 7, -9, -23, -20,
					-- layer=2 filter=240 channel=67
					29, 15, -2, 4, -25, -10, -32, -84, -13,
					-- layer=2 filter=240 channel=68
					0, 1, -7, 9, 10, 0, -4, -1, -8,
					-- layer=2 filter=240 channel=69
					11, -1, -16, 24, -11, -18, -5, -35, -11,
					-- layer=2 filter=240 channel=70
					5, -25, 9, 6, 9, 14, 14, 38, 32,
					-- layer=2 filter=240 channel=71
					-6, 23, -28, -48, -41, -23, -31, -8, 8,
					-- layer=2 filter=240 channel=72
					-17, -18, 44, 26, 6, 54, 34, 45, 32,
					-- layer=2 filter=240 channel=73
					59, 69, 45, 9, 42, 15, -21, -5, 7,
					-- layer=2 filter=240 channel=74
					3, 10, 3, -7, -24, -14, -6, -25, 17,
					-- layer=2 filter=240 channel=75
					47, 4, 6, 32, 28, -7, -25, -45, 4,
					-- layer=2 filter=240 channel=76
					11, 43, -22, -5, 30, 17, -68, -12, -5,
					-- layer=2 filter=240 channel=77
					3, -9, 6, 10, 11, -8, 2, 2, 6,
					-- layer=2 filter=240 channel=78
					1, 23, -8, -8, -6, 23, -12, 2, 10,
					-- layer=2 filter=240 channel=79
					-3, 1, -3, -7, 0, 7, -1, 4, 0,
					-- layer=2 filter=240 channel=80
					12, 8, -19, 34, -12, -5, 21, -18, -8,
					-- layer=2 filter=240 channel=81
					-7, 0, -2, -9, 0, 1, -7, -9, 6,
					-- layer=2 filter=240 channel=82
					-8, 11, -1, -7, 3, 2, -1, 8, 8,
					-- layer=2 filter=240 channel=83
					10, -7, -59, 7, -3, -28, 64, 16, 33,
					-- layer=2 filter=240 channel=84
					0, 0, 0, 0, 0, -3, -1, -1, -3,
					-- layer=2 filter=240 channel=85
					-3, 0, -23, 0, -11, 1, -8, 2, 3,
					-- layer=2 filter=240 channel=86
					-8, -9, -10, -9, -17, -14, -1, -9, 9,
					-- layer=2 filter=240 channel=87
					-10, 14, 22, -6, 0, 1, -12, 0, -76,
					-- layer=2 filter=240 channel=88
					14, 12, -10, 20, 5, -35, 25, -23, 1,
					-- layer=2 filter=240 channel=89
					-33, 11, 10, 0, -6, -14, 22, -10, -16,
					-- layer=2 filter=240 channel=90
					6, -2, 7, -2, 3, 0, 1, -4, -8,
					-- layer=2 filter=240 channel=91
					-23, 5, -1, 0, 30, 6, -25, -13, 23,
					-- layer=2 filter=240 channel=92
					-37, -9, -9, -15, 4, -16, 17, -4, 2,
					-- layer=2 filter=240 channel=93
					10, -2, 55, -10, -47, 40, -57, -18, -9,
					-- layer=2 filter=240 channel=94
					35, -29, -5, -55, -24, -3, -9, -3, -21,
					-- layer=2 filter=240 channel=95
					-2, -3, 0, -10, 0, -1, -14, -17, -5,
					-- layer=2 filter=240 channel=96
					-24, 20, 37, 18, 26, 28, 16, 13, 20,
					-- layer=2 filter=240 channel=97
					24, 35, -27, 28, -25, 0, 12, 8, -2,
					-- layer=2 filter=240 channel=98
					0, -7, 4, 20, 20, 16, -5, 40, 8,
					-- layer=2 filter=240 channel=99
					15, 47, 46, 17, -52, 29, -48, 35, -22,
					-- layer=2 filter=240 channel=100
					-39, -24, -25, 14, 17, 31, 29, 11, 25,
					-- layer=2 filter=240 channel=101
					15, 26, -10, 5, 21, -23, -8, 9, 5,
					-- layer=2 filter=240 channel=102
					-12, 13, 16, 17, -33, -12, 10, -30, -36,
					-- layer=2 filter=240 channel=103
					9, 24, 23, 5, -37, -31, -43, 23, 51,
					-- layer=2 filter=240 channel=104
					11, -16, -19, -45, 20, -44, 2, -100, -65,
					-- layer=2 filter=240 channel=105
					8, 68, 11, 7, 3, -18, -11, -3, 22,
					-- layer=2 filter=240 channel=106
					25, 13, -11, 38, 3, 4, -28, -22, -16,
					-- layer=2 filter=240 channel=107
					56, 56, 30, 25, 43, -40, 0, 48, -19,
					-- layer=2 filter=240 channel=108
					-51, -17, -27, -11, -76, -41, -23, -18, -32,
					-- layer=2 filter=240 channel=109
					-13, -7, -4, -4, 4, 2, 8, -13, -2,
					-- layer=2 filter=240 channel=110
					45, 7, -36, 32, 0, -44, -17, -43, -73,
					-- layer=2 filter=240 channel=111
					-10, -4, -2, 2, 2, -10, -5, 8, -3,
					-- layer=2 filter=240 channel=112
					12, 4, -11, -13, -18, -27, -33, -56, -42,
					-- layer=2 filter=240 channel=113
					4, -22, -21, -14, -2, -27, -32, -4, -17,
					-- layer=2 filter=240 channel=114
					1, 6, 15, 3, 7, -7, 1, 0, 20,
					-- layer=2 filter=240 channel=115
					6, 10, -8, 0, -5, 9, 7, 7, 3,
					-- layer=2 filter=240 channel=116
					-14, 0, 12, 2, -26, -6, -16, -29, -82,
					-- layer=2 filter=240 channel=117
					12, 3, 27, 7, -2, -12, -22, 21, -13,
					-- layer=2 filter=240 channel=118
					3, 29, 31, 17, 7, 21, -10, 7, 32,
					-- layer=2 filter=240 channel=119
					20, -19, -9, -2, 12, -21, 12, -17, -47,
					-- layer=2 filter=240 channel=120
					-5, -7, 1, -3, -7, -1, -7, -6, 5,
					-- layer=2 filter=240 channel=121
					0, -3, -7, -7, -3, 2, -1, -2, -1,
					-- layer=2 filter=240 channel=122
					2, 10, -2, -18, 0, -7, -7, 15, -8,
					-- layer=2 filter=240 channel=123
					-34, -6, 6, 15, 0, 28, -3, 6, 8,
					-- layer=2 filter=240 channel=124
					-15, -26, -23, 3, 7, -27, 1, -37, 13,
					-- layer=2 filter=240 channel=125
					8, 1, -10, -3, 6, 6, 6, 6, 2,
					-- layer=2 filter=240 channel=126
					16, -9, 26, -38, -63, 2, -9, -12, -51,
					-- layer=2 filter=240 channel=127
					-19, -9, -1, 34, 0, -3, 14, -39, 30,
					-- layer=2 filter=241 channel=0
					4, -12, -11, -3, -13, -10, 0, -10, -10,
					-- layer=2 filter=241 channel=1
					5, 1, -9, 6, 6, -3, -7, -10, 1,
					-- layer=2 filter=241 channel=2
					1, -5, -9, 5, -9, -2, 9, 6, 0,
					-- layer=2 filter=241 channel=3
					-4, -8, -13, 7, -13, -1, -10, 1, -10,
					-- layer=2 filter=241 channel=4
					-5, 2, 5, -1, -9, 5, 4, -3, -8,
					-- layer=2 filter=241 channel=5
					-8, 0, -8, 5, -8, -11, 0, -3, 5,
					-- layer=2 filter=241 channel=6
					2, -3, 3, -5, -13, -3, 6, -2, 0,
					-- layer=2 filter=241 channel=7
					-10, -5, -1, -11, 5, 6, 0, 4, 3,
					-- layer=2 filter=241 channel=8
					-6, 2, 0, 5, 9, -7, -1, 9, -6,
					-- layer=2 filter=241 channel=9
					-3, -4, -1, 7, -1, -12, 7, -5, -11,
					-- layer=2 filter=241 channel=10
					-16, -3, -1, 1, -13, -1, -10, 4, -8,
					-- layer=2 filter=241 channel=11
					0, 8, 6, -5, -11, -12, -8, -12, -6,
					-- layer=2 filter=241 channel=12
					0, 0, -2, 6, 3, -9, -14, -14, 0,
					-- layer=2 filter=241 channel=13
					-4, -10, -3, 0, 3, 0, -5, 5, 5,
					-- layer=2 filter=241 channel=14
					-5, 1, 0, -11, -3, -10, -13, -5, 6,
					-- layer=2 filter=241 channel=15
					0, -10, 3, 1, -2, -6, -5, 2, -3,
					-- layer=2 filter=241 channel=16
					3, 5, -1, 4, 3, -3, 7, -8, -2,
					-- layer=2 filter=241 channel=17
					6, 2, 8, 2, 9, 2, -8, -3, 4,
					-- layer=2 filter=241 channel=18
					-5, 7, -9, -4, -15, 2, -7, -12, -11,
					-- layer=2 filter=241 channel=19
					-8, -3, 2, -6, -10, 1, -7, -4, -14,
					-- layer=2 filter=241 channel=20
					4, 3, -6, 7, -8, -2, -3, 4, 2,
					-- layer=2 filter=241 channel=21
					7, 2, 4, 0, 8, -10, -3, -8, -1,
					-- layer=2 filter=241 channel=22
					-5, -4, 1, -8, -5, -2, -2, 5, 11,
					-- layer=2 filter=241 channel=23
					-11, -11, -6, 4, -9, 2, -6, -7, -5,
					-- layer=2 filter=241 channel=24
					0, 2, 2, -7, -12, -6, 1, -9, -3,
					-- layer=2 filter=241 channel=25
					3, -11, 5, -8, -4, -9, 0, -13, 0,
					-- layer=2 filter=241 channel=26
					-1, 5, -4, -3, 2, 0, 9, 3, -2,
					-- layer=2 filter=241 channel=27
					4, 1, -4, 9, -7, -8, 5, 3, 2,
					-- layer=2 filter=241 channel=28
					0, 8, -5, -9, -6, 0, 10, -8, -2,
					-- layer=2 filter=241 channel=29
					5, 7, 0, 2, -4, 3, -4, -4, 8,
					-- layer=2 filter=241 channel=30
					2, -2, -6, 0, 1, -7, -15, -2, -9,
					-- layer=2 filter=241 channel=31
					-6, 0, -10, 3, 1, 5, 3, 8, -8,
					-- layer=2 filter=241 channel=32
					-8, 0, 3, 3, -9, -7, 1, 3, -8,
					-- layer=2 filter=241 channel=33
					-9, -6, 2, 2, 3, 0, 0, -6, -11,
					-- layer=2 filter=241 channel=34
					-9, -4, 3, 0, 0, -6, -6, 3, 1,
					-- layer=2 filter=241 channel=35
					3, -5, -3, 0, 3, 1, 4, 0, -5,
					-- layer=2 filter=241 channel=36
					-9, -11, -10, 6, -6, 3, 3, 5, -2,
					-- layer=2 filter=241 channel=37
					-8, -7, -8, -3, 5, -10, 0, 0, 0,
					-- layer=2 filter=241 channel=38
					-10, -2, 4, 3, -12, -12, -15, -7, 5,
					-- layer=2 filter=241 channel=39
					8, -7, 0, 1, -9, -7, 6, -8, -7,
					-- layer=2 filter=241 channel=40
					-8, -4, -5, 5, 6, -8, -10, -9, -6,
					-- layer=2 filter=241 channel=41
					0, -11, 0, 0, 0, -6, 0, -7, 9,
					-- layer=2 filter=241 channel=42
					0, -14, 0, -12, -10, -15, 5, 5, -12,
					-- layer=2 filter=241 channel=43
					-5, 1, -11, -6, 2, -12, 7, -2, -9,
					-- layer=2 filter=241 channel=44
					-2, -5, 4, -3, 0, -4, 8, 3, 3,
					-- layer=2 filter=241 channel=45
					2, -6, -10, -3, 8, -9, -1, -5, -11,
					-- layer=2 filter=241 channel=46
					0, -6, 2, -9, 3, 3, -3, -1, 4,
					-- layer=2 filter=241 channel=47
					-3, -13, -8, -1, 7, -15, 4, -11, -2,
					-- layer=2 filter=241 channel=48
					-7, 2, -1, -9, 6, 0, 5, -6, -7,
					-- layer=2 filter=241 channel=49
					9, 6, -13, 10, -6, -1, -6, 5, -17,
					-- layer=2 filter=241 channel=50
					0, 0, -10, -7, 5, -3, -2, 0, -10,
					-- layer=2 filter=241 channel=51
					-4, -12, -7, -15, -2, -3, -16, 0, 1,
					-- layer=2 filter=241 channel=52
					10, 2, 1, 4, -10, 0, -13, 0, -8,
					-- layer=2 filter=241 channel=53
					5, 0, -6, -6, -5, -9, 8, 0, 5,
					-- layer=2 filter=241 channel=54
					-5, -15, -12, -9, 7, -8, -11, -2, -5,
					-- layer=2 filter=241 channel=55
					1, 3, 0, -2, 8, -8, 5, -6, 9,
					-- layer=2 filter=241 channel=56
					5, 7, 5, -12, 5, -13, -13, -1, 2,
					-- layer=2 filter=241 channel=57
					-2, 2, -7, -10, -3, 11, 7, -2, -1,
					-- layer=2 filter=241 channel=58
					-4, -11, -9, 0, 7, -3, -11, 3, -3,
					-- layer=2 filter=241 channel=59
					1, -3, -7, -5, -12, -11, 0, -1, 2,
					-- layer=2 filter=241 channel=60
					-7, -2, -9, -6, -10, -4, -3, 2, -12,
					-- layer=2 filter=241 channel=61
					-11, -11, -12, -9, -3, -6, 1, -12, -5,
					-- layer=2 filter=241 channel=62
					4, 7, 1, 3, -16, -5, 5, -2, -4,
					-- layer=2 filter=241 channel=63
					-10, -8, -6, -16, 1, 0, 5, 1, 1,
					-- layer=2 filter=241 channel=64
					-5, -2, -12, 2, -12, 4, 1, -12, 0,
					-- layer=2 filter=241 channel=65
					1, -12, -5, -11, 0, 8, -10, -3, 1,
					-- layer=2 filter=241 channel=66
					-5, -1, -5, -3, 0, -1, -6, -1, -2,
					-- layer=2 filter=241 channel=67
					8, 6, -12, 4, -15, 6, -13, 6, -4,
					-- layer=2 filter=241 channel=68
					2, -11, -6, -7, -2, -2, -2, 8, 9,
					-- layer=2 filter=241 channel=69
					0, -19, -5, -9, -4, 1, 2, -10, 4,
					-- layer=2 filter=241 channel=70
					-2, 0, -4, 0, -14, -10, -13, 5, -8,
					-- layer=2 filter=241 channel=71
					4, 0, -7, 6, 0, 0, 1, 7, 0,
					-- layer=2 filter=241 channel=72
					0, -7, -3, -6, -4, -8, -6, 3, -9,
					-- layer=2 filter=241 channel=73
					2, -8, 0, 5, 6, -2, -8, -10, 1,
					-- layer=2 filter=241 channel=74
					-3, 7, -10, -11, -6, -9, -5, 3, 3,
					-- layer=2 filter=241 channel=75
					-3, 4, -9, 7, -1, 2, 5, 3, 0,
					-- layer=2 filter=241 channel=76
					-2, -2, -1, 3, -6, 4, 2, 7, 0,
					-- layer=2 filter=241 channel=77
					-7, -3, 4, 4, -3, -9, 0, -1, -6,
					-- layer=2 filter=241 channel=78
					5, 0, 0, 2, -5, 1, 5, -8, 0,
					-- layer=2 filter=241 channel=79
					6, -9, -8, -8, 3, -11, -8, -6, -7,
					-- layer=2 filter=241 channel=80
					0, 1, -8, 7, -1, 7, -3, -3, -9,
					-- layer=2 filter=241 channel=81
					6, 0, 5, -1, 0, 8, 4, -9, 8,
					-- layer=2 filter=241 channel=82
					6, -4, 2, -4, 7, 0, 7, 8, -9,
					-- layer=2 filter=241 channel=83
					0, -11, -6, -8, -8, 6, -10, 0, 1,
					-- layer=2 filter=241 channel=84
					6, -4, -10, 1, 2, -3, -1, -11, -7,
					-- layer=2 filter=241 channel=85
					0, 7, 5, 5, -7, -5, 8, -6, 2,
					-- layer=2 filter=241 channel=86
					-4, 0, -4, -10, 1, 8, 6, 8, 2,
					-- layer=2 filter=241 channel=87
					-11, 0, 0, -1, -3, -3, -9, -10, 8,
					-- layer=2 filter=241 channel=88
					4, 7, 2, 3, -8, 6, -6, -12, 4,
					-- layer=2 filter=241 channel=89
					-11, -8, -4, 2, 5, -10, 4, -11, -5,
					-- layer=2 filter=241 channel=90
					2, -6, 5, -7, 7, 9, 4, 4, 8,
					-- layer=2 filter=241 channel=91
					-7, 3, -3, -1, 0, -3, -2, -10, 8,
					-- layer=2 filter=241 channel=92
					5, 6, -9, 4, 3, 2, -10, -5, -3,
					-- layer=2 filter=241 channel=93
					-2, 1, 0, -12, -1, 0, 4, -4, -14,
					-- layer=2 filter=241 channel=94
					-6, -1, -4, 11, -3, 3, -11, -7, 0,
					-- layer=2 filter=241 channel=95
					8, 1, -3, -7, -12, -5, -5, 0, 6,
					-- layer=2 filter=241 channel=96
					-6, -11, 7, -13, -5, -10, 3, 0, -11,
					-- layer=2 filter=241 channel=97
					-5, 0, -13, -8, -6, -12, -10, 8, -8,
					-- layer=2 filter=241 channel=98
					-13, 0, -14, -13, -16, -12, -9, 6, -15,
					-- layer=2 filter=241 channel=99
					-1, 0, -10, 0, -1, 0, 0, -6, -3,
					-- layer=2 filter=241 channel=100
					-6, -13, 7, 4, -4, -9, -9, 4, -9,
					-- layer=2 filter=241 channel=101
					1, 8, -12, 2, -10, -8, -15, -8, -13,
					-- layer=2 filter=241 channel=102
					-7, -9, -7, 0, 6, -5, -5, -10, -7,
					-- layer=2 filter=241 channel=103
					1, -4, 8, 3, 0, 3, -10, -5, 0,
					-- layer=2 filter=241 channel=104
					-8, -9, 0, 5, -8, -13, -7, -12, 4,
					-- layer=2 filter=241 channel=105
					-5, -7, 7, -4, -6, 9, 7, 2, -9,
					-- layer=2 filter=241 channel=106
					-9, 0, 6, -9, -13, 6, 0, 0, -8,
					-- layer=2 filter=241 channel=107
					6, 9, -7, -6, -6, -10, 0, -9, 0,
					-- layer=2 filter=241 channel=108
					0, 0, 3, -1, -2, 5, -4, 7, -11,
					-- layer=2 filter=241 channel=109
					-8, -1, 7, 7, 1, -5, 8, -8, -4,
					-- layer=2 filter=241 channel=110
					-11, -8, -16, -4, 3, -7, -7, -10, -8,
					-- layer=2 filter=241 channel=111
					6, 2, 7, -5, 8, -6, 8, 4, 8,
					-- layer=2 filter=241 channel=112
					-13, 0, 0, -4, -3, -6, 0, 3, -1,
					-- layer=2 filter=241 channel=113
					-2, -9, -11, 0, -9, 7, 2, -18, 7,
					-- layer=2 filter=241 channel=114
					-9, 5, -11, -2, 12, 5, -1, -2, -2,
					-- layer=2 filter=241 channel=115
					-5, -7, 3, 2, -3, 2, -4, 8, -8,
					-- layer=2 filter=241 channel=116
					5, -3, -10, 0, -2, -15, 1, 6, -7,
					-- layer=2 filter=241 channel=117
					1, -4, 2, -13, -9, -4, 5, -3, 3,
					-- layer=2 filter=241 channel=118
					5, -10, -14, -7, 3, 1, -1, -9, -5,
					-- layer=2 filter=241 channel=119
					-6, 4, -12, 4, -1, 7, -4, 0, -12,
					-- layer=2 filter=241 channel=120
					-8, -1, -4, -1, 2, -2, 0, -10, 0,
					-- layer=2 filter=241 channel=121
					4, -3, -6, -3, -1, -5, -6, -8, -8,
					-- layer=2 filter=241 channel=122
					4, 4, -11, -3, -6, -8, 2, -10, -4,
					-- layer=2 filter=241 channel=123
					-9, -5, -4, -16, -11, 5, 6, -14, 6,
					-- layer=2 filter=241 channel=124
					-9, 0, 1, -5, -4, -15, 4, -2, -9,
					-- layer=2 filter=241 channel=125
					5, 3, 4, -10, 3, -7, 6, 3, -9,
					-- layer=2 filter=241 channel=126
					0, -14, -3, 1, 8, -10, 5, 3, 5,
					-- layer=2 filter=241 channel=127
					0, 0, 2, -3, -14, -10, 1, -16, -8,
					-- layer=2 filter=242 channel=0
					-15, -8, -30, -1, -3, -32, -2, -3, 13,
					-- layer=2 filter=242 channel=1
					-18, -13, -23, -11, -33, -8, -14, 0, -14,
					-- layer=2 filter=242 channel=2
					-3, -3, 6, 0, 0, 2, 11, 4, -3,
					-- layer=2 filter=242 channel=3
					-6, -20, -11, 16, -19, -7, 0, -10, -7,
					-- layer=2 filter=242 channel=4
					0, -12, -1, 5, -11, 0, -8, -40, -14,
					-- layer=2 filter=242 channel=5
					8, 7, 0, 3, -11, 10, -3, 8, -5,
					-- layer=2 filter=242 channel=6
					-27, 23, 14, -18, 24, 3, -15, 25, -26,
					-- layer=2 filter=242 channel=7
					32, -4, -19, 0, -3, -9, -28, 0, -8,
					-- layer=2 filter=242 channel=8
					5, 3, 1, 0, 5, 0, 1, 8, 7,
					-- layer=2 filter=242 channel=9
					9, -21, 4, -17, -20, 5, -11, -21, -5,
					-- layer=2 filter=242 channel=10
					-23, -20, -23, 0, -32, -13, 5, 4, 0,
					-- layer=2 filter=242 channel=11
					3, 1, -17, -2, -12, -10, -5, -11, -9,
					-- layer=2 filter=242 channel=12
					-22, 4, -4, -22, -30, -41, 17, 2, 1,
					-- layer=2 filter=242 channel=13
					-1, 0, -9, 6, -8, -5, 4, 3, -5,
					-- layer=2 filter=242 channel=14
					-3, -31, -32, -19, -27, -34, 4, -33, -19,
					-- layer=2 filter=242 channel=15
					6, -31, -2, -7, 23, -24, -22, -34, -35,
					-- layer=2 filter=242 channel=16
					43, -4, -27, -23, -23, 1, -16, -14, -11,
					-- layer=2 filter=242 channel=17
					1, 10, 1, -3, 4, 4, 1, 8, 11,
					-- layer=2 filter=242 channel=18
					-11, -9, 8, 8, 0, -4, 0, -28, -9,
					-- layer=2 filter=242 channel=19
					-10, 31, 20, -16, -33, 12, -23, -4, 1,
					-- layer=2 filter=242 channel=20
					9, 9, 1, 8, 12, 1, 4, 9, 3,
					-- layer=2 filter=242 channel=21
					-10, 1, 0, 0, -1, -11, 0, -2, 7,
					-- layer=2 filter=242 channel=22
					9, 0, -10, 7, -4, -2, 10, -5, -10,
					-- layer=2 filter=242 channel=23
					-26, -33, -36, -1, -28, -34, -30, -25, -29,
					-- layer=2 filter=242 channel=24
					5, 6, -10, -4, -4, -9, -3, -8, -4,
					-- layer=2 filter=242 channel=25
					17, 1, -20, -2, -2, -9, 3, -4, 10,
					-- layer=2 filter=242 channel=26
					5, 9, 8, 6, 7, 1, -5, 6, 10,
					-- layer=2 filter=242 channel=27
					-26, 4, 17, -34, -18, -5, -20, -19, 1,
					-- layer=2 filter=242 channel=28
					35, 3, 16, -10, 0, 6, 21, -11, -37,
					-- layer=2 filter=242 channel=29
					-7, 4, 2, -5, -9, -10, 4, 8, 0,
					-- layer=2 filter=242 channel=30
					-17, -9, -14, -2, -3, 0, -15, 16, -22,
					-- layer=2 filter=242 channel=31
					-16, 9, 19, 0, 8, -18, -10, -2, -21,
					-- layer=2 filter=242 channel=32
					5, -5, 2, -1, 5, 1, -5, 2, 6,
					-- layer=2 filter=242 channel=33
					0, -25, -19, 0, -16, -5, -20, -34, -26,
					-- layer=2 filter=242 channel=34
					4, 1, 20, -7, 7, 3, 0, 0, -6,
					-- layer=2 filter=242 channel=35
					22, -11, -5, -4, -5, -10, -17, 0, -25,
					-- layer=2 filter=242 channel=36
					6, -10, 8, -2, -8, -1, 7, -4, 5,
					-- layer=2 filter=242 channel=37
					-2, -10, 0, -20, 0, 19, -15, 0, 4,
					-- layer=2 filter=242 channel=38
					-49, -5, -8, 7, -17, -15, -9, 15, -20,
					-- layer=2 filter=242 channel=39
					22, -26, -25, -8, -14, -39, -36, -18, 19,
					-- layer=2 filter=242 channel=40
					29, -6, 27, 13, 8, 10, -29, -32, -25,
					-- layer=2 filter=242 channel=41
					1, 0, -7, 8, 7, -10, 0, -2, 0,
					-- layer=2 filter=242 channel=42
					-38, 5, 13, -14, 0, -28, -27, -32, -1,
					-- layer=2 filter=242 channel=43
					3, -46, 29, -4, -21, 25, 18, 0, -20,
					-- layer=2 filter=242 channel=44
					9, 0, -8, -5, -4, -1, -2, -6, 1,
					-- layer=2 filter=242 channel=45
					-1, 12, 11, -7, -13, -5, -28, -33, -12,
					-- layer=2 filter=242 channel=46
					-9, -6, -22, 20, 4, -19, 10, 17, -32,
					-- layer=2 filter=242 channel=47
					39, 18, -6, -34, 5, 3, -15, -30, -34,
					-- layer=2 filter=242 channel=48
					-3, 0, -7, -1, 8, -6, -2, 5, -6,
					-- layer=2 filter=242 channel=49
					-17, -2, -1, -12, -11, -9, -12, -23, -12,
					-- layer=2 filter=242 channel=50
					-9, 2, 7, -5, -3, -3, 3, 0, 7,
					-- layer=2 filter=242 channel=51
					8, -4, -17, 5, 3, -14, 12, 8, -10,
					-- layer=2 filter=242 channel=52
					0, -16, 0, -21, 16, -6, -23, -12, 7,
					-- layer=2 filter=242 channel=53
					24, 17, 25, 6, -4, -3, -16, -19, -4,
					-- layer=2 filter=242 channel=54
					-21, 6, -18, -5, 0, -10, -19, -4, -23,
					-- layer=2 filter=242 channel=55
					9, 4, -1, 0, 1, 5, -6, 1, 3,
					-- layer=2 filter=242 channel=56
					0, -13, -1, -6, -22, -15, -4, 0, -3,
					-- layer=2 filter=242 channel=57
					-10, 5, 6, -3, 6, -7, -5, -3, -7,
					-- layer=2 filter=242 channel=58
					-44, -2, 11, -1, -20, -41, 4, -2, 0,
					-- layer=2 filter=242 channel=59
					0, -22, -2, 16, -19, -27, -12, 4, -4,
					-- layer=2 filter=242 channel=60
					-2, 41, -42, -14, -8, -9, -27, -1, 7,
					-- layer=2 filter=242 channel=61
					-7, 19, -37, 4, 11, -22, -49, 25, -5,
					-- layer=2 filter=242 channel=62
					-22, -2, 13, -8, 16, 16, -26, 10, -5,
					-- layer=2 filter=242 channel=63
					2, -17, -1, -12, -22, -23, -35, -1, -4,
					-- layer=2 filter=242 channel=64
					-29, -24, -25, -9, -6, 4, -29, -17, 0,
					-- layer=2 filter=242 channel=65
					-46, 10, -5, 14, 20, -8, -5, 36, -28,
					-- layer=2 filter=242 channel=66
					23, -16, -6, -21, -4, -4, -10, 11, -16,
					-- layer=2 filter=242 channel=67
					-15, -4, -28, -4, -13, -8, 5, -8, 0,
					-- layer=2 filter=242 channel=68
					1, -3, -11, 3, 3, -8, -11, 1, 0,
					-- layer=2 filter=242 channel=69
					-28, -37, -26, -19, -24, -14, -30, -8, -3,
					-- layer=2 filter=242 channel=70
					14, -6, 0, -14, -3, -17, -8, 6, -31,
					-- layer=2 filter=242 channel=71
					-24, -2, 2, -33, -16, -8, -9, -29, 4,
					-- layer=2 filter=242 channel=72
					19, -3, -26, 26, 2, -21, -35, -12, -38,
					-- layer=2 filter=242 channel=73
					6, -4, 9, -18, -12, 10, -33, -54, 6,
					-- layer=2 filter=242 channel=74
					-13, -18, -13, -4, -24, 5, -5, -5, -3,
					-- layer=2 filter=242 channel=75
					37, 32, -16, -25, -8, -14, 27, 26, 7,
					-- layer=2 filter=242 channel=76
					16, 13, 22, -16, 3, -7, 3, -7, 8,
					-- layer=2 filter=242 channel=77
					8, -7, -2, -10, -11, 2, 1, -8, 4,
					-- layer=2 filter=242 channel=78
					-2, -15, -9, 0, -1, 17, -6, -5, -10,
					-- layer=2 filter=242 channel=79
					-9, 2, 1, -2, -9, -6, 0, -9, 8,
					-- layer=2 filter=242 channel=80
					-18, 5, -19, -21, -10, -9, -1, -43, -7,
					-- layer=2 filter=242 channel=81
					3, 0, 1, -10, 0, -5, -5, 3, 1,
					-- layer=2 filter=242 channel=82
					10, -3, 5, 6, 2, 0, 1, 1, -6,
					-- layer=2 filter=242 channel=83
					-30, -10, 2, -3, -16, -24, -43, 12, -18,
					-- layer=2 filter=242 channel=84
					0, 0, 11, 10, 6, 1, 0, 0, -11,
					-- layer=2 filter=242 channel=85
					0, 6, 0, 0, 0, -11, 3, 5, -9,
					-- layer=2 filter=242 channel=86
					-2, 0, 8, 6, -5, 3, 9, 9, 4,
					-- layer=2 filter=242 channel=87
					-11, -23, 12, -32, 9, -8, -11, -33, -23,
					-- layer=2 filter=242 channel=88
					-11, -27, -21, -29, -11, -23, -23, 0, -23,
					-- layer=2 filter=242 channel=89
					18, 4, -19, -4, -18, -29, -6, -17, -31,
					-- layer=2 filter=242 channel=90
					-4, 5, 8, 2, -10, -1, -9, 0, -3,
					-- layer=2 filter=242 channel=91
					8, 10, 7, -17, -46, -12, -7, -15, 11,
					-- layer=2 filter=242 channel=92
					-34, -22, -1, -5, -2, -24, -2, 7, -2,
					-- layer=2 filter=242 channel=93
					-48, 39, 22, -28, 24, 27, -15, 48, 7,
					-- layer=2 filter=242 channel=94
					-30, 9, 3, -6, 1, 1, -5, 13, -1,
					-- layer=2 filter=242 channel=95
					1, 2, -8, 0, 0, -1, -1, -1, -10,
					-- layer=2 filter=242 channel=96
					4, -26, -12, -12, 9, -21, -18, -36, -3,
					-- layer=2 filter=242 channel=97
					-10, -20, -14, 0, -5, -5, 3, -28, -8,
					-- layer=2 filter=242 channel=98
					28, 10, -9, -25, 11, 15, -19, -5, -20,
					-- layer=2 filter=242 channel=99
					-17, 5, 22, -4, 7, 34, -23, -8, -2,
					-- layer=2 filter=242 channel=100
					-24, 30, 1, -16, -56, 15, -10, 19, -7,
					-- layer=2 filter=242 channel=101
					-8, -10, -14, -25, -47, -20, -12, -12, -10,
					-- layer=2 filter=242 channel=102
					-7, -46, -20, -15, 3, -12, -11, -9, 22,
					-- layer=2 filter=242 channel=103
					-14, 17, -7, 2, -7, 10, 4, 9, -4,
					-- layer=2 filter=242 channel=104
					-9, -11, 1, -3, -2, -15, 9, -23, 1,
					-- layer=2 filter=242 channel=105
					56, 31, 13, -4, 15, 4, -2, -1, 11,
					-- layer=2 filter=242 channel=106
					11, 0, -22, -17, -34, -40, -33, -18, -4,
					-- layer=2 filter=242 channel=107
					0, 5, -18, -4, -13, 4, 1, 6, 13,
					-- layer=2 filter=242 channel=108
					-9, -14, -6, -43, -17, -10, -21, -22, 0,
					-- layer=2 filter=242 channel=109
					-2, 0, 1, 3, 6, 7, -5, -6, 3,
					-- layer=2 filter=242 channel=110
					3, -17, -17, 1, -4, -38, -35, -7, 2,
					-- layer=2 filter=242 channel=111
					-4, -4, -7, -7, -7, -2, -5, -3, 7,
					-- layer=2 filter=242 channel=112
					3, 18, -45, 30, 9, -38, -3, 40, -2,
					-- layer=2 filter=242 channel=113
					-23, -27, 0, 21, 9, -21, -23, 24, -11,
					-- layer=2 filter=242 channel=114
					5, 3, 2, -2, -1, 4, 0, -1, 2,
					-- layer=2 filter=242 channel=115
					2, 0, -2, -7, 0, 9, -4, -8, 8,
					-- layer=2 filter=242 channel=116
					-8, -27, 0, -23, 24, -5, -24, -26, -4,
					-- layer=2 filter=242 channel=117
					28, 17, -23, -15, 3, -2, -42, -20, -22,
					-- layer=2 filter=242 channel=118
					-6, -34, -8, -1, -6, 24, -10, -36, -4,
					-- layer=2 filter=242 channel=119
					-17, -7, -6, -13, 0, -8, 0, -24, -19,
					-- layer=2 filter=242 channel=120
					0, -8, 9, 6, -9, 3, -2, -6, 10,
					-- layer=2 filter=242 channel=121
					-6, -9, 8, -11, 0, -7, -8, 0, 5,
					-- layer=2 filter=242 channel=122
					-4, 2, -2, -4, -7, 0, 4, -2, 6,
					-- layer=2 filter=242 channel=123
					29, -13, -6, 7, 19, -17, -43, -23, -19,
					-- layer=2 filter=242 channel=124
					9, -2, 18, 28, 13, -12, -12, -35, -2,
					-- layer=2 filter=242 channel=125
					11, -6, 3, 0, 9, -9, -8, -9, -4,
					-- layer=2 filter=242 channel=126
					1, -3, 8, 8, 15, -10, -9, -9, 10,
					-- layer=2 filter=242 channel=127
					-7, -33, 14, 0, 13, -20, 1, -2, -26,
					-- layer=2 filter=243 channel=0
					2, 4, -10, 0, -4, -13, -6, -6, 0,
					-- layer=2 filter=243 channel=1
					4, -1, 3, 0, -11, -1, -6, -14, -12,
					-- layer=2 filter=243 channel=2
					0, 5, 9, -3, 0, 2, 7, 2, 0,
					-- layer=2 filter=243 channel=3
					0, -10, 0, -5, -2, -8, 1, -10, 2,
					-- layer=2 filter=243 channel=4
					1, -12, 6, -7, 4, 8, -1, -5, 6,
					-- layer=2 filter=243 channel=5
					5, 2, -11, -4, -11, -7, -6, 0, 4,
					-- layer=2 filter=243 channel=6
					-11, 3, -10, 0, 6, -13, 0, 1, -9,
					-- layer=2 filter=243 channel=7
					-11, -5, 5, 5, -4, -1, -6, 10, 1,
					-- layer=2 filter=243 channel=8
					7, 0, -6, 0, -9, 5, 5, -9, 4,
					-- layer=2 filter=243 channel=9
					-5, -5, 7, -8, 3, 7, -8, -7, -6,
					-- layer=2 filter=243 channel=10
					-7, 6, 1, 5, 1, -1, -4, -7, -2,
					-- layer=2 filter=243 channel=11
					-3, 3, -7, 6, -1, 5, -2, -6, 6,
					-- layer=2 filter=243 channel=12
					-10, -4, -7, -1, 0, 2, -4, 3, 3,
					-- layer=2 filter=243 channel=13
					-7, 5, -3, -3, 4, -8, -7, 8, 6,
					-- layer=2 filter=243 channel=14
					-13, -8, 9, -5, -9, 5, -5, -4, 3,
					-- layer=2 filter=243 channel=15
					4, -10, 3, 0, -2, -3, 5, -6, -2,
					-- layer=2 filter=243 channel=16
					-6, 3, 1, -13, 2, 6, 0, 8, -8,
					-- layer=2 filter=243 channel=17
					10, 7, 0, -4, -3, -4, -8, 0, 4,
					-- layer=2 filter=243 channel=18
					-5, 2, -12, -9, 6, -10, 0, 1, 0,
					-- layer=2 filter=243 channel=19
					10, -7, -5, -7, -10, -6, -4, -4, 0,
					-- layer=2 filter=243 channel=20
					6, -4, -6, -7, 4, -4, -10, 6, 2,
					-- layer=2 filter=243 channel=21
					1, 7, -10, -1, 2, -2, -9, 3, -8,
					-- layer=2 filter=243 channel=22
					4, -9, 0, 0, 7, -2, 0, -1, -8,
					-- layer=2 filter=243 channel=23
					-6, 7, 9, 3, 4, 5, -7, -1, 8,
					-- layer=2 filter=243 channel=24
					6, -8, -11, 1, -2, 6, 0, -5, -1,
					-- layer=2 filter=243 channel=25
					-5, -5, 3, 7, -7, 3, -7, 7, 0,
					-- layer=2 filter=243 channel=26
					3, 9, 3, 0, 6, -9, -1, 8, 4,
					-- layer=2 filter=243 channel=27
					-3, 1, -6, 1, -2, -9, 0, -7, -5,
					-- layer=2 filter=243 channel=28
					-9, 0, -7, 1, -3, -3, -13, 6, -7,
					-- layer=2 filter=243 channel=29
					3, -8, -4, 10, 3, 8, -2, -12, -1,
					-- layer=2 filter=243 channel=30
					-7, -11, 7, 2, -10, -10, -4, 4, -5,
					-- layer=2 filter=243 channel=31
					6, 0, 1, 6, -8, -5, -4, -2, 7,
					-- layer=2 filter=243 channel=32
					1, -3, 0, 6, 0, 7, -9, -8, 9,
					-- layer=2 filter=243 channel=33
					2, -2, 3, 4, 3, -7, 4, -2, -6,
					-- layer=2 filter=243 channel=34
					3, 9, -6, -10, -6, -12, 0, -7, -11,
					-- layer=2 filter=243 channel=35
					9, -6, 5, 3, 6, -7, 2, -8, -9,
					-- layer=2 filter=243 channel=36
					-8, 3, -3, 0, -10, 7, 5, 7, -6,
					-- layer=2 filter=243 channel=37
					-1, 7, -1, 1, 0, -10, -10, -4, -3,
					-- layer=2 filter=243 channel=38
					8, 1, 1, 4, -10, 5, -12, -2, 0,
					-- layer=2 filter=243 channel=39
					4, 3, -10, 0, -8, 0, -5, -1, 8,
					-- layer=2 filter=243 channel=40
					4, 7, -12, 4, -6, 1, -5, 5, 6,
					-- layer=2 filter=243 channel=41
					0, -6, 9, 7, 2, 6, 5, 0, -6,
					-- layer=2 filter=243 channel=42
					-7, 3, 1, 6, -7, -5, 5, 6, -4,
					-- layer=2 filter=243 channel=43
					0, 2, -8, -2, -12, -14, 1, 1, -4,
					-- layer=2 filter=243 channel=44
					5, -10, -9, -6, -5, 4, -7, -4, 2,
					-- layer=2 filter=243 channel=45
					-10, -5, 9, -9, -1, 0, -4, 4, 0,
					-- layer=2 filter=243 channel=46
					-9, 3, 6, 0, 2, 0, -5, -8, 2,
					-- layer=2 filter=243 channel=47
					3, 0, -1, -3, 1, -12, -5, -5, -1,
					-- layer=2 filter=243 channel=48
					0, 2, 9, -5, 11, -9, 4, -8, 9,
					-- layer=2 filter=243 channel=49
					-1, -11, -8, 1, 3, 0, -1, -6, 8,
					-- layer=2 filter=243 channel=50
					11, -8, 3, 6, 11, 4, -1, -3, -1,
					-- layer=2 filter=243 channel=51
					10, -5, -4, 2, 0, -9, -2, -11, 4,
					-- layer=2 filter=243 channel=52
					8, -2, -12, -5, 1, -8, -9, -9, -11,
					-- layer=2 filter=243 channel=53
					-3, -5, 1, 5, -10, -6, 0, 4, -11,
					-- layer=2 filter=243 channel=54
					-8, -1, -1, 0, 0, 0, 3, 4, -4,
					-- layer=2 filter=243 channel=55
					9, -9, 8, -5, -6, 8, 3, -3, 1,
					-- layer=2 filter=243 channel=56
					3, -10, -7, -6, -9, -7, -12, -8, 3,
					-- layer=2 filter=243 channel=57
					0, 3, 4, -10, 0, 5, 5, 2, 0,
					-- layer=2 filter=243 channel=58
					-10, 8, 6, -9, 7, -10, 0, -4, -3,
					-- layer=2 filter=243 channel=59
					-2, 10, -11, -7, -4, 4, -7, -10, 6,
					-- layer=2 filter=243 channel=60
					-5, 3, -11, 4, -4, -4, 6, -1, 2,
					-- layer=2 filter=243 channel=61
					4, -10, 3, -3, 6, 1, -3, 4, 9,
					-- layer=2 filter=243 channel=62
					-6, -4, -4, 9, -10, 8, -14, -10, -9,
					-- layer=2 filter=243 channel=63
					0, -10, 0, -15, 7, 2, -14, 1, -4,
					-- layer=2 filter=243 channel=64
					6, -5, -8, -7, -9, 5, -8, -7, 7,
					-- layer=2 filter=243 channel=65
					7, -9, 0, -10, 8, 4, -8, -7, -9,
					-- layer=2 filter=243 channel=66
					-9, 3, -1, 6, -4, 5, 10, -8, -3,
					-- layer=2 filter=243 channel=67
					-4, -3, 0, -2, -1, -3, -7, -5, 7,
					-- layer=2 filter=243 channel=68
					-5, -6, -6, -4, 8, -6, -2, 2, 1,
					-- layer=2 filter=243 channel=69
					-8, 0, 0, -3, 7, -7, -9, 2, 10,
					-- layer=2 filter=243 channel=70
					-3, -6, -3, -8, 5, 2, -1, -12, -9,
					-- layer=2 filter=243 channel=71
					2, 0, 0, -4, 0, -4, -4, -8, -5,
					-- layer=2 filter=243 channel=72
					0, -9, -9, 0, -5, 0, 0, -2, -10,
					-- layer=2 filter=243 channel=73
					-2, -7, 5, 5, 0, -8, -5, 2, -5,
					-- layer=2 filter=243 channel=74
					-1, 5, -5, 4, -3, -11, -1, -5, -6,
					-- layer=2 filter=243 channel=75
					0, -6, 1, 8, -5, -3, 5, 2, -9,
					-- layer=2 filter=243 channel=76
					-10, 7, 0, 1, 0, -4, 8, 2, 8,
					-- layer=2 filter=243 channel=77
					-3, -1, 6, -4, 3, -4, -2, -8, -1,
					-- layer=2 filter=243 channel=78
					3, -3, 1, -1, -6, -7, 0, -2, -12,
					-- layer=2 filter=243 channel=79
					-4, -8, -5, -2, -5, -9, 5, -3, -4,
					-- layer=2 filter=243 channel=80
					6, -1, -11, 3, -8, 1, -14, -14, -4,
					-- layer=2 filter=243 channel=81
					4, -4, -8, -6, 0, -2, 6, 0, -6,
					-- layer=2 filter=243 channel=82
					-3, -3, 10, -4, 4, 0, 6, 5, 0,
					-- layer=2 filter=243 channel=83
					-16, -3, 2, 5, -7, -8, 4, -13, 7,
					-- layer=2 filter=243 channel=84
					9, 5, 3, 8, -4, 10, 5, -4, -2,
					-- layer=2 filter=243 channel=85
					0, -7, 3, 9, -4, -3, 0, 10, 0,
					-- layer=2 filter=243 channel=86
					-10, -5, -8, 0, -9, -4, -4, 10, 6,
					-- layer=2 filter=243 channel=87
					-3, -3, -8, -11, -16, 0, -7, -8, 6,
					-- layer=2 filter=243 channel=88
					-13, -11, 5, 1, 0, 0, -8, -3, -3,
					-- layer=2 filter=243 channel=89
					-15, 1, -6, 7, 10, -8, -7, 8, -2,
					-- layer=2 filter=243 channel=90
					-4, -9, 1, 5, -6, -2, 5, -9, 0,
					-- layer=2 filter=243 channel=91
					4, -12, -2, -8, -5, 0, 1, -9, 7,
					-- layer=2 filter=243 channel=92
					1, 11, -6, 0, 5, 4, -12, -8, -11,
					-- layer=2 filter=243 channel=93
					8, -10, -3, 0, 7, -4, -5, 8, -7,
					-- layer=2 filter=243 channel=94
					1, 12, -14, 7, -2, 1, -10, -3, 5,
					-- layer=2 filter=243 channel=95
					-10, -8, -5, 3, -8, 0, 2, 1, 6,
					-- layer=2 filter=243 channel=96
					0, -6, -11, 4, 3, 1, -8, 0, -5,
					-- layer=2 filter=243 channel=97
					-13, -3, -9, 0, -9, -6, 5, 2, -3,
					-- layer=2 filter=243 channel=98
					-6, 9, -9, 3, 2, 0, 6, 6, -4,
					-- layer=2 filter=243 channel=99
					0, -1, -4, 3, -6, -12, 6, 3, -11,
					-- layer=2 filter=243 channel=100
					-2, -11, -3, -9, 1, 4, -7, -3, 8,
					-- layer=2 filter=243 channel=101
					-1, -6, -10, -6, -2, -5, 0, 1, -4,
					-- layer=2 filter=243 channel=102
					1, -4, 1, -2, 2, -7, 2, -5, 4,
					-- layer=2 filter=243 channel=103
					-8, -7, 0, 0, -8, -9, -4, -2, -10,
					-- layer=2 filter=243 channel=104
					-3, 1, -2, -9, -4, -5, 0, -5, -2,
					-- layer=2 filter=243 channel=105
					3, 0, 3, -1, -6, -5, -1, 6, -9,
					-- layer=2 filter=243 channel=106
					3, -6, -2, 1, -9, 5, -11, -4, -9,
					-- layer=2 filter=243 channel=107
					10, -3, 1, -2, 6, 0, -7, -6, 4,
					-- layer=2 filter=243 channel=108
					1, 12, 0, 1, 6, -7, 2, 10, -7,
					-- layer=2 filter=243 channel=109
					-2, -8, -9, -9, -2, 0, -3, 4, 5,
					-- layer=2 filter=243 channel=110
					-18, -9, 3, -4, -8, 9, -2, -11, -5,
					-- layer=2 filter=243 channel=111
					-5, -6, 2, 0, -8, -1, 6, 5, -8,
					-- layer=2 filter=243 channel=112
					-12, 0, 1, -2, 6, -11, -2, -4, 3,
					-- layer=2 filter=243 channel=113
					2, -11, -1, -7, -10, -6, -10, -6, -4,
					-- layer=2 filter=243 channel=114
					-8, 0, -4, -5, -8, 2, 9, 5, 7,
					-- layer=2 filter=243 channel=115
					5, 1, 0, 10, 1, -6, -8, 0, 6,
					-- layer=2 filter=243 channel=116
					-8, -6, 0, 7, 3, 3, 0, 6, -8,
					-- layer=2 filter=243 channel=117
					4, 3, -3, 0, -16, 1, -3, -1, 0,
					-- layer=2 filter=243 channel=118
					6, 0, 4, 4, 4, 0, 6, 1, 4,
					-- layer=2 filter=243 channel=119
					-2, 4, 4, -7, -2, 2, -10, -10, 3,
					-- layer=2 filter=243 channel=120
					2, 9, 10, 8, -1, 2, 7, 7, 0,
					-- layer=2 filter=243 channel=121
					11, 1, 4, 9, -3, 1, 2, -4, 10,
					-- layer=2 filter=243 channel=122
					0, 7, -9, 0, 3, 1, 5, -2, -9,
					-- layer=2 filter=243 channel=123
					-7, 4, 4, -5, 2, -14, 5, 2, -3,
					-- layer=2 filter=243 channel=124
					-3, -7, -1, -11, 6, -8, -6, -2, 3,
					-- layer=2 filter=243 channel=125
					0, 4, 0, -8, 5, 1, 5, -6, -9,
					-- layer=2 filter=243 channel=126
					-9, 7, -3, -1, -10, -3, 6, 3, 5,
					-- layer=2 filter=243 channel=127
					-16, -4, 0, -11, -12, 3, -2, 2, -1,
					-- layer=2 filter=244 channel=0
					-10, -10, -37, -3, 16, -29, 17, 34, 5,
					-- layer=2 filter=244 channel=1
					-5, -14, 28, 30, 12, 7, 24, -9, 5,
					-- layer=2 filter=244 channel=2
					-6, -5, -9, -5, -4, 8, 7, -1, -11,
					-- layer=2 filter=244 channel=3
					-9, 10, 29, -3, -11, -23, 21, 10, -15,
					-- layer=2 filter=244 channel=4
					45, 35, 5, -27, -34, 31, -42, -67, -15,
					-- layer=2 filter=244 channel=5
					28, -10, -34, 9, 7, -14, -1, 18, -4,
					-- layer=2 filter=244 channel=6
					-12, 4, -42, -42, -18, 7, -35, -48, 0,
					-- layer=2 filter=244 channel=7
					-4, -5, -44, -71, -56, -28, 15, -34, -5,
					-- layer=2 filter=244 channel=8
					-1, -4, 7, 2, 3, -7, 9, -10, 0,
					-- layer=2 filter=244 channel=9
					-20, 22, 35, -1, 1, 9, -3, -11, -30,
					-- layer=2 filter=244 channel=10
					-22, -7, -2, -7, 9, 1, 9, 32, -3,
					-- layer=2 filter=244 channel=11
					15, 2, -12, 27, 13, 4, 24, 8, -1,
					-- layer=2 filter=244 channel=12
					9, 33, 38, 7, 15, 2, 0, -15, -21,
					-- layer=2 filter=244 channel=13
					0, -1, -1, -12, -8, 1, 1, 0, 1,
					-- layer=2 filter=244 channel=14
					8, 4, 29, 35, 23, -3, -7, -21, -23,
					-- layer=2 filter=244 channel=15
					26, 15, -37, 59, 33, -1, 49, 45, 18,
					-- layer=2 filter=244 channel=16
					37, 26, 47, -29, -37, -3, -77, -89, -7,
					-- layer=2 filter=244 channel=17
					4, 3, 4, -9, -5, -4, 9, 5, 1,
					-- layer=2 filter=244 channel=18
					27, 14, -6, 18, -39, 22, -8, -50, -24,
					-- layer=2 filter=244 channel=19
					-11, -39, -23, 17, -24, 4, -4, -27, -16,
					-- layer=2 filter=244 channel=20
					3, 7, 0, -9, -3, 2, 9, -1, -5,
					-- layer=2 filter=244 channel=21
					13, 12, 13, 7, 0, 20, -6, -1, 10,
					-- layer=2 filter=244 channel=22
					8, 3, 9, 7, 7, -5, 7, -9, 0,
					-- layer=2 filter=244 channel=23
					48, 29, 44, -18, -10, -16, -34, -50, -28,
					-- layer=2 filter=244 channel=24
					0, 17, 42, -39, 30, 43, -30, 7, 16,
					-- layer=2 filter=244 channel=25
					16, 27, 36, -10, 15, 19, 0, 9, 6,
					-- layer=2 filter=244 channel=26
					11, -2, -1, -8, -3, 0, -3, -7, -4,
					-- layer=2 filter=244 channel=27
					1, 19, 10, 20, 15, -4, 23, 14, 1,
					-- layer=2 filter=244 channel=28
					15, 0, -19, 35, -39, -89, -37, -27, -33,
					-- layer=2 filter=244 channel=29
					8, 2, -11, -6, 7, 6, -4, 0, 5,
					-- layer=2 filter=244 channel=30
					7, -4, 35, 28, -18, 0, -34, -38, -12,
					-- layer=2 filter=244 channel=31
					44, 12, -50, -48, -2, -23, -30, -32, -47,
					-- layer=2 filter=244 channel=32
					7, -3, 1, -4, 4, -10, -3, 9, 9,
					-- layer=2 filter=244 channel=33
					8, 35, -37, 38, 10, -39, 24, -40, 0,
					-- layer=2 filter=244 channel=34
					47, 35, 3, 59, -7, -19, 33, -35, -16,
					-- layer=2 filter=244 channel=35
					33, -7, -29, 15, -18, -76, -17, -19, -6,
					-- layer=2 filter=244 channel=36
					-3, 1, 3, -5, -1, -19, 1, -8, -6,
					-- layer=2 filter=244 channel=37
					-6, -3, -33, 26, 20, -3, 31, 18, -9,
					-- layer=2 filter=244 channel=38
					4, 1, 0, 23, 10, -15, 9, -17, -25,
					-- layer=2 filter=244 channel=39
					37, 43, 40, 16, -15, -44, 7, -44, -21,
					-- layer=2 filter=244 channel=40
					48, 54, -11, 37, -2, -52, 31, 19, 46,
					-- layer=2 filter=244 channel=41
					4, 8, -9, 9, 3, 0, -8, -8, 12,
					-- layer=2 filter=244 channel=42
					47, 18, 27, -17, 6, 21, -64, -43, 1,
					-- layer=2 filter=244 channel=43
					-13, -2, -50, 17, 14, -68, 32, 0, -37,
					-- layer=2 filter=244 channel=44
					-6, 1, 5, -1, 6, 6, -2, -3, -2,
					-- layer=2 filter=244 channel=45
					2, -8, -22, -18, -11, 19, -3, -33, -23,
					-- layer=2 filter=244 channel=46
					-2, -47, -24, -12, -42, -24, 12, 1, -3,
					-- layer=2 filter=244 channel=47
					38, 40, -15, 4, -40, -52, -18, -1, -27,
					-- layer=2 filter=244 channel=48
					-8, 8, 0, 2, 4, -7, 4, -5, -6,
					-- layer=2 filter=244 channel=49
					12, -31, 9, 22, -27, 48, -26, -29, -15,
					-- layer=2 filter=244 channel=50
					-3, -7, -11, -8, 0, -12, 16, -5, -3,
					-- layer=2 filter=244 channel=51
					0, -2, -21, 24, 19, -24, 26, 10, 7,
					-- layer=2 filter=244 channel=52
					-12, -23, -27, 24, 9, -3, 33, -8, -2,
					-- layer=2 filter=244 channel=53
					-29, -39, -104, 15, -11, 11, -36, 7, 5,
					-- layer=2 filter=244 channel=54
					27, -6, -33, 3, -24, 8, -2, -17, 22,
					-- layer=2 filter=244 channel=55
					6, 13, 0, 6, -3, 12, -10, -2, 1,
					-- layer=2 filter=244 channel=56
					-10, 1, 0, 33, 12, -9, 14, 11, -3,
					-- layer=2 filter=244 channel=57
					8, 0, 8, -2, -10, 12, 1, 1, 6,
					-- layer=2 filter=244 channel=58
					31, 2, 37, 0, 12, -33, -8, -17, -36,
					-- layer=2 filter=244 channel=59
					-15, 0, -9, 31, 37, -35, 25, -7, 5,
					-- layer=2 filter=244 channel=60
					2, 17, -29, 14, 10, 5, -12, -30, 44,
					-- layer=2 filter=244 channel=61
					-53, -21, -53, -30, 3, -26, -34, -26, 5,
					-- layer=2 filter=244 channel=62
					19, -4, -40, -22, -39, 3, 9, -64, 15,
					-- layer=2 filter=244 channel=63
					6, 51, 18, 17, -15, -32, -25, -4, -31,
					-- layer=2 filter=244 channel=64
					-3, 18, 56, -18, -36, -30, -75, -73, -34,
					-- layer=2 filter=244 channel=65
					-44, -25, -21, -32, -1, -7, -36, -29, 11,
					-- layer=2 filter=244 channel=66
					14, -62, -13, -8, -38, -28, 2, -58, 46,
					-- layer=2 filter=244 channel=67
					7, 1, 7, 15, -22, -17, 11, -22, -29,
					-- layer=2 filter=244 channel=68
					-3, -11, -11, -11, -6, -8, -7, 0, -3,
					-- layer=2 filter=244 channel=69
					16, 27, 54, 0, 7, 3, -72, -39, -13,
					-- layer=2 filter=244 channel=70
					13, -28, -19, 30, -16, -46, 0, -19, -20,
					-- layer=2 filter=244 channel=71
					-5, 23, -27, 25, 11, 6, 31, 16, -22,
					-- layer=2 filter=244 channel=72
					8, -8, 2, 39, 25, 35, 43, -1, -2,
					-- layer=2 filter=244 channel=73
					34, 17, 5, -27, -23, 56, 4, -4, 4,
					-- layer=2 filter=244 channel=74
					17, 29, 27, -1, -43, -49, -42, -51, -32,
					-- layer=2 filter=244 channel=75
					13, -26, -10, -11, -28, -7, -10, -37, 35,
					-- layer=2 filter=244 channel=76
					51, 5, 14, 9, 17, 20, -75, -27, 11,
					-- layer=2 filter=244 channel=77
					-3, -2, 7, -7, 1, 6, 8, -4, 6,
					-- layer=2 filter=244 channel=78
					1, 3, -6, -11, 14, 23, -6, 9, 0,
					-- layer=2 filter=244 channel=79
					-10, 0, -5, -6, 0, -7, 0, 3, 1,
					-- layer=2 filter=244 channel=80
					26, 2, 2, -47, -50, -11, -57, -32, -33,
					-- layer=2 filter=244 channel=81
					8, -10, -3, -8, 5, 1, -6, -2, -5,
					-- layer=2 filter=244 channel=82
					8, 5, 5, 8, 3, 6, 6, 2, 4,
					-- layer=2 filter=244 channel=83
					46, 13, 29, -11, 0, 9, -46, 6, -16,
					-- layer=2 filter=244 channel=84
					5, 4, 9, -3, -4, 7, 7, -6, 0,
					-- layer=2 filter=244 channel=85
					0, -7, -1, -8, -6, 6, 11, 3, -7,
					-- layer=2 filter=244 channel=86
					-6, -10, -2, -14, -1, 5, 0, 3, 0,
					-- layer=2 filter=244 channel=87
					6, 7, 12, 7, 8, -20, -33, -7, 40,
					-- layer=2 filter=244 channel=88
					5, 45, 28, 22, -11, -11, -51, -72, -27,
					-- layer=2 filter=244 channel=89
					6, 1, 24, 21, 40, -3, 16, -2, 0,
					-- layer=2 filter=244 channel=90
					1, 10, 10, 0, -8, 6, 3, 0, -4,
					-- layer=2 filter=244 channel=91
					29, 26, -3, 19, 18, -2, -8, -23, 34,
					-- layer=2 filter=244 channel=92
					-3, 21, 11, 31, 40, 23, 12, 5, 20,
					-- layer=2 filter=244 channel=93
					-51, 72, -7, -84, -13, -71, 1, 2, -40,
					-- layer=2 filter=244 channel=94
					-32, -44, -50, -24, -37, 59, -25, 0, 1,
					-- layer=2 filter=244 channel=95
					-5, -2, -12, -8, -7, -16, -7, -4, -4,
					-- layer=2 filter=244 channel=96
					-12, -9, -56, -44, -22, -27, -3, -15, -35,
					-- layer=2 filter=244 channel=97
					23, 30, 11, -32, -14, -19, -33, -25, -29,
					-- layer=2 filter=244 channel=98
					17, 5, -7, 41, -6, -32, 5, 13, -16,
					-- layer=2 filter=244 channel=99
					4, -39, -42, -5, 4, -36, -1, 26, 7,
					-- layer=2 filter=244 channel=100
					47, 35, 34, -14, 25, -5, -31, -23, 4,
					-- layer=2 filter=244 channel=101
					4, 14, -2, 31, 25, -33, 12, 31, -2,
					-- layer=2 filter=244 channel=102
					-1, 10, -11, 4, -36, 9, 18, -32, -31,
					-- layer=2 filter=244 channel=103
					-15, 6, -16, -33, -49, 0, -17, 2, 15,
					-- layer=2 filter=244 channel=104
					-1, -67, -39, 5, -48, 79, -19, 3, 4,
					-- layer=2 filter=244 channel=105
					-32, -22, -36, -29, 9, -5, -48, -47, -9,
					-- layer=2 filter=244 channel=106
					-6, -9, 27, -7, 25, -16, -9, 7, 4,
					-- layer=2 filter=244 channel=107
					25, -29, 26, -6, 16, 19, -17, 7, 4,
					-- layer=2 filter=244 channel=108
					-24, 13, -3, 13, 10, -2, 16, 0, 8,
					-- layer=2 filter=244 channel=109
					-5, 8, 7, -10, -8, -3, -3, -6, 0,
					-- layer=2 filter=244 channel=110
					12, 19, 59, -1, -6, 11, -59, -38, -28,
					-- layer=2 filter=244 channel=111
					-8, 4, -4, -7, -9, 5, 0, 8, 6,
					-- layer=2 filter=244 channel=112
					6, -19, -32, 3, 50, -23, 27, 13, 27,
					-- layer=2 filter=244 channel=113
					-22, -11, 34, -21, -26, -35, -39, -10, -9,
					-- layer=2 filter=244 channel=114
					23, -7, 2, 0, 12, 5, 12, 4, 2,
					-- layer=2 filter=244 channel=115
					6, 2, 8, 9, 14, 0, 1, -8, 0,
					-- layer=2 filter=244 channel=116
					32, 22, -12, 45, -14, -31, -21, -8, -2,
					-- layer=2 filter=244 channel=117
					6, 23, -22, -18, 9, 21, 44, -16, 0,
					-- layer=2 filter=244 channel=118
					-18, -32, -33, -27, -4, 9, 12, -22, -18,
					-- layer=2 filter=244 channel=119
					58, -1, 33, -6, -77, -13, -31, -68, -47,
					-- layer=2 filter=244 channel=120
					-2, -3, 7, -8, 8, -3, -9, 0, -9,
					-- layer=2 filter=244 channel=121
					7, 3, 1, 0, -4, 5, -4, 7, 4,
					-- layer=2 filter=244 channel=122
					-4, 1, 1, -14, 13, 8, 13, 5, -3,
					-- layer=2 filter=244 channel=123
					16, 1, -23, -4, 11, -40, 22, -15, -14,
					-- layer=2 filter=244 channel=124
					50, 4, -2, -14, 9, -34, 26, -15, 5,
					-- layer=2 filter=244 channel=125
					-8, -4, 2, 3, 1, -13, -4, 1, 0,
					-- layer=2 filter=244 channel=126
					-10, -64, -11, -49, -6, -32, 17, -5, -28,
					-- layer=2 filter=244 channel=127
					16, -9, 55, 6, 70, -14, -9, -37, 0,
					-- layer=2 filter=245 channel=0
					-22, -21, -32, -6, -13, -22, -7, -19, -7,
					-- layer=2 filter=245 channel=1
					28, 1, 9, -4, 34, 13, -18, -18, 4,
					-- layer=2 filter=245 channel=2
					-2, -1, -9, 6, 0, 6, -11, 0, 8,
					-- layer=2 filter=245 channel=3
					-34, -22, -42, -39, -42, -20, -21, 23, -26,
					-- layer=2 filter=245 channel=4
					14, 7, -5, -16, 9, -4, -30, 4, -2,
					-- layer=2 filter=245 channel=5
					-45, -14, -36, 8, -24, 1, -48, -7, -36,
					-- layer=2 filter=245 channel=6
					41, 12, -54, 30, 8, -38, 28, 54, 28,
					-- layer=2 filter=245 channel=7
					-6, 19, 5, -51, 4, -52, -65, -69, -1,
					-- layer=2 filter=245 channel=8
					-8, 0, 0, 6, -8, 4, 1, -8, -5,
					-- layer=2 filter=245 channel=9
					14, -16, -8, 22, -1, -10, 17, 15, 4,
					-- layer=2 filter=245 channel=10
					0, -19, -9, -36, 5, -19, -40, 1, -16,
					-- layer=2 filter=245 channel=11
					-9, -17, -69, -20, -16, -47, -36, -41, -40,
					-- layer=2 filter=245 channel=12
					17, 0, 12, 12, 20, -8, -53, -18, 8,
					-- layer=2 filter=245 channel=13
					-1, -5, 0, -7, -7, -10, -2, 8, 5,
					-- layer=2 filter=245 channel=14
					6, -5, 17, 2, 21, -2, -20, -19, -23,
					-- layer=2 filter=245 channel=15
					-33, -31, 2, -1, -17, -21, 11, -33, 13,
					-- layer=2 filter=245 channel=16
					12, 9, 1, 15, 12, 32, 18, -2, -2,
					-- layer=2 filter=245 channel=17
					-10, 3, -9, -7, -4, 4, 1, -4, 3,
					-- layer=2 filter=245 channel=18
					-3, -24, -28, -1, -2, -13, -9, -53, -9,
					-- layer=2 filter=245 channel=19
					-6, 17, 0, 43, 18, 11, 15, 41, 19,
					-- layer=2 filter=245 channel=20
					-2, 4, -3, 8, -2, -7, -1, 7, -10,
					-- layer=2 filter=245 channel=21
					5, 9, 14, 1, -4, -9, -3, 1, -1,
					-- layer=2 filter=245 channel=22
					-11, -2, -2, -3, 3, 8, 3, -3, 5,
					-- layer=2 filter=245 channel=23
					1, -3, -16, 11, 10, 9, -9, -14, -15,
					-- layer=2 filter=245 channel=24
					-8, 26, -37, -58, -40, -26, -11, -2, 27,
					-- layer=2 filter=245 channel=25
					-25, 21, -15, -63, -15, -76, -31, -26, 25,
					-- layer=2 filter=245 channel=26
					8, 0, 2, 0, 9, 0, -8, 7, 5,
					-- layer=2 filter=245 channel=27
					10, 16, 21, -5, 7, -12, -16, -23, -13,
					-- layer=2 filter=245 channel=28
					18, 28, -1, 30, 33, -6, -59, -6, -22,
					-- layer=2 filter=245 channel=29
					-8, 5, 10, 4, 2, -8, 0, -7, -8,
					-- layer=2 filter=245 channel=30
					7, -4, 18, -13, 0, 22, 19, -6, -20,
					-- layer=2 filter=245 channel=31
					39, 72, 66, 22, -14, -16, 32, 3, 60,
					-- layer=2 filter=245 channel=32
					-3, -11, 2, -3, 4, 4, 5, 5, 0,
					-- layer=2 filter=245 channel=33
					2, -32, -7, -14, -10, -26, -55, -13, -21,
					-- layer=2 filter=245 channel=34
					-32, 33, 15, 18, 13, 11, -8, 5, 6,
					-- layer=2 filter=245 channel=35
					-10, 9, 11, -15, -3, -19, -67, -23, -54,
					-- layer=2 filter=245 channel=36
					0, -5, 7, 11, -3, 13, -13, -9, 0,
					-- layer=2 filter=245 channel=37
					1, -27, -32, -23, -32, -41, -29, -36, -8,
					-- layer=2 filter=245 channel=38
					16, -19, 21, -6, 7, 19, -27, -9, 3,
					-- layer=2 filter=245 channel=39
					0, 29, 24, -9, -12, 17, -3, -3, 1,
					-- layer=2 filter=245 channel=40
					-3, 11, -39, -14, 37, -30, -3, 14, 35,
					-- layer=2 filter=245 channel=41
					-4, -5, 2, 2, -9, 8, 2, -4, -11,
					-- layer=2 filter=245 channel=42
					3, -2, 22, -12, 20, -1, -4, -6, 8,
					-- layer=2 filter=245 channel=43
					-24, -39, -73, -36, -49, -23, -35, -10, 0,
					-- layer=2 filter=245 channel=44
					-7, 8, 8, 9, 5, -4, 4, -6, -7,
					-- layer=2 filter=245 channel=45
					8, 37, 32, -2, 11, -5, 5, 25, 2,
					-- layer=2 filter=245 channel=46
					1, -2, 13, 7, -15, -8, 11, -6, -8,
					-- layer=2 filter=245 channel=47
					11, 19, -33, -16, 8, -40, -37, -41, -38,
					-- layer=2 filter=245 channel=48
					-11, -9, 1, -8, 8, -8, -8, -8, 9,
					-- layer=2 filter=245 channel=49
					-17, -37, -9, -2, -8, -35, -28, 0, 18,
					-- layer=2 filter=245 channel=50
					14, 10, 11, 1, 7, -9, 10, 2, -13,
					-- layer=2 filter=245 channel=51
					-22, -38, -40, -28, -19, -7, -47, -36, -10,
					-- layer=2 filter=245 channel=52
					36, 1, 42, 27, 31, -22, 14, -20, -21,
					-- layer=2 filter=245 channel=53
					-46, 27, -13, -33, -3, -37, -31, -6, -31,
					-- layer=2 filter=245 channel=54
					22, -5, -19, -3, 17, -11, -4, -44, -6,
					-- layer=2 filter=245 channel=55
					0, -5, -2, -2, 3, 7, -3, 5, 1,
					-- layer=2 filter=245 channel=56
					-24, -2, -58, -22, -16, -76, -35, -46, -38,
					-- layer=2 filter=245 channel=57
					7, -1, -2, -2, -3, 1, 18, 24, 13,
					-- layer=2 filter=245 channel=58
					1, -7, 18, 5, 37, -10, -37, -26, -17,
					-- layer=2 filter=245 channel=59
					35, -11, 24, -9, 31, 23, -35, 26, -16,
					-- layer=2 filter=245 channel=60
					19, -7, 15, 20, 38, 40, -39, -1, 9,
					-- layer=2 filter=245 channel=61
					2, -17, 5, -19, -36, -9, -68, -22, 8,
					-- layer=2 filter=245 channel=62
					18, 29, -14, -8, 18, 0, 1, 15, 15,
					-- layer=2 filter=245 channel=63
					20, 1, -25, 11, 8, 14, -21, -9, 24,
					-- layer=2 filter=245 channel=64
					5, 18, 27, 27, 7, 5, 32, -6, -27,
					-- layer=2 filter=245 channel=65
					2, -23, 29, 16, 10, -30, -31, -6, 26,
					-- layer=2 filter=245 channel=66
					-13, 7, -28, 28, -2, -31, -21, 30, 0,
					-- layer=2 filter=245 channel=67
					11, 3, -26, -14, -10, -32, 4, 31, -17,
					-- layer=2 filter=245 channel=68
					0, 7, 4, 0, -2, 3, -8, 8, -10,
					-- layer=2 filter=245 channel=69
					3, 6, 0, 7, 0, 27, 24, 7, -23,
					-- layer=2 filter=245 channel=70
					4, 6, 13, 6, -1, -36, -49, -39, -38,
					-- layer=2 filter=245 channel=71
					-1, -2, 29, -2, 17, 2, 7, 10, -7,
					-- layer=2 filter=245 channel=72
					-9, 5, 19, 11, 14, 0, -1, -1, 20,
					-- layer=2 filter=245 channel=73
					-2, 22, 7, -27, -55, -37, 2, 50, 44,
					-- layer=2 filter=245 channel=74
					35, 12, 16, -5, 9, 23, -12, 11, -48,
					-- layer=2 filter=245 channel=75
					6, -7, -28, 7, 8, 0, 45, 25, 19,
					-- layer=2 filter=245 channel=76
					11, 13, -41, 1, -57, -59, -2, -38, -67,
					-- layer=2 filter=245 channel=77
					-11, -4, -1, -6, -3, -2, 1, -5, 7,
					-- layer=2 filter=245 channel=78
					1, -2, -42, -33, -19, -55, -19, -24, -19,
					-- layer=2 filter=245 channel=79
					11, 4, -1, 4, -1, -6, -7, -8, 5,
					-- layer=2 filter=245 channel=80
					12, -2, -3, -1, -18, 8, -7, 16, -2,
					-- layer=2 filter=245 channel=81
					-7, -24, -7, -19, -19, -14, -4, -18, -11,
					-- layer=2 filter=245 channel=82
					-12, 0, 0, -2, -1, 2, 11, -2, -2,
					-- layer=2 filter=245 channel=83
					-7, 13, 27, 7, 17, 1, -22, 4, -40,
					-- layer=2 filter=245 channel=84
					2, -1, 8, -8, 7, -6, -3, -1, 7,
					-- layer=2 filter=245 channel=85
					-2, 3, -9, -1, 5, 6, -6, -4, 15,
					-- layer=2 filter=245 channel=86
					2, -7, 0, 16, 6, 6, 13, 16, -10,
					-- layer=2 filter=245 channel=87
					27, 16, -7, 46, 61, -25, 74, 5, 43,
					-- layer=2 filter=245 channel=88
					19, 14, 3, 0, 19, 7, -17, 9, -29,
					-- layer=2 filter=245 channel=89
					17, 17, 22, 13, 40, 8, -21, -5, 2,
					-- layer=2 filter=245 channel=90
					-8, -9, 7, -5, -8, 4, -9, -11, -1,
					-- layer=2 filter=245 channel=91
					-9, 10, 12, 17, 24, 17, -33, -5, 37,
					-- layer=2 filter=245 channel=92
					-4, 4, 18, 7, 33, 12, -35, -11, 17,
					-- layer=2 filter=245 channel=93
					33, 19, 28, 41, 39, -48, 4, 54, 32,
					-- layer=2 filter=245 channel=94
					21, 6, -52, -43, -2, -8, -13, 46, 34,
					-- layer=2 filter=245 channel=95
					-10, -3, 9, -3, 3, 8, -5, 5, 2,
					-- layer=2 filter=245 channel=96
					-5, -17, -28, 24, 8, 7, 18, 38, -4,
					-- layer=2 filter=245 channel=97
					20, -3, -20, 12, -19, -12, 18, -5, -33,
					-- layer=2 filter=245 channel=98
					1, 19, -17, 13, 16, -33, -67, -51, 1,
					-- layer=2 filter=245 channel=99
					32, -18, 7, 66, 25, -33, 8, 26, -61,
					-- layer=2 filter=245 channel=100
					25, -20, 26, 19, 24, 12, -21, -1, -23,
					-- layer=2 filter=245 channel=101
					-16, 10, 36, -35, -32, -59, -31, 0, -14,
					-- layer=2 filter=245 channel=102
					-14, -24, -21, 0, 11, -8, 9, 4, 26,
					-- layer=2 filter=245 channel=103
					-42, -6, 13, -29, 24, -15, -54, -20, -1,
					-- layer=2 filter=245 channel=104
					-3, -2, -51, -38, -5, -59, -22, 13, -20,
					-- layer=2 filter=245 channel=105
					0, 7, -2, 14, 51, -29, 13, -18, -10,
					-- layer=2 filter=245 channel=106
					-15, -23, -39, -33, -42, -43, -35, -19, 2,
					-- layer=2 filter=245 channel=107
					-13, 20, 20, 5, 9, -17, 20, 33, 58,
					-- layer=2 filter=245 channel=108
					0, 0, -5, 27, 28, -6, 10, 15, 9,
					-- layer=2 filter=245 channel=109
					27, -15, -9, 6, -6, -2, 17, 12, -2,
					-- layer=2 filter=245 channel=110
					0, 19, 21, 11, -2, -20, 32, 30, -12,
					-- layer=2 filter=245 channel=111
					-6, -6, -11, -5, -10, -7, -1, -8, -4,
					-- layer=2 filter=245 channel=112
					-56, -70, -30, -63, -66, -21, -25, -51, -8,
					-- layer=2 filter=245 channel=113
					-8, -14, 47, 6, 5, 12, 18, -18, 0,
					-- layer=2 filter=245 channel=114
					12, 6, -2, -2, 0, 6, -12, 16, 9,
					-- layer=2 filter=245 channel=115
					-4, -3, -2, -1, 1, -1, -3, 2, -4,
					-- layer=2 filter=245 channel=116
					3, -12, -8, 43, 65, -9, 42, 18, 17,
					-- layer=2 filter=245 channel=117
					-12, -7, -49, -43, -11, -49, 0, -24, 15,
					-- layer=2 filter=245 channel=118
					-14, -27, -54, -25, -61, -9, -4, -29, -6,
					-- layer=2 filter=245 channel=119
					-5, -11, -38, -17, 0, 13, 6, -30, -29,
					-- layer=2 filter=245 channel=120
					-1, 8, 7, -4, 10, -2, -9, -4, -4,
					-- layer=2 filter=245 channel=121
					-7, -6, -8, -7, 0, 5, 3, 8, 3,
					-- layer=2 filter=245 channel=122
					-16, -13, -3, -6, -8, 11, 1, 5, -6,
					-- layer=2 filter=245 channel=123
					28, 26, 1, -3, 23, 4, -2, -20, -3,
					-- layer=2 filter=245 channel=124
					10, -29, 7, -27, -6, -25, 11, -8, 12,
					-- layer=2 filter=245 channel=125
					4, 8, 10, 8, -7, -8, 13, 4, -5,
					-- layer=2 filter=245 channel=126
					-2, 0, 19, -50, -20, -9, -26, 100, -17,
					-- layer=2 filter=245 channel=127
					32, 0, 32, 20, 6, 3, -10, 9, -3,
					-- layer=2 filter=246 channel=0
					-3, -24, 14, -17, 11, 29, -25, 0, 12,
					-- layer=2 filter=246 channel=1
					4, 0, -3, 14, 35, 3, 0, -32, -37,
					-- layer=2 filter=246 channel=2
					-6, 2, -10, -9, 1, -10, 2, -4, -9,
					-- layer=2 filter=246 channel=3
					-10, 14, 34, -5, 8, 24, 52, 66, 48,
					-- layer=2 filter=246 channel=4
					18, -61, -32, 1, -1, -41, -24, -42, -57,
					-- layer=2 filter=246 channel=5
					-37, -23, -14, 2, -10, 12, 8, 12, 14,
					-- layer=2 filter=246 channel=6
					-12, 19, 61, -17, -24, 24, -54, -97, -14,
					-- layer=2 filter=246 channel=7
					-22, -33, -2, 9, -6, -6, -22, -41, -60,
					-- layer=2 filter=246 channel=8
					-7, -4, 3, 5, -13, -6, -3, 2, -1,
					-- layer=2 filter=246 channel=9
					-43, -35, -58, -5, 7, -29, 10, 3, -4,
					-- layer=2 filter=246 channel=10
					-1, 13, 0, 23, 10, 43, 15, 34, 41,
					-- layer=2 filter=246 channel=11
					-12, -8, 6, -27, 16, 12, -12, 12, 7,
					-- layer=2 filter=246 channel=12
					-13, -38, -57, -1, -13, -22, -19, 13, 16,
					-- layer=2 filter=246 channel=13
					8, -8, 10, 1, 2, -3, 1, -1, -6,
					-- layer=2 filter=246 channel=14
					-17, -33, -25, 11, -1, 9, -20, 7, -1,
					-- layer=2 filter=246 channel=15
					92, 25, 48, 13, 38, 62, 50, 19, 45,
					-- layer=2 filter=246 channel=16
					28, 29, -6, 14, 6, -30, -17, -36, -14,
					-- layer=2 filter=246 channel=17
					-4, 7, -3, -6, 4, -1, 0, -7, 3,
					-- layer=2 filter=246 channel=18
					30, -6, 19, 1, 24, 20, 21, 19, 8,
					-- layer=2 filter=246 channel=19
					51, 21, 27, 2, 24, -12, 4, -19, -34,
					-- layer=2 filter=246 channel=20
					4, 1, -3, -10, 0, 2, -8, -7, -4,
					-- layer=2 filter=246 channel=21
					-7, -1, -12, 20, 15, -2, 19, 7, 5,
					-- layer=2 filter=246 channel=22
					1, -3, -2, -3, 5, 3, 7, 5, -2,
					-- layer=2 filter=246 channel=23
					26, -2, -8, 41, 7, -4, 0, -26, -46,
					-- layer=2 filter=246 channel=24
					-11, -12, 20, -23, -2, 4, 8, 17, 39,
					-- layer=2 filter=246 channel=25
					-23, 6, 39, -15, -9, -3, -17, -3, 21,
					-- layer=2 filter=246 channel=26
					-10, -1, 1, 1, -9, 9, -8, 4, 11,
					-- layer=2 filter=246 channel=27
					18, -31, -48, 32, -28, -39, 32, 20, 16,
					-- layer=2 filter=246 channel=28
					-9, 14, -7, 12, 11, -1, -12, 16, 2,
					-- layer=2 filter=246 channel=29
					-8, 3, -2, 6, -7, -8, 7, -9, -9,
					-- layer=2 filter=246 channel=30
					-6, -19, -20, -16, -51, -84, -3, -3, -7,
					-- layer=2 filter=246 channel=31
					-21, -42, -33, 8, -33, 26, -30, -12, 15,
					-- layer=2 filter=246 channel=32
					9, -3, -2, 2, 6, 3, 10, -1, 5,
					-- layer=2 filter=246 channel=33
					-18, -45, -13, 0, 24, 8, 20, 28, 0,
					-- layer=2 filter=246 channel=34
					25, -16, -2, -25, -11, -1, -21, -39, -50,
					-- layer=2 filter=246 channel=35
					13, 21, -4, 8, 4, -4, 3, 8, 4,
					-- layer=2 filter=246 channel=36
					-11, 11, 8, 13, 10, -8, 11, 6, 19,
					-- layer=2 filter=246 channel=37
					7, 7, 9, -14, -13, -11, 10, 18, 2,
					-- layer=2 filter=246 channel=38
					0, -44, -57, 11, -29, -33, 3, 9, 8,
					-- layer=2 filter=246 channel=39
					31, -19, -30, 42, -21, -32, -12, -31, -15,
					-- layer=2 filter=246 channel=40
					22, 21, 9, 14, -18, 22, 1, 50, 33,
					-- layer=2 filter=246 channel=41
					9, -2, 1, -7, 6, 7, 8, -3, 0,
					-- layer=2 filter=246 channel=42
					37, -4, 14, 18, -20, -22, 13, 10, 36,
					-- layer=2 filter=246 channel=43
					20, 27, 10, 5, 36, 27, 21, 38, 29,
					-- layer=2 filter=246 channel=44
					10, 2, -4, -8, -7, 5, 6, -2, -9,
					-- layer=2 filter=246 channel=45
					-3, -14, -26, 27, 16, -34, 71, 26, 29,
					-- layer=2 filter=246 channel=46
					-12, -22, -41, 0, -6, -20, -33, -10, -21,
					-- layer=2 filter=246 channel=47
					-46, -22, -2, 25, 16, 1, 1, 10, -8,
					-- layer=2 filter=246 channel=48
					8, 6, -4, 6, 8, 10, -2, -9, -5,
					-- layer=2 filter=246 channel=49
					45, -16, 36, -11, 5, 18, 32, -11, 37,
					-- layer=2 filter=246 channel=50
					31, 28, 42, 10, 19, 33, 15, 24, 27,
					-- layer=2 filter=246 channel=51
					-17, 9, 23, -21, -4, 14, -28, -4, -5,
					-- layer=2 filter=246 channel=52
					20, 19, 54, -29, -4, -26, 18, 16, -13,
					-- layer=2 filter=246 channel=53
					31, -24, 16, 5, -4, 4, -51, 18, -30,
					-- layer=2 filter=246 channel=54
					16, 20, 35, 28, 20, 33, -30, -17, -1,
					-- layer=2 filter=246 channel=55
					0, 6, -6, -2, 2, -6, -10, -6, 1,
					-- layer=2 filter=246 channel=56
					-11, -15, -12, -9, -9, 14, -14, 21, 20,
					-- layer=2 filter=246 channel=57
					-15, 0, -3, -9, 4, 4, 1, -2, 5,
					-- layer=2 filter=246 channel=58
					-16, -29, -36, 12, -27, -38, -37, -2, -6,
					-- layer=2 filter=246 channel=59
					13, 2, 27, 16, -32, -44, 33, -47, -1,
					-- layer=2 filter=246 channel=60
					5, 3, 2, 0, -14, -33, -72, -76, -16,
					-- layer=2 filter=246 channel=61
					18, -4, 25, 29, 12, -6, -12, -39, 32,
					-- layer=2 filter=246 channel=62
					0, -17, 25, -16, -37, 19, -33, -81, -11,
					-- layer=2 filter=246 channel=63
					-29, -15, -13, 38, -3, 6, -3, -18, -7,
					-- layer=2 filter=246 channel=64
					24, 18, 7, 23, 9, -2, 36, -6, 31,
					-- layer=2 filter=246 channel=65
					2, 0, 28, 2, -18, 1, -50, -45, -20,
					-- layer=2 filter=246 channel=66
					-26, 19, 12, 40, 26, 2, 23, 37, 22,
					-- layer=2 filter=246 channel=67
					-22, -16, -16, 39, 0, -12, -16, -22, -29,
					-- layer=2 filter=246 channel=68
					-7, 2, -5, -7, 3, 5, 10, -6, 0,
					-- layer=2 filter=246 channel=69
					25, 14, 5, 29, 5, -17, 2, 6, 41,
					-- layer=2 filter=246 channel=70
					-2, -3, -2, 5, 9, 15, -7, 10, -13,
					-- layer=2 filter=246 channel=71
					-12, -15, -24, 0, -13, -6, 30, -12, -7,
					-- layer=2 filter=246 channel=72
					-38, -30, 2, -12, -22, -14, -21, -22, -16,
					-- layer=2 filter=246 channel=73
					60, 55, 22, 52, 63, 32, 9, 34, 38,
					-- layer=2 filter=246 channel=74
					-22, -23, -44, 3, 18, -7, -22, 5, -13,
					-- layer=2 filter=246 channel=75
					5, 0, -7, 11, -12, 11, -58, -55, -61,
					-- layer=2 filter=246 channel=76
					69, -17, 0, 16, -13, -10, -36, -40, -14,
					-- layer=2 filter=246 channel=77
					3, 1, 4, 9, -6, 2, 0, -9, -7,
					-- layer=2 filter=246 channel=78
					-10, 28, 33, -19, 10, 17, 6, 0, 16,
					-- layer=2 filter=246 channel=79
					-3, 0, -4, 2, 3, -11, 7, 1, 6,
					-- layer=2 filter=246 channel=80
					8, -1, -9, -5, -17, -5, 17, 0, -6,
					-- layer=2 filter=246 channel=81
					18, 9, -1, 0, 19, -5, 10, 4, 11,
					-- layer=2 filter=246 channel=82
					8, 9, -3, 1, 4, -13, -3, 11, 12,
					-- layer=2 filter=246 channel=83
					6, -4, -16, 32, -25, -52, 6, -3, -33,
					-- layer=2 filter=246 channel=84
					5, -7, -4, 1, -1, -5, -8, 5, 9,
					-- layer=2 filter=246 channel=85
					16, 8, -7, 21, 4, -1, -14, -6, -5,
					-- layer=2 filter=246 channel=86
					1, 1, 12, -11, 12, -3, 20, -10, 10,
					-- layer=2 filter=246 channel=87
					10, -3, 11, -14, -18, 6, -32, -24, -27,
					-- layer=2 filter=246 channel=88
					-21, -6, -13, 9, -16, -37, 13, 5, 23,
					-- layer=2 filter=246 channel=89
					16, -10, 8, -12, -20, -20, -26, -30, -16,
					-- layer=2 filter=246 channel=90
					8, 5, -2, 8, -11, -3, -8, -7, 1,
					-- layer=2 filter=246 channel=91
					23, 13, -10, 4, -11, -30, -16, -2, -4,
					-- layer=2 filter=246 channel=92
					4, -3, -34, -22, -6, -35, 4, 16, 0,
					-- layer=2 filter=246 channel=93
					37, 14, -4, 55, 2, -27, -46, -46, -32,
					-- layer=2 filter=246 channel=94
					21, 7, 56, 11, 14, -27, -20, -46, 4,
					-- layer=2 filter=246 channel=95
					15, 19, 8, -6, -1, -5, 8, 15, 9,
					-- layer=2 filter=246 channel=96
					0, 19, 25, 15, -24, -20, -48, -39, -116,
					-- layer=2 filter=246 channel=97
					-27, -24, -4, -13, 6, -18, 10, 22, 22,
					-- layer=2 filter=246 channel=98
					-24, 2, 3, 5, 1, 3, -4, 14, 12,
					-- layer=2 filter=246 channel=99
					97, 43, 29, 16, 25, -41, 20, -18, -8,
					-- layer=2 filter=246 channel=100
					8, -24, -33, 32, -55, -44, 16, -4, -8,
					-- layer=2 filter=246 channel=101
					-18, 23, 16, -36, -9, 14, -13, 1, 10,
					-- layer=2 filter=246 channel=102
					-2, 39, -1, 34, 11, -23, 10, -11, -52,
					-- layer=2 filter=246 channel=103
					19, 46, -39, -28, -1, 30, -35, 19, -40,
					-- layer=2 filter=246 channel=104
					13, -3, 36, 30, 8, 14, 5, 9, 1,
					-- layer=2 filter=246 channel=105
					31, -12, -47, -24, -55, -39, -2, -85, 25,
					-- layer=2 filter=246 channel=106
					2, -11, 3, -3, -14, 10, -10, 0, 12,
					-- layer=2 filter=246 channel=107
					71, -9, 4, 41, 18, 61, 31, 25, 30,
					-- layer=2 filter=246 channel=108
					-8, 10, -13, 0, -30, -32, 34, 5, -6,
					-- layer=2 filter=246 channel=109
					1, 12, 19, -1, -4, 0, 3, -16, 11,
					-- layer=2 filter=246 channel=110
					35, 0, 18, 28, -11, -12, 25, -16, 15,
					-- layer=2 filter=246 channel=111
					-10, 12, 0, -8, 1, -7, 0, -6, -9,
					-- layer=2 filter=246 channel=112
					-5, 0, -1, -4, -7, 18, -18, -12, 41,
					-- layer=2 filter=246 channel=113
					-25, -42, -19, 8, -27, -53, 1, 3, 6,
					-- layer=2 filter=246 channel=114
					17, 9, 1, -8, 13, 0, -8, -7, 6,
					-- layer=2 filter=246 channel=115
					0, -3, 4, -4, -5, 3, 6, -13, 2,
					-- layer=2 filter=246 channel=116
					36, 6, 3, 7, 1, -5, -5, -22, -52,
					-- layer=2 filter=246 channel=117
					13, 30, 29, 59, 51, 25, 23, -8, -2,
					-- layer=2 filter=246 channel=118
					2, 31, 26, -1, 24, 28, 34, 20, 24,
					-- layer=2 filter=246 channel=119
					37, -37, -40, 19, -38, -26, 21, -18, -10,
					-- layer=2 filter=246 channel=120
					-4, 8, -5, 0, 2, 1, -7, -7, -9,
					-- layer=2 filter=246 channel=121
					3, 6, -6, -8, 8, -2, 0, -9, 0,
					-- layer=2 filter=246 channel=122
					6, 4, 11, 2, 15, -2, -6, 10, 6,
					-- layer=2 filter=246 channel=123
					-7, -8, 15, 26, 15, -10, -29, -61, -49,
					-- layer=2 filter=246 channel=124
					66, 20, 17, 46, 73, 57, 19, -11, -2,
					-- layer=2 filter=246 channel=125
					1, 1, -5, -4, -4, 2, -5, 3, 6,
					-- layer=2 filter=246 channel=126
					15, -12, -10, -39, 0, 41, -31, 24, -24,
					-- layer=2 filter=246 channel=127
					-15, -14, -17, -8, -7, -26, 27, 2, -18,
					-- layer=2 filter=247 channel=0
					1, -11, 3, -19, 5, -9, -9, -10, -1,
					-- layer=2 filter=247 channel=1
					-52, 35, 17, -10, 4, 28, 23, 11, -23,
					-- layer=2 filter=247 channel=2
					9, 0, 7, 7, -8, 0, 12, 8, 0,
					-- layer=2 filter=247 channel=3
					26, 16, 1, 13, -8, -44, 2, 4, 30,
					-- layer=2 filter=247 channel=4
					-13, 28, -3, 0, 47, -59, -16, -8, -40,
					-- layer=2 filter=247 channel=5
					-22, -23, -5, -52, -16, 13, -11, -25, 5,
					-- layer=2 filter=247 channel=6
					-42, -10, -68, -9, 6, -7, 6, -28, 31,
					-- layer=2 filter=247 channel=7
					7, 29, 6, 6, -23, -2, -15, 11, 8,
					-- layer=2 filter=247 channel=8
					0, 0, 0, -7, 0, -1, 9, -5, -4,
					-- layer=2 filter=247 channel=9
					30, 33, -5, -4, 5, -28, 28, -23, -26,
					-- layer=2 filter=247 channel=10
					-6, 8, -2, 20, 6, -46, -13, -19, -4,
					-- layer=2 filter=247 channel=11
					4, -14, -18, -15, -26, -9, 1, -8, 10,
					-- layer=2 filter=247 channel=12
					-25, 15, -5, 0, 5, 34, 0, 19, -13,
					-- layer=2 filter=247 channel=13
					2, 5, 2, -1, 0, -2, -1, -2, 3,
					-- layer=2 filter=247 channel=14
					-36, -9, 1, -36, -20, -11, 5, -12, -25,
					-- layer=2 filter=247 channel=15
					-14, 19, 18, 9, 40, 42, 56, 23, -16,
					-- layer=2 filter=247 channel=16
					4, 49, -32, -27, -48, -84, -48, -55, -24,
					-- layer=2 filter=247 channel=17
					-6, 1, 8, 0, -6, 2, -6, -4, -7,
					-- layer=2 filter=247 channel=18
					19, 29, -5, 4, 40, -11, -11, 6, 19,
					-- layer=2 filter=247 channel=19
					-42, 22, -21, -1, 22, 36, 3, -4, -8,
					-- layer=2 filter=247 channel=20
					-7, 0, 2, -7, 8, 12, 7, -7, -7,
					-- layer=2 filter=247 channel=21
					-6, 0, 19, 0, 0, -7, 19, 10, 8,
					-- layer=2 filter=247 channel=22
					-9, -4, -7, -1, 0, -2, 0, -10, 0,
					-- layer=2 filter=247 channel=23
					-41, 10, -23, 0, 18, 6, -9, -21, -21,
					-- layer=2 filter=247 channel=24
					42, 16, 6, 24, -12, -14, -10, -1, 13,
					-- layer=2 filter=247 channel=25
					22, -9, -7, -6, -13, -24, 13, -14, 14,
					-- layer=2 filter=247 channel=26
					-8, -8, 3, 7, -8, -3, -14, -2, 0,
					-- layer=2 filter=247 channel=27
					-63, -51, 6, -92, -48, 28, -63, 16, 30,
					-- layer=2 filter=247 channel=28
					-45, 6, -4, 12, 34, 2, 28, 20, 24,
					-- layer=2 filter=247 channel=29
					-3, -10, 0, 9, 6, 12, 11, -2, -1,
					-- layer=2 filter=247 channel=30
					10, 13, 6, 0, 11, 9, -40, -14, -40,
					-- layer=2 filter=247 channel=31
					-11, 20, 29, -31, 13, 80, 16, 37, -16,
					-- layer=2 filter=247 channel=32
					0, 11, -7, -7, -6, -5, 3, -3, 8,
					-- layer=2 filter=247 channel=33
					-27, 37, 87, -44, -21, -3, -13, 23, 28,
					-- layer=2 filter=247 channel=34
					0, 23, 29, -24, 36, 24, 5, 12, 0,
					-- layer=2 filter=247 channel=35
					-2, -13, -11, 13, 27, 3, 6, -3, 27,
					-- layer=2 filter=247 channel=36
					7, -3, -6, -2, -9, -3, -1, 2, -2,
					-- layer=2 filter=247 channel=37
					-19, -14, -2, -28, -15, 17, 0, 13, 8,
					-- layer=2 filter=247 channel=38
					-55, -40, 20, -59, -2, 47, -43, 10, 13,
					-- layer=2 filter=247 channel=39
					3, 34, -15, -11, 7, -10, -18, -17, 29,
					-- layer=2 filter=247 channel=40
					18, -81, 23, 25, 58, 57, 5, 31, 12,
					-- layer=2 filter=247 channel=41
					-2, 9, 0, -8, -2, -2, 1, 4, 0,
					-- layer=2 filter=247 channel=42
					14, 8, -29, 27, 9, 5, 22, -23, -26,
					-- layer=2 filter=247 channel=43
					0, 6, -40, 17, -25, 3, -24, -17, 44,
					-- layer=2 filter=247 channel=44
					0, -6, -5, -1, 2, -10, 9, -4, 0,
					-- layer=2 filter=247 channel=45
					-5, 41, -3, 1, 8, 10, 27, 41, 43,
					-- layer=2 filter=247 channel=46
					-1, 10, 17, 41, 21, 3, -41, -33, -39,
					-- layer=2 filter=247 channel=47
					-26, 8, 15, -1, -1, -28, 27, 35, -22,
					-- layer=2 filter=247 channel=48
					5, -3, 1, 12, 1, 0, -8, 8, 8,
					-- layer=2 filter=247 channel=49
					55, 46, -52, 41, 5, -10, -6, -22, -4,
					-- layer=2 filter=247 channel=50
					10, -10, 1, -13, 6, -5, -5, 2, -5,
					-- layer=2 filter=247 channel=51
					-9, -22, -2, -18, -40, -26, 0, -10, 20,
					-- layer=2 filter=247 channel=52
					-10, -16, 0, -19, 9, 17, -10, 27, 23,
					-- layer=2 filter=247 channel=53
					10, -36, -6, 3, 6, -18, -11, -38, 0,
					-- layer=2 filter=247 channel=54
					-37, 1, -7, -15, 24, 5, 4, 19, 18,
					-- layer=2 filter=247 channel=55
					11, 8, 0, 5, 1, 5, 2, 7, 5,
					-- layer=2 filter=247 channel=56
					0, -5, -28, -26, -36, -17, -12, 9, 12,
					-- layer=2 filter=247 channel=57
					3, -7, 8, 3, 10, 0, -6, 0, -5,
					-- layer=2 filter=247 channel=58
					-44, -28, 25, -22, 7, 43, 3, 18, 1,
					-- layer=2 filter=247 channel=59
					-53, -3, 34, -60, 12, 39, -37, -1, 46,
					-- layer=2 filter=247 channel=60
					-48, -13, 0, -45, 23, 73, -43, -11, 22,
					-- layer=2 filter=247 channel=61
					-88, -23, -8, -45, -28, -5, -22, -7, 40,
					-- layer=2 filter=247 channel=62
					21, 13, -40, -22, -6, -5, -7, -10, -27,
					-- layer=2 filter=247 channel=63
					-50, -15, -14, -36, 3, 8, -29, -7, 3,
					-- layer=2 filter=247 channel=64
					-2, 21, 9, -9, 23, -4, -8, -26, -27,
					-- layer=2 filter=247 channel=65
					-97, -26, -20, -47, -69, 28, -59, -12, 30,
					-- layer=2 filter=247 channel=66
					-18, -10, -22, 24, 24, 40, -9, -34, -30,
					-- layer=2 filter=247 channel=67
					-3, 21, 2, -6, 50, -8, -52, -13, -59,
					-- layer=2 filter=247 channel=68
					-2, -8, -7, 3, -1, 4, -4, -4, -9,
					-- layer=2 filter=247 channel=69
					8, 38, -10, 7, -10, -24, 26, -19, -18,
					-- layer=2 filter=247 channel=70
					-31, 14, 2, 15, 24, -12, -5, 6, 29,
					-- layer=2 filter=247 channel=71
					3, -5, -45, -42, -12, 2, -30, -14, 13,
					-- layer=2 filter=247 channel=72
					-26, 35, 65, -35, 9, -16, -10, 6, 7,
					-- layer=2 filter=247 channel=73
					53, 9, 34, 69, 51, 1, 71, 21, 12,
					-- layer=2 filter=247 channel=74
					-43, 1, 2, 3, 26, 6, -50, 9, -27,
					-- layer=2 filter=247 channel=75
					-40, -32, -53, 20, -28, 38, -52, 0, 7,
					-- layer=2 filter=247 channel=76
					-28, 41, 57, 0, 70, -50, 28, -6, 0,
					-- layer=2 filter=247 channel=77
					10, -7, -10, -5, 6, 5, -10, -10, -2,
					-- layer=2 filter=247 channel=78
					38, 14, -20, 10, -22, 0, 11, 11, 26,
					-- layer=2 filter=247 channel=79
					-5, 0, 6, -7, 6, -1, 12, -1, 2,
					-- layer=2 filter=247 channel=80
					-3, 41, -20, 52, 45, -40, -40, -33, -71,
					-- layer=2 filter=247 channel=81
					-4, 7, -3, 12, -2, 0, -8, 1, -1,
					-- layer=2 filter=247 channel=82
					9, -5, -9, 7, -9, -6, -8, 1, 5,
					-- layer=2 filter=247 channel=83
					-34, 1, -34, 0, 34, -2, -48, -11, -44,
					-- layer=2 filter=247 channel=84
					2, 1, -10, 6, 0, 2, -7, -5, 1,
					-- layer=2 filter=247 channel=85
					-5, -10, 5, -12, 9, 0, -5, 5, 5,
					-- layer=2 filter=247 channel=86
					-2, 0, -17, 3, 2, -12, 10, -2, -22,
					-- layer=2 filter=247 channel=87
					0, 30, 26, -13, 44, 36, 30, 64, 33,
					-- layer=2 filter=247 channel=88
					-63, 26, -1, -57, 0, -2, 4, 21, 1,
					-- layer=2 filter=247 channel=89
					-26, 21, 6, -47, -28, -8, 6, -22, -33,
					-- layer=2 filter=247 channel=90
					8, 2, 10, 0, 6, 3, 3, 9, -3,
					-- layer=2 filter=247 channel=91
					-20, -1, -26, -27, -17, 26, -8, 12, -3,
					-- layer=2 filter=247 channel=92
					-24, 16, 4, -6, 3, 40, 0, 24, -3,
					-- layer=2 filter=247 channel=93
					-22, 0, -45, 16, -54, 27, -46, -11, -37,
					-- layer=2 filter=247 channel=94
					-12, -21, -26, -9, -36, 8, -13, -50, 8,
					-- layer=2 filter=247 channel=95
					-13, -7, 0, 2, 0, 10, -11, -14, -8,
					-- layer=2 filter=247 channel=96
					-48, -33, -4, -13, -11, -1, 63, -5, -28,
					-- layer=2 filter=247 channel=97
					39, 37, 14, 24, 18, -15, 4, 10, -18,
					-- layer=2 filter=247 channel=98
					-22, -7, 16, 5, 5, 16, 13, 52, 29,
					-- layer=2 filter=247 channel=99
					-19, -20, -31, 12, -30, 10, 25, 23, 7,
					-- layer=2 filter=247 channel=100
					-26, -20, -17, 13, 1, 21, -59, -53, 6,
					-- layer=2 filter=247 channel=101
					25, -43, 5, -36, -40, -17, -53, -56, -8,
					-- layer=2 filter=247 channel=102
					7, -15, -15, 18, -7, -2, 36, -2, -9,
					-- layer=2 filter=247 channel=103
					27, 22, 4, 56, 12, 27, 21, -8, 16,
					-- layer=2 filter=247 channel=104
					33, 48, -64, 15, 17, 11, -15, 3, -8,
					-- layer=2 filter=247 channel=105
					22, 28, 11, -28, 56, -23, 11, 38, 40,
					-- layer=2 filter=247 channel=106
					-8, -23, 4, -40, -63, -27, -26, -47, -29,
					-- layer=2 filter=247 channel=107
					32, -1, -10, 68, 37, 23, 5, -26, -23,
					-- layer=2 filter=247 channel=108
					-19, -4, -25, -13, -9, -35, 4, 3, -11,
					-- layer=2 filter=247 channel=109
					7, -10, 10, 8, 5, 12, 2, 0, 12,
					-- layer=2 filter=247 channel=110
					-20, 10, -22, -43, -8, 0, -50, -19, -18,
					-- layer=2 filter=247 channel=111
					-3, 6, 7, -6, 5, -9, -4, 10, -1,
					-- layer=2 filter=247 channel=112
					-21, -13, -6, -11, -38, -23, -21, -7, 20,
					-- layer=2 filter=247 channel=113
					-5, -14, -17, 33, 11, 24, -31, -20, -10,
					-- layer=2 filter=247 channel=114
					-1, -6, -13, -1, -1, -10, -1, -4, -7,
					-- layer=2 filter=247 channel=115
					-9, -8, -11, 2, 7, 12, -9, 9, -5,
					-- layer=2 filter=247 channel=116
					-67, -11, 22, -15, 67, 34, 22, 49, 20,
					-- layer=2 filter=247 channel=117
					12, -3, -22, 16, -29, -35, 33, 19, 0,
					-- layer=2 filter=247 channel=118
					27, 38, 4, 30, 6, -31, -5, 14, 17,
					-- layer=2 filter=247 channel=119
					0, 17, -48, 0, -1, -55, -9, -27, -5,
					-- layer=2 filter=247 channel=120
					-3, 0, -5, 2, 1, 4, 6, -3, 8,
					-- layer=2 filter=247 channel=121
					-1, -1, -9, -7, 1, -8, -5, 0, -1,
					-- layer=2 filter=247 channel=122
					-6, 2, -12, 14, 5, -4, -14, 7, -1,
					-- layer=2 filter=247 channel=123
					-17, 27, 46, -6, -5, -9, 11, 40, 15,
					-- layer=2 filter=247 channel=124
					-3, 56, 27, 5, 23, 17, 45, 14, 5,
					-- layer=2 filter=247 channel=125
					8, -8, 2, 3, 3, -7, -8, -2, 3,
					-- layer=2 filter=247 channel=126
					9, -9, 116, 12, 46, 14, -14, -74, -1,
					-- layer=2 filter=247 channel=127
					-32, 4, -14, 0, 27, 9, 4, 2, 22,
					-- layer=2 filter=248 channel=0
					18, 8, 14, -46, -31, -23, -21, -19, 4,
					-- layer=2 filter=248 channel=1
					9, 10, 11, -18, -21, -5, -18, -36, 11,
					-- layer=2 filter=248 channel=2
					5, -1, 11, -5, -9, 2, 7, -6, -8,
					-- layer=2 filter=248 channel=3
					-51, -8, -3, -64, -12, -3, 48, 55, 55,
					-- layer=2 filter=248 channel=4
					8, -12, -6, -21, -37, -18, -3, 12, 22,
					-- layer=2 filter=248 channel=5
					1, 35, 17, 33, -14, 16, -18, -20, 2,
					-- layer=2 filter=248 channel=6
					95, 41, 24, 52, 47, 18, 17, 13, 16,
					-- layer=2 filter=248 channel=7
					-4, -35, -26, 0, -20, 6, 30, 24, 34,
					-- layer=2 filter=248 channel=8
					-3, -6, -5, 0, 0, -6, 4, -9, 8,
					-- layer=2 filter=248 channel=9
					-1, 18, 6, -18, 5, 22, -45, -16, 16,
					-- layer=2 filter=248 channel=10
					-15, 13, 18, -58, -38, -13, -10, 22, 19,
					-- layer=2 filter=248 channel=11
					36, 18, 1, 9, 4, 6, -7, -32, -23,
					-- layer=2 filter=248 channel=12
					17, 2, 25, 18, 12, 20, 16, -11, 4,
					-- layer=2 filter=248 channel=13
					-8, 0, -7, -2, -6, -6, 8, -1, 4,
					-- layer=2 filter=248 channel=14
					33, 11, 17, 3, -9, -9, -22, -42, -24,
					-- layer=2 filter=248 channel=15
					2, -10, 50, -12, -23, 22, -11, -25, -11,
					-- layer=2 filter=248 channel=16
					36, 9, 0, -35, -39, -11, -19, 19, 5,
					-- layer=2 filter=248 channel=17
					-7, -9, -1, -8, -9, 3, -8, -5, -2,
					-- layer=2 filter=248 channel=18
					5, -2, -29, 13, -9, -19, 30, 3, 14,
					-- layer=2 filter=248 channel=19
					-10, 33, 12, -3, -8, 3, 4, -47, -39,
					-- layer=2 filter=248 channel=20
					7, -5, 0, -10, -3, -7, -4, 7, 3,
					-- layer=2 filter=248 channel=21
					7, 0, 6, 10, -5, -7, -2, 4, -1,
					-- layer=2 filter=248 channel=22
					9, -7, 7, -7, -1, -5, -9, -9, 6,
					-- layer=2 filter=248 channel=23
					1, -42, 15, -50, -22, 2, 0, -10, 17,
					-- layer=2 filter=248 channel=24
					10, 24, -6, -55, -16, -24, 2, 6, -10,
					-- layer=2 filter=248 channel=25
					28, 43, -2, -12, 3, 25, -11, -9, -14,
					-- layer=2 filter=248 channel=26
					7, -9, 2, -4, 10, -7, 3, 3, 2,
					-- layer=2 filter=248 channel=27
					61, 37, 30, -1, -47, -38, -26, -68, -30,
					-- layer=2 filter=248 channel=28
					-96, -55, -11, -95, -46, 0, 12, 15, 27,
					-- layer=2 filter=248 channel=29
					6, -8, -4, -6, 6, -2, -5, 2, 1,
					-- layer=2 filter=248 channel=30
					2, 8, 19, -15, -20, 5, -4, -28, -11,
					-- layer=2 filter=248 channel=31
					-48, -59, -18, -88, -80, -11, -56, 14, 2,
					-- layer=2 filter=248 channel=32
					5, 7, -7, 6, 1, -7, -8, -5, -2,
					-- layer=2 filter=248 channel=33
					-27, -17, -8, -23, -28, -4, 9, 28, 22,
					-- layer=2 filter=248 channel=34
					-33, 40, -2, 41, -6, -5, -5, 29, -6,
					-- layer=2 filter=248 channel=35
					-82, -62, -7, -18, -59, -4, 17, 16, 18,
					-- layer=2 filter=248 channel=36
					0, 2, 0, 6, -7, 0, 5, 2, 16,
					-- layer=2 filter=248 channel=37
					39, 25, 9, 30, -12, 12, -14, -25, -27,
					-- layer=2 filter=248 channel=38
					42, 45, 48, 24, -30, -20, -17, -31, -27,
					-- layer=2 filter=248 channel=39
					-6, -1, 2, -27, -14, -15, 35, -19, -33,
					-- layer=2 filter=248 channel=40
					-8, 7, 29, -13, -12, -35, -23, 29, 0,
					-- layer=2 filter=248 channel=41
					0, -6, 5, -1, -8, 6, 9, 6, 4,
					-- layer=2 filter=248 channel=42
					-12, -14, 1, -3, -20, -26, 20, 30, 19,
					-- layer=2 filter=248 channel=43
					4, 32, 31, -22, -33, 15, 19, 17, 90,
					-- layer=2 filter=248 channel=44
					7, -8, 3, -5, 4, 0, -6, -11, -4,
					-- layer=2 filter=248 channel=45
					56, -8, 14, 14, -70, -29, 6, -26, 0,
					-- layer=2 filter=248 channel=46
					30, 31, 1, 4, -19, 14, -51, -5, 5,
					-- layer=2 filter=248 channel=47
					-22, 1, 18, -67, -68, -11, -20, 0, 21,
					-- layer=2 filter=248 channel=48
					-9, 7, -1, 3, 3, 1, 10, -6, 2,
					-- layer=2 filter=248 channel=49
					17, 25, -7, 24, -9, -8, -28, -33, -7,
					-- layer=2 filter=248 channel=50
					12, 0, 10, -4, -6, 1, -2, 6, -3,
					-- layer=2 filter=248 channel=51
					9, 2, -4, 7, -6, 8, -24, -20, -27,
					-- layer=2 filter=248 channel=52
					-5, -5, 0, 34, 7, 9, 58, -5, -8,
					-- layer=2 filter=248 channel=53
					30, 34, -10, -11, 16, -58, 5, 3, -43,
					-- layer=2 filter=248 channel=54
					-24, -34, -32, -3, -31, 26, -9, -11, -7,
					-- layer=2 filter=248 channel=55
					-6, -8, 9, -5, 2, 9, -11, -4, -11,
					-- layer=2 filter=248 channel=56
					51, 32, 14, 7, -3, -3, -8, -29, -16,
					-- layer=2 filter=248 channel=57
					14, 12, 10, -1, 9, 4, 1, -3, 9,
					-- layer=2 filter=248 channel=58
					34, -11, 45, 8, 7, 38, 31, -36, -7,
					-- layer=2 filter=248 channel=59
					38, -3, 27, -37, -22, -12, 17, -24, -20,
					-- layer=2 filter=248 channel=60
					22, 13, 7, 11, 3, -4, 4, -41, -51,
					-- layer=2 filter=248 channel=61
					29, -77, -40, -25, -36, -31, -10, -73, -96,
					-- layer=2 filter=248 channel=62
					32, -8, 5, 31, 40, 16, 5, -10, -7,
					-- layer=2 filter=248 channel=63
					8, -16, -7, -40, -48, -15, 5, -34, -17,
					-- layer=2 filter=248 channel=64
					-14, 18, 0, -13, 5, 5, 0, 11, 4,
					-- layer=2 filter=248 channel=65
					37, -29, 2, -1, -36, 9, -7, -26, -22,
					-- layer=2 filter=248 channel=66
					17, -4, -47, -6, 10, 37, 21, -20, -45,
					-- layer=2 filter=248 channel=67
					39, 36, 23, -10, -14, -1, -44, 16, 1,
					-- layer=2 filter=248 channel=68
					-1, 7, 5, 7, -7, -2, 9, -7, 5,
					-- layer=2 filter=248 channel=69
					33, 12, 12, -14, 0, -1, 5, 6, 16,
					-- layer=2 filter=248 channel=70
					-60, -2, -5, -7, -45, -15, 2, 0, -11,
					-- layer=2 filter=248 channel=71
					54, 46, 27, 0, -32, -51, -14, -43, -33,
					-- layer=2 filter=248 channel=72
					-13, 0, -4, 3, -11, 1, 25, 16, 28,
					-- layer=2 filter=248 channel=73
					-19, 46, -50, -48, -23, -27, -3, -8, -50,
					-- layer=2 filter=248 channel=74
					-12, 26, 12, -9, -12, -14, -31, -8, -12,
					-- layer=2 filter=248 channel=75
					-2, -18, 7, -19, 17, 27, -20, -33, 2,
					-- layer=2 filter=248 channel=76
					-32, -13, -32, 4, 43, 54, -38, -47, -29,
					-- layer=2 filter=248 channel=77
					-7, 3, 1, 0, 4, 2, 1, 4, 6,
					-- layer=2 filter=248 channel=78
					11, 1, 26, 17, 17, 21, 11, -6, 0,
					-- layer=2 filter=248 channel=79
					0, 2, -5, 0, 9, 2, 4, 8, -8,
					-- layer=2 filter=248 channel=80
					-9, 31, 10, -15, -17, 2, -23, 29, 41,
					-- layer=2 filter=248 channel=81
					8, 7, 3, 12, -2, 6, 12, -3, 4,
					-- layer=2 filter=248 channel=82
					-3, 11, 9, 4, 4, 8, 0, 4, -10,
					-- layer=2 filter=248 channel=83
					10, 9, -6, -40, -51, -40, -2, -12, -8,
					-- layer=2 filter=248 channel=84
					3, 1, 5, 4, -2, -6, 6, 5, -3,
					-- layer=2 filter=248 channel=85
					-3, 0, 10, 4, 11, 14, -9, 14, 11,
					-- layer=2 filter=248 channel=86
					7, 11, -8, 17, -6, -11, -12, 5, -14,
					-- layer=2 filter=248 channel=87
					34, -5, 33, 14, 52, -11, 5, -12, 50,
					-- layer=2 filter=248 channel=88
					12, 26, 16, -8, -3, 8, -36, -15, -6,
					-- layer=2 filter=248 channel=89
					25, 14, 34, 13, 16, 32, 12, -51, 9,
					-- layer=2 filter=248 channel=90
					-9, 5, 4, -8, -8, 0, 8, 3, 5,
					-- layer=2 filter=248 channel=91
					-10, 8, 28, 13, 13, 42, 7, -9, -4,
					-- layer=2 filter=248 channel=92
					26, 14, 9, 17, 8, 4, -2, -26, 12,
					-- layer=2 filter=248 channel=93
					-64, -36, -32, 3, -11, 18, 12, 35, 44,
					-- layer=2 filter=248 channel=94
					35, -13, -7, -12, 18, -3, 32, -16, -1,
					-- layer=2 filter=248 channel=95
					17, 16, 17, 0, 1, 11, 12, 14, -4,
					-- layer=2 filter=248 channel=96
					8, 8, -25, 17, 44, 20, -6, -16, 46,
					-- layer=2 filter=248 channel=97
					-10, 24, 7, -32, 2, 3, -11, 11, 3,
					-- layer=2 filter=248 channel=98
					-82, -60, -18, -44, -33, 3, -2, 8, -1,
					-- layer=2 filter=248 channel=99
					9, 16, -26, 52, 6, 6, 16, -64, -39,
					-- layer=2 filter=248 channel=100
					20, 18, 42, 2, -8, -2, 7, 4, 23,
					-- layer=2 filter=248 channel=101
					26, 19, -16, -14, 4, 31, -8, -27, 0,
					-- layer=2 filter=248 channel=102
					17, 6, -22, 37, 5, 6, 14, -7, -4,
					-- layer=2 filter=248 channel=103
					-7, 0, -6, 2, 18, -8, 0, -35, 27,
					-- layer=2 filter=248 channel=104
					56, -9, -5, -11, 16, -44, -18, -31, 3,
					-- layer=2 filter=248 channel=105
					-2, -17, 6, -62, 90, 34, -3, -65, -32,
					-- layer=2 filter=248 channel=106
					7, 10, 24, -46, -21, 40, -44, -37, 5,
					-- layer=2 filter=248 channel=107
					-17, -2, -34, 42, -10, -25, 12, -15, 57,
					-- layer=2 filter=248 channel=108
					28, 20, 4, 34, -26, -47, -4, -66, -7,
					-- layer=2 filter=248 channel=109
					9, 1, 8, 5, 9, -3, 10, -2, -12,
					-- layer=2 filter=248 channel=110
					4, 9, -8, -17, 21, -12, -3, 11, 4,
					-- layer=2 filter=248 channel=111
					-1, 9, 2, -1, -9, -5, 0, -7, 4,
					-- layer=2 filter=248 channel=112
					47, -21, 37, -13, -51, -1, -30, 20, 1,
					-- layer=2 filter=248 channel=113
					6, -31, 0, -47, -21, -20, -10, -33, -35,
					-- layer=2 filter=248 channel=114
					4, 1, -9, -3, 6, -8, -12, -6, 5,
					-- layer=2 filter=248 channel=115
					-4, -6, 10, 4, 9, -4, 5, 0, 3,
					-- layer=2 filter=248 channel=116
					39, 34, 43, 30, -2, 8, 17, -19, 48,
					-- layer=2 filter=248 channel=117
					-14, -12, -50, 8, -41, -9, 29, -14, -12,
					-- layer=2 filter=248 channel=118
					-13, 14, 21, -42, -30, -2, -2, 18, 37,
					-- layer=2 filter=248 channel=119
					20, 22, 6, 6, -73, -24, -23, 8, 34,
					-- layer=2 filter=248 channel=120
					-3, 8, 0, 4, 8, 10, -5, 1, 5,
					-- layer=2 filter=248 channel=121
					-3, -1, 0, 4, -3, -5, -3, -10, 0,
					-- layer=2 filter=248 channel=122
					0, -7, 4, 2, -13, 3, 3, -2, -7,
					-- layer=2 filter=248 channel=123
					7, -28, -26, -43, -25, -1, 27, 16, 4,
					-- layer=2 filter=248 channel=124
					-35, -28, 1, 13, 0, 35, 13, 40, 16,
					-- layer=2 filter=248 channel=125
					11, -2, -1, 0, -10, 4, -12, -2, -6,
					-- layer=2 filter=248 channel=126
					-4, -10, -34, -22, 49, 11, 34, 18, 42,
					-- layer=2 filter=248 channel=127
					22, -15, -2, -42, -26, -2, -23, -22, -8,
					-- layer=2 filter=249 channel=0
					8, 1, 0, -16, -2, 14, -14, 0, 1,
					-- layer=2 filter=249 channel=1
					10, 25, 6, -3, -4, 14, 10, -15, -18,
					-- layer=2 filter=249 channel=2
					3, -5, 0, -6, -2, 0, -4, -9, -2,
					-- layer=2 filter=249 channel=3
					-33, -14, 11, 0, 26, 14, 0, 20, 19,
					-- layer=2 filter=249 channel=4
					-2, 5, 13, -13, -46, -19, -26, -25, -7,
					-- layer=2 filter=249 channel=5
					12, 16, 7, -17, 9, -2, 3, 20, 2,
					-- layer=2 filter=249 channel=6
					-66, -1, -34, -50, -87, -77, -37, -50, -33,
					-- layer=2 filter=249 channel=7
					-41, 19, 2, -4, 5, -38, -14, -32, -14,
					-- layer=2 filter=249 channel=8
					-7, -1, -2, -1, 5, 4, -8, -7, 0,
					-- layer=2 filter=249 channel=9
					0, 3, 19, 12, -17, 6, 10, -1, -36,
					-- layer=2 filter=249 channel=10
					-9, -1, -4, -20, 31, 18, -24, 20, 10,
					-- layer=2 filter=249 channel=11
					2, 29, 14, 15, 10, 16, -4, 5, -2,
					-- layer=2 filter=249 channel=12
					10, 21, 3, 23, 22, 19, -6, -16, -1,
					-- layer=2 filter=249 channel=13
					-2, 4, 1, 8, -4, 5, -3, -3, -8,
					-- layer=2 filter=249 channel=14
					23, 9, 18, 6, 15, 32, 10, -6, 8,
					-- layer=2 filter=249 channel=15
					34, 40, 30, -8, 18, -23, -36, 4, 25,
					-- layer=2 filter=249 channel=16
					-15, -3, -27, -21, -16, -21, 30, 37, 10,
					-- layer=2 filter=249 channel=17
					-7, 9, 8, -5, -2, -1, -9, 8, 9,
					-- layer=2 filter=249 channel=18
					10, 20, 10, 10, -1, 22, 31, 1, 43,
					-- layer=2 filter=249 channel=19
					14, 7, 0, -5, -1, -9, -14, -36, -39,
					-- layer=2 filter=249 channel=20
					-6, 1, 8, 6, 3, 3, 6, 8, -5,
					-- layer=2 filter=249 channel=21
					4, -10, -11, -4, -9, -5, 15, 2, 8,
					-- layer=2 filter=249 channel=22
					-9, 6, 5, -7, -2, -9, -5, 3, -7,
					-- layer=2 filter=249 channel=23
					7, -7, -5, -3, -20, -12, 12, 8, 4,
					-- layer=2 filter=249 channel=24
					-8, -5, -2, 4, 36, 27, 24, 35, 22,
					-- layer=2 filter=249 channel=25
					-9, -3, 2, -10, 20, 13, -9, 15, 4,
					-- layer=2 filter=249 channel=26
					2, -4, 2, -9, 3, 10, 4, -8, -9,
					-- layer=2 filter=249 channel=27
					0, 7, 0, 6, 25, 0, -32, 1, 12,
					-- layer=2 filter=249 channel=28
					27, -17, 40, -9, -4, -15, -34, -53, 0,
					-- layer=2 filter=249 channel=29
					8, 7, 2, -7, 2, -6, -7, 6, 10,
					-- layer=2 filter=249 channel=30
					5, -11, -6, 5, -14, 0, 6, -1, -24,
					-- layer=2 filter=249 channel=31
					14, 23, -59, -7, 24, 1, 8, 39, -3,
					-- layer=2 filter=249 channel=32
					4, 1, -10, -5, -6, -9, 1, 0, 0,
					-- layer=2 filter=249 channel=33
					-34, -10, 1, 1, -5, -22, -36, -31, -11,
					-- layer=2 filter=249 channel=34
					16, -39, 3, 22, -13, -78, 46, -107, -24,
					-- layer=2 filter=249 channel=35
					7, 14, 3, -25, 2, -3, -14, -30, 0,
					-- layer=2 filter=249 channel=36
					0, 7, -6, 2, 5, -5, 0, -9, -1,
					-- layer=2 filter=249 channel=37
					-2, 1, 18, -15, 7, 5, 4, 14, 17,
					-- layer=2 filter=249 channel=38
					22, 25, 13, -3, -4, -4, -33, -15, -23,
					-- layer=2 filter=249 channel=39
					2, -5, -1, 23, 8, -18, 15, 28, 26,
					-- layer=2 filter=249 channel=40
					16, 32, 64, 8, -21, 10, -17, -8, 29,
					-- layer=2 filter=249 channel=41
					7, -7, 5, -4, 0, 3, -6, 4, -8,
					-- layer=2 filter=249 channel=42
					-17, -5, -19, -24, 10, 8, 16, 1, 22,
					-- layer=2 filter=249 channel=43
					-26, -32, -31, -5, -1, -4, -17, -3, 14,
					-- layer=2 filter=249 channel=44
					-10, 2, 5, -10, 4, -5, 6, -1, 2,
					-- layer=2 filter=249 channel=45
					13, 34, -2, -2, 19, 10, -20, 3, 18,
					-- layer=2 filter=249 channel=46
					7, -51, -10, -11, 10, -10, -13, -5, 0,
					-- layer=2 filter=249 channel=47
					37, 28, 26, 3, 1, 7, -19, 15, 42,
					-- layer=2 filter=249 channel=48
					-9, -6, 7, 0, -7, -9, 0, -10, -4,
					-- layer=2 filter=249 channel=49
					-16, 20, -25, 8, -15, 50, 55, 29, 47,
					-- layer=2 filter=249 channel=50
					-15, 3, 3, -4, -8, -3, 0, -1, 14,
					-- layer=2 filter=249 channel=51
					8, 25, 18, -4, 16, -11, 4, -1, 4,
					-- layer=2 filter=249 channel=52
					14, 35, 56, 3, 13, 2, -3, -37, -19,
					-- layer=2 filter=249 channel=53
					29, -9, -11, -10, -74, -50, -24, -52, -8,
					-- layer=2 filter=249 channel=54
					-12, 43, 14, -6, 21, -39, -30, -38, -33,
					-- layer=2 filter=249 channel=55
					9, 0, 10, 8, 2, 11, -1, -4, -10,
					-- layer=2 filter=249 channel=56
					-7, 13, 1, 6, 0, 16, -4, 8, 17,
					-- layer=2 filter=249 channel=57
					-13, -2, 4, -17, -7, 2, 3, 4, -3,
					-- layer=2 filter=249 channel=58
					1, 52, 4, 6, -2, 14, -4, -14, -12,
					-- layer=2 filter=249 channel=59
					6, 31, 7, 47, -15, -10, -21, -30, -19,
					-- layer=2 filter=249 channel=60
					46, 53, 14, 44, 30, -12, -15, 9, -2,
					-- layer=2 filter=249 channel=61
					18, 5, 27, 23, 14, -2, 26, 41, 35,
					-- layer=2 filter=249 channel=62
					-1, 1, 0, -2, -71, -25, 32, -69, 18,
					-- layer=2 filter=249 channel=63
					13, 2, 25, 10, 5, -31, -10, 17, 27,
					-- layer=2 filter=249 channel=64
					6, -7, -13, 11, 0, -11, 15, -2, -3,
					-- layer=2 filter=249 channel=65
					-2, 1, 0, -32, -24, -49, -22, -14, 10,
					-- layer=2 filter=249 channel=66
					-41, -14, 0, -20, -36, -7, 2, 7, 53,
					-- layer=2 filter=249 channel=67
					-2, -26, -36, -8, -25, -21, 2, -10, -59,
					-- layer=2 filter=249 channel=68
					7, -6, 8, 2, -10, 10, 4, 3, 4,
					-- layer=2 filter=249 channel=69
					-16, -9, 0, -1, -16, -3, 16, 12, 0,
					-- layer=2 filter=249 channel=70
					0, -1, 32, -7, 9, -12, -21, -20, -8,
					-- layer=2 filter=249 channel=71
					6, -16, -6, -8, 23, 0, -12, 28, -13,
					-- layer=2 filter=249 channel=72
					14, 0, 25, 13, 5, 5, -5, -42, 44,
					-- layer=2 filter=249 channel=73
					50, 7, 0, 20, 28, 17, 60, 71, 29,
					-- layer=2 filter=249 channel=74
					3, 25, -35, 5, -7, 14, -22, 8, -16,
					-- layer=2 filter=249 channel=75
					-6, -11, 0, -13, -26, 8, 6, 0, -5,
					-- layer=2 filter=249 channel=76
					42, 8, -7, 7, -65, -33, -37, -64, -25,
					-- layer=2 filter=249 channel=77
					2, 1, -6, 7, -2, 0, -1, 6, 6,
					-- layer=2 filter=249 channel=78
					4, 20, 13, 21, 6, 3, 0, -1, -3,
					-- layer=2 filter=249 channel=79
					-9, 3, 6, -3, 2, -1, -10, 8, 4,
					-- layer=2 filter=249 channel=80
					7, -21, -15, -7, 23, 15, 22, 25, 12,
					-- layer=2 filter=249 channel=81
					15, -3, 18, 17, 8, -1, 5, 6, -1,
					-- layer=2 filter=249 channel=82
					-11, -4, -5, 3, -2, -8, 7, -12, 4,
					-- layer=2 filter=249 channel=83
					14, -8, 25, 2, 6, -15, 5, 12, 0,
					-- layer=2 filter=249 channel=84
					1, -1, 5, 5, 5, 7, 2, -7, 0,
					-- layer=2 filter=249 channel=85
					10, -2, 4, -6, 7, 0, 7, 5, 4,
					-- layer=2 filter=249 channel=86
					-12, -9, -20, -7, -4, 2, -3, 4, 4,
					-- layer=2 filter=249 channel=87
					10, 46, 34, 5, -42, -62, -10, -96, 10,
					-- layer=2 filter=249 channel=88
					3, 6, 0, 1, 5, -19, -10, 0, -25,
					-- layer=2 filter=249 channel=89
					28, 13, 3, 36, 3, 17, 15, -14, -6,
					-- layer=2 filter=249 channel=90
					6, 5, 8, -8, 5, 0, 5, 2, -4,
					-- layer=2 filter=249 channel=91
					17, 4, -15, 11, -7, 9, -4, -12, -16,
					-- layer=2 filter=249 channel=92
					18, 5, 24, 16, 9, 6, 1, -9, -3,
					-- layer=2 filter=249 channel=93
					-11, 0, 8, -3, -40, -48, 36, -55, 27,
					-- layer=2 filter=249 channel=94
					-24, 3, -10, 23, -22, -22, -1, -33, 13,
					-- layer=2 filter=249 channel=95
					-4, 4, 1, -3, 4, -5, 1, 4, 1,
					-- layer=2 filter=249 channel=96
					-30, -17, -30, -51, -91, -89, 2, -80, -72,
					-- layer=2 filter=249 channel=97
					-5, -19, -10, 0, -11, 21, -8, 0, 0,
					-- layer=2 filter=249 channel=98
					4, 10, 22, 14, -6, -13, 0, -8, 45,
					-- layer=2 filter=249 channel=99
					28, 8, 32, 7, 0, 4, 20, 3, 19,
					-- layer=2 filter=249 channel=100
					17, 35, -4, 31, 40, 8, -28, 2, -18,
					-- layer=2 filter=249 channel=101
					-38, -22, -12, -34, 8, 16, 20, 16, 9,
					-- layer=2 filter=249 channel=102
					-4, -32, -6, -12, -78, -38, 10, -82, -26,
					-- layer=2 filter=249 channel=103
					-23, -5, 13, -62, -1, 2, -28, -1, -29,
					-- layer=2 filter=249 channel=104
					-24, 27, -48, -41, -55, 3, 7, -32, 7,
					-- layer=2 filter=249 channel=105
					17, -19, 10, -29, -67, -31, -76, -23, -2,
					-- layer=2 filter=249 channel=106
					1, 0, -9, 0, 2, -6, 4, 12, -5,
					-- layer=2 filter=249 channel=107
					-24, -12, -44, -9, 33, 27, 20, 8, -18,
					-- layer=2 filter=249 channel=108
					23, -11, 7, -18, -9, -9, 7, -7, -30,
					-- layer=2 filter=249 channel=109
					17, 0, -13, -11, -1, 1, 10, 5, 10,
					-- layer=2 filter=249 channel=110
					2, -21, 3, 8, 3, -14, 39, 12, -2,
					-- layer=2 filter=249 channel=111
					7, 0, -4, -1, 5, -5, 2, 0, -9,
					-- layer=2 filter=249 channel=112
					0, -6, -11, -11, 10, -19, -8, 23, 12,
					-- layer=2 filter=249 channel=113
					0, -15, 26, 10, 7, -12, 15, 6, 12,
					-- layer=2 filter=249 channel=114
					2, 0, 3, 8, -10, -3, -10, -18, -9,
					-- layer=2 filter=249 channel=115
					5, 8, 5, 0, 0, -11, 3, -3, 7,
					-- layer=2 filter=249 channel=116
					-2, 52, 15, 24, -7, -92, 0, -77, -9,
					-- layer=2 filter=249 channel=117
					-8, 26, -4, 30, 23, 11, 27, -6, -5,
					-- layer=2 filter=249 channel=118
					-10, -18, -11, -11, 3, 2, 0, 27, 18,
					-- layer=2 filter=249 channel=119
					0, 24, -5, -2, 9, 3, -2, -26, 0,
					-- layer=2 filter=249 channel=120
					-4, -5, -10, -3, 9, 9, 3, -5, -8,
					-- layer=2 filter=249 channel=121
					-10, 8, -5, 7, 7, -3, -1, -10, -8,
					-- layer=2 filter=249 channel=122
					-13, -12, -10, 7, -7, 0, 6, 8, 4,
					-- layer=2 filter=249 channel=123
					15, 12, 28, 19, -29, -17, -31, -45, 5,
					-- layer=2 filter=249 channel=124
					12, 17, -9, -13, -18, -26, -23, -17, 0,
					-- layer=2 filter=249 channel=125
					-8, -9, 3, -7, 3, -8, 0, 2, 2,
					-- layer=2 filter=249 channel=126
					49, 20, 14, -5, -22, 32, 21, 38, -41,
					-- layer=2 filter=249 channel=127
					15, 17, 29, 5, -17, 7, -23, -28, -3,
					-- layer=2 filter=250 channel=0
					-13, 0, -15, -24, -34, -14, -6, 3, -6,
					-- layer=2 filter=250 channel=1
					2, 10, -11, 9, 2, -5, -10, -11, -22,
					-- layer=2 filter=250 channel=2
					-4, 1, -6, 0, -3, 0, -8, 3, 5,
					-- layer=2 filter=250 channel=3
					-19, -9, 0, 2, 6, 3, 0, -6, -1,
					-- layer=2 filter=250 channel=4
					-7, -17, -7, -5, -26, -4, -22, 19, -8,
					-- layer=2 filter=250 channel=5
					0, 3, 1, -12, -7, -4, -2, -13, 2,
					-- layer=2 filter=250 channel=6
					-9, 10, 6, 10, 4, -29, 3, 7, -19,
					-- layer=2 filter=250 channel=7
					-3, -5, -13, -15, -6, 5, 0, 0, -19,
					-- layer=2 filter=250 channel=8
					-10, 0, -4, -1, 0, 2, 8, 1, 1,
					-- layer=2 filter=250 channel=9
					-13, -8, -12, -9, -16, -14, -6, -3, 3,
					-- layer=2 filter=250 channel=10
					-31, -12, -6, -2, -8, 0, -4, -9, 2,
					-- layer=2 filter=250 channel=11
					-10, -23, -3, -14, -17, -16, 5, -22, -29,
					-- layer=2 filter=250 channel=12
					10, -8, 5, 6, -11, -1, -23, -21, -14,
					-- layer=2 filter=250 channel=13
					10, 0, -8, 4, 1, 4, 2, -6, 0,
					-- layer=2 filter=250 channel=14
					-2, -11, -18, 6, -6, -3, -13, -9, -15,
					-- layer=2 filter=250 channel=15
					-10, -12, 27, 3, 1, -7, -3, -7, 0,
					-- layer=2 filter=250 channel=16
					-12, -10, 2, -16, -8, -9, 2, 13, 6,
					-- layer=2 filter=250 channel=17
					-1, -4, -7, -6, 2, 6, -1, 6, 6,
					-- layer=2 filter=250 channel=18
					5, -24, 4, -7, -1, 3, -13, 10, -10,
					-- layer=2 filter=250 channel=19
					-8, -15, -14, -18, 0, -15, 0, -2, 0,
					-- layer=2 filter=250 channel=20
					-11, -4, -6, -5, 4, -5, 0, 1, 5,
					-- layer=2 filter=250 channel=21
					-4, 0, 8, -1, 0, -9, 7, 8, 11,
					-- layer=2 filter=250 channel=22
					7, 9, -4, 2, 1, -2, 9, -5, -1,
					-- layer=2 filter=250 channel=23
					-26, -9, -12, -20, -14, -15, -1, -14, -8,
					-- layer=2 filter=250 channel=24
					-33, 3, -7, -24, -16, -1, -27, -23, -7,
					-- layer=2 filter=250 channel=25
					-2, -9, -3, -7, -21, -1, -22, -18, -3,
					-- layer=2 filter=250 channel=26
					-4, 1, 4, -2, 4, -5, -4, 9, 5,
					-- layer=2 filter=250 channel=27
					-7, -15, -4, 3, 2, 0, 4, -6, -3,
					-- layer=2 filter=250 channel=28
					-7, -23, -18, -22, -7, -12, -13, -7, 4,
					-- layer=2 filter=250 channel=29
					-8, -4, 4, 0, -8, 6, -5, -8, -6,
					-- layer=2 filter=250 channel=30
					-5, -11, -15, 4, -13, -16, -3, -18, 1,
					-- layer=2 filter=250 channel=31
					-9, -16, -3, -10, 3, -3, -10, -2, 4,
					-- layer=2 filter=250 channel=32
					0, -8, -2, 2, 0, 1, -9, 4, 2,
					-- layer=2 filter=250 channel=33
					-17, -8, -36, -11, -8, 0, 1, -11, -29,
					-- layer=2 filter=250 channel=34
					6, 6, -15, 17, -10, 1, -1, 16, 1,
					-- layer=2 filter=250 channel=35
					0, 2, -7, -14, -4, 5, -17, 14, 11,
					-- layer=2 filter=250 channel=36
					6, -10, 0, 0, 1, 6, -9, -9, -8,
					-- layer=2 filter=250 channel=37
					-16, -27, -19, -8, -2, -11, -1, -22, -17,
					-- layer=2 filter=250 channel=38
					-20, -11, 1, 16, -16, 9, -7, -29, 5,
					-- layer=2 filter=250 channel=39
					0, 13, -2, -17, 6, 6, -11, -11, -13,
					-- layer=2 filter=250 channel=40
					-3, 5, 0, -3, 9, -10, -18, -4, -13,
					-- layer=2 filter=250 channel=41
					-4, -3, -3, 10, -10, 4, -6, 10, -6,
					-- layer=2 filter=250 channel=42
					-18, -12, -13, 8, -1, -17, 1, 0, -6,
					-- layer=2 filter=250 channel=43
					10, -9, -1, 8, 6, -15, 0, 8, 0,
					-- layer=2 filter=250 channel=44
					5, 2, -7, -8, 3, -5, 10, 1, -2,
					-- layer=2 filter=250 channel=45
					-13, -26, -6, -2, -1, 2, 2, 2, 2,
					-- layer=2 filter=250 channel=46
					4, -21, -8, -7, -19, -16, -11, -13, 12,
					-- layer=2 filter=250 channel=47
					-21, -14, -7, -16, -16, 10, 0, 9, 1,
					-- layer=2 filter=250 channel=48
					-2, 3, -6, 3, -5, 6, -6, -8, -3,
					-- layer=2 filter=250 channel=49
					8, -9, -7, 6, -12, -10, -9, 0, -14,
					-- layer=2 filter=250 channel=50
					3, -4, 10, 14, 3, 2, -1, 0, 3,
					-- layer=2 filter=250 channel=51
					-25, -31, -26, -12, -18, -19, -13, -30, -15,
					-- layer=2 filter=250 channel=52
					-4, 1, 3, 8, 3, 1, -17, 13, -23,
					-- layer=2 filter=250 channel=53
					-13, -6, -12, -11, -4, -24, -10, -7, -5,
					-- layer=2 filter=250 channel=54
					11, 11, -13, -11, -5, -3, -3, -3, -5,
					-- layer=2 filter=250 channel=55
					10, 4, 1, -6, -8, -4, 3, -9, -5,
					-- layer=2 filter=250 channel=56
					-16, -8, 9, -25, -12, -20, -1, 1, -4,
					-- layer=2 filter=250 channel=57
					3, 0, -6, 0, -9, 8, -5, -2, 8,
					-- layer=2 filter=250 channel=58
					1, 1, 7, 3, -5, -16, -6, -21, -3,
					-- layer=2 filter=250 channel=59
					-4, 10, -4, 7, -8, -16, -7, -4, -20,
					-- layer=2 filter=250 channel=60
					-5, 5, -3, -13, -15, -14, -13, -28, 1,
					-- layer=2 filter=250 channel=61
					-12, -5, -8, -19, 6, 5, 6, -17, -19,
					-- layer=2 filter=250 channel=62
					12, 6, -2, 6, -8, -15, -7, 1, -2,
					-- layer=2 filter=250 channel=63
					-3, -7, -18, -12, -7, -2, -16, -17, 2,
					-- layer=2 filter=250 channel=64
					-3, -6, -1, -17, -9, -8, -7, 0, -16,
					-- layer=2 filter=250 channel=65
					4, 6, -13, 14, 9, 4, -5, -1, -29,
					-- layer=2 filter=250 channel=66
					6, 0, 16, 18, -11, 15, -9, 12, 14,
					-- layer=2 filter=250 channel=67
					-7, 3, -17, -2, -20, -19, -5, -4, -15,
					-- layer=2 filter=250 channel=68
					-10, -5, -7, 0, 4, 4, -5, -10, -8,
					-- layer=2 filter=250 channel=69
					0, -4, 2, 0, 8, -4, -17, 6, -12,
					-- layer=2 filter=250 channel=70
					-1, -4, 8, -18, -20, 4, 3, 15, 20,
					-- layer=2 filter=250 channel=71
					-10, -7, -12, -19, -18, 5, -2, -8, -16,
					-- layer=2 filter=250 channel=72
					-9, -3, -10, -1, -11, 5, -4, -9, -19,
					-- layer=2 filter=250 channel=73
					-13, -3, 17, 13, -10, 7, 10, -10, -1,
					-- layer=2 filter=250 channel=74
					-9, 11, -18, 0, -8, -1, -14, -9, -9,
					-- layer=2 filter=250 channel=75
					-11, 2, -3, -11, -17, -10, -7, 5, -6,
					-- layer=2 filter=250 channel=76
					4, -19, -5, 7, 9, -3, -10, 1, -23,
					-- layer=2 filter=250 channel=77
					5, -4, 8, -8, 1, -1, -8, 7, -9,
					-- layer=2 filter=250 channel=78
					-5, -2, 0, -9, -11, -12, -8, -16, -6,
					-- layer=2 filter=250 channel=79
					7, 8, -2, -11, 4, -3, -10, 0, 0,
					-- layer=2 filter=250 channel=80
					-25, -19, -7, -11, -3, -19, -18, 3, -4,
					-- layer=2 filter=250 channel=81
					-3, -6, -9, -12, 6, 2, 6, -10, 7,
					-- layer=2 filter=250 channel=82
					0, 4, 10, 5, -1, 1, 9, -8, 2,
					-- layer=2 filter=250 channel=83
					-12, 0, -10, -11, -23, -15, -2, -23, -2,
					-- layer=2 filter=250 channel=84
					4, -8, -7, -2, -7, -2, 0, -8, 8,
					-- layer=2 filter=250 channel=85
					0, -10, 9, -4, -2, -3, 5, -9, -6,
					-- layer=2 filter=250 channel=86
					5, 1, 3, -2, -11, 10, 4, -10, -7,
					-- layer=2 filter=250 channel=87
					-10, -24, -11, -8, -25, -22, -16, 1, -12,
					-- layer=2 filter=250 channel=88
					-2, -10, -21, -4, 10, -2, -28, -11, -13,
					-- layer=2 filter=250 channel=89
					0, -24, 6, 9, -10, -9, -9, -15, -19,
					-- layer=2 filter=250 channel=90
					0, 8, 1, -9, -3, 6, -7, -5, -7,
					-- layer=2 filter=250 channel=91
					-10, -1, -11, 1, -11, -4, -14, 2, -6,
					-- layer=2 filter=250 channel=92
					8, 0, -12, 10, -5, 4, -23, -4, -12,
					-- layer=2 filter=250 channel=93
					19, 5, 4, 12, 16, 0, 2, -7, -12,
					-- layer=2 filter=250 channel=94
					-6, -10, -15, -6, -11, -20, -6, -21, -16,
					-- layer=2 filter=250 channel=95
					-6, -7, -11, 0, 3, 0, -5, -9, -2,
					-- layer=2 filter=250 channel=96
					6, -20, 8, -1, -28, 0, -14, 5, -5,
					-- layer=2 filter=250 channel=97
					-2, -32, -18, -6, -16, -9, -5, -10, 5,
					-- layer=2 filter=250 channel=98
					-21, -28, 0, -4, -13, 16, 6, 11, -5,
					-- layer=2 filter=250 channel=99
					-2, -13, 8, -20, 1, -13, -7, -9, -10,
					-- layer=2 filter=250 channel=100
					-12, 10, -26, -16, -1, -3, 4, -13, 11,
					-- layer=2 filter=250 channel=101
					-4, -1, 2, -11, -26, -23, -24, -14, -17,
					-- layer=2 filter=250 channel=102
					-5, -6, -4, -16, -9, 7, -21, 3, 1,
					-- layer=2 filter=250 channel=103
					0, -1, -3, 7, 7, -11, -3, -1, 14,
					-- layer=2 filter=250 channel=104
					-6, -12, -14, 4, -15, -9, -23, 2, -21,
					-- layer=2 filter=250 channel=105
					-5, -22, 0, -2, 7, 11, -4, -6, -8,
					-- layer=2 filter=250 channel=106
					-13, 0, -8, -11, 0, 3, -6, -27, -7,
					-- layer=2 filter=250 channel=107
					7, -11, -12, 10, -12, -8, 10, 1, -4,
					-- layer=2 filter=250 channel=108
					-9, -26, -10, -3, -21, 1, 3, -2, -25,
					-- layer=2 filter=250 channel=109
					-8, -11, -10, -1, 8, -1, 8, -2, -6,
					-- layer=2 filter=250 channel=110
					-8, 1, 0, -12, 3, 2, -27, 1, 3,
					-- layer=2 filter=250 channel=111
					0, 4, -1, -1, 1, -5, -4, -9, -9,
					-- layer=2 filter=250 channel=112
					-24, -11, -15, -1, -14, 11, -6, -14, -13,
					-- layer=2 filter=250 channel=113
					3, -15, 2, -15, -13, -5, -23, -22, 3,
					-- layer=2 filter=250 channel=114
					-3, 4, -4, 7, 10, 0, 10, 4, 3,
					-- layer=2 filter=250 channel=115
					5, 3, -9, 0, 0, -10, -6, 6, 7,
					-- layer=2 filter=250 channel=116
					-24, -7, 1, -19, -3, 5, -22, 12, -14,
					-- layer=2 filter=250 channel=117
					1, 1, -16, -6, -15, 1, -4, -4, 3,
					-- layer=2 filter=250 channel=118
					-9, 4, 8, 1, -2, -5, -1, 0, -21,
					-- layer=2 filter=250 channel=119
					3, -10, -14, -14, -20, 1, -11, 2, 8,
					-- layer=2 filter=250 channel=120
					9, 0, 9, 0, 9, 6, -3, -6, -2,
					-- layer=2 filter=250 channel=121
					-7, -4, 0, -5, -2, 1, 8, 0, -4,
					-- layer=2 filter=250 channel=122
					-1, 3, 5, -2, -10, 1, -6, -7, 2,
					-- layer=2 filter=250 channel=123
					7, -7, -2, 3, 15, 24, 0, 0, -14,
					-- layer=2 filter=250 channel=124
					11, -3, 1, 13, 19, -16, -13, 4, -15,
					-- layer=2 filter=250 channel=125
					7, 2, -4, 2, 0, -6, 7, -8, 7,
					-- layer=2 filter=250 channel=126
					-2, -6, 8, -12, 0, 0, -21, -16, -17,
					-- layer=2 filter=250 channel=127
					7, -15, 0, -1, 11, -15, -23, -11, -6,
					-- layer=2 filter=251 channel=0
					5, -9, -6, -8, -1, -2, 0, 7, -7,
					-- layer=2 filter=251 channel=1
					-8, 3, -10, 0, 5, -12, 5, -1, 0,
					-- layer=2 filter=251 channel=2
					-4, -3, 6, 9, 5, 2, -10, -4, -8,
					-- layer=2 filter=251 channel=3
					-2, -10, -4, -2, 3, -11, 0, -10, -11,
					-- layer=2 filter=251 channel=4
					3, 6, -11, 2, -7, 3, -3, -7, -8,
					-- layer=2 filter=251 channel=5
					-12, -5, 4, -9, 3, -3, -7, 0, -7,
					-- layer=2 filter=251 channel=6
					1, -5, -4, -2, 5, -5, -3, -11, 8,
					-- layer=2 filter=251 channel=7
					-1, -5, 2, -9, 0, -16, 4, -6, -8,
					-- layer=2 filter=251 channel=8
					2, 6, -2, 6, -7, 9, 0, 2, 4,
					-- layer=2 filter=251 channel=9
					-8, -2, 1, -3, 0, 0, 4, -12, 5,
					-- layer=2 filter=251 channel=10
					-13, 7, -8, -17, -3, 2, -9, 4, -1,
					-- layer=2 filter=251 channel=11
					1, 7, -4, -6, -4, -7, 5, 0, -14,
					-- layer=2 filter=251 channel=12
					-7, -1, -9, 3, 0, 4, 0, 0, -5,
					-- layer=2 filter=251 channel=13
					1, 7, 0, -3, -8, 2, -12, 6, -3,
					-- layer=2 filter=251 channel=14
					-3, 0, -3, 0, 5, -7, -7, 0, -6,
					-- layer=2 filter=251 channel=15
					-11, 1, -2, -1, 4, 8, -1, 5, -1,
					-- layer=2 filter=251 channel=16
					6, 7, -8, 4, -6, -12, -2, 7, -10,
					-- layer=2 filter=251 channel=17
					-11, 9, -1, 10, 6, 7, -6, -9, -11,
					-- layer=2 filter=251 channel=18
					0, -11, 1, -9, 5, 1, 3, 5, -8,
					-- layer=2 filter=251 channel=19
					-8, 3, -4, 2, -11, 0, -2, 2, -7,
					-- layer=2 filter=251 channel=20
					0, -4, -7, -6, -9, -10, -6, 1, -3,
					-- layer=2 filter=251 channel=21
					5, -6, -6, -1, -3, 6, 6, -4, -11,
					-- layer=2 filter=251 channel=22
					-1, -2, 0, -5, 3, -3, -1, 9, 3,
					-- layer=2 filter=251 channel=23
					-8, 8, 3, -8, -10, 5, 0, 10, -13,
					-- layer=2 filter=251 channel=24
					2, -10, -8, -8, -4, -2, 2, 6, 3,
					-- layer=2 filter=251 channel=25
					0, 1, -4, 3, 1, -12, 1, 2, 5,
					-- layer=2 filter=251 channel=26
					-5, 5, -5, -6, -7, -7, 6, -7, 9,
					-- layer=2 filter=251 channel=27
					0, 0, -9, 0, -9, -8, -7, 2, 4,
					-- layer=2 filter=251 channel=28
					-15, 1, -18, -5, 4, -9, -2, 5, 0,
					-- layer=2 filter=251 channel=29
					7, -9, -7, 0, -2, 1, -6, 4, -3,
					-- layer=2 filter=251 channel=30
					-11, -1, -5, 7, -4, 0, -3, -11, -12,
					-- layer=2 filter=251 channel=31
					-1, -4, -6, 0, 0, 4, 7, -6, 8,
					-- layer=2 filter=251 channel=32
					-5, 5, 1, -4, 3, -4, -1, 5, -11,
					-- layer=2 filter=251 channel=33
					-10, -1, 5, -6, 5, 7, -1, -5, 5,
					-- layer=2 filter=251 channel=34
					-8, 0, 5, -8, -2, -4, -5, 5, -7,
					-- layer=2 filter=251 channel=35
					-7, -8, -14, -12, -8, -10, -2, 3, 0,
					-- layer=2 filter=251 channel=36
					6, -8, 0, 5, 8, -8, -4, -8, 2,
					-- layer=2 filter=251 channel=37
					-1, 3, -13, 6, -8, 3, -13, -13, -5,
					-- layer=2 filter=251 channel=38
					8, 6, 1, 0, -2, -8, -4, 4, -10,
					-- layer=2 filter=251 channel=39
					8, 8, 2, -5, 6, -4, 6, 3, -7,
					-- layer=2 filter=251 channel=40
					5, 1, -7, 5, -1, 6, 5, 8, 0,
					-- layer=2 filter=251 channel=41
					7, 3, -2, -8, -9, -2, 4, -6, -10,
					-- layer=2 filter=251 channel=42
					-10, -5, 1, -10, -11, 8, -9, -7, -14,
					-- layer=2 filter=251 channel=43
					4, 4, -7, 5, 6, -6, 7, 7, -1,
					-- layer=2 filter=251 channel=44
					7, 1, 2, 0, 0, 8, -9, 0, -6,
					-- layer=2 filter=251 channel=45
					1, 5, -3, 0, -5, -7, 0, -1, 4,
					-- layer=2 filter=251 channel=46
					-7, 0, 2, 5, 0, -10, -2, -2, 5,
					-- layer=2 filter=251 channel=47
					0, 1, -13, -8, -6, 5, -1, -6, -7,
					-- layer=2 filter=251 channel=48
					-6, -5, -7, 5, -8, 0, 0, -10, 1,
					-- layer=2 filter=251 channel=49
					-20, -12, -13, 0, 0, -6, 0, -8, 2,
					-- layer=2 filter=251 channel=50
					-5, 3, 0, 8, -8, -5, 0, 0, -3,
					-- layer=2 filter=251 channel=51
					1, 0, -6, 1, -2, 0, 7, -1, -6,
					-- layer=2 filter=251 channel=52
					6, -4, 0, 1, -12, -8, 4, 2, -13,
					-- layer=2 filter=251 channel=53
					4, 0, -6, -2, -11, 0, -2, 4, 3,
					-- layer=2 filter=251 channel=54
					-6, -4, -5, -2, -12, 4, 3, -12, -4,
					-- layer=2 filter=251 channel=55
					3, 4, 0, -7, 7, -5, 7, 3, -2,
					-- layer=2 filter=251 channel=56
					0, 6, -12, 4, -4, -5, -1, -7, -2,
					-- layer=2 filter=251 channel=57
					-9, -4, -7, -1, -3, -6, -9, -9, -9,
					-- layer=2 filter=251 channel=58
					5, 0, -2, -9, -9, -9, -3, -2, -7,
					-- layer=2 filter=251 channel=59
					-5, 1, 3, 3, -7, 7, 0, -1, 7,
					-- layer=2 filter=251 channel=60
					5, -3, -11, -5, -6, -9, -9, -14, -11,
					-- layer=2 filter=251 channel=61
					4, 0, -3, -7, 4, -12, -4, -1, 0,
					-- layer=2 filter=251 channel=62
					-8, -4, -3, 4, -5, -10, 5, 1, -4,
					-- layer=2 filter=251 channel=63
					2, -6, -7, -1, 2, -12, -13, -6, -6,
					-- layer=2 filter=251 channel=64
					-4, -3, -11, -6, 0, -11, 1, 5, -8,
					-- layer=2 filter=251 channel=65
					4, -1, -6, -6, -6, 4, 8, -11, -12,
					-- layer=2 filter=251 channel=66
					-7, 6, 8, 2, 6, -4, -8, 6, 0,
					-- layer=2 filter=251 channel=67
					-1, -3, -4, -6, -4, -7, 1, 0, 6,
					-- layer=2 filter=251 channel=68
					5, 7, -10, 3, 2, -8, -1, -8, -1,
					-- layer=2 filter=251 channel=69
					-7, -6, -9, -9, 2, -4, 2, 4, 0,
					-- layer=2 filter=251 channel=70
					-1, -10, 0, -7, -2, 5, -6, 4, 2,
					-- layer=2 filter=251 channel=71
					-6, 6, 0, -10, -6, -10, -13, 6, 3,
					-- layer=2 filter=251 channel=72
					-7, 11, 0, -2, -2, -4, -2, -3, 7,
					-- layer=2 filter=251 channel=73
					5, -1, -9, 0, -6, -3, -3, -7, -6,
					-- layer=2 filter=251 channel=74
					-3, -8, 5, 0, -6, -12, 1, 6, 3,
					-- layer=2 filter=251 channel=75
					-6, -8, 4, -1, -11, -7, 4, 11, 8,
					-- layer=2 filter=251 channel=76
					-6, -11, -3, 5, -6, 1, -9, -9, 6,
					-- layer=2 filter=251 channel=77
					-1, -6, 7, -11, -11, -7, -9, 2, 5,
					-- layer=2 filter=251 channel=78
					0, -8, 0, 5, -4, 1, -8, 3, 5,
					-- layer=2 filter=251 channel=79
					4, -7, -4, -11, -9, -4, -4, -11, 5,
					-- layer=2 filter=251 channel=80
					-11, -5, -7, 1, -1, -1, -4, 4, -11,
					-- layer=2 filter=251 channel=81
					2, 7, 0, 8, -1, 4, -6, -8, -9,
					-- layer=2 filter=251 channel=82
					-5, -5, 9, 3, -3, -9, -7, -9, 9,
					-- layer=2 filter=251 channel=83
					0, -6, -11, -3, 5, -8, -8, 3, 7,
					-- layer=2 filter=251 channel=84
					8, 7, 8, -2, -5, 0, -2, 3, 6,
					-- layer=2 filter=251 channel=85
					6, 3, 7, -10, -7, 8, -7, 2, 2,
					-- layer=2 filter=251 channel=86
					0, -5, -4, -4, 1, 3, 11, -5, -2,
					-- layer=2 filter=251 channel=87
					6, 4, 2, -3, 6, 7, -6, -5, 7,
					-- layer=2 filter=251 channel=88
					-4, -1, -5, 3, -8, 7, -9, 3, -6,
					-- layer=2 filter=251 channel=89
					-7, -6, 3, -9, 7, -7, 5, 4, 2,
					-- layer=2 filter=251 channel=90
					4, 4, -6, -8, 6, -6, -1, -4, 10,
					-- layer=2 filter=251 channel=91
					-10, 2, 2, -8, -12, -9, 4, 0, 1,
					-- layer=2 filter=251 channel=92
					-4, -3, 1, -6, 6, -6, 9, 2, -1,
					-- layer=2 filter=251 channel=93
					0, 2, -5, 8, 0, -11, -6, -8, 2,
					-- layer=2 filter=251 channel=94
					-15, 0, 1, 4, -3, 10, -8, -6, -8,
					-- layer=2 filter=251 channel=95
					4, 2, -2, -9, 9, -8, -11, -3, 7,
					-- layer=2 filter=251 channel=96
					-3, 8, -5, -9, -10, -3, -5, -5, -3,
					-- layer=2 filter=251 channel=97
					0, -5, -1, -2, 1, 0, 1, 0, -10,
					-- layer=2 filter=251 channel=98
					-12, 7, -10, 2, -5, -4, 4, -10, 2,
					-- layer=2 filter=251 channel=99
					6, -2, -3, -9, 0, -3, -11, -1, -10,
					-- layer=2 filter=251 channel=100
					-2, -12, 3, -2, 5, 6, 2, 5, 0,
					-- layer=2 filter=251 channel=101
					5, 0, 0, 3, 4, -1, 6, 6, -5,
					-- layer=2 filter=251 channel=102
					6, -7, 0, -11, -6, -4, 1, -4, -2,
					-- layer=2 filter=251 channel=103
					-8, 4, 8, 4, 2, -4, -11, -7, 9,
					-- layer=2 filter=251 channel=104
					-4, 6, 4, -3, 0, -2, -8, 4, -2,
					-- layer=2 filter=251 channel=105
					-8, -7, 8, 3, -8, -4, -5, -9, -3,
					-- layer=2 filter=251 channel=106
					2, -11, -7, -8, 9, -8, -11, 0, -12,
					-- layer=2 filter=251 channel=107
					2, 5, 2, 11, -4, 6, -4, 1, 8,
					-- layer=2 filter=251 channel=108
					-6, -1, -3, -8, -3, -7, 0, 3, 3,
					-- layer=2 filter=251 channel=109
					5, -4, -1, -6, -7, -10, -1, -3, -5,
					-- layer=2 filter=251 channel=110
					-3, -10, -8, -4, -6, 3, 7, 3, 3,
					-- layer=2 filter=251 channel=111
					-3, -2, 3, -3, 4, -5, 9, 11, -10,
					-- layer=2 filter=251 channel=112
					-8, 7, -5, 4, 4, -11, -1, 2, -6,
					-- layer=2 filter=251 channel=113
					-9, 4, -1, 0, -8, -3, 7, -1, -3,
					-- layer=2 filter=251 channel=114
					-5, 9, 0, -9, 1, -7, -9, -4, -10,
					-- layer=2 filter=251 channel=115
					-9, -9, 1, 1, 0, 0, 0, -8, 4,
					-- layer=2 filter=251 channel=116
					-5, -12, -7, -9, 2, -1, 3, -2, -3,
					-- layer=2 filter=251 channel=117
					6, 4, -11, 3, -6, -10, -8, -6, -12,
					-- layer=2 filter=251 channel=118
					7, -4, 1, -9, 4, -7, 2, -5, -11,
					-- layer=2 filter=251 channel=119
					-6, -9, -6, -6, -8, -9, -10, -10, -1,
					-- layer=2 filter=251 channel=120
					-9, 8, -6, -8, -9, 7, -2, 5, 1,
					-- layer=2 filter=251 channel=121
					-1, 1, 1, -8, -8, 4, 4, -4, -9,
					-- layer=2 filter=251 channel=122
					-4, -5, -7, 0, -1, 4, 1, -9, 9,
					-- layer=2 filter=251 channel=123
					4, -2, -8, 2, -7, -11, -3, 4, -10,
					-- layer=2 filter=251 channel=124
					1, -6, -8, -1, 5, -6, -3, -7, -2,
					-- layer=2 filter=251 channel=125
					-9, 6, -7, 8, -11, -6, -7, -8, -8,
					-- layer=2 filter=251 channel=126
					7, -8, -7, -10, -5, -5, 3, -7, -2,
					-- layer=2 filter=251 channel=127
					-4, 0, 2, 4, 6, -4, 2, -1, -4,
					-- layer=2 filter=252 channel=0
					0, 18, 11, 32, 9, 16, 22, 8, 13,
					-- layer=2 filter=252 channel=1
					-27, -24, -26, -17, -58, -4, 16, -14, -45,
					-- layer=2 filter=252 channel=2
					1, -9, 0, -3, 0, -7, 0, 8, -3,
					-- layer=2 filter=252 channel=3
					-15, 17, 1, -5, 40, -22, -16, 14, 14,
					-- layer=2 filter=252 channel=4
					10, -34, -44, -24, -20, 17, 9, 4, -36,
					-- layer=2 filter=252 channel=5
					2, -27, -3, 0, 8, 15, 10, 0, 22,
					-- layer=2 filter=252 channel=6
					48, 53, 1, 3, 19, 0, 3, 6, 35,
					-- layer=2 filter=252 channel=7
					-29, -20, 17, 33, -22, -13, 14, -9, 33,
					-- layer=2 filter=252 channel=8
					-9, 6, 1, -1, 1, 3, -3, -5, 4,
					-- layer=2 filter=252 channel=9
					-27, -28, -56, -29, -34, -50, -30, -32, -39,
					-- layer=2 filter=252 channel=10
					13, 1, 14, 0, -3, 2, 17, 35, 25,
					-- layer=2 filter=252 channel=11
					11, 6, 0, 0, 21, 18, -4, 5, 13,
					-- layer=2 filter=252 channel=12
					0, 19, -53, 6, 3, 8, 8, -27, -7,
					-- layer=2 filter=252 channel=13
					-2, 4, 8, 9, 2, 8, 1, -7, -5,
					-- layer=2 filter=252 channel=14
					4, -1, -20, 1, 0, 33, 22, -8, -25,
					-- layer=2 filter=252 channel=15
					-16, -27, -23, 4, -2, -20, 17, 0, 20,
					-- layer=2 filter=252 channel=16
					-13, -14, -3, 11, 31, -11, 2, 3, -34,
					-- layer=2 filter=252 channel=17
					4, 6, 0, -6, 1, -10, -4, -8, 6,
					-- layer=2 filter=252 channel=18
					-29, -2, -10, -15, -18, 0, -2, 9, -9,
					-- layer=2 filter=252 channel=19
					-30, -34, 0, -20, -51, -43, 39, -25, -50,
					-- layer=2 filter=252 channel=20
					0, 4, -8, 7, 4, -5, 0, 9, -7,
					-- layer=2 filter=252 channel=21
					6, -13, 2, 0, -10, 0, -20, 1, -6,
					-- layer=2 filter=252 channel=22
					-7, 6, 2, 9, 2, -9, -7, -5, -1,
					-- layer=2 filter=252 channel=23
					-17, 8, 25, -3, 19, -1, -44, 14, -16,
					-- layer=2 filter=252 channel=24
					-26, 4, -36, 33, 39, 11, -2, 10, -3,
					-- layer=2 filter=252 channel=25
					16, 23, -5, 29, 55, 13, 4, 7, 34,
					-- layer=2 filter=252 channel=26
					-6, 0, 1, 6, -8, 10, 9, 3, -9,
					-- layer=2 filter=252 channel=27
					-9, -26, 2, 7, -35, -8, 25, -9, -15,
					-- layer=2 filter=252 channel=28
					-1, 4, -10, -13, -30, -32, 16, 9, 5,
					-- layer=2 filter=252 channel=29
					4, -4, 0, 7, 0, -7, -7, 2, 7,
					-- layer=2 filter=252 channel=30
					-13, -76, -5, -40, -68, -39, 10, -39, -5,
					-- layer=2 filter=252 channel=31
					-10, -24, -56, 17, 45, -5, -70, -20, -74,
					-- layer=2 filter=252 channel=32
					-4, -8, -8, -6, 3, 0, 5, 0, 2,
					-- layer=2 filter=252 channel=33
					-20, 36, 28, 41, -4, -13, 26, -11, 21,
					-- layer=2 filter=252 channel=34
					11, 6, 23, 5, 0, -3, -12, -30, -33,
					-- layer=2 filter=252 channel=35
					33, 51, 11, -23, -7, -52, 5, -19, 16,
					-- layer=2 filter=252 channel=36
					-3, -1, 1, -1, -6, -10, -8, 2, -13,
					-- layer=2 filter=252 channel=37
					5, -17, -8, 5, -10, 16, 17, 0, 7,
					-- layer=2 filter=252 channel=38
					-16, -45, -28, -5, -65, -38, 38, -26, -2,
					-- layer=2 filter=252 channel=39
					0, -6, -18, -1, -18, -39, 29, 0, 22,
					-- layer=2 filter=252 channel=40
					23, 11, -64, -16, 14, -30, -3, 43, 46,
					-- layer=2 filter=252 channel=41
					-5, 3, -3, -2, 8, -4, -1, 8, -3,
					-- layer=2 filter=252 channel=42
					30, 34, 8, 31, 44, -7, 0, 1, 3,
					-- layer=2 filter=252 channel=43
					-50, -14, 9, -1, -22, -6, 0, 22, -17,
					-- layer=2 filter=252 channel=44
					0, 0, -4, 8, 0, 0, 0, 5, 0,
					-- layer=2 filter=252 channel=45
					-56, 3, -1, -26, -25, -26, -4, -57, -58,
					-- layer=2 filter=252 channel=46
					-24, -1, -23, -20, 5, -39, 17, -8, -8,
					-- layer=2 filter=252 channel=47
					-2, 9, 18, -20, -49, -67, 29, 8, -5,
					-- layer=2 filter=252 channel=48
					4, 0, -6, -2, -10, -5, 0, 7, 0,
					-- layer=2 filter=252 channel=49
					-41, -11, 21, -37, 15, -9, -4, 20, -3,
					-- layer=2 filter=252 channel=50
					-13, 12, 13, -2, -11, -13, 0, -15, 4,
					-- layer=2 filter=252 channel=51
					8, -5, 12, 24, 20, 13, 4, 15, 17,
					-- layer=2 filter=252 channel=52
					-21, 7, 51, 35, -34, -28, 24, 20, -7,
					-- layer=2 filter=252 channel=53
					-23, -10, 1, -9, -114, -27, -1, 7, 17,
					-- layer=2 filter=252 channel=54
					29, 44, 31, 32, 29, 29, 23, 22, 21,
					-- layer=2 filter=252 channel=55
					5, -8, -2, 4, -7, -7, 2, 0, -4,
					-- layer=2 filter=252 channel=56
					26, -6, -3, 6, -9, 9, 7, 0, 14,
					-- layer=2 filter=252 channel=57
					0, -6, -5, 6, -3, -6, -1, -5, -4,
					-- layer=2 filter=252 channel=58
					9, 29, -9, 19, 3, 18, 16, -8, -22,
					-- layer=2 filter=252 channel=59
					-43, -9, 3, -1, -79, -25, -2, 8, -21,
					-- layer=2 filter=252 channel=60
					23, -28, 51, -7, 4, -1, 12, -7, 0,
					-- layer=2 filter=252 channel=61
					10, 9, 44, 1, -32, -6, 2, 12, 16,
					-- layer=2 filter=252 channel=62
					26, 34, 13, 20, 49, 15, 20, -7, 0,
					-- layer=2 filter=252 channel=63
					-17, -42, -51, -30, -38, -8, -8, -3, -15,
					-- layer=2 filter=252 channel=64
					8, 19, 22, 44, 36, 6, -12, 16, -5,
					-- layer=2 filter=252 channel=65
					29, 8, 21, -18, -21, -10, -2, 35, 0,
					-- layer=2 filter=252 channel=66
					46, 15, 5, 5, -44, 25, 18, -30, -9,
					-- layer=2 filter=252 channel=67
					-37, -81, -66, -27, -31, -64, -25, -45, -28,
					-- layer=2 filter=252 channel=68
					-6, -8, -2, -8, 3, 8, 3, 0, 6,
					-- layer=2 filter=252 channel=69
					-8, 23, 24, 35, 17, 11, 10, 5, -24,
					-- layer=2 filter=252 channel=70
					28, 28, -1, -43, -23, -24, 4, -28, 1,
					-- layer=2 filter=252 channel=71
					-16, -22, 16, -1, -38, 15, 7, -17, -19,
					-- layer=2 filter=252 channel=72
					40, -3, -9, 34, 25, -13, 53, 12, 36,
					-- layer=2 filter=252 channel=73
					-38, -34, 18, -21, -96, -18, -48, -24, -21,
					-- layer=2 filter=252 channel=74
					-20, 0, -33, 0, -62, -15, 30, 11, -2,
					-- layer=2 filter=252 channel=75
					30, 46, -57, 26, -6, 10, 10, 12, -13,
					-- layer=2 filter=252 channel=76
					50, -21, -28, 1, -43, -26, 33, -19, -77,
					-- layer=2 filter=252 channel=77
					-6, -5, -9, -3, 7, 11, 0, -6, -3,
					-- layer=2 filter=252 channel=78
					-4, 17, -8, 13, 23, 6, -33, 19, 0,
					-- layer=2 filter=252 channel=79
					9, 2, -5, 0, 8, 0, 9, -4, -1,
					-- layer=2 filter=252 channel=80
					-52, -21, -26, -8, 23, -24, -4, -2, -24,
					-- layer=2 filter=252 channel=81
					-11, -3, 3, -9, -13, -3, -4, -9, 0,
					-- layer=2 filter=252 channel=82
					4, 8, 1, -7, 9, -5, -10, -9, -7,
					-- layer=2 filter=252 channel=83
					-3, -19, -19, -29, 2, 0, -33, -3, -41,
					-- layer=2 filter=252 channel=84
					2, 2, -3, -8, 1, -8, -5, -4, 2,
					-- layer=2 filter=252 channel=85
					-8, 13, 12, 7, 9, 17, 0, 13, 11,
					-- layer=2 filter=252 channel=86
					6, 0, 10, -8, 7, -9, -1, 2, 17,
					-- layer=2 filter=252 channel=87
					0, 0, 12, -12, -13, -3, -22, -32, 0,
					-- layer=2 filter=252 channel=88
					4, -20, -18, -50, -48, 4, -3, -18, -12,
					-- layer=2 filter=252 channel=89
					20, 18, -28, 13, 5, -13, 10, -3, -38,
					-- layer=2 filter=252 channel=90
					-4, 0, -9, -5, -5, -11, 3, 4, 10,
					-- layer=2 filter=252 channel=91
					25, 38, -27, 41, 22, -14, 39, -9, -27,
					-- layer=2 filter=252 channel=92
					2, -10, -13, 0, -15, -7, 36, -25, -40,
					-- layer=2 filter=252 channel=93
					54, -26, 19, -10, 35, -9, 8, 23, -35,
					-- layer=2 filter=252 channel=94
					-4, -18, -23, -19, -25, -21, 15, 0, -3,
					-- layer=2 filter=252 channel=95
					6, -11, -12, 5, -2, -1, -6, 4, 6,
					-- layer=2 filter=252 channel=96
					39, 13, 48, 26, 70, 33, 27, 35, 3,
					-- layer=2 filter=252 channel=97
					-20, -4, -65, -8, 0, -28, -22, 17, -38,
					-- layer=2 filter=252 channel=98
					3, 33, 12, 7, -32, -36, 2, 6, -3,
					-- layer=2 filter=252 channel=99
					-10, 14, -2, 5, -8, 2, 3, 28, -4,
					-- layer=2 filter=252 channel=100
					0, -49, -47, -17, -37, -65, -2, -64, -22,
					-- layer=2 filter=252 channel=101
					5, 9, -20, 37, 32, 11, 36, 13, -5,
					-- layer=2 filter=252 channel=102
					7, -11, 5, -13, 8, -16, 30, 8, -60,
					-- layer=2 filter=252 channel=103
					-15, 4, -6, 26, -44, 23, 14, 8, 16,
					-- layer=2 filter=252 channel=104
					-36, -29, 19, -6, -55, 9, -15, 8, -22,
					-- layer=2 filter=252 channel=105
					0, -19, 0, 5, 0, 4, -16, 3, 6,
					-- layer=2 filter=252 channel=106
					15, 23, -26, 39, 43, 20, 25, 13, 14,
					-- layer=2 filter=252 channel=107
					8, -2, -29, -7, -12, -12, -14, -11, -7,
					-- layer=2 filter=252 channel=108
					-14, -72, -25, -39, -70, -57, 24, -11, -61,
					-- layer=2 filter=252 channel=109
					5, -21, 21, 7, -13, 5, 11, 0, -14,
					-- layer=2 filter=252 channel=110
					27, 31, -7, 36, 31, 14, -1, -21, 10,
					-- layer=2 filter=252 channel=111
					4, 10, 0, -10, -6, 4, -3, 0, -9,
					-- layer=2 filter=252 channel=112
					-7, 23, 28, -10, 10, 18, 14, 22, 45,
					-- layer=2 filter=252 channel=113
					-20, -38, 6, -24, -65, -10, -24, 9, 11,
					-- layer=2 filter=252 channel=114
					-4, -9, 11, 9, -10, -11, 10, -5, 0,
					-- layer=2 filter=252 channel=115
					2, -6, -3, -2, 9, -4, -2, 0, 3,
					-- layer=2 filter=252 channel=116
					-14, -22, -3, -30, -35, -12, -20, -6, 9,
					-- layer=2 filter=252 channel=117
					-3, -20, 8, -6, -26, -19, 33, 9, 20,
					-- layer=2 filter=252 channel=118
					-36, 3, 24, 5, -2, 4, 7, 28, -3,
					-- layer=2 filter=252 channel=119
					11, -4, 1, -4, 7, -25, 55, 16, -33,
					-- layer=2 filter=252 channel=120
					8, 5, -5, 1, 3, -2, -9, 1, 8,
					-- layer=2 filter=252 channel=121
					2, -6, 12, -7, -6, -5, -6, -2, 3,
					-- layer=2 filter=252 channel=122
					0, 5, -12, -11, -3, 0, 7, -8, 9,
					-- layer=2 filter=252 channel=123
					2, 36, 14, 53, -14, 15, 10, 17, 18,
					-- layer=2 filter=252 channel=124
					25, 32, -18, 61, -7, -23, 10, 29, -1,
					-- layer=2 filter=252 channel=125
					-1, 0, 4, 13, 3, -5, 13, 7, -6,
					-- layer=2 filter=252 channel=126
					35, 0, 26, 27, -1, 15, 28, 17, 18,
					-- layer=2 filter=252 channel=127
					-27, -19, -18, -17, -39, -14, -13, 14, -38,
					-- layer=2 filter=253 channel=0
					-18, -21, 29, -24, 7, 26, 6, 11, 45,
					-- layer=2 filter=253 channel=1
					20, 17, 19, -19, -18, 0, -24, 10, 5,
					-- layer=2 filter=253 channel=2
					2, -2, 4, 5, 11, 0, -5, 10, 2,
					-- layer=2 filter=253 channel=3
					-11, -27, 19, 3, 13, 26, -17, -20, 26,
					-- layer=2 filter=253 channel=4
					-48, -10, -20, -19, -3, 5, -13, 25, 2,
					-- layer=2 filter=253 channel=5
					0, 11, 2, -23, -23, -7, -15, 2, 3,
					-- layer=2 filter=253 channel=6
					4, 8, 25, 21, -25, -82, -16, 16, 26,
					-- layer=2 filter=253 channel=7
					-25, -48, -13, -48, -3, -8, -7, -27, -8,
					-- layer=2 filter=253 channel=8
					-4, 10, -1, 3, 5, -8, -8, 5, 0,
					-- layer=2 filter=253 channel=9
					-29, -36, 5, -23, 20, 3, -23, 5, 28,
					-- layer=2 filter=253 channel=10
					-7, -3, 26, 0, -7, 50, 7, 15, 46,
					-- layer=2 filter=253 channel=11
					-6, -8, 0, -20, -23, -30, 0, -2, -13,
					-- layer=2 filter=253 channel=12
					-46, -35, 3, -88, -53, -27, -71, -15, -32,
					-- layer=2 filter=253 channel=13
					7, -9, 8, -1, -6, -1, 3, -4, -6,
					-- layer=2 filter=253 channel=14
					1, 1, -7, -33, -36, -29, -30, 4, -3,
					-- layer=2 filter=253 channel=15
					14, 43, 9, -44, -36, 20, 6, -13, 13,
					-- layer=2 filter=253 channel=16
					-26, -42, 26, -26, -19, 46, 10, -18, 8,
					-- layer=2 filter=253 channel=17
					-7, 2, -9, -9, 7, 10, 7, -3, -5,
					-- layer=2 filter=253 channel=18
					42, 7, -8, 50, 16, -9, 42, 19, -17,
					-- layer=2 filter=253 channel=19
					29, 35, -9, -19, 28, -4, -15, 34, 27,
					-- layer=2 filter=253 channel=20
					2, 0, 9, -3, -7, 11, -8, 4, -3,
					-- layer=2 filter=253 channel=21
					-6, -9, -12, -14, -8, 2, 0, -2, 4,
					-- layer=2 filter=253 channel=22
					8, -1, 0, -11, -7, 3, -3, -5, -2,
					-- layer=2 filter=253 channel=23
					-26, 7, -4, -3, 8, 6, 19, 30, 20,
					-- layer=2 filter=253 channel=24
					35, -24, 26, 0, -18, 31, 5, -38, 7,
					-- layer=2 filter=253 channel=25
					-49, -37, 9, -6, -54, -2, -20, -73, -68,
					-- layer=2 filter=253 channel=26
					9, 8, 0, 7, 0, -9, -1, 5, -7,
					-- layer=2 filter=253 channel=27
					-2, 9, -7, 7, 20, -7, -5, 14, 6,
					-- layer=2 filter=253 channel=28
					-34, -95, -19, -21, -13, 7, 14, 0, 19,
					-- layer=2 filter=253 channel=29
					-10, 5, 6, -3, -5, -4, 0, 6, -9,
					-- layer=2 filter=253 channel=30
					-6, 10, -26, 22, 31, 5, 10, 22, -8,
					-- layer=2 filter=253 channel=31
					-20, 26, 2, 44, -4, 5, -33, -1, 12,
					-- layer=2 filter=253 channel=32
					-6, -3, -2, -1, 6, 0, -4, -4, -5,
					-- layer=2 filter=253 channel=33
					-5, 23, -15, -40, -45, -5, -34, -38, -11,
					-- layer=2 filter=253 channel=34
					81, -10, -5, 44, -49, -10, 41, -15, 20,
					-- layer=2 filter=253 channel=35
					-14, -32, -23, -36, 1, 4, 16, 17, 14,
					-- layer=2 filter=253 channel=36
					-5, -3, -5, -14, -7, -9, -8, 1, -11,
					-- layer=2 filter=253 channel=37
					16, 4, -10, -14, 11, -17, -15, 4, -7,
					-- layer=2 filter=253 channel=38
					2, 4, -18, -6, -8, -14, -8, 10, -10,
					-- layer=2 filter=253 channel=39
					-43, -13, 24, -38, -18, 28, 1, -28, 15,
					-- layer=2 filter=253 channel=40
					-43, 4, -5, 11, -41, -24, 0, 6, -8,
					-- layer=2 filter=253 channel=41
					-1, -1, -6, 4, -3, 0, 0, -2, 0,
					-- layer=2 filter=253 channel=42
					-28, -8, 36, -18, -13, 23, -10, 13, -1,
					-- layer=2 filter=253 channel=43
					4, -15, -17, -17, 15, -1, -44, -16, 28,
					-- layer=2 filter=253 channel=44
					5, 8, -8, 7, -8, -3, 9, -7, 10,
					-- layer=2 filter=253 channel=45
					6, 7, 3, 34, 37, 45, 15, 11, 14,
					-- layer=2 filter=253 channel=46
					-24, -6, -7, -11, -8, 9, -1, 15, 19,
					-- layer=2 filter=253 channel=47
					-14, -41, -10, -42, 0, 3, -14, -20, -8,
					-- layer=2 filter=253 channel=48
					4, 9, 4, 0, -2, 8, 8, -3, 8,
					-- layer=2 filter=253 channel=49
					62, 30, -10, 48, 25, -1, 63, 38, -20,
					-- layer=2 filter=253 channel=50
					0, 3, -8, 17, 21, -13, 14, 7, -1,
					-- layer=2 filter=253 channel=51
					-1, -4, 0, -9, 2, 4, -6, 1, -15,
					-- layer=2 filter=253 channel=52
					44, 9, 34, 7, 7, -3, -9, -9, -15,
					-- layer=2 filter=253 channel=53
					-21, 52, -6, -7, -37, -20, -21, 26, -20,
					-- layer=2 filter=253 channel=54
					10, -2, -25, -22, -38, 7, -6, 14, 7,
					-- layer=2 filter=253 channel=55
					12, -11, 5, 9, -8, -8, -5, 9, 4,
					-- layer=2 filter=253 channel=56
					-18, -8, 4, 10, -9, -17, -21, 0, 1,
					-- layer=2 filter=253 channel=57
					-8, 6, 1, -3, 16, 11, -1, 10, -5,
					-- layer=2 filter=253 channel=58
					-45, -52, 1, -124, -61, -57, -52, -16, -21,
					-- layer=2 filter=253 channel=59
					22, -24, 13, -24, 2, 11, 3, 0, -8,
					-- layer=2 filter=253 channel=60
					53, 3, -23, -19, 11, -22, -1, 14, -16,
					-- layer=2 filter=253 channel=61
					19, 3, 16, 27, 20, -10, 44, 21, 18,
					-- layer=2 filter=253 channel=62
					58, 14, 44, 2, -14, -33, 7, 4, 8,
					-- layer=2 filter=253 channel=63
					-23, -43, 8, -27, 2, 18, 5, -6, 28,
					-- layer=2 filter=253 channel=64
					14, 9, 32, 18, 23, 13, 44, 22, 22,
					-- layer=2 filter=253 channel=65
					25, 6, -10, 20, 20, -30, 33, 23, -5,
					-- layer=2 filter=253 channel=66
					35, 26, 4, 1, -18, -5, -13, 30, 51,
					-- layer=2 filter=253 channel=67
					3, -12, -18, 9, 7, 14, -8, -12, 16,
					-- layer=2 filter=253 channel=68
					0, 6, 6, 6, 3, -4, -5, -4, -1,
					-- layer=2 filter=253 channel=69
					0, -11, 28, -9, 16, 12, 22, 30, 21,
					-- layer=2 filter=253 channel=70
					-34, -48, -34, -16, -16, 2, 12, 19, 16,
					-- layer=2 filter=253 channel=71
					-10, 7, 13, 16, 42, -6, 15, 22, 6,
					-- layer=2 filter=253 channel=72
					-19, -12, -27, -71, -64, -48, -46, -56, -18,
					-- layer=2 filter=253 channel=73
					-17, -3, -19, 36, 53, 52, 41, 74, 61,
					-- layer=2 filter=253 channel=74
					-24, -29, -7, -19, -44, 23, -1, 5, 36,
					-- layer=2 filter=253 channel=75
					-39, -75, -23, -54, -60, -46, 28, 22, 5,
					-- layer=2 filter=253 channel=76
					19, 27, -12, -5, -35, 10, -37, 21, -9,
					-- layer=2 filter=253 channel=77
					0, -3, -9, -5, -8, 0, 10, 3, 10,
					-- layer=2 filter=253 channel=78
					15, 3, -3, 23, -24, -17, 16, -20, -10,
					-- layer=2 filter=253 channel=79
					5, -1, 0, 0, -7, 10, 7, 6, 0,
					-- layer=2 filter=253 channel=80
					-20, -13, 15, -11, -16, 48, 3, -10, 32,
					-- layer=2 filter=253 channel=81
					-2, -2, 6, 0, 0, 9, -1, 10, 5,
					-- layer=2 filter=253 channel=82
					-8, -2, -5, -3, 8, -1, -5, -7, -5,
					-- layer=2 filter=253 channel=83
					-22, 13, -2, -1, -10, -1, 29, 16, 9,
					-- layer=2 filter=253 channel=84
					-3, 5, 12, 10, 8, 4, -7, 5, 0,
					-- layer=2 filter=253 channel=85
					2, -8, -17, 7, -7, 6, -12, -13, -4,
					-- layer=2 filter=253 channel=86
					7, 6, 8, -11, 25, -3, 9, 8, 3,
					-- layer=2 filter=253 channel=87
					31, 32, 7, 12, -15, 15, 19, 14, -33,
					-- layer=2 filter=253 channel=88
					-17, -17, -29, -1, -12, 5, 7, 4, 7,
					-- layer=2 filter=253 channel=89
					-25, 4, 4, -73, -54, -15, -30, 7, -35,
					-- layer=2 filter=253 channel=90
					0, -6, -9, -2, 7, 6, -2, 6, -3,
					-- layer=2 filter=253 channel=91
					-68, -28, -17, -118, -42, -37, -37, -14, -40,
					-- layer=2 filter=253 channel=92
					-22, 16, 18, -65, -51, -12, -64, 0, -28,
					-- layer=2 filter=253 channel=93
					9, 65, 55, -26, 16, 20, -73, 33, -20,
					-- layer=2 filter=253 channel=94
					23, 7, 22, 11, 13, -15, -15, 34, -26,
					-- layer=2 filter=253 channel=95
					13, -3, -11, 3, 5, 4, -2, -3, -7,
					-- layer=2 filter=253 channel=96
					2, 0, 17, 21, 11, 21, 33, 40, -29,
					-- layer=2 filter=253 channel=97
					-1, -12, 7, 4, 12, 8, 14, 16, 32,
					-- layer=2 filter=253 channel=98
					-36, -66, -22, -20, 4, 19, 16, 12, 15,
					-- layer=2 filter=253 channel=99
					38, 32, -20, -4, -2, 14, -10, 23, -28,
					-- layer=2 filter=253 channel=100
					-12, -33, -5, -32, -40, 12, 9, 30, 3,
					-- layer=2 filter=253 channel=101
					-30, -51, 33, -37, 0, 10, 6, -24, -48,
					-- layer=2 filter=253 channel=102
					41, 24, -10, 55, 45, 22, 65, 51, -33,
					-- layer=2 filter=253 channel=103
					30, 0, 30, -13, 10, -13, -35, 4, -9,
					-- layer=2 filter=253 channel=104
					16, 59, 7, 30, 23, -13, 27, 20, -22,
					-- layer=2 filter=253 channel=105
					11, -16, 10, -64, -72, 41, -22, 35, -5,
					-- layer=2 filter=253 channel=106
					-65, -59, 21, -34, -53, -5, -11, -36, -21,
					-- layer=2 filter=253 channel=107
					4, 14, 9, 28, 24, 16, -6, 49, -25,
					-- layer=2 filter=253 channel=108
					39, 24, 17, 37, 20, 26, 30, 36, 8,
					-- layer=2 filter=253 channel=109
					11, -3, 3, 14, -5, -6, -8, 6, 1,
					-- layer=2 filter=253 channel=110
					-15, 8, 24, -5, -18, -8, 14, -30, -8,
					-- layer=2 filter=253 channel=111
					8, 1, -11, -6, -1, 2, -1, 9, -7,
					-- layer=2 filter=253 channel=112
					-11, 6, -10, -14, -4, 8, 6, -16, -35,
					-- layer=2 filter=253 channel=113
					-12, 4, -13, 13, 33, 22, 31, 3, 0,
					-- layer=2 filter=253 channel=114
					-11, 12, 14, 7, 1, 11, 9, 5, 5,
					-- layer=2 filter=253 channel=115
					-4, -8, 6, -1, -8, -1, -4, 7, 0,
					-- layer=2 filter=253 channel=116
					14, 16, -24, 18, -25, 17, 2, 18, -21,
					-- layer=2 filter=253 channel=117
					13, -15, -36, -26, 3, -28, 0, -1, -12,
					-- layer=2 filter=253 channel=118
					21, 10, 0, 4, 1, 17, 1, 13, 28,
					-- layer=2 filter=253 channel=119
					5, -30, 17, 28, -3, -5, 18, 21, 8,
					-- layer=2 filter=253 channel=120
					8, 8, -8, 9, -7, 3, 4, 2, -8,
					-- layer=2 filter=253 channel=121
					-5, -1, -6, 1, -6, 3, 8, -7, 1,
					-- layer=2 filter=253 channel=122
					-3, 0, 2, 0, -1, 0, -5, 3, -8,
					-- layer=2 filter=253 channel=123
					-20, -14, -34, -49, -1, 16, -15, -5, -10,
					-- layer=2 filter=253 channel=124
					13, 49, 17, -27, -29, 20, -10, 19, -6,
					-- layer=2 filter=253 channel=125
					3, 9, 0, 5, -8, -5, 6, 8, -2,
					-- layer=2 filter=253 channel=126
					-8, 14, 37, -4, 17, 21, 11, 2, 31,
					-- layer=2 filter=253 channel=127
					-2, 25, -9, 1, 7, 18, -13, 5, 23,
					-- layer=2 filter=254 channel=0
					-13, -5, -6, 0, 0, 2, 24, 31, 29,
					-- layer=2 filter=254 channel=1
					21, 29, 2, 13, 20, 7, -21, 2, 12,
					-- layer=2 filter=254 channel=2
					-6, -5, 2, 9, 3, 8, 10, 5, -3,
					-- layer=2 filter=254 channel=3
					-31, -30, -57, 3, -30, 5, 62, 21, 40,
					-- layer=2 filter=254 channel=4
					32, 34, 33, 12, 4, -37, -54, -22, -41,
					-- layer=2 filter=254 channel=5
					-1, -54, -6, 1, 3, -6, 46, -12, 38,
					-- layer=2 filter=254 channel=6
					13, -19, -5, 42, 14, -24, 5, 64, 22,
					-- layer=2 filter=254 channel=7
					4, 18, -4, 8, 34, 38, 14, 41, 3,
					-- layer=2 filter=254 channel=8
					-3, -3, 9, 12, -5, -9, -8, -2, 10,
					-- layer=2 filter=254 channel=9
					0, 31, -2, -13, -6, 15, 49, 10, 31,
					-- layer=2 filter=254 channel=10
					-24, -4, 10, -7, 12, 3, 43, 4, 26,
					-- layer=2 filter=254 channel=11
					-15, -35, 0, 17, -11, -21, 40, 19, 19,
					-- layer=2 filter=254 channel=12
					1, 0, -10, 11, 17, 28, 7, 9, 4,
					-- layer=2 filter=254 channel=13
					0, -8, -3, -6, 1, -7, 10, -11, 1,
					-- layer=2 filter=254 channel=14
					19, -10, 2, 9, 7, 6, -19, -8, 9,
					-- layer=2 filter=254 channel=15
					-53, -24, 35, -26, -46, -21, -59, 28, 11,
					-- layer=2 filter=254 channel=16
					34, 40, 3, -36, -25, 28, -58, -83, -39,
					-- layer=2 filter=254 channel=17
					4, -1, 1, -4, 7, -1, 5, -6, 0,
					-- layer=2 filter=254 channel=18
					-9, 0, 21, -29, -16, -17, -42, -30, -12,
					-- layer=2 filter=254 channel=19
					18, 15, -40, -10, 17, -16, 0, 21, -24,
					-- layer=2 filter=254 channel=20
					-3, 6, -1, 2, -6, -1, -7, 7, 3,
					-- layer=2 filter=254 channel=21
					-13, -11, -18, -9, 9, -2, 4, -8, 1,
					-- layer=2 filter=254 channel=22
					3, -9, 6, 7, 0, 4, -1, -8, 0,
					-- layer=2 filter=254 channel=23
					42, 45, 16, -34, 14, 14, -6, -21, -34,
					-- layer=2 filter=254 channel=24
					-38, -16, -35, 0, -15, -42, 48, 23, 15,
					-- layer=2 filter=254 channel=25
					-48, -43, 0, 8, -29, -40, 66, 22, 25,
					-- layer=2 filter=254 channel=26
					6, 4, 2, 0, -8, -6, 2, -3, -1,
					-- layer=2 filter=254 channel=27
					43, 29, 14, 16, -20, -24, -8, -25, -23,
					-- layer=2 filter=254 channel=28
					-17, -14, -8, 30, 21, 39, 20, 32, -2,
					-- layer=2 filter=254 channel=29
					0, 1, 2, -4, -1, 6, 5, 5, 7,
					-- layer=2 filter=254 channel=30
					7, 33, 26, -27, 8, 23, -41, -25, -26,
					-- layer=2 filter=254 channel=31
					15, 7, 34, -37, -46, -2, 30, 28, 26,
					-- layer=2 filter=254 channel=32
					-7, 7, -1, 6, 9, -11, -1, -3, 8,
					-- layer=2 filter=254 channel=33
					8, -29, -11, 18, -36, -6, -26, -22, 18,
					-- layer=2 filter=254 channel=34
					52, 9, -44, 36, -21, 4, -8, -23, -69,
					-- layer=2 filter=254 channel=35
					5, -38, -50, 16, 15, -8, 21, 7, -47,
					-- layer=2 filter=254 channel=36
					-7, -4, 0, 4, 2, 2, 7, -4, -11,
					-- layer=2 filter=254 channel=37
					0, -24, 14, 26, -22, 0, 2, -5, 17,
					-- layer=2 filter=254 channel=38
					33, 5, -1, -14, -12, -24, -6, -5, -27,
					-- layer=2 filter=254 channel=39
					21, 0, 3, -5, 14, 18, -6, -79, -64,
					-- layer=2 filter=254 channel=40
					-16, -63, 19, 29, -3, 45, -23, -30, -7,
					-- layer=2 filter=254 channel=41
					-10, 0, -11, -9, 6, 2, 9, 8, 3,
					-- layer=2 filter=254 channel=42
					23, 31, 0, -16, 32, -4, -44, -22, -56,
					-- layer=2 filter=254 channel=43
					-16, -41, -9, 6, -34, -9, 53, 1, 26,
					-- layer=2 filter=254 channel=44
					-4, -3, 3, 1, -1, 9, -1, -6, 0,
					-- layer=2 filter=254 channel=45
					4, -27, -31, -34, 8, -15, -55, -51, -45,
					-- layer=2 filter=254 channel=46
					20, 1, 6, 14, -7, -2, -6, -6, -26,
					-- layer=2 filter=254 channel=47
					38, 25, -2, 69, 7, 58, -16, 25, 18,
					-- layer=2 filter=254 channel=48
					-4, -7, 0, -2, -1, -6, 0, 4, 0,
					-- layer=2 filter=254 channel=49
					-9, -18, 2, -29, 11, -4, -45, -27, -4,
					-- layer=2 filter=254 channel=50
					19, 8, 9, -5, 2, 8, 5, 13, 11,
					-- layer=2 filter=254 channel=51
					-23, -47, -1, 11, -13, -19, 43, 13, 14,
					-- layer=2 filter=254 channel=52
					5, -20, -6, 1, -8, -26, 36, 7, 14,
					-- layer=2 filter=254 channel=53
					-5, -2, 16, 31, 10, -28, -3, 4, 15,
					-- layer=2 filter=254 channel=54
					10, -28, -18, 7, 42, -22, -2, 17, 15,
					-- layer=2 filter=254 channel=55
					6, -5, 10, 1, -4, 3, -5, 3, -8,
					-- layer=2 filter=254 channel=56
					-13, -25, -4, 17, -21, -16, 40, 26, 39,
					-- layer=2 filter=254 channel=57
					0, 8, 10, 3, -8, -5, 3, 14, 7,
					-- layer=2 filter=254 channel=58
					8, -6, -21, 0, -1, 23, -19, 10, -11,
					-- layer=2 filter=254 channel=59
					-8, 33, -19, -25, -9, -2, -18, -10, -61,
					-- layer=2 filter=254 channel=60
					0, -19, 0, -17, 22, -4, -11, -12, -43,
					-- layer=2 filter=254 channel=61
					-10, -8, 18, -22, -5, 30, -18, -17, -26,
					-- layer=2 filter=254 channel=62
					-7, -36, -43, 4, 6, -27, -7, 24, -25,
					-- layer=2 filter=254 channel=63
					7, 25, 20, -36, -1, 27, -26, 0, -21,
					-- layer=2 filter=254 channel=64
					0, 40, -3, -31, 8, 21, -53, -34, -27,
					-- layer=2 filter=254 channel=65
					5, -13, 11, -4, 18, -21, -11, 13, 18,
					-- layer=2 filter=254 channel=66
					-1, 14, 23, -27, 24, -48, 18, 38, 11,
					-- layer=2 filter=254 channel=67
					3, 1, -4, 19, -2, -7, 28, -24, 0,
					-- layer=2 filter=254 channel=68
					9, -3, 10, 0, 5, -7, 0, -3, -4,
					-- layer=2 filter=254 channel=69
					35, 63, 14, -15, 38, 13, -79, -26, -30,
					-- layer=2 filter=254 channel=70
					6, -23, -3, 9, 12, 8, 13, 5, -10,
					-- layer=2 filter=254 channel=71
					26, 17, -23, 12, -24, -27, 35, -7, 18,
					-- layer=2 filter=254 channel=72
					3, -14, 11, -7, -14, -20, -12, 21, 11,
					-- layer=2 filter=254 channel=73
					12, 17, -32, -22, 8, 10, 9, -35, 8,
					-- layer=2 filter=254 channel=74
					6, -1, 21, 8, -11, 1, -15, -58, -51,
					-- layer=2 filter=254 channel=75
					-31, -15, 1, 2, -25, 40, -10, -37, -22,
					-- layer=2 filter=254 channel=76
					-21, -12, 1, 18, -4, 0, -37, -19, 18,
					-- layer=2 filter=254 channel=77
					12, 2, -7, 1, 2, 5, 1, -2, 1,
					-- layer=2 filter=254 channel=78
					-42, -41, -16, 17, 0, -1, 45, 9, 22,
					-- layer=2 filter=254 channel=79
					9, -7, 0, 8, 3, 0, -3, -7, 1,
					-- layer=2 filter=254 channel=80
					24, 30, 15, -25, -18, -16, -15, -68, -71,
					-- layer=2 filter=254 channel=81
					0, 4, -14, -17, -17, -1, 0, -7, -14,
					-- layer=2 filter=254 channel=82
					5, 0, 3, -7, -7, -6, 9, -1, 2,
					-- layer=2 filter=254 channel=83
					32, 38, 54, -47, -9, 6, -33, -43, -54,
					-- layer=2 filter=254 channel=84
					10, 0, 4, 1, 3, 3, -2, -1, -4,
					-- layer=2 filter=254 channel=85
					3, -5, 18, -6, 14, -16, -13, 9, 10,
					-- layer=2 filter=254 channel=86
					-6, 18, -5, -4, 6, 0, 0, 1, -3,
					-- layer=2 filter=254 channel=87
					12, -16, -26, -14, -12, -22, -34, 33, -45,
					-- layer=2 filter=254 channel=88
					18, 18, 21, -13, -1, 36, -71, -28, -17,
					-- layer=2 filter=254 channel=89
					1, -2, -13, 1, 9, 0, -20, 18, -14,
					-- layer=2 filter=254 channel=90
					5, -2, -7, -1, -6, -3, 1, -2, 0,
					-- layer=2 filter=254 channel=91
					-16, -38, -14, -3, -3, 10, -2, -16, -32,
					-- layer=2 filter=254 channel=92
					21, 14, 0, 12, 6, 3, -9, 4, -5,
					-- layer=2 filter=254 channel=93
					-32, 3, -31, 26, -22, -32, 17, 11, 37,
					-- layer=2 filter=254 channel=94
					21, 50, 44, -10, 67, 12, 6, 50, 26,
					-- layer=2 filter=254 channel=95
					1, -1, 5, 12, 0, -11, 8, -2, -1,
					-- layer=2 filter=254 channel=96
					13, -17, -30, 27, 49, 40, 21, 25, 32,
					-- layer=2 filter=254 channel=97
					-10, 16, -29, -15, 7, 10, 12, 19, -16,
					-- layer=2 filter=254 channel=98
					8, -18, -12, 43, 12, 37, 13, 40, -3,
					-- layer=2 filter=254 channel=99
					11, -21, 3, 8, -11, -1, 5, -24, -3,
					-- layer=2 filter=254 channel=100
					51, 16, 2, -11, 16, 2, -61, -43, -39,
					-- layer=2 filter=254 channel=101
					-14, -12, -26, 3, -15, -31, 60, 0, -3,
					-- layer=2 filter=254 channel=102
					-1, -9, -26, -5, 47, 0, 16, 22, -9,
					-- layer=2 filter=254 channel=103
					-17, -18, 3, -3, -1, 8, -24, -25, -25,
					-- layer=2 filter=254 channel=104
					5, -41, -8, -22, 5, -21, -42, 12, 17,
					-- layer=2 filter=254 channel=105
					-3, -6, 28, 0, 2, 3, -32, 11, 29,
					-- layer=2 filter=254 channel=106
					-64, -41, -37, -10, -42, -38, 59, 0, -3,
					-- layer=2 filter=254 channel=107
					25, -12, 2, -29, 20, -28, 43, 24, -31,
					-- layer=2 filter=254 channel=108
					11, 4, -11, 12, -2, 15, -18, -26, -15,
					-- layer=2 filter=254 channel=109
					0, 0, -1, 7, -5, -1, 8, -18, -6,
					-- layer=2 filter=254 channel=110
					0, -8, 13, -6, -17, -5, -21, -3, 23,
					-- layer=2 filter=254 channel=111
					-11, 8, 5, -12, -7, 5, 0, -3, 1,
					-- layer=2 filter=254 channel=112
					-17, -39, 3, 15, 15, -42, 52, 10, -2,
					-- layer=2 filter=254 channel=113
					-17, -8, 42, -31, 15, 28, -17, -20, -4,
					-- layer=2 filter=254 channel=114
					-7, 4, 13, -9, -6, 2, -10, -7, -4,
					-- layer=2 filter=254 channel=115
					-7, -10, -12, 5, -3, 10, -5, 3, -1,
					-- layer=2 filter=254 channel=116
					-3, -16, 16, -21, -20, 19, -19, 16, -14,
					-- layer=2 filter=254 channel=117
					0, -14, -77, 52, 37, 3, 40, 40, 9,
					-- layer=2 filter=254 channel=118
					-2, -17, -19, 7, -21, 13, 27, -11, 0,
					-- layer=2 filter=254 channel=119
					47, 42, -33, -36, 5, -18, -36, -56, -15,
					-- layer=2 filter=254 channel=120
					-6, -2, 2, 5, 7, 1, 6, 2, -3,
					-- layer=2 filter=254 channel=121
					8, -8, 4, -3, 9, -2, -6, 9, 4,
					-- layer=2 filter=254 channel=122
					-13, 1, 6, -9, -7, -5, -13, -5, -8,
					-- layer=2 filter=254 channel=123
					19, 17, -2, 7, 29, 0, -12, 28, 7,
					-- layer=2 filter=254 channel=124
					-77, -12, -52, -32, 35, -4, -15, 25, -8,
					-- layer=2 filter=254 channel=125
					-6, -7, 10, -1, 6, 4, -7, -3, -8,
					-- layer=2 filter=254 channel=126
					11, 7, -12, -14, -40, 47, 29, -3, -2,
					-- layer=2 filter=254 channel=127
					17, 16, 3, -4, 19, 7, -32, -13, 17,
					-- layer=2 filter=255 channel=0
					5, -2, 1, -11, -12, -8, 6, -8, -3,
					-- layer=2 filter=255 channel=1
					-20, -11, -16, -2, -14, -18, -5, -7, -7,
					-- layer=2 filter=255 channel=2
					3, -8, -9, 5, -6, -8, -11, 7, 3,
					-- layer=2 filter=255 channel=3
					-2, -3, -14, -1, -18, 12, 1, -9, 6,
					-- layer=2 filter=255 channel=4
					-8, -6, -1, -9, -6, -13, 3, -8, -11,
					-- layer=2 filter=255 channel=5
					-7, 5, -7, -9, -11, -13, -1, -11, -11,
					-- layer=2 filter=255 channel=6
					-1, -4, 0, 6, -13, -1, 14, 2, -7,
					-- layer=2 filter=255 channel=7
					12, -9, -12, -10, -2, 4, 5, 0, -15,
					-- layer=2 filter=255 channel=8
					11, -8, 3, 0, -2, -8, -9, 0, 3,
					-- layer=2 filter=255 channel=9
					-12, -8, -4, 4, 0, -7, -2, 0, -5,
					-- layer=2 filter=255 channel=10
					0, -15, -5, 0, -9, 1, -7, -2, -5,
					-- layer=2 filter=255 channel=11
					-9, -5, -8, 0, -11, -7, 5, -11, -4,
					-- layer=2 filter=255 channel=12
					-16, -1, -8, -6, 0, -18, -12, -10, 5,
					-- layer=2 filter=255 channel=13
					-4, -10, 5, 6, -1, -10, -1, -3, -7,
					-- layer=2 filter=255 channel=14
					-4, 1, -2, -9, -1, 0, -12, -5, 0,
					-- layer=2 filter=255 channel=15
					0, 3, 6, -2, 5, -9, 5, 0, -10,
					-- layer=2 filter=255 channel=16
					10, 10, 7, -3, -12, -12, -1, -4, -1,
					-- layer=2 filter=255 channel=17
					0, 6, -5, 9, 6, 9, -7, 3, -2,
					-- layer=2 filter=255 channel=18
					-2, 10, -6, -18, -3, -13, 8, 7, -4,
					-- layer=2 filter=255 channel=19
					4, 3, 0, -12, -1, -14, -1, -9, -7,
					-- layer=2 filter=255 channel=20
					2, -4, 5, 0, -9, -1, 1, 6, 8,
					-- layer=2 filter=255 channel=21
					-7, 6, 7, 0, 0, 0, 2, 0, -8,
					-- layer=2 filter=255 channel=22
					4, 0, 5, 3, 5, -1, 0, 11, 10,
					-- layer=2 filter=255 channel=23
					-4, -7, 0, -19, 4, 9, 5, -7, 0,
					-- layer=2 filter=255 channel=24
					0, -6, -8, 1, -3, -5, -9, -1, -6,
					-- layer=2 filter=255 channel=25
					-15, -11, -1, -1, -15, -12, -13, -2, -7,
					-- layer=2 filter=255 channel=26
					3, 5, 3, 9, -9, -9, 0, -9, 8,
					-- layer=2 filter=255 channel=27
					-15, -4, -13, -13, -8, -10, -9, -16, -9,
					-- layer=2 filter=255 channel=28
					-5, -2, 1, -4, 10, 0, -2, 5, -15,
					-- layer=2 filter=255 channel=29
					2, -6, -7, -11, 5, -6, -4, -9, -1,
					-- layer=2 filter=255 channel=30
					-4, -10, 3, -2, -1, -13, -2, -14, -12,
					-- layer=2 filter=255 channel=31
					-5, 8, -10, 8, -11, -7, -5, 3, -4,
					-- layer=2 filter=255 channel=32
					-7, 1, -11, 7, -5, 7, -11, 0, -9,
					-- layer=2 filter=255 channel=33
					3, 1, 1, -17, -4, 0, -10, -15, -14,
					-- layer=2 filter=255 channel=34
					-6, -8, -9, -2, -8, -6, -7, -6, 2,
					-- layer=2 filter=255 channel=35
					-1, -5, -16, 8, 4, -13, -10, 3, -4,
					-- layer=2 filter=255 channel=36
					5, 6, -8, -2, 0, -4, -11, 2, -4,
					-- layer=2 filter=255 channel=37
					5, -5, -15, -12, -12, -8, 7, -7, -9,
					-- layer=2 filter=255 channel=38
					3, 3, 0, 0, -7, -18, -4, 0, -5,
					-- layer=2 filter=255 channel=39
					1, 7, 0, -1, -6, -18, 0, -19, -9,
					-- layer=2 filter=255 channel=40
					-12, -12, 4, -16, 9, -5, -7, -15, -11,
					-- layer=2 filter=255 channel=41
					-3, 5, -4, 1, -1, -4, 1, 6, -6,
					-- layer=2 filter=255 channel=42
					-2, -4, 0, 1, -10, -2, -11, -13, 12,
					-- layer=2 filter=255 channel=43
					-10, -3, 3, -8, 4, 5, 0, 3, -10,
					-- layer=2 filter=255 channel=44
					-6, -8, -1, -2, -9, -2, -9, 3, 6,
					-- layer=2 filter=255 channel=45
					0, 8, -8, -12, 7, 0, 3, 0, 0,
					-- layer=2 filter=255 channel=46
					6, -12, -7, 4, -11, -8, 3, -9, -7,
					-- layer=2 filter=255 channel=47
					4, -12, -15, 8, -5, -17, -2, 2, -20,
					-- layer=2 filter=255 channel=48
					-9, -11, -8, -7, -9, -3, 10, -7, 2,
					-- layer=2 filter=255 channel=49
					-6, 0, 0, -11, -11, -12, -2, 1, 0,
					-- layer=2 filter=255 channel=50
					-1, 8, -1, 4, 7, 1, -1, 4, -1,
					-- layer=2 filter=255 channel=51
					-4, -1, -14, -10, -10, -3, -2, -8, -9,
					-- layer=2 filter=255 channel=52
					0, -7, -7, -4, -12, -9, 9, 9, -8,
					-- layer=2 filter=255 channel=53
					-15, 3, -8, 0, -6, -11, 13, 11, -1,
					-- layer=2 filter=255 channel=54
					-2, -13, -11, 3, 1, 0, -8, -10, 1,
					-- layer=2 filter=255 channel=55
					5, 7, 3, 5, 10, 7, 0, -6, 6,
					-- layer=2 filter=255 channel=56
					0, -3, 2, -3, -5, -1, 1, 0, 6,
					-- layer=2 filter=255 channel=57
					1, -9, -11, -11, 1, 7, -8, -4, 8,
					-- layer=2 filter=255 channel=58
					-13, -8, 3, 9, -7, -16, -5, -7, -15,
					-- layer=2 filter=255 channel=59
					5, -14, 0, 11, -9, -15, 0, 1, -14,
					-- layer=2 filter=255 channel=60
					-5, -4, -2, 0, -7, -2, -14, 5, -3,
					-- layer=2 filter=255 channel=61
					3, -15, -14, -12, -11, 4, -4, -3, 4,
					-- layer=2 filter=255 channel=62
					-12, -8, 5, -21, -16, 8, 3, 5, 6,
					-- layer=2 filter=255 channel=63
					3, -14, -2, -6, -7, 0, -15, -8, 0,
					-- layer=2 filter=255 channel=64
					-8, -4, -9, -6, 1, 3, -4, -4, 4,
					-- layer=2 filter=255 channel=65
					-1, -10, -7, -4, 0, -2, -2, -11, 0,
					-- layer=2 filter=255 channel=66
					0, -7, 0, -10, -6, 0, 1, 0, -9,
					-- layer=2 filter=255 channel=67
					-5, -4, 0, 5, 6, -1, 6, 5, 1,
					-- layer=2 filter=255 channel=68
					5, -10, -5, 2, -9, 0, 0, -11, 2,
					-- layer=2 filter=255 channel=69
					-9, -12, -1, -1, 0, 0, -18, -6, -3,
					-- layer=2 filter=255 channel=70
					-1, -21, -4, 2, 3, -11, -9, -7, -13,
					-- layer=2 filter=255 channel=71
					4, -11, -10, -2, -12, 0, 7, -6, -3,
					-- layer=2 filter=255 channel=72
					10, 7, 1, -5, 9, 9, 7, -2, 2,
					-- layer=2 filter=255 channel=73
					5, 20, 1, -4, -10, 1, -2, 8, 0,
					-- layer=2 filter=255 channel=74
					-10, -4, 4, 3, 4, -3, -10, -3, -7,
					-- layer=2 filter=255 channel=75
					-18, 2, 6, 1, 11, -15, -23, -15, 1,
					-- layer=2 filter=255 channel=76
					-3, 2, -4, -16, -4, 6, 11, 3, -1,
					-- layer=2 filter=255 channel=77
					2, -7, -4, -11, -9, -4, -3, 3, 6,
					-- layer=2 filter=255 channel=78
					-7, -2, 7, -4, -12, -5, 6, -13, -14,
					-- layer=2 filter=255 channel=79
					2, -7, -3, 8, -1, -2, -3, 2, 4,
					-- layer=2 filter=255 channel=80
					-13, 5, -10, 4, 0, -6, -9, -3, 3,
					-- layer=2 filter=255 channel=81
					7, -6, 5, 1, -11, 7, 2, 6, 4,
					-- layer=2 filter=255 channel=82
					4, 3, -4, -3, 8, -6, 3, 3, -1,
					-- layer=2 filter=255 channel=83
					-12, 5, -10, -13, 1, 2, 4, -10, -12,
					-- layer=2 filter=255 channel=84
					-3, -6, -10, 4, 0, 5, -9, -2, -11,
					-- layer=2 filter=255 channel=85
					-3, -8, 0, -9, 6, -4, -5, -2, 2,
					-- layer=2 filter=255 channel=86
					2, 2, -3, 9, 0, 3, -2, -8, 11,
					-- layer=2 filter=255 channel=87
					-10, 0, 5, 1, -1, 7, 9, -15, -5,
					-- layer=2 filter=255 channel=88
					-1, -8, -12, 6, -13, -4, -7, -22, -15,
					-- layer=2 filter=255 channel=89
					-14, -7, 3, -3, -6, -14, -9, 7, -14,
					-- layer=2 filter=255 channel=90
					-9, 2, -1, -1, 5, 9, -9, 0, 3,
					-- layer=2 filter=255 channel=91
					-14, 0, -5, 4, -4, -7, -2, -10, -3,
					-- layer=2 filter=255 channel=92
					-15, -5, -9, 9, -13, -14, 4, 2, 1,
					-- layer=2 filter=255 channel=93
					-1, -5, -4, -1, -9, -13, 8, -7, -7,
					-- layer=2 filter=255 channel=94
					16, 3, -10, -11, -7, 0, 9, 7, -9,
					-- layer=2 filter=255 channel=95
					-4, -9, 0, -8, -8, -9, 6, 2, -5,
					-- layer=2 filter=255 channel=96
					-1, -7, 0, 2, 11, -13, 4, 0, 0,
					-- layer=2 filter=255 channel=97
					4, 2, -1, -12, -14, -7, -5, 0, -1,
					-- layer=2 filter=255 channel=98
					0, -21, -5, 7, 9, 6, 2, -12, -2,
					-- layer=2 filter=255 channel=99
					16, -7, -10, 1, -11, -9, 11, -9, -18,
					-- layer=2 filter=255 channel=100
					0, -4, 2, 0, -4, -12, 4, -9, -10,
					-- layer=2 filter=255 channel=101
					1, -8, -5, -4, -4, -10, -4, -2, 1,
					-- layer=2 filter=255 channel=102
					-23, -5, -19, -2, -2, -6, 5, 2, 1,
					-- layer=2 filter=255 channel=103
					6, -4, -1, 0, -8, -1, 4, -9, 1,
					-- layer=2 filter=255 channel=104
					0, 0, 2, -9, -15, 3, -1, -13, 5,
					-- layer=2 filter=255 channel=105
					12, 5, -3, -4, -4, -10, 12, 12, 6,
					-- layer=2 filter=255 channel=106
					-13, -9, -7, 9, -7, -4, -4, -8, -3,
					-- layer=2 filter=255 channel=107
					-4, 5, 1, 3, -1, 2, -6, 6, -10,
					-- layer=2 filter=255 channel=108
					-14, -4, -7, -13, 5, -6, -10, -8, -7,
					-- layer=2 filter=255 channel=109
					0, -9, -7, 7, -7, -8, 8, -7, -8,
					-- layer=2 filter=255 channel=110
					-1, -9, -12, -14, -7, -2, -8, -5, 3,
					-- layer=2 filter=255 channel=111
					-3, -5, -9, 7, -6, 7, 4, 9, 0,
					-- layer=2 filter=255 channel=112
					-8, 4, 1, 0, 4, -9, -4, -3, 2,
					-- layer=2 filter=255 channel=113
					8, -4, -13, 0, -6, -15, -8, -18, -12,
					-- layer=2 filter=255 channel=114
					8, 0, 1, 7, 2, 3, 8, 4, 5,
					-- layer=2 filter=255 channel=115
					0, 2, 5, -1, -1, -1, -3, -10, 0,
					-- layer=2 filter=255 channel=116
					-20, 5, -12, -12, 11, 1, 12, -11, 10,
					-- layer=2 filter=255 channel=117
					0, -3, -8, -2, -9, -9, 3, 7, -17,
					-- layer=2 filter=255 channel=118
					-10, 7, -13, -4, -5, -6, 0, -3, -2,
					-- layer=2 filter=255 channel=119
					-9, -8, -12, 2, -5, -10, -2, -11, 3,
					-- layer=2 filter=255 channel=120
					1, 9, -9, -4, 0, -6, -9, 3, -7,
					-- layer=2 filter=255 channel=121
					3, 5, 2, 3, -2, 3, 0, 10, -3,
					-- layer=2 filter=255 channel=122
					-3, 0, -3, -3, -5, 6, 1, 3, 0,
					-- layer=2 filter=255 channel=123
					2, -6, -12, -7, 10, -9, 12, -1, -9,
					-- layer=2 filter=255 channel=124
					-1, -7, 4, -8, -14, 2, 10, -1, -2,
					-- layer=2 filter=255 channel=125
					2, -10, 2, 1, 3, 0, -8, -3, 8,
					-- layer=2 filter=255 channel=126
					5, -8, -2, -2, -11, -5, -5, 5, -8,
					-- layer=2 filter=255 channel=127
					1, 2, -1, 5, -11, 0, 1, -10, -5,

			0, 0, 0, 0, 0, 0, 0, 
			23, 0, 0, 58, 0, 119, 14, 
			98, 86, 0, 114, 0, 110, 0, 
			76, 34, 0, 71, 43, 68, 0, 
			39, 158, 192, 0, 0, 0, 0, 
			0, 6, 8, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 3, 
			0, 0, 0, 0, 13, 0, 0, 
			0, 0, 6, 0, 0, 0, 0, 
			0, 0, 57, 0, 38, 0, 0, 
			0, 0, 0, 0, 10, 0, 0, 
			114, 0, 40, 27, 0, 0, 0, 
			0, 195, 0, 0, 0, 2, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 5, 
			0, 0, 0, 0, 0, 15, 0, 
			0, 0, 0, 29, 47, 50, 51, 
			0, 0, 0, 32, 57, 36, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			9, 0, 0, 0, 63, 0, 0, 
			0, 0, 0, 0, 146, 0, 0, 
			0, 0, 0, 0, 21, 0, 0, 
			0, 128, 126, 0, 0, 0, 0, 
			0, 111, 0, 0, 0, 80, 44, 
			232, 0, 0, 11, 84, 89, 124, 
			

			0, 0, 4, 49, 0, 24, 0, 
			0, 0, 0, 56, 59, 84, 40, 
			111, 132, 0, 62, 50, 56, 0, 
			0, 0, 146, 57, 171, 92, 57, 
			14, 71, 15, 0, 42, 0, 58, 
			0, 148, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 36, 0, 0, 0, 0, 0, 
			0, 0, 0, 61, 0, 0, 236, 
			0, 277, 0, 0, 0, 216, 0, 
			0, 131, 0, 0, 0, 268, 0, 
			0, 0, 90, 0, 0, 70, 0, 
			0, 0, 104, 0, 37, 0, 0, 
			186, 0, 0, 2, 0, 0, 0, 
			

			0, 0, 0, 0, 70, 198, 0, 
			179, 0, 209, 29, 0, 70, 43, 
			0, 0, 0, 0, 0, 0, 0, 
			7, 23, 0, 0, 0, 0, 0, 
			0, 43, 274, 0, 3, 80, 0, 
			0, 0, 0, 151, 26, 0, 42, 
			25, 0, 0, 0, 32, 12, 42, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			45, 62, 0, 0, 0, 0, 34, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 22, 0, 0, 0, 44, 
			2, 0, 0, 0, 0, 0, 0, 
			75, 0, 0, 68, 0, 0, 0, 
			0, 90, 0, 29, 32, 2, 0, 
			

			0, 0, 0, 0, 0, 20, 0, 
			0, 0, 0, 82, 0, 111, 0, 
			0, 0, 0, 101, 0, 50, 56, 
			0, 0, 0, 78, 0, 0, 53, 
			77, 0, 33, 0, 4, 0, 0, 
			0, 0, 0, 0, 21, 45, 11, 
			0, 0, 0, 21, 39, 18, 0, 
			

			80, 65, 51, 44, 45, 31, 47, 
			41, 89, 62, 8, 53, 2, 50, 
			0, 98, 86, 12, 35, 31, 25, 
			0, 52, 26, 0, 32, 48, 68, 
			0, 14, 13, 0, 0, 0, 8, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 106, 18, 0, 71, 
			0, 0, 0, 0, 8, 0, 21, 
			13, 59, 0, 0, 0, 5, 0, 
			0, 0, 99, 68, 13, 3, 0, 
			0, 0, 0, 0, 70, 13, 36, 
			125, 20, 204, 121, 0, 0, 0, 
			13, 167, 0, 0, 0, 8, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			73, 33, 77, 52, 0, 0, 42, 
			0, 0, 0, 0, 31, 0, 3, 
			0, 55, 104, 0, 51, 1, 0, 
			0, 8, 113, 33, 57, 56, 27, 
			0, 0, 0, 0, 0, 2, 21, 
			122, 0, 90, 13, 0, 0, 0, 
			0, 113, 15, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 40, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 34, 
			0, 0, 0, 0, 0, 7, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 88, 145, 265, 281, 
			158, 60, 233, 238, 271, 304, 316, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 4, 0, 0, 0, 0, 
			0, 0, 0, 0, 35, 0, 0, 
			0, 40, 0, 0, 33, 0, 0, 
			0, 0, 87, 0, 0, 0, 11, 
			0, 0, 0, 0, 0, 0, 88, 
			0, 35, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 46, 33, 77, 2, 
			6, 0, 0, 18, 15, 0, 65, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 54, 4, 0, 60, 21, 0, 
			0, 0, 53, 0, 56, 34, 0, 
			39, 0, 0, 31, 0, 0, 0, 
			0, 124, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 10, 0, 0, 
			8, 0, 0, 0, 59, 0, 0, 
			17, 0, 0, 0, 0, 0, 0, 
			0, 175, 57, 0, 0, 15, 0, 
			124, 103, 149, 98, 136, 118, 145, 
			186, 145, 123, 68, 59, 95, 70, 
			

			7, 31, 11, 63, 12, 55, 28, 
			32, 0, 13, 60, 0, 86, 54, 
			0, 0, 0, 30, 0, 5, 41, 
			0, 0, 0, 40, 0, 62, 41, 
			16, 0, 36, 0, 0, 55, 65, 
			0, 0, 0, 0, 66, 30, 36, 
			14, 0, 88, 80, 82, 57, 60, 
			

			109, 79, 96, 107, 39, 46, 89, 
			111, 117, 0, 25, 54, 0, 50, 
			0, 63, 0, 0, 22, 0, 5, 
			0, 35, 13, 0, 0, 5, 53, 
			0, 17, 0, 0, 0, 0, 29, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			193, 199, 182, 234, 140, 121, 128, 
			92, 229, 209, 73, 5, 45, 10, 
			0, 131, 103, 62, 0, 41, 0, 
			0, 43, 56, 29, 24, 10, 0, 
			21, 1, 71, 0, 64, 57, 76, 
			0, 0, 36, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			20, 7, 55, 0, 0, 0, 0, 
			0, 0, 0, 44, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 123, 0, 0, 111, 
			0, 0, 0, 0, 3, 63, 28, 
			0, 0, 32, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			6, 9, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 21, 0, 0, 
			178, 0, 56, 0, 0, 0, 15, 
			109, 0, 14, 0, 0, 0, 77, 
			173, 0, 0, 0, 0, 0, 63, 
			130, 174, 0, 0, 0, 19, 0, 
			0, 175, 0, 4, 0, 0, 12, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 55, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 94, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 39, 139, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			140, 16, 0, 0, 0, 0, 0, 
			48, 0, 234, 0, 141, 0, 39, 
			28, 0, 0, 405, 0, 0, 181, 
			0, 487, 0, 0, 0, 46, 0, 
			0, 165, 42, 0, 31, 0, 117, 
			

			0, 0, 0, 27, 140, 132, 3, 
			109, 0, 184, 95, 0, 0, 0, 
			9, 0, 0, 0, 73, 0, 8, 
			0, 55, 0, 0, 0, 0, 0, 
			0, 0, 95, 142, 11, 33, 146, 
			0, 171, 54, 0, 130, 224, 117, 
			0, 0, 0, 0, 37, 0, 22, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			40, 21, 11, 21, 13, 47, 52, 
			16, 57, 7, 45, 51, 18, 2, 
			4, 0, 84, 45, 11, 30, 25, 
			0, 49, 47, 16, 12, 15, 65, 
			2, 4, 0, 0, 23, 0, 35, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			37, 63, 53, 102, 0, 10, 0, 
			0, 44, 53, 44, 0, 0, 0, 
			0, 112, 107, 68, 0, 51, 0, 
			89, 66, 52, 64, 0, 3, 0, 
			70, 0, 0, 0, 65, 0, 0, 
			0, 0, 66, 0, 0, 0, 0, 
			0, 81, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 48, 0, 
			0, 0, 0, 0, 0, 23, 0, 
			0, 0, 0, 18, 0, 36, 0, 
			0, 0, 245, 0, 0, 144, 0, 
			7, 0, 163, 190, 213, 138, 189, 
			59, 0, 218, 159, 190, 213, 233, 
			

			0, 50, 74, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 7, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 37, 0, 
			62, 0, 266, 156, 123, 137, 108, 
			206, 10, 151, 82, 96, 117, 72, 
			

			52, 189, 1, 0, 0, 0, 0, 
			0, 31, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 69, 
			0, 0, 0, 0, 0, 0, 78, 
			0, 0, 0, 0, 0, 77, 0, 
			0, 0, 0, 0, 12, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 118, 16, 0, 0, 0, 0, 
			0, 68, 21, 0, 0, 29, 0, 
			0, 0, 0, 15, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			38, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 5, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 24, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 44, 
			0, 18, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 3, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			59, 35, 0, 0, 0, 0, 64, 
			0, 15, 0, 0, 82, 0, 0, 
			0, 113, 0, 0, 7, 0, 0, 
			0, 19, 128, 0, 0, 0, 25, 
			0, 0, 0, 0, 0, 0, 42, 
			106, 0, 0, 0, 0, 84, 30, 
			165, 0, 0, 46, 90, 124, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			98, 81, 67, 51, 31, 39, 84, 
			70, 114, 75, 38, 79, 52, 44, 
			121, 79, 102, 79, 65, 49, 31, 
			84, 103, 81, 45, 72, 26, 83, 
			49, 110, 88, 0, 8, 0, 27, 
			9, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 40, 0, 19, 
			97, 0, 34, 0, 63, 0, 0, 
			24, 0, 26, 0, 130, 0, 72, 
			152, 201, 0, 0, 0, 0, 17, 
			0, 97, 0, 0, 0, 63, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			54, 0, 0, 1, 0, 21, 133, 
			165, 90, 0, 0, 0, 0, 165, 
			0, 97, 0, 0, 0, 0, 0, 
			0, 147, 0, 0, 0, 0, 0, 
			0, 0, 28, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			12, 0, 0, 47, 120, 62, 26, 
			55, 141, 0, 0, 112, 38, 6, 
			0, 0, 73, 43, 104, 0, 81, 
			0, 66, 142, 0, 101, 0, 0, 
			0, 100, 64, 0, 0, 22, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			67, 45, 89, 67, 42, 0, 20, 
			8, 38, 24, 0, 0, 0, 32, 
			0, 147, 80, 0, 0, 0, 0, 
			0, 2, 18, 0, 51, 24, 7, 
			0, 0, 0, 0, 0, 0, 7, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			1, 0, 0, 190, 115, 3, 81, 
			0, 71, 0, 0, 36, 0, 0, 
			5, 26, 155, 0, 0, 59, 0, 
			0, 0, 0, 95, 0, 0, 0, 
			0, 0, 0, 0, 110, 15, 0, 
			93, 0, 412, 126, 48, 52, 19, 
			0, 122, 0, 0, 0, 45, 0, 
			

			100, 94, 0, 206, 258, 64, 87, 
			127, 245, 171, 0, 0, 47, 30, 
			0, 0, 82, 5, 0, 191, 38, 
			45, 137, 0, 246, 0, 53, 0, 
			0, 174, 161, 0, 65, 217, 0, 
			0, 0, 245, 86, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 42, 323, 0, 122, 20, 
			3, 64, 81, 207, 57, 186, 11, 
			127, 125, 0, 261, 48, 306, 0, 
			165, 89, 242, 147, 109, 145, 0, 
			0, 109, 118, 20, 402, 0, 0, 
			0, 58, 335, 48, 0, 0, 0, 
			0, 299, 0, 0, 0, 14, 0, 
			

			0, 0, 0, 33, 0, 148, 0, 
			151, 0, 52, 182, 0, 191, 184, 
			178, 0, 0, 344, 0, 286, 83, 
			202, 172, 0, 112, 0, 209, 0, 
			63, 106, 202, 89, 60, 30, 0, 
			0, 0, 228, 0, 3, 0, 0, 
			6, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 37, 0, 0, 42, 
			44, 190, 29, 0, 0, 79, 0, 
			85, 140, 0, 0, 3, 105, 0, 
			0, 0, 104, 58, 40, 32, 0, 
			0, 0, 0, 0, 41, 4, 0, 
			0, 182, 21, 0, 0, 4, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 33, 0, 
			29, 0, 0, 104, 0, 78, 0, 
			52, 0, 0, 63, 0, 113, 0, 
			81, 183, 9, 0, 0, 0, 0, 
			0, 50, 222, 0, 77, 0, 38, 
			0, 0, 149, 55, 35, 66, 75, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 34, 0, 0, 
			32, 0, 0, 0, 97, 0, 10, 
			32, 0, 0, 0, 0, 0, 0, 
			122, 126, 0, 59, 0, 1, 0, 
			231, 134, 0, 106, 112, 134, 151, 
			170, 142, 144, 134, 142, 166, 198, 
			

			0, 2, 0, 0, 0, 46, 0, 
			0, 0, 0, 37, 0, 0, 53, 
			0, 0, 13, 134, 0, 106, 149, 
			234, 171, 0, 0, 0, 79, 0, 
			21, 0, 0, 163, 1, 5, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			62, 69, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 22, 0, 0, 
			0, 0, 6, 0, 0, 0, 0, 
			

			240, 315, 71, 167, 0, 0, 136, 
			0, 47, 0, 0, 0, 70, 0, 
			0, 0, 0, 20, 0, 39, 0, 
			0, 0, 0, 66, 0, 14, 0, 
			105, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 55, 
			0, 0, 0, 138, 91, 94, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 1, 0, 
			0, 0, 0, 0, 0, 36, 0, 
			0, 0, 0, 0, 0, 11, 0, 
			173, 0, 141, 93, 87, 118, 104, 
			71, 110, 155, 133, 128, 173, 137, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 18, 24, 0, 0, 0, 
			0, 0, 17, 0, 0, 0, 0, 
			0, 0, 30, 0, 0, 0, 0, 
			0, 0, 58, 64, 20, 0, 68, 
			0, 94, 80, 0, 69, 81, 44, 
			0, 0, 0, 0, 0, 0, 0, 
			

			327, 330, 201, 343, 142, 124, 240, 
			184, 252, 108, 0, 0, 0, 32, 
			0, 139, 0, 0, 0, 0, 0, 
			0, 21, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 125, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 12, 0, 30, 119, 0, 
			156, 0, 142, 51, 0, 0, 93, 
			0, 77, 0, 30, 55, 0, 0, 
			14, 35, 0, 0, 83, 47, 0, 
			0, 0, 79, 32, 0, 102, 9, 
			0, 29, 0, 68, 0, 0, 0, 
			40, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 15, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 15, 0, 
			0, 0, 0, 0, 0, 70, 0, 
			0, 0, 0, 72, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 172, 12, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			149, 0, 123, 212, 0, 0, 91, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 8, 0, 
			0, 0, 0, 0, 0, 0, 169, 
			74, 0, 0, 0, 0, 0, 0, 
			8, 83, 53, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			150, 26, 0, 0, 60, 0, 0, 
			0, 0, 0, 0, 212, 0, 0, 
			0, 123, 0, 0, 0, 0, 0, 
			0, 368, 82, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			10, 0, 0, 0, 26, 43, 8, 
			53, 41, 0, 32, 82, 0, 78, 
			0, 54, 37, 0, 105, 20, 41, 
			0, 89, 22, 0, 12, 27, 60, 
			0, 68, 27, 0, 0, 0, 29, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 3, 145, 134, 
			124, 0, 0, 142, 162, 166, 105, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			4, 0, 0, 0, 35, 0, 39, 
			67, 0, 2, 0, 38, 0, 0, 
			0, 0, 0, 0, 82, 0, 0, 
			92, 89, 0, 0, 0, 0, 111, 
			137, 242, 138, 84, 95, 130, 129, 
			240, 19, 83, 96, 89, 132, 102, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 203, 0, 0, 
			200, 41, 103, 0, 0, 0, 0, 
			0, 8, 0, 0, 227, 0, 6, 
			0, 61, 0, 0, 0, 0, 0, 
			0, 99, 24, 0, 0, 247, 0, 
			0, 129, 0, 0, 188, 20, 0, 
			132, 0, 33, 0, 43, 0, 117, 
			

			0, 0, 0, 0, 0, 0, 0, 
			46, 0, 0, 0, 0, 10, 24, 
			196, 0, 0, 0, 0, 19, 0, 
			68, 0, 0, 69, 3, 19, 139, 
			90, 9, 0, 0, 0, 0, 0, 
			164, 17, 44, 29, 0, 0, 0, 
			43, 133, 38, 31, 11, 40, 59, 
			

			59, 0, 0, 95, 132, 68, 89, 
			108, 25, 0, 0, 2, 0, 44, 
			0, 0, 18, 0, 0, 0, 0, 
			0, 91, 0, 44, 0, 11, 0, 
			0, 0, 0, 0, 0, 98, 0, 
			58, 0, 120, 78, 0, 0, 0, 
			0, 38, 5, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			6, 0, 50, 209, 141, 116, 53, 
			0, 0, 41, 41, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 18, 2, 0, 0, 0, 
			0, 0, 0, 0, 49, 21, 0, 
			0, 0, 174, 157, 11, 0, 0, 
			0, 85, 59, 0, 0, 0, 0, 
			

			0, 0, 0, 87, 36, 31, 41, 
			0, 0, 0, 0, 0, 0, 29, 
			0, 48, 0, 0, 0, 15, 0, 
			0, 0, 30, 61, 19, 0, 0, 
			0, 0, 0, 0, 32, 34, 0, 
			20, 0, 138, 134, 0, 0, 0, 
			0, 77, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 1, 
			0, 0, 0, 0, 0, 61, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 2, 0, 
			0, 232, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 21, 0, 
			0, 0, 0, 109, 0, 33, 277, 
			0, 301, 0, 76, 0, 178, 0, 
			0, 0, 0, 0, 89, 237, 0, 
			0, 0, 216, 0, 0, 23, 0, 
			0, 0, 203, 0, 0, 0, 0, 
			111, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			77, 0, 30, 38, 101, 0, 91, 
			578, 198, 25, 7, 393, 20, 0, 
			394, 89, 0, 19, 850, 0, 0, 
			163, 102, 68, 121, 314, 0, 0, 
			88, 826, 171, 0, 3, 0, 0, 
			0, 430, 252, 0, 16, 0, 0, 
			42, 0, 177, 0, 0, 2, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 51, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 39, 
			4, 0, 0, 58, 51, 79, 0, 
			

			0, 0, 117, 0, 0, 2, 0, 
			40, 31, 80, 95, 0, 0, 0, 
			0, 0, 0, 139, 61, 0, 30, 
			0, 0, 0, 0, 0, 39, 0, 
			0, 94, 91, 219, 0, 0, 64, 
			0, 58, 0, 0, 1, 15, 10, 
			0, 0, 2, 25, 26, 0, 73, 
			

			116, 61, 148, 99, 131, 66, 102, 
			121, 212, 0, 68, 99, 0, 34, 
			0, 0, 0, 64, 184, 24, 120, 
			0, 161, 0, 0, 0, 10, 8, 
			0, 216, 0, 0, 42, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 137, 0, 39, 0, 
			0, 0, 0, 50, 0, 0, 0, 
			0, 0, 0, 0, 0, 27, 0, 
			0, 0, 10, 3, 0, 0, 0, 
			0, 0, 0, 0, 126, 0, 75, 
			0, 0, 176, 87, 48, 95, 131, 
			28, 261, 61, 86, 40, 94, 0, 
			

			269, 270, 251, 249, 214, 63, 238, 
			199, 295, 155, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 20, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 5, 0, 108, 0, 27, 
			141, 83, 14, 0, 260, 0, 0, 
			88, 0, 0, 0, 420, 0, 0, 
			0, 0, 206, 0, 233, 0, 4, 
			47, 283, 0, 0, 0, 0, 0, 
			2, 261, 0, 0, 0, 0, 0, 
			0, 0, 79, 0, 0, 0, 1, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			56, 0, 0, 0, 0, 0, 95, 
			0, 304, 0, 0, 14, 0, 0, 
			0, 0, 0, 0, 35, 0, 0, 
			0, 0, 76, 0, 0, 9, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			55, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 42, 0, 0, 
			25, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 66, 0, 0, 0, 0, 0, 
			0, 3, 26, 0, 0, 116, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			168, 131, 141, 175, 62, 40, 68, 
			0, 151, 51, 19, 0, 0, 0, 
			0, 5, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 27, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			166, 77, 77, 83, 19, 0, 142, 
			22, 132, 0, 0, 116, 0, 0, 
			0, 0, 0, 0, 135, 0, 0, 
			0, 45, 173, 0, 50, 0, 23, 
			62, 81, 0, 0, 0, 0, 42, 
			150, 0, 0, 0, 0, 0, 0, 
			0, 70, 33, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			45, 0, 0, 150, 58, 174, 189, 
			297, 57, 0, 0, 5, 0, 116, 
			144, 0, 0, 0, 19, 0, 45, 
			25, 68, 0, 0, 0, 8, 0, 
			0, 87, 0, 14, 107, 129, 299, 
			157, 24, 70, 160, 189, 105, 148, 
			152, 207, 194, 115, 97, 108, 159, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			1, 83, 65, 65, 0, 42, 4, 
			0, 49, 130, 64, 0, 149, 0, 
			81, 0, 35, 252, 0, 95, 50, 
			33, 0, 0, 75, 0, 29, 0, 
			84, 0, 11, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 13, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			146, 0, 205, 103, 0, 0, 82, 
			149, 0, 0, 13, 0, 24, 0, 
			155, 95, 0, 78, 0, 0, 6, 
			57, 45, 203, 71, 139, 41, 59, 
			0, 230, 140, 39, 11, 18, 15, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			197, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 325, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 29, 0, 0, 0, 30, 30, 
			0, 212, 0, 0, 85, 0, 0, 
			15, 0, 39, 0, 0, 0, 72, 
			

			0, 6, 0, 0, 0, 89, 0, 
			251, 0, 176, 78, 0, 46, 81, 
			0, 66, 0, 67, 143, 0, 0, 
			42, 2, 0, 0, 46, 0, 0, 
			0, 119, 192, 0, 0, 0, 0, 
			0, 64, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 4, 0, 0, 0, 7, 0, 
			0, 0, 0, 0, 7, 0, 42, 
			0, 0, 0, 0, 0, 12, 62, 
			35, 82, 0, 0, 0, 0, 26, 
			0, 0, 56, 0, 0, 35, 0, 
			0, 0, 0, 0, 33, 76, 67, 
			75, 0, 0, 56, 79, 54, 3, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 43, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 132, 80, 
			0, 0, 6, 26, 88, 88, 77, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 1, 0, 
			0, 0, 0, 55, 32, 12, 24, 
			41, 0, 0, 3, 0, 59, 0, 
			0, 153, 106, 7, 0, 96, 0, 
			0, 0, 0, 12, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 39, 
			0, 0, 0, 0, 0, 0, 61, 
			0, 0, 0, 0, 0, 193, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			49, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			76, 0, 0, 65, 0, 0, 0, 
			0, 0, 0, 0, 0, 162, 0, 
			0, 24, 0, 60, 0, 17, 0, 
			0, 189, 0, 0, 0, 0, 0, 
			0, 0, 229, 0, 42, 0, 0, 
			0, 0, 175, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 37, 0, 0, 
			71, 0, 88, 0, 79, 0, 0, 
			0, 5, 70, 22, 75, 0, 0, 
			0, 14, 0, 0, 25, 0, 0, 
			128, 23, 148, 13, 0, 0, 0, 
			71, 205, 59, 0, 0, 18, 0, 
			
		others=>0 );
END inmem_package;
