library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    588, 408, 450, 
    449, 458, 153, 
    35, 13, 0, 
    
    -- channel=1
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=2
    114, 147, 83, 
    0, 0, 40, 
    222, 208, 308, 
    
    -- channel=3
    196, 123, 136, 
    113, 230, 129, 
    0, 14, 24, 
    
    -- channel=4
    0, 0, 85, 
    0, 53, 230, 
    0, 0, 202, 
    
    -- channel=5
    0, 0, 0, 
    234, 0, 0, 
    0, 0, 0, 
    
    -- channel=6
    59, 0, 0, 
    0, 156, 189, 
    471, 173, 52, 
    
    -- channel=7
    272, 234, 253, 
    0, 270, 242, 
    0, 210, 203, 
    
    -- channel=8
    360, 301, 0, 
    0, 184, 76, 
    141, 192, 0, 
    
    -- channel=9
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=12
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 
    0, 0, 0, 
    91, 0, 0, 
    
    -- channel=14
    0, 0, 0, 
    0, 0, 0, 
    297, 235, 231, 
    
    -- channel=15
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=16
    0, 20, 110, 
    0, 0, 26, 
    0, 0, 0, 
    
    -- channel=17
    112, 152, 0, 
    0, 0, 14, 
    209, 259, 182, 
    
    -- channel=18
    7, 28, 0, 
    0, 0, 18, 
    0, 47, 0, 
    
    -- channel=19
    97, 215, 13, 
    0, 190, 239, 
    210, 332, 374, 
    
    -- channel=20
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=21
    417, 62, 266, 
    82, 528, 429, 
    110, 287, 339, 
    
    -- channel=22
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=23
    0, 198, 0, 
    158, 0, 21, 
    138, 191, 119, 
    
    -- channel=24
    44, 0, 297, 
    142, 136, 253, 
    0, 0, 0, 
    
    -- channel=25
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=26
    351, 297, 308, 
    129, 416, 358, 
    0, 19, 0, 
    
    -- channel=27
    0, 87, 99, 
    110, 0, 0, 
    0, 0, 0, 
    
    -- channel=28
    310, 83, 80, 
    0, 0, 158, 
    0, 41, 132, 
    
    -- channel=29
    0, 91, 0, 
    0, 0, 0, 
    599, 811, 1065, 
    
    -- channel=30
    476, 417, 214, 
    60, 27, 0, 
    0, 0, 0, 
    
    -- channel=31
    47, 274, 173, 
    241, 191, 15, 
    167, 98, 174, 
    
    -- channel=32
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=33
    0, 0, 100, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=34
    240, 360, 444, 
    0, 353, 264, 
    0, 0, 194, 
    
    -- channel=35
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=36
    0, 9, 90, 
    21, 299, 156, 
    0, 0, 0, 
    
    -- channel=37
    164, 0, 28, 
    168, 0, 49, 
    0, 103, 0, 
    
    -- channel=38
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=39
    0, 97, 0, 
    243, 287, 310, 
    701, 71, 156, 
    
    -- channel=40
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=41
    0, 0, 224, 
    140, 0, 0, 
    235, 0, 328, 
    
    -- channel=42
    56, 577, 463, 
    280, 249, 245, 
    0, 0, 0, 
    
    -- channel=43
    199, 35, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=44
    153, 214, 85, 
    173, 106, 22, 
    0, 69, 0, 
    
    -- channel=45
    89, 82, 86, 
    562, 209, 68, 
    428, 338, 192, 
    
    -- channel=46
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 
    0, 0, 0, 
    27, 0, 0, 
    
    -- channel=48
    47, 0, 0, 
    0, 0, 58, 
    0, 0, 0, 
    
    -- channel=49
    0, 399, 49, 
    261, 73, 13, 
    0, 0, 0, 
    
    -- channel=50
    539, 632, 592, 
    290, 578, 329, 
    144, 100, 141, 
    
    -- channel=51
    28, 175, 58, 
    0, 0, 0, 
    53, 0, 0, 
    
    -- channel=52
    192, 0, 0, 
    0, 171, 40, 
    236, 0, 0, 
    
    -- channel=53
    0, 0, 0, 
    0, 0, 0, 
    70, 166, 0, 
    
    -- channel=54
    585, 486, 455, 
    407, 330, 364, 
    0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 
    24, 0, 0, 
    295, 177, 80, 
    
    -- channel=56
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=57
    0, 0, 113, 
    9, 40, 2, 
    0, 0, 0, 
    
    -- channel=58
    525, 303, 140, 
    361, 106, 0, 
    171, 0, 182, 
    
    -- channel=59
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=60
    0, 0, 193, 
    0, 0, 146, 
    0, 0, 0, 
    
    -- channel=61
    398, 423, 487, 
    454, 237, 226, 
    195, 0, 0, 
    
    -- channel=62
    285, 179, 204, 
    474, 322, 225, 
    95, 173, 166, 
    
    -- channel=63
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
