library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_36k_layer0_entity13 is
    generic (
        DEVICE: string := "7SERIES"
        );
  
    port (reset   : in std_logic;
          clock   : in std_logic;
          chip_en : in std_logic;
          wr_en   : in std_logic;
          data_in : in std_logic_vector(INPUT_SIZE-1 downto 0);
          address : in std_logic_vector(11-1 downto 0);
  
          data_av  : out std_logic;
          data_out : out std_logic_vector(INPUT_SIZE-1 downto 0);
  
          n_read  : out std_logic_vector(31 downto 0);
          n_write : out std_logic_vector(31 downto 0)
          );
  end ifmap_36k_layer0_entity13;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,             -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"0017001c0013002800710073006d007400710067006a0069006900690069006b",
       INIT_01 => X"006a0063004c003a0054005600720089007c007d007c007d007f007d007a0078",
       INIT_02 => X"0018001b0014001a006a00820076007c007d0072006d00750078007600720079",
       INIT_03 => X"00850083006a0044003e0051008c0096008a008c008900880088008500810080",
       INIT_04 => X"0018001a00170012005800830074007b008b008d007400740081007f007d0084",
       INIT_05 => X"008e009a0098006900370059009f009e009700970092008e008e008b00880084",
       INIT_06 => X"00180019001900120045007c006a0073009c00a6009200780089009400950097",
       INIT_07 => X"0096009c0094006d004a007a00b100a900a1009d00980095009600940091008e",
       INIT_08 => X"00190018001900170033006d0060006800a100b800b2008d007c008000860093",
       INIT_09 => X"009700960089006c0060009800b700b500b300ae00a800a400a0009c00980093",
       INIT_0A => X"001a001a001b001c00230059005f0066009600c100c7009f0074006600620076",
       INIT_0B => X"008200830077007a008400a700a600aa00b200b700b300b700b700b100af00a9",
       INIT_0C => X"001a00160019001a001d005c0080007b009300c300c700ab007e005e0063006a",
       INIT_0D => X"0060006d0065007a00ac00c000aa00b000c300c400c500ca00c500bf00bf00c2",
       INIT_0E => X"004d0021001100190058009a009b007e008c00be00c100b900a30081007b0071",
       INIT_0F => X"005800670068007900b100c600a500bd00e400db00e000da00ba00bb00c400cd",
       INIT_10 => X"0095008000560060009b00a700990077006f00a800bf00bf00b700aa0094007f",
       INIT_11 => X"007000700074007c00a300bb00a200c100df00d500cf00bb009d00a600c400d2",
       INIT_12 => X"00a1009e0092009b00a700a9009f00750068009b00b300b500b600b4009f0087",
       INIT_13 => X"0064007400750079009e00b200b200cc00d800d600cb00a70093009600b000cf",
       INIT_14 => X"00aa00a5009e00a500af00b000a00070007b00a400b100b400b600ac00950079",
       INIT_15 => X"006a007400750076009c00a600af00d100de00d800cd00a900910093009f00ba",
       INIT_16 => X"00ac00ae00a900a600b000b0009d007a008d00b100b900b600b6009d007f0068",
       INIT_17 => X"00730084007b007d009f00a400a300ce00e000d900cd00b50092008e0093009c",
       INIT_18 => X"00a700a700a500a000a500a40099008f009100a300ae00a400a3009f00850076",
       INIT_19 => X"0086009f0087009200a300a300a800cd00df00dc00d600c700a3009000900098",
       INIT_1A => X"00a900a200a0009b00a30088008300a40092008800840085009f009e00870092",
       INIT_1B => X"00a700a20090009e0098009800b000cb00d700d800dd00da00c5009f00a200b6",
       INIT_1C => X"00ae00a400a2009d00a80078006d00b200a600a700a100a300b600ab00840078",
       INIT_1D => X"00a900a3008c009500a600a400aa00cc00d300d500da00e400d600b000bb00c7",
       INIT_1E => X"00af00a000a1009f00aa0084006800b700bc00b600b800b000a200a800a3008d",
       INIT_1F => X"009100a50092008500af00a5009600a900ca00d400d900dd00c400ba00c700c7",
       INIT_20 => X"00b3009f0092009400a10097006d00a800c700b500a400ae00a5009c00aa00a6",
       INIT_21 => X"00690088009f0077008f009e007e0050007600b700d100cd00af00b700c900c5",
       INIT_22 => X"00b500a400850083009500a50097009f00c200c700c400cd00b900a800ac00a2",
       INIT_23 => X"00680069009b0077008600ad0088005c004b006f0098009e009800b000cb00c8",
       INIT_24 => X"00b700ac008e0085009f00b000b100aa00b100c500cf00d900d900c600bb00aa",
       INIT_25 => X"0083005a0085007e008b00a20082007e006f006000760084007c009200b800c7",
       INIT_26 => X"00b900b000a1009500af00b700b600bc00aa00aa00b900c200c900d000ca00af",
       INIT_27 => X"00a4007b00710091009d008c0071007b007700700086008e007f0079008400a6",
       INIT_28 => X"00bd00b700ad009b00ab00ba00b100b200b400ac00b200b100a400bc00c300bd",
       INIT_29 => X"00c900b60088009d00930078006a007c0080008a0094008a00780077007a0082",
       INIT_2A => X"00bd00bc00b700a1009e00b700bb00b000b800bf00c000a4008b00a600ad00b1",
       INIT_2B => X"00c000bc00a200960076006b00790085008e0096008d007d0075007c007d006c",
       INIT_2C => X"00ba00ba00bb00a6009400b400c700c500c100c300c000a80091009f00a900aa",
       INIT_2D => X"00af00ac00a30086005d006c0086008b008d0097008e007c007c00720065005b",
       INIT_2E => X"00ba00b500b700ac008f00b000c900cf00ce00cb00bd00af00a500ab00ae00ac",
       INIT_2F => X"00b200ab009e007500610078008a0088008a00a1009200840082006d00640068",
       INIT_30 => X"00b800b200af00a9009200aa00c600ca00c800c500ab008800a100b400ab00aa",
       INIT_31 => X"00ad00a800900073006c007c0086007e0082009900910087007700750074006f",
       INIT_32 => X"00b800b000a8009d009300a200c000c800bf00b900810052008d00b300a6009f",
       INIT_33 => X"009f0096008400740069007a007f007a007f00840080007a00770077006b0062",
       INIT_34 => X"00b800ac00a300940086009200ba00ca00c000b200820058008c00ac00980090",
       INIT_35 => X"00910084007a00690064007700790070007a00710064006c007c007a00750072",
       INIT_36 => X"00b700a9009e008e007e008400b200cc00c300af009d009000a4009800870083",
       INIT_37 => X"007c0074006f0054006100730071006d00720066005f0064007400820082007b",
       INIT_38 => X"00b100a10099008e0077007a00b200cc00c500b400aa00a8009d0087007a007b",
       INIT_39 => X"0077006d005e004b0068006f0070007100700064005c006600770082007e0073",
       INIT_3A => X"00a30090008d00910074006b00a900c800c200b700ac00a30096008100730079",
       INIT_3B => X"00700064004e005100680065006a00720072006300630070007600750074006e",
       INIT_3C => X"008e007e0083008f007c005f009100c000be00b700b200a800820062005c0065",
       INIT_3D => X"0068005c004b005f00630061006a0074006d006c0071006e0067006c00740077",
       INIT_3E => X"007b00680070007800740057007600ae00b500ae00a4008d0063004500390046",
       INIT_3F => X"0057005100580060005d005e006b0070006b006c0061005d00650076007b0076",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INIT_40 => X"00d900d200cd00c700da00d600cf00bd00bb00ae00a600a90096009a008c008f",
       INIT_41 => X"00a700bf00db00df00db00d700e200e100db00be00af00bb00c800aa00a100a2",
       INIT_42 => X"00de00dd00dc00d700d800e100d300b300b400c000be00bc00c700ce00d100db",
       INIT_43 => X"00e500eb00ec00ec00e900e200e100e500e700d400d000cd00d800b700ba00c8",
       INIT_44 => X"00ea00e900e700e800e900ef00d900ad00a400b400ad00b700be00bc00d400e0",
       INIT_45 => X"00da00eb00e300e100e500df00d600e100ea00e800e600d800d100ca00d000d3",
       INIT_46 => X"00f500f400f400f200f400f300e4009e0092009d0083009f0091008800a2009f",
       INIT_47 => X"00a900cb00c300d300d100cb00d000e200e600e900e400d500c700db00e000d4",
       INIT_48 => X"00f500f300f400f400f500f100cf00750063006c0059006b0064005b0064005c",
       INIT_49 => X"0066007c007c009500b600b900ca00e900e100e200e300cd00c200d500e200de",
       INIT_4A => X"00f500f400f400f300f500ed00d8007e0048005a005b006600650067006b0063",
       INIT_4B => X"00590059005b005d007e00be00d800eb00e700df00d800c400ae00bd00d900ec",
       INIT_4C => X"00f500f300f300f400f100db00d9009e0050007200840097008c0084008f008a",
       INIT_4D => X"0082007a00720078006e009b00dd00e900eb00e000c600c000a700ab00cc00eb",
       INIT_4E => X"00f400f300f300f600e300c700d700990051009200bb00ca00cf009e00830083",
       INIT_4F => X"0081008d00830084009f0084009f00d700e500d700d400d100c500ab00b200dd",
       INIT_50 => X"00f400f300f400f500e300ce00da0082005100820080008100b800910074007d",
       INIT_51 => X"007c0089008e007d00990093009000c600d600db00e900dc00b800a400a900c9",
       INIT_52 => X"00f300f300f400f200e400be00a8006e005300860077006e008f008000730078",
       INIT_53 => X"007d00830092007d0095009b008c00c400e900f000f000e900c800c800d700dc",
       INIT_54 => X"00ef00f100f400f500dc00850082005f004e00740074006c006d006b006d006c",
       INIT_55 => X"007300780078007300880096008f00a700d000e400f500f300f400f500f500f4",
       INIT_56 => X"00de00e900f200f400d800a900a50059003d0043005b0064005f005f00620060",
       INIT_57 => X"0060005f005a0061006900790081007e009b00d800f800f300f400f400f400f4",
       INIT_58 => X"00d000df00ec00e300bf00b700b500640037003800580065006f006300560054",
       INIT_59 => X"00520054005d0071006d00620070008100ae00e200f500f400f400f400f400f4",
       INIT_5A => X"00c800cc00db00c300aa009a009c006600680063006c006600730075005e0055",
       INIT_5B => X"005a006a007a008c00800068006c007c009600b300c300d400ef00f500f400f4",
       INIT_5C => X"00c800d200cf00a900a400940093008a0081005c006a005d0059005d0054004d",
       INIT_5D => X"004c005100510051004f004a004b00520065007b008c008f00bf00f400f400f4",
       INIT_5E => X"00d200e200c400770070009600ba00c0006c004d004d0037002d002f003c003f",
       INIT_5F => X"003b003f003b003600310032003d00400047004b005b0067008700e100f600f4",
       INIT_60 => X"00c700c100b40060005d009100c000a100560049005c00620068004f004f0047",
       INIT_61 => X"0025001c001e001b003400320016001c00180035005b0068008000ce00f700f3",
       INIT_62 => X"00d300c700c200710078009d009f00470044005a0074007c0095007900800066",
       INIT_63 => X"004e00620070006400940093005c0063005e006c0087008e009c00b700f200f5",
       INIT_64 => X"00dc00ca00b70066006e00a50084001e00390062006b00530052006500810064",
       INIT_65 => X"009900ae009e009f00ac00a800a200a300a000af009c00770072008700e400f7",
       INIT_66 => X"00db00cf00bc00620053008d006f002a003a0048004c003e003500380040005d",
       INIT_67 => X"00a0007c005b00650074006b006700670063009b007e00430051007600d900f8",
       INIT_68 => X"00d900d200c7006500380058005d003c0038002e003f0046003c003600400041",
       INIT_69 => X"006300720069006700640060005d00610066006f006400490052007200d400f9",
       INIT_6A => X"00d100cd00ca0075005300460051004400320023002b00330044004d0057003f",
       INIT_6B => X"003400470052004800400043003e005d0058003c0053006c0070006c00cc00fa",
       INIT_6C => X"00cd00ca00c50068005d006f00470049003f002900260022004b0063008e004f",
       INIT_6D => X"001e005600930076006300720066009900b2003f004a008d0077005a00c300f6",
       INIT_6E => X"00c600c200b900570031006c00610063005f0033002700240028003200570037",
       INIT_6F => X"0020004f0097007f007a00880074009c009f00370035004a003e004e00c200f0",
       INIT_70 => X"00b600b400a9004d0025003b006c0090006a003c002b0020001d001c001e0021",
       INIT_71 => X"0027002a003a0058006a0079007a00750043002f003300320033005000ba00e1",
       INIT_72 => X"00a800a500a4007d005b0060006f008d0060004a00370024001e001e001d001f",
       INIT_73 => X"00230018004000ae00cd00cb00b300b500570026002b00300042005b00ae00d3",
       INIT_74 => X"00a200a300af00b400980076006c008d005b0053004e0030001900180019001d",
       INIT_75 => X"00270026004700a400b800b100a900a60051001e001e0031004e005f00a900ce",
       INIT_76 => X"009a00ac00b300a6009200750067009200570055005200360020001e00210025",
       INIT_77 => X"0036004d00560065006b0079008e0089003c001e00210036004e005b00a500c7",
       INIT_78 => X"00a600a9009e0094008f008500670071004f0051004b003c002a0027002a002c",
       INIT_79 => X"003000360041004d005a006e0083008b0035001d002600360046005b00a900c4",
       INIT_7A => X"00a200970093008d00890085006b004e0048004e0046003c0032002a002e0030",
       INIT_7B => X"00310033003b0042004c0059006500710045001d00230034003f006200ae00ba",
       INIT_7C => X"0094008d008e008c008f008c006a003c0042004a00420037003900340036003a",
       INIT_7D => X"003a003a00410046004900500057005d004d002500260037004a008300b300b4",
       INIT_7E => X"0090009500a000a2009e0092007e003d00390039003a00430046004500490048",
       INIT_7F => X"0044004900590062005e0061006300610052004500400047007700a400b600ba",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
