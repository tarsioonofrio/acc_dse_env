library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 7, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    55, 56, 57, 59, 57, 54, 58, 62, 58, 47, 37, 38, 44, 51, 53, 
    54, 60, 60, 60, 59, 47, 55, 46, 33, 19, 15, 15, 18, 35, 50, 
    35, 34, 58, 61, 59, 45, 26, 21, 18, 9, 17, 16, 15, 17, 35, 
    32, 15, 55, 57, 47, 35, 30, 21, 10, 10, 16, 12, 10, 11, 21, 
    23, 17, 51, 50, 43, 32, 23, 16, 9, 0, 22, 22, 14, 17, 11, 
    7, 3, 47, 30, 0, 14, 19, 26, 19, 0, 17, 14, 13, 16, 15, 
    11, 0, 23, 54, 15, 9, 20, 17, 24, 0, 14, 13, 6, 10, 21, 
    3, 10, 15, 35, 31, 18, 18, 6, 20, 13, 11, 14, 7, 14, 32, 
    2, 0, 5, 2, 19, 4, 15, 13, 15, 18, 14, 11, 6, 26, 46, 
    2, 1, 10, 0, 20, 11, 8, 21, 12, 16, 9, 7, 10, 31, 42, 
    0, 1, 9, 0, 18, 21, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    25, 25, 26, 26, 25, 21, 27, 27, 23, 19, 16, 19, 21, 23, 25, 
    26, 24, 27, 26, 27, 21, 17, 16, 12, 6, 3, 0, 4, 21, 25, 
    10, 26, 26, 26, 26, 9, 5, 0, 10, 14, 10, 15, 11, 11, 25, 
    3, 15, 24, 24, 13, 10, 12, 13, 14, 16, 8, 8, 10, 12, 22, 
    8, 16, 21, 22, 20, 6, 0, 6, 8, 12, 4, 8, 13, 17, 8, 
    0, 6, 20, 3, 0, 2, 6, 9, 9, 20, 0, 3, 13, 14, 14, 
    0, 0, 10, 21, 11, 6, 7, 6, 10, 13, 0, 3, 6, 12, 16, 
    0, 1, 0, 13, 19, 19, 2, 5, 14, 16, 5, 0, 11, 14, 24, 
    0, 0, 0, 12, 1, 0, 1, 5, 15, 0, 3, 6, 10, 25, 29, 
    0, 0, 0, 0, 5, 7, 6, 9, 0, 16, 10, 11, 21, 25, 18, 
    0, 0, 0, 11, 12, 9, 12, 4, 7, 0, 2, 10, 0, 0, 0, 
    0, 0, 9, 5, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 6, 5, 0, 0, 0, 4, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 5, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 3, 16, 0, 4, 0, 1, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 2, 16, 1, 0, 2, 0, 7, 
    13, 8, 0, 0, 14, 0, 0, 0, 0, 32, 0, 0, 7, 0, 0, 
    9, 8, 0, 0, 9, 5, 0, 0, 0, 31, 0, 1, 9, 9, 0, 
    12, 0, 6, 0, 4, 13, 0, 0, 0, 15, 0, 1, 12, 2, 0, 
    10, 16, 3, 4, 1, 5, 0, 5, 4, 0, 13, 0, 7, 0, 0, 
    8, 17, 0, 26, 2, 2, 5, 0, 14, 0, 0, 5, 7, 0, 0, 
    25, 14, 0, 38, 0, 14, 22, 4, 0, 5, 25, 26, 32, 28, 25, 
    56, 20, 1, 33, 10, 25, 40, 37, 34, 36, 38, 42, 43, 46, 43, 
    48, 53, 28, 20, 9, 35, 35, 35, 37, 41, 45, 47, 45, 45, 49, 
    48, 47, 65, 0, 25, 39, 35, 38, 39, 43, 49, 49, 46, 59, 49, 
    44, 49, 48, 36, 38, 44, 38, 33, 38, 41, 44, 45, 50, 50, 37, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 2, 
    0, 15, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 43, 0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 29, 9, 9, 0, 0, 62, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 45, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 20, 0, 10, 0, 3, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    11, 18, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 12, 0, 55, 0, 0, 36, 14, 0, 0, 0, 0, 6, 7, 0, 
    60, 34, 0, 72, 3, 0, 13, 9, 0, 4, 9, 13, 13, 16, 9, 
    10, 49, 31, 38, 0, 5, 6, 6, 5, 8, 14, 15, 19, 18, 18, 
    7, 15, 66, 10, 0, 11, 1, 6, 10, 13, 17, 20, 13, 26, 26, 
    5, 18, 20, 18, 2, 17, 15, 7, 12, 11, 8, 12, 27, 18, 0, 
    
    -- channel=6
    2, 0, 1, 4, 3, 0, 2, 3, 3, 4, 5, 0, 2, 6, 8, 
    1, 0, 0, 5, 0, 0, 22, 4, 16, 0, 6, 3, 0, 0, 4, 
    9, 0, 1, 4, 0, 0, 26, 10, 0, 0, 8, 7, 20, 0, 0, 
    51, 0, 3, 0, 6, 0, 1, 18, 4, 0, 26, 0, 18, 15, 0, 
    57, 0, 32, 0, 0, 16, 25, 24, 9, 0, 1, 36, 0, 22, 0, 
    48, 0, 42, 4, 0, 16, 17, 19, 28, 0, 36, 43, 0, 13, 18, 
    50, 0, 9, 30, 0, 0, 0, 25, 34, 0, 44, 25, 0, 0, 17, 
    34, 4, 27, 17, 0, 0, 50, 0, 23, 0, 22, 26, 0, 0, 11, 
    27, 0, 64, 0, 19, 0, 9, 0, 0, 9, 0, 36, 0, 0, 0, 
    0, 0, 56, 0, 27, 11, 0, 0, 8, 5, 34, 3, 0, 0, 8, 
    0, 0, 49, 0, 56, 19, 0, 3, 46, 22, 0, 0, 0, 0, 6, 
    0, 0, 21, 0, 52, 32, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 18, 18, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 8, 9, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 8, 9, 0, 1, 2, 4, 0, 0, 
    27, 7, 0, 0, 0, 9, 1, 3, 4, 1, 4, 8, 3, 6, 0, 
    35, 7, 0, 0, 0, 0, 0, 3, 7, 3, 12, 5, 3, 9, 7, 
    33, 20, 0, 0, 0, 0, 1, 6, 6, 10, 13, 9, 9, 10, 4, 
    32, 20, 12, 0, 0, 0, 8, 0, 0, 0, 6, 7, 7, 1, 0, 
    35, 30, 30, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    19, 29, 25, 25, 9, 3, 1, 16, 12, 0, 2, 6, 1, 0, 0, 
    20, 23, 25, 19, 45, 37, 34, 23, 25, 23, 33, 46, 47, 32, 32, 
    53, 31, 28, 29, 42, 41, 46, 46, 52, 59, 65, 69, 74, 76, 75, 
    89, 51, 28, 30, 42, 62, 64, 61, 64, 69, 76, 78, 77, 79, 84, 
    91, 78, 50, 31, 55, 66, 68, 64, 67, 72, 82, 80, 84, 89, 89, 
    91, 83, 76, 46, 62, 62, 63, 63, 70, 75, 79, 77, 83, 95, 87, 
    
    -- channel=10
    31, 33, 31, 28, 29, 28, 33, 35, 31, 30, 27, 31, 23, 19, 21, 
    28, 31, 34, 30, 33, 19, 8, 31, 31, 15, 0, 0, 17, 30, 21, 
    26, 54, 32, 31, 36, 69, 11, 6, 0, 16, 0, 0, 0, 12, 31, 
    0, 18, 26, 36, 23, 21, 0, 0, 0, 42, 0, 2, 0, 0, 43, 
    0, 0, 0, 46, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 6, 
    0, 12, 0, 26, 84, 8, 0, 0, 0, 57, 0, 0, 5, 0, 0, 
    0, 0, 16, 8, 57, 22, 18, 0, 0, 62, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 57, 0, 14, 0, 51, 0, 0, 7, 5, 0, 
    0, 4, 0, 19, 0, 28, 0, 0, 4, 0, 35, 0, 8, 12, 16, 
    8, 3, 0, 16, 0, 0, 7, 0, 0, 23, 0, 0, 1, 26, 21, 
    44, 0, 0, 41, 0, 0, 15, 13, 0, 0, 0, 0, 0, 5, 0, 
    44, 26, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 23, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 47, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 19, 14, 7, 0, 0, 
    10, 0, 0, 0, 0, 0, 1, 15, 13, 2, 10, 9, 15, 13, 0, 
    30, 0, 0, 0, 0, 0, 8, 16, 11, 4, 9, 15, 10, 14, 0, 
    40, 12, 0, 0, 1, 11, 9, 9, 11, 3, 16, 20, 10, 14, 14, 
    44, 9, 0, 0, 0, 7, 7, 13, 15, 0, 21, 20, 12, 16, 13, 
    42, 18, 15, 0, 0, 5, 12, 7, 16, 0, 16, 18, 14, 8, 0, 
    37, 25, 40, 8, 13, 0, 10, 11, 8, 0, 13, 11, 8, 0, 0, 
    26, 25, 34, 9, 28, 10, 7, 12, 17, 11, 8, 15, 5, 0, 0, 
    18, 23, 28, 19, 34, 36, 23, 25, 33, 18, 34, 38, 32, 23, 30, 
    38, 31, 31, 2, 36, 56, 41, 44, 53, 49, 53, 53, 59, 57, 63, 
    67, 40, 33, 18, 59, 53, 51, 50, 52, 56, 59, 62, 59, 62, 66, 
    74, 61, 41, 31, 56, 51, 54, 53, 54, 58, 61, 65, 65, 74, 65, 
    71, 66, 56, 39, 52, 55, 55, 53, 53, 56, 62, 60, 63, 68, 70, 
    
    -- channel=12
    19, 15, 17, 17, 18, 11, 21, 27, 20, 10, 6, 8, 8, 13, 14, 
    19, 18, 18, 19, 16, 0, 7, 10, 1, 0, 0, 0, 0, 9, 11, 
    2, 24, 22, 22, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 17, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    11, 4, 0, 0, 13, 0, 0, 0, 0, 1, 0, 3, 3, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 6, 0, 0, 
    4, 6, 0, 1, 0, 7, 0, 0, 5, 0, 0, 9, 5, 0, 0, 
    7, 7, 0, 3, 1, 2, 4, 0, 0, 5, 6, 7, 0, 0, 0, 
    8, 2, 0, 9, 0, 0, 1, 15, 12, 3, 10, 9, 14, 17, 13, 
    45, 27, 8, 0, 4, 41, 31, 32, 33, 29, 32, 33, 35, 35, 36, 
    39, 40, 31, 0, 41, 30, 28, 29, 30, 32, 36, 35, 36, 39, 40, 
    46, 38, 42, 20, 30, 32, 28, 29, 32, 35, 38, 43, 42, 44, 42, 
    41, 42, 32, 42, 33, 38, 40, 34, 28, 30, 33, 40, 36, 33, 41, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 0, 0, 
    2, 0, 0, 0, 0, 24, 0, 13, 0, 0, 0, 0, 0, 19, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 
    0, 0, 0, 40, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 15, 24, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 0, 0, 0, 0, 0, 41, 33, 0, 0, 0, 0, 0, 0, 0, 
    0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 19, 20, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 2, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 
    1, 13, 0, 0, 18, 0, 0, 0, 0, 10, 0, 0, 1, 0, 0, 
    0, 24, 0, 0, 28, 0, 15, 0, 0, 35, 0, 0, 0, 0, 0, 
    0, 23, 0, 0, 4, 18, 11, 3, 0, 37, 0, 0, 0, 7, 0, 
    8, 26, 0, 0, 0, 24, 0, 1, 0, 13, 7, 0, 3, 0, 0, 
    22, 33, 0, 21, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    30, 26, 8, 29, 0, 0, 10, 18, 0, 0, 0, 0, 3, 0, 0, 
    50, 21, 5, 51, 38, 5, 36, 28, 9, 3, 11, 26, 26, 19, 12, 
    38, 47, 15, 53, 12, 17, 24, 23, 27, 30, 36, 39, 45, 41, 40, 
    42, 33, 40, 36, 6, 36, 33, 33, 32, 36, 43, 45, 43, 46, 55, 
    46, 43, 36, 45, 28, 36, 35, 32, 38, 41, 45, 45, 47, 57, 47, 
    45, 50, 42, 24, 24, 34, 36, 37, 42, 45, 38, 41, 57, 53, 38, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 16, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 8, 1, 0, 0, 10, 0, 0, 0, 0, 4, 0, 0, 
    5, 2, 0, 30, 28, 25, 11, 2, 0, 0, 12, 21, 14, 0, 0, 
    19, 8, 16, 19, 0, 0, 0, 3, 14, 19, 27, 27, 34, 34, 33, 
    38, 17, 11, 0, 0, 27, 27, 25, 26, 31, 36, 40, 36, 33, 46, 
    41, 35, 18, 0, 11, 30, 29, 29, 29, 33, 32, 35, 35, 46, 31, 
    40, 41, 24, 16, 14, 22, 25, 30, 35, 37, 35, 36, 50, 49, 41, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 3, 0, 0, 
    7, 11, 0, 0, 0, 11, 18, 10, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 12, 39, 11, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 14, 4, 0, 5, 1, 0, 0, 0, 
    0, 0, 1, 0, 0, 25, 6, 0, 0, 0, 17, 29, 10, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 20, 18, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 0, 0, 32, 61, 28, 27, 12, 0, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 30, 10, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 
    0, 0, 0, 23, 9, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 2, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 7, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 14, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 7, 9, 13, 13, 13, 11, 10, 9, 
    13, 0, 0, 0, 0, 10, 10, 14, 17, 18, 16, 11, 3, 4, 4, 
    11, 16, 0, 0, 0, 10, 11, 15, 13, 12, 13, 9, 13, 11, 0, 
    8, 17, 11, 0, 17, 16, 7, 8, 8, 8, 11, 16, 5, 0, 12, 
    
    -- channel=19
    5, 7, 7, 5, 7, 7, 6, 8, 11, 12, 14, 12, 10, 9, 10, 
    7, 7, 8, 5, 6, 0, 10, 14, 24, 13, 6, 11, 14, 7, 6, 
    17, 6, 6, 7, 7, 10, 21, 22, 12, 0, 0, 0, 5, 7, 3, 
    6, 0, 0, 9, 14, 11, 0, 5, 2, 0, 2, 7, 10, 8, 3, 
    0, 0, 1, 7, 0, 1, 4, 8, 8, 5, 0, 5, 1, 3, 14, 
    6, 0, 0, 29, 0, 12, 0, 2, 3, 0, 0, 11, 0, 3, 5, 
    5, 0, 2, 14, 3, 0, 0, 0, 1, 0, 2, 6, 5, 0, 0, 
    3, 0, 2, 0, 1, 0, 3, 6, 0, 0, 2, 7, 2, 0, 0, 
    0, 0, 7, 0, 9, 14, 6, 2, 0, 14, 2, 17, 9, 0, 0, 
    0, 0, 0, 0, 0, 14, 4, 0, 2, 6, 15, 14, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 3, 0, 0, 0, 6, 
    0, 0, 0, 0, 6, 15, 10, 10, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    18, 14, 15, 17, 18, 11, 18, 20, 18, 13, 8, 6, 6, 17, 18, 
    17, 14, 17, 17, 14, 0, 19, 10, 3, 0, 0, 1, 4, 3, 13, 
    13, 0, 16, 17, 20, 10, 0, 1, 0, 0, 0, 0, 3, 11, 0, 
    0, 0, 14, 14, 8, 0, 0, 4, 0, 0, 0, 3, 0, 13, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 5, 0, 0, 3, 0, 1, 23, 
    0, 0, 12, 32, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 
    0, 0, 2, 0, 10, 0, 0, 0, 0, 4, 0, 6, 1, 0, 16, 
    0, 0, 0, 0, 0, 10, 0, 0, 17, 0, 0, 0, 0, 2, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    4, 7, 2, 6, 5, 3, 6, 4, 3, 8, 7, 2, 4, 6, 6, 
    2, 3, 1, 8, 0, 20, 17, 9, 13, 5, 27, 19, 3, 0, 7, 
    22, 0, 4, 6, 2, 23, 32, 13, 0, 6, 48, 32, 41, 0, 4, 
    71, 0, 13, 0, 19, 0, 38, 23, 25, 0, 61, 26, 37, 20, 0, 
    71, 31, 30, 0, 55, 24, 62, 41, 35, 0, 47, 47, 24, 37, 0, 
    47, 56, 38, 0, 30, 29, 79, 45, 61, 0, 73, 50, 17, 31, 18, 
    36, 96, 19, 41, 0, 10, 76, 52, 67, 0, 79, 45, 18, 19, 35, 
    45, 86, 22, 43, 0, 26, 79, 42, 46, 1, 62, 53, 9, 28, 20, 
    72, 63, 72, 29, 23, 23, 42, 41, 8, 43, 26, 44, 4, 11, 8, 
    68, 59, 102, 14, 60, 0, 1, 73, 25, 29, 45, 8, 0, 4, 15, 
    46, 55, 100, 0, 114, 48, 25, 71, 67, 35, 16, 16, 22, 30, 36, 
    32, 43, 61, 33, 143, 68, 43, 43, 46, 36, 41, 41, 46, 48, 52, 
    62, 20, 0, 111, 94, 43, 45, 41, 42, 39, 41, 45, 53, 48, 48, 
    68, 45, 0, 144, 54, 40, 51, 42, 38, 42, 49, 54, 54, 42, 78, 
    73, 51, 44, 68, 46, 35, 42, 42, 40, 51, 57, 42, 34, 81, 79, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 3, 
    25, 9, 0, 0, 5, 0, 0, 0, 0, 3, 5, 2, 3, 0, 0, 
    24, 6, 0, 0, 0, 0, 0, 0, 0, 7, 3, 3, 5, 0, 2, 
    21, 5, 5, 0, 0, 0, 10, 4, 0, 3, 0, 5, 6, 7, 0, 
    18, 18, 18, 0, 0, 8, 0, 0, 0, 0, 0, 4, 10, 0, 0, 
    12, 20, 6, 13, 6, 8, 0, 0, 20, 0, 0, 0, 0, 0, 0, 
    10, 16, 11, 16, 0, 6, 13, 13, 8, 4, 13, 13, 22, 11, 5, 
    53, 24, 10, 9, 23, 38, 41, 40, 34, 33, 37, 42, 45, 47, 47, 
    55, 53, 27, 15, 34, 38, 39, 39, 39, 41, 44, 48, 48, 47, 50, 
    56, 49, 59, 15, 29, 42, 39, 41, 41, 45, 51, 53, 50, 56, 62, 
    57, 53, 50, 40, 40, 45, 42, 39, 39, 44, 49, 49, 47, 55, 50, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 15, 0, 0, 0, 4, 0, 0, 
    19, 13, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 4, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 14, 47, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 11, 15, 0, 6, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 23, 17, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 21, 0, 0, 0, 0, 0, 0, 0, 
    44, 13, 0, 0, 33, 25, 18, 16, 2, 0, 0, 0, 0, 0, 0, 
    0, 34, 0, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 38, 28, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 20, 
    0, 0, 1, 22, 3, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 3, 0, 0, 11, 20, 14, 9, 2, 0, 
    0, 5, 0, 0, 0, 17, 0, 6, 12, 41, 40, 32, 21, 13, 3, 
    15, 21, 1, 0, 0, 11, 25, 24, 22, 48, 25, 26, 14, 7, 16, 
    41, 57, 9, 27, 54, 51, 35, 19, 15, 33, 42, 23, 24, 13, 13, 
    51, 59, 10, 0, 47, 40, 34, 30, 14, 57, 45, 20, 32, 24, 15, 
    51, 51, 16, 0, 38, 40, 58, 34, 24, 66, 38, 22, 25, 31, 25, 
    54, 58, 39, 15, 36, 73, 43, 32, 20, 49, 31, 21, 31, 33, 12, 
    63, 74, 31, 41, 21, 34, 22, 24, 37, 21, 26, 10, 17, 17, 10, 
    60, 71, 36, 57, 41, 27, 39, 48, 38, 23, 13, 12, 30, 20, 6, 
    68, 66, 40, 83, 61, 60, 73, 64, 39, 23, 31, 40, 50, 47, 37, 
    85, 71, 64, 99, 64, 35, 46, 45, 43, 49, 54, 58, 61, 64, 61, 
    66, 73, 72, 81, 39, 53, 54, 51, 51, 54, 62, 67, 68, 68, 75, 
    67, 61, 88, 59, 45, 59, 54, 53, 55, 60, 65, 66, 63, 75, 73, 
    67, 64, 58, 58, 47, 53, 57, 55, 60, 63, 62, 62, 77, 82, 60, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 3, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 4, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 9, 1, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 0, 4, 5, 0, 
    3, 14, 0, 0, 24, 0, 0, 0, 4, 0, 0, 4, 7, 5, 0, 
    1, 13, 0, 0, 0, 0, 6, 0, 10, 2, 8, 4, 5, 9, 0, 
    0, 22, 0, 0, 0, 0, 0, 2, 9, 0, 6, 8, 8, 0, 0, 
    8, 18, 1, 13, 0, 6, 8, 3, 5, 0, 11, 4, 7, 0, 0, 
    15, 13, 18, 16, 10, 0, 0, 10, 0, 0, 6, 14, 7, 0, 0, 
    33, 8, 20, 9, 4, 0, 0, 17, 15, 11, 26, 23, 23, 28, 28, 
    50, 31, 17, 0, 25, 51, 47, 47, 49, 43, 47, 48, 54, 50, 53, 
    55, 41, 19, 11, 44, 44, 44, 43, 46, 48, 53, 51, 50, 54, 58, 
    65, 54, 26, 48, 42, 44, 45, 44, 46, 49, 53, 60, 60, 61, 59, 
    58, 60, 47, 64, 46, 50, 50, 45, 43, 48, 52, 54, 54, 57, 62, 
    
    -- channel=29
    3, 5, 6, 7, 6, 6, 8, 8, 8, 5, 4, 4, 6, 7, 5, 
    7, 9, 8, 7, 5, 8, 14, 12, 0, 0, 0, 0, 0, 0, 6, 
    8, 0, 6, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 6, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 5, 0, 0, 1, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 3, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 2, 5, 0, 
    3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 1, 16, 0, 0, 1, 12, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 2, 21, 20, 14, 1, 0, 0, 8, 22, 25, 16, 8, 8, 
    11, 5, 7, 10, 0, 5, 18, 17, 20, 25, 28, 31, 37, 33, 32, 
    36, 14, 8, 0, 1, 28, 28, 27, 28, 32, 36, 37, 31, 32, 43, 
    38, 35, 10, 0, 18, 30, 31, 29, 29, 32, 34, 33, 37, 42, 28, 
    38, 38, 30, 16, 23, 23, 21, 27, 33, 37, 34, 36, 45, 43, 36, 
    
    -- channel=31
    8, 7, 7, 9, 7, 3, 9, 5, 3, 3, 2, 0, 4, 7, 5, 
    3, 2, 4, 10, 4, 17, 24, 5, 4, 0, 18, 8, 0, 0, 5, 
    10, 0, 6, 8, 3, 0, 34, 2, 0, 0, 48, 37, 30, 0, 0, 
    53, 0, 10, 0, 14, 0, 30, 31, 21, 0, 64, 21, 32, 13, 0, 
    84, 13, 42, 0, 57, 53, 66, 48, 23, 0, 44, 53, 16, 28, 0, 
    85, 47, 61, 20, 8, 63, 81, 45, 45, 0, 89, 61, 8, 29, 20, 
    90, 69, 23, 36, 0, 26, 62, 68, 54, 0, 88, 48, 12, 14, 37, 
    91, 77, 41, 29, 0, 17, 103, 40, 47, 0, 69, 49, 3, 24, 29, 
    103, 64, 102, 16, 45, 17, 37, 29, 7, 26, 6, 46, 0, 9, 11, 
    80, 68, 108, 0, 61, 28, 14, 56, 37, 32, 37, 0, 0, 0, 12, 
    21, 66, 98, 0, 138, 60, 31, 72, 76, 28, 4, 11, 12, 9, 21, 
    0, 48, 79, 24, 131, 71, 24, 27, 36, 25, 28, 29, 36, 37, 43, 
    52, 2, 27, 92, 114, 37, 36, 31, 30, 28, 30, 36, 42, 40, 44, 
    59, 33, 0, 114, 57, 32, 44, 31, 29, 34, 38, 39, 44, 35, 59, 
    69, 39, 33, 25, 32, 21, 31, 38, 34, 43, 46, 34, 30, 69, 68, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 14, 0, 0, 0, 0, 8, 0, 0, 
    44, 0, 0, 0, 3, 0, 3, 0, 0, 0, 18, 0, 17, 2, 0, 
    38, 0, 5, 0, 0, 0, 13, 12, 5, 0, 2, 18, 0, 15, 0, 
    11, 0, 12, 0, 0, 0, 18, 13, 28, 0, 9, 26, 0, 6, 4, 
    13, 0, 0, 32, 0, 0, 0, 10, 28, 0, 30, 17, 0, 0, 0, 
    3, 10, 0, 16, 0, 0, 15, 0, 15, 0, 18, 23, 0, 0, 0, 
    6, 0, 31, 0, 0, 0, 15, 3, 0, 16, 0, 23, 0, 0, 0, 
    0, 0, 44, 0, 4, 0, 0, 8, 0, 0, 19, 2, 0, 0, 0, 
    0, 0, 42, 0, 36, 0, 0, 0, 11, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 40, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 11, 14, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 24, 16, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    4, 0, 10, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 13, 5, 0, 6, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 33, 6, 0, 0, 0, 0, 31, 6, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 18, 28, 9, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 15, 11, 0, 0, 0, 0, 0, 1, 
    14, 16, 0, 0, 29, 56, 22, 22, 11, 0, 0, 0, 0, 0, 0, 
    0, 8, 9, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    3, 0, 0, 32, 14, 0, 0, 0, 0, 0, 0, 4, 6, 0, 9, 
    0, 0, 0, 30, 10, 8, 12, 2, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 11, 0, 0, 
    7, 7, 0, 0, 0, 35, 17, 28, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 10, 4, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 12, 
    23, 0, 0, 26, 25, 16, 0, 0, 0, 0, 2, 14, 0, 0, 0, 
    9, 0, 16, 0, 2, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 19, 0, 0, 3, 11, 0, 0, 0, 
    0, 0, 8, 0, 0, 45, 14, 0, 0, 18, 21, 29, 10, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 6, 11, 19, 7, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 6, 
    34, 0, 0, 0, 59, 59, 42, 39, 13, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 15, 5, 0, 0, 0, 0, 0, 0, 5, 2, 0, 18, 
    0, 0, 9, 39, 16, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    17, 19, 19, 18, 18, 18, 22, 24, 18, 11, 8, 10, 12, 16, 14, 
    18, 23, 21, 20, 18, 9, 16, 15, 8, 0, 0, 0, 0, 8, 12, 
    5, 10, 21, 22, 21, 9, 2, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 18, 20, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    4, 3, 2, 1, 2, 31, 17, 0, 0, 0, 21, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 9, 8, 15, 0, 0, 
    24, 25, 5, 0, 0, 0, 23, 16, 5, 0, 1, 0, 0, 3, 0, 
    34, 48, 18, 4, 62, 59, 6, 8, 0, 3, 21, 25, 6, 16, 0, 
    8, 0, 17, 0, 0, 0, 18, 18, 20, 14, 4, 0, 0, 9, 29, 
    26, 0, 0, 0, 0, 9, 0, 15, 4, 0, 0, 10, 4, 10, 20, 
    25, 3, 34, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 21, 0, 21, 0, 0, 5, 6, 4, 0, 0, 0, 0, 19, 
    0, 0, 10, 4, 3, 2, 3, 34, 15, 0, 0, 0, 16, 15, 0, 
    0, 0, 0, 24, 95, 71, 7, 0, 0, 7, 19, 34, 11, 0, 0, 
    0, 0, 17, 22, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 12, 0, 0, 14, 
    0, 2, 0, 0, 0, 1, 10, 2, 0, 1, 0, 0, 0, 5, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 12, 15, 6, 1, 23, 21, 7, 
    
    -- channel=38
    34, 31, 33, 33, 34, 30, 35, 36, 34, 31, 29, 29, 28, 32, 31, 
    36, 31, 32, 33, 31, 24, 32, 32, 23, 18, 16, 23, 28, 30, 31, 
    32, 30, 35, 34, 36, 20, 27, 20, 21, 8, 10, 10, 17, 31, 27, 
    10, 33, 35, 33, 32, 18, 13, 17, 19, 14, 12, 19, 16, 29, 27, 
    0, 14, 32, 17, 0, 7, 7, 16, 19, 19, 7, 16, 15, 16, 34, 
    11, 11, 31, 38, 7, 9, 5, 9, 15, 16, 10, 15, 14, 12, 20, 
    10, 8, 32, 22, 11, 16, 0, 10, 8, 9, 8, 16, 18, 14, 20, 
    12, 0, 24, 16, 14, 3, 6, 15, 14, 15, 12, 16, 15, 18, 24, 
    2, 0, 19, 12, 28, 12, 16, 16, 15, 18, 21, 17, 21, 22, 31, 
    1, 2, 6, 4, 12, 21, 9, 0, 25, 18, 14, 15, 19, 28, 30, 
    0, 4, 3, 1, 0, 7, 5, 0, 6, 9, 11, 9, 10, 11, 12, 
    4, 0, 0, 0, 1, 11, 8, 7, 8, 5, 5, 2, 1, 4, 3, 
    6, 12, 7, 1, 0, 3, 3, 5, 5, 5, 1, 1, 1, 0, 0, 
    0, 5, 14, 0, 5, 2, 4, 5, 3, 2, 2, 1, 0, 1, 3, 
    0, 1, 11, 0, 9, 9, 5, 3, 1, 0, 2, 2, 0, 0, 0, 
    
    -- channel=39
    44, 44, 44, 45, 46, 42, 47, 50, 45, 39, 35, 36, 36, 38, 37, 
    44, 45, 46, 47, 45, 39, 43, 43, 32, 19, 10, 17, 27, 34, 38, 
    37, 42, 48, 47, 48, 47, 26, 20, 8, 7, 0, 0, 4, 20, 33, 
    8, 28, 47, 47, 43, 29, 15, 2, 1, 10, 6, 5, 0, 1, 28, 
    0, 16, 40, 36, 21, 15, 10, 2, 2, 6, 9, 2, 3, 0, 16, 
    0, 13, 35, 26, 18, 9, 8, 5, 0, 9, 9, 1, 5, 0, 0, 
    0, 9, 31, 31, 21, 14, 16, 7, 1, 13, 4, 0, 2, 0, 2, 
    0, 3, 11, 28, 15, 17, 11, 10, 3, 18, 4, 2, 1, 7, 16, 
    0, 3, 0, 10, 12, 13, 9, 6, 9, 25, 12, 4, 3, 15, 32, 
    2, 2, 0, 4, 3, 7, 9, 4, 7, 10, 4, 0, 5, 30, 37, 
    7, 5, 0, 3, 0, 0, 1, 3, 0, 0, 0, 0, 0, 11, 9, 
    0, 0, 0, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 4, 15, 27, 16, 5, 0, 0, 
    9, 0, 0, 0, 0, 3, 21, 13, 10, 18, 37, 30, 28, 2, 1, 
    44, 0, 0, 0, 6, 5, 29, 22, 24, 5, 42, 20, 31, 18, 0, 
    57, 28, 9, 0, 44, 17, 40, 31, 25, 0, 37, 32, 23, 27, 0, 
    46, 50, 17, 0, 33, 27, 54, 32, 38, 0, 50, 38, 21, 28, 18, 
    43, 63, 15, 13, 4, 25, 53, 42, 43, 7, 56, 36, 22, 26, 27, 
    48, 66, 23, 27, 0, 30, 52, 31, 37, 7, 47, 38, 18, 23, 13, 
    64, 57, 56, 34, 21, 19, 34, 34, 20, 21, 26, 30, 12, 12, 0, 
    62, 54, 72, 26, 45, 9, 18, 54, 22, 25, 30, 15, 10, 0, 4, 
    54, 51, 69, 21, 87, 44, 34, 58, 55, 33, 32, 34, 39, 45, 50, 
    46, 55, 56, 39, 93, 69, 49, 50, 56, 49, 52, 54, 59, 58, 62, 
    69, 38, 35, 78, 81, 53, 51, 50, 52, 53, 57, 60, 61, 62, 68, 
    76, 58, 20, 103, 62, 51, 57, 50, 50, 55, 61, 65, 66, 66, 74, 
    75, 63, 54, 63, 53, 50, 54, 53, 52, 60, 62, 57, 58, 80, 76, 
    
    -- channel=41
    36, 35, 35, 37, 37, 34, 37, 42, 40, 33, 29, 28, 30, 34, 35, 
    36, 38, 35, 38, 35, 16, 41, 34, 27, 11, 6, 13, 18, 25, 33, 
    29, 25, 39, 40, 37, 23, 31, 26, 13, 0, 1, 3, 5, 15, 19, 
    25, 0, 36, 37, 34, 22, 8, 9, 1, 0, 11, 4, 10, 11, 4, 
    14, 0, 39, 17, 0, 3, 12, 12, 6, 0, 4, 14, 1, 9, 9, 
    15, 0, 42, 23, 0, 11, 4, 13, 11, 0, 12, 21, 0, 5, 8, 
    18, 0, 29, 40, 0, 0, 0, 10, 14, 0, 16, 13, 0, 0, 10, 
    7, 0, 14, 24, 0, 0, 19, 3, 17, 0, 6, 16, 0, 1, 21, 
    0, 0, 18, 0, 18, 5, 14, 1, 0, 13, 6, 22, 2, 5, 18, 
    0, 0, 12, 0, 12, 11, 0, 0, 8, 11, 14, 5, 0, 8, 33, 
    0, 0, 12, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    63, 73, 67, 68, 65, 68, 69, 72, 68, 61, 54, 54, 57, 55, 53, 
    62, 71, 69, 71, 68, 90, 60, 68, 55, 44, 32, 27, 35, 47, 53, 
    61, 55, 68, 72, 69, 98, 63, 34, 18, 46, 50, 36, 24, 17, 52, 
    36, 21, 63, 71, 72, 51, 58, 25, 25, 46, 62, 41, 32, 8, 32, 
    48, 54, 57, 59, 96, 55, 71, 40, 28, 24, 63, 35, 31, 16, 3, 
    47, 86, 64, 65, 127, 83, 92, 47, 30, 46, 77, 42, 34, 26, 5, 
    44, 91, 56, 69, 70, 81, 106, 61, 45, 65, 72, 36, 26, 35, 27, 
    64, 91, 23, 56, 40, 103, 80, 64, 47, 70, 75, 42, 31, 44, 41, 
    87, 91, 45, 65, 43, 61, 58, 53, 35, 51, 66, 37, 23, 43, 53, 
    106, 91, 69, 53, 56, 24, 47, 74, 32, 58, 31, 5, 16, 51, 60, 
    98, 88, 72, 75, 83, 35, 63, 88, 44, 13, 0, 0, 9, 27, 24, 
    49, 82, 67, 115, 123, 49, 35, 33, 19, 9, 8, 11, 13, 14, 14, 
    1, 35, 64, 137, 56, 14, 11, 9, 7, 4, 6, 10, 16, 16, 17, 
    7, 3, 38, 119, 25, 13, 11, 8, 9, 10, 11, 16, 10, 13, 24, 
    10, 9, 10, 43, 8, 12, 16, 12, 13, 16, 11, 6, 16, 28, 3, 
    
    -- channel=43
    5, 4, 7, 2, 3, 5, 4, 4, 3, 2, 2, 7, 4, 0, 0, 
    4, 4, 8, 1, 9, 0, 0, 0, 4, 9, 0, 0, 5, 9, 0, 
    0, 25, 4, 2, 10, 10, 0, 0, 7, 23, 0, 0, 0, 9, 9, 
    0, 31, 0, 8, 0, 14, 0, 0, 0, 39, 0, 0, 0, 0, 34, 
    0, 0, 0, 47, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 17, 
    0, 0, 0, 22, 33, 1, 0, 0, 0, 84, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 39, 23, 0, 0, 0, 66, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 30, 27, 0, 0, 0, 40, 0, 0, 10, 0, 0, 
    0, 0, 0, 5, 0, 11, 0, 0, 6, 0, 6, 0, 13, 6, 5, 
    0, 0, 0, 25, 0, 5, 17, 0, 0, 0, 0, 0, 13, 11, 0, 
    17, 0, 0, 62, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 9, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 1, 5, 0, 0, 0, 0, 9, 6, 0, 0, 0, 
    21, 6, 0, 0, 0, 0, 1, 0, 0, 0, 12, 0, 0, 0, 0, 
    20, 4, 0, 0, 0, 0, 15, 4, 0, 0, 4, 3, 0, 0, 0, 
    21, 13, 22, 0, 0, 3, 0, 0, 0, 0, 1, 6, 0, 0, 0, 
    12, 13, 18, 0, 11, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 
    4, 12, 17, 0, 0, 2, 8, 23, 17, 0, 1, 4, 10, 15, 21, 
    35, 23, 11, 0, 51, 48, 32, 33, 31, 27, 28, 30, 32, 31, 34, 
    39, 32, 10, 23, 50, 26, 27, 25, 25, 26, 27, 30, 34, 36, 31, 
    44, 35, 29, 38, 30, 25, 26, 27, 27, 30, 35, 40, 39, 37, 52, 
    44, 38, 35, 33, 31, 31, 32, 27, 24, 26, 34, 31, 24, 38, 42, 
    
    -- channel=45
    0, 5, 1, 5, 4, 2, 2, 5, 3, 0, 3, 0, 6, 6, 7, 
    4, 2, 0, 6, 0, 9, 12, 3, 9, 1, 13, 2, 0, 0, 7, 
    5, 0, 3, 7, 0, 0, 29, 7, 0, 0, 7, 14, 19, 0, 0, 
    55, 0, 3, 0, 11, 0, 11, 9, 6, 0, 36, 0, 24, 11, 0, 
    61, 0, 21, 0, 26, 0, 28, 24, 11, 0, 10, 29, 2, 28, 0, 
    20, 0, 36, 0, 0, 7, 41, 21, 39, 0, 29, 39, 0, 16, 17, 
    26, 17, 9, 35, 0, 0, 8, 31, 41, 0, 46, 25, 0, 0, 15, 
    17, 31, 7, 30, 0, 0, 43, 2, 32, 0, 31, 27, 0, 0, 18, 
    25, 0, 48, 0, 0, 0, 18, 4, 0, 6, 0, 34, 0, 0, 0, 
    10, 0, 67, 0, 20, 0, 0, 22, 0, 1, 34, 3, 0, 0, 7, 
    0, 0, 58, 0, 82, 6, 0, 9, 47, 23, 0, 0, 0, 0, 5, 
    0, 0, 27, 0, 40, 34, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 56, 21, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 
    
    -- channel=46
    0, 6, 8, 10, 8, 7, 6, 6, 9, 0, 0, 0, 4, 6, 8, 
    9, 10, 9, 9, 11, 49, 13, 2, 0, 2, 20, 0, 0, 0, 7, 
    0, 0, 5, 8, 5, 0, 0, 0, 0, 17, 15, 17, 17, 0, 0, 
    30, 8, 5, 9, 13, 5, 34, 17, 9, 0, 14, 0, 0, 0, 0, 
    40, 42, 12, 14, 88, 49, 15, 13, 0, 0, 25, 23, 13, 22, 0, 
    0, 6, 10, 0, 0, 0, 37, 21, 27, 17, 10, 0, 0, 16, 21, 
    7, 13, 0, 17, 0, 18, 12, 20, 19, 5, 4, 9, 1, 15, 16, 
    13, 26, 9, 19, 11, 12, 0, 0, 0, 0, 6, 0, 0, 0, 2, 
    20, 9, 9, 9, 8, 0, 0, 17, 6, 0, 0, 0, 0, 5, 21, 
    2, 5, 24, 5, 8, 0, 5, 51, 0, 0, 0, 0, 12, 15, 2, 
    0, 5, 8, 31, 108, 61, 22, 0, 8, 8, 13, 32, 8, 0, 0, 
    0, 0, 23, 38, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 
    3, 0, 0, 4, 0, 3, 2, 0, 1, 6, 8, 11, 2, 0, 15, 
    1, 0, 0, 0, 0, 2, 9, 1, 2, 4, 0, 0, 0, 8, 0, 
    6, 2, 0, 0, 0, 0, 0, 3, 15, 15, 4, 0, 25, 25, 8, 
    
    -- channel=47
    0, 5, 2, 3, 0, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 3, 2, 26, 4, 1, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 2, 3, 0, 10, 5, 0, 0, 9, 18, 9, 0, 0, 0, 
    5, 0, 3, 2, 6, 0, 14, 0, 0, 4, 24, 2, 0, 0, 0, 
    28, 28, 9, 2, 52, 29, 30, 8, 0, 0, 26, 8, 0, 0, 0, 
    28, 47, 19, 1, 45, 37, 46, 13, 1, 10, 38, 10, 0, 0, 0, 
    31, 48, 10, 1, 9, 34, 48, 29, 11, 20, 35, 8, 0, 5, 3, 
    44, 52, 10, 9, 0, 42, 37, 17, 10, 17, 32, 8, 0, 7, 5, 
    57, 53, 27, 27, 8, 12, 16, 12, 8, 6, 8, 0, 0, 4, 3, 
    57, 52, 39, 22, 22, 0, 15, 37, 8, 7, 0, 0, 0, 3, 2, 
    47, 50, 38, 41, 73, 24, 32, 44, 22, 0, 0, 0, 1, 3, 1, 
    15, 45, 43, 66, 64, 20, 8, 6, 5, 0, 2, 4, 10, 11, 10, 
    9, 11, 39, 74, 26, 7, 5, 3, 1, 2, 6, 10, 13, 11, 19, 
    13, 6, 14, 61, 10, 7, 8, 3, 4, 7, 8, 10, 9, 14, 17, 
    15, 10, 8, 9, 0, 0, 4, 7, 9, 13, 9, 6, 18, 28, 11, 
    
    -- channel=48
    45, 44, 42, 43, 42, 42, 45, 46, 41, 41, 40, 41, 37, 35, 33, 
    41, 41, 43, 44, 43, 38, 39, 41, 41, 31, 19, 24, 35, 40, 35, 
    40, 54, 46, 44, 47, 74, 46, 33, 18, 34, 35, 25, 15, 30, 38, 
    11, 25, 45, 45, 40, 38, 28, 18, 22, 50, 40, 35, 25, 10, 36, 
    26, 34, 43, 44, 35, 30, 44, 24, 23, 34, 40, 20, 21, 6, 19, 
    51, 66, 48, 51, 98, 67, 48, 28, 10, 41, 56, 35, 30, 17, 2, 
    45, 59, 57, 34, 53, 57, 70, 42, 24, 57, 54, 27, 26, 27, 20, 
    54, 56, 29, 36, 35, 72, 63, 57, 36, 58, 54, 33, 30, 41, 34, 
    62, 71, 38, 47, 38, 65, 47, 32, 33, 44, 56, 35, 29, 32, 32, 
    79, 73, 42, 47, 41, 29, 42, 36, 35, 48, 29, 11, 14, 36, 43, 
    80, 71, 51, 58, 27, 15, 49, 70, 33, 15, 5, 1, 16, 42, 37, 
    76, 81, 53, 84, 102, 66, 53, 51, 32, 24, 24, 27, 27, 29, 28, 
    24, 64, 74, 99, 61, 24, 22, 23, 21, 20, 21, 23, 30, 32, 29, 
    26, 24, 73, 90, 34, 26, 21, 21, 22, 23, 28, 35, 29, 29, 46, 
    27, 23, 33, 59, 29, 33, 33, 24, 21, 24, 25, 25, 26, 31, 19, 
    
    -- channel=49
    35, 36, 40, 42, 41, 40, 41, 40, 40, 31, 21, 24, 34, 35, 32, 
    41, 43, 42, 42, 45, 80, 56, 35, 8, 30, 47, 30, 14, 23, 35, 
    15, 13, 40, 41, 37, 15, 16, 12, 24, 46, 46, 44, 33, 8, 27, 
    54, 43, 45, 44, 43, 43, 62, 36, 25, 22, 44, 18, 16, 7, 13, 
    78, 86, 56, 63, 134, 93, 57, 35, 10, 26, 70, 48, 34, 32, 2, 
    47, 60, 58, 0, 1, 38, 74, 57, 40, 50, 58, 27, 28, 36, 35, 
    63, 52, 28, 38, 19, 59, 66, 59, 44, 44, 51, 38, 26, 39, 40, 
    66, 80, 58, 62, 41, 62, 42, 17, 30, 31, 38, 29, 21, 23, 30, 
    75, 72, 44, 46, 41, 1, 30, 39, 46, 35, 6, 0, 0, 27, 45, 
    56, 63, 59, 47, 53, 26, 50, 87, 36, 9, 3, 6, 34, 50, 43, 
    51, 67, 52, 89, 144, 102, 59, 46, 43, 33, 37, 46, 36, 31, 28, 
    5, 40, 80, 99, 29, 0, 0, 0, 10, 19, 23, 22, 29, 30, 29, 
    30, 2, 51, 67, 14, 27, 24, 21, 23, 26, 33, 40, 31, 27, 51, 
    29, 23, 9, 33, 22, 30, 33, 24, 22, 28, 22, 18, 22, 37, 8, 
    32, 22, 9, 6, 7, 3, 10, 26, 36, 42, 29, 26, 55, 58, 31, 
    
    -- channel=50
    2, 3, 3, 3, 1, 3, 6, 1, 0, 11, 16, 13, 8, 4, 0, 
    1, 4, 4, 5, 2, 1, 13, 17, 16, 0, 4, 2, 1, 9, 7, 
    19, 15, 3, 0, 0, 0, 0, 0, 0, 2, 9, 4, 12, 8, 8, 
    7, 2, 9, 1, 6, 0, 10, 13, 9, 11, 3, 4, 0, 4, 8, 
    12, 28, 18, 4, 45, 33, 6, 0, 1, 0, 0, 12, 1, 8, 7, 
    4, 12, 17, 0, 0, 2, 2, 0, 2, 8, 18, 0, 4, 6, 7, 
    0, 14, 9, 2, 0, 0, 26, 9, 7, 10, 1, 0, 0, 0, 10, 
    6, 1, 15, 14, 8, 40, 16, 0, 0, 0, 0, 0, 1, 12, 0, 
    5, 10, 4, 9, 9, 0, 0, 0, 7, 0, 0, 0, 0, 0, 9, 
    0, 2, 5, 0, 22, 14, 0, 13, 8, 20, 12, 0, 23, 22, 13, 
    5, 6, 0, 0, 31, 42, 55, 38, 36, 4, 0, 21, 20, 17, 14, 
    16, 14, 17, 24, 14, 0, 0, 0, 0, 4, 8, 3, 0, 0, 2, 
    10, 7, 0, 24, 0, 2, 7, 2, 0, 1, 1, 6, 14, 8, 1, 
    2, 7, 16, 14, 0, 1, 1, 3, 5, 5, 1, 1, 0, 3, 19, 
    7, 1, 2, 0, 0, 0, 8, 7, 8, 0, 1, 0, 0, 8, 7, 
    
    -- channel=51
    23, 20, 22, 24, 25, 19, 25, 26, 24, 19, 13, 11, 17, 24, 26, 
    24, 24, 23, 25, 21, 16, 29, 17, 17, 4, 15, 13, 6, 13, 23, 
    12, 7, 25, 26, 25, 2, 18, 12, 7, 0, 1, 0, 19, 5, 12, 
    34, 0, 28, 21, 22, 8, 14, 9, 6, 0, 9, 2, 9, 13, 0, 
    16, 0, 32, 0, 7, 7, 7, 9, 7, 0, 5, 18, 4, 17, 3, 
    0, 0, 27, 15, 0, 0, 10, 11, 24, 0, 4, 8, 0, 8, 15, 
    0, 3, 6, 34, 0, 0, 0, 7, 16, 0, 9, 10, 2, 0, 12, 
    0, 0, 8, 25, 1, 0, 0, 0, 7, 0, 3, 11, 0, 0, 10, 
    0, 0, 12, 0, 11, 0, 5, 6, 0, 25, 0, 5, 0, 6, 20, 
    0, 0, 14, 0, 2, 0, 0, 11, 0, 0, 8, 3, 0, 8, 17, 
    0, 0, 12, 0, 24, 7, 0, 0, 0, 10, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 2, 0, 0, 
    15, 0, 0, 0, 1, 0, 2, 3, 1, 0, 0, 5, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 10, 5, 19, 0, 0, 1, 0, 3, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 16, 0, 4, 2, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 5, 0, 1, 0, 3, 5, 0, 0, 0, 
    1, 0, 6, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 34, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 1, 5, 5, 7, 
    9, 0, 0, 0, 16, 4, 5, 3, 5, 5, 6, 5, 4, 2, 5, 
    14, 0, 0, 18, 6, 3, 9, 5, 3, 5, 6, 4, 8, 3, 7, 
    18, 9, 0, 0, 3, 0, 0, 5, 6, 10, 11, 6, 4, 22, 21, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 38, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 11, 4, 0, 0, 0, 29, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 4, 0, 5, 0, 20, 0, 0, 0, 0, 0, 
    6, 20, 0, 3, 0, 18, 1, 0, 0, 0, 6, 0, 3, 0, 0, 
    18, 22, 0, 26, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 16, 0, 34, 0, 0, 0, 3, 0, 0, 0, 0, 5, 10, 0, 
    53, 30, 0, 34, 20, 32, 40, 39, 20, 15, 17, 24, 26, 28, 23, 
    25, 48, 35, 26, 12, 17, 16, 18, 19, 20, 24, 24, 24, 27, 30, 
    28, 26, 55, 19, 9, 23, 17, 18, 19, 22, 30, 33, 31, 35, 34, 
    24, 29, 34, 42, 21, 29, 23, 16, 18, 24, 24, 29, 32, 29, 17, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 19, 0, 6, 0, 11, 8, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 19, 9, 0, 0, 13, 6, 32, 0, 0, 
    77, 0, 0, 0, 10, 0, 13, 9, 2, 0, 32, 0, 18, 13, 0, 
    56, 0, 24, 0, 11, 4, 35, 23, 16, 0, 13, 37, 0, 30, 0, 
    20, 0, 27, 0, 0, 0, 33, 28, 53, 0, 37, 36, 0, 14, 13, 
    11, 37, 0, 36, 0, 0, 18, 19, 54, 0, 48, 27, 0, 0, 16, 
    4, 32, 16, 27, 0, 0, 45, 0, 18, 0, 20, 34, 0, 0, 1, 
    18, 0, 51, 0, 0, 0, 13, 8, 0, 28, 0, 33, 0, 0, 0, 
    0, 0, 71, 0, 31, 0, 0, 29, 2, 0, 34, 0, 0, 0, 6, 
    0, 0, 68, 0, 72, 23, 0, 8, 42, 28, 0, 0, 0, 0, 6, 
    0, 0, 13, 0, 82, 22, 0, 0, 3, 0, 0, 0, 0, 0, 2, 
    14, 0, 0, 17, 68, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 64, 12, 0, 9, 0, 0, 0, 0, 0, 2, 0, 13, 
    24, 0, 0, 13, 6, 0, 0, 0, 0, 0, 10, 0, 0, 21, 41, 
    
    -- channel=55
    23, 23, 22, 24, 24, 20, 20, 25, 27, 23, 20, 16, 17, 20, 25, 
    22, 20, 20, 24, 21, 19, 19, 21, 17, 12, 10, 9, 12, 16, 22, 
    28, 14, 24, 25, 23, 18, 31, 18, 12, 0, 12, 12, 13, 8, 13, 
    28, 0, 19, 22, 26, 12, 12, 13, 10, 0, 22, 9, 20, 18, 0, 
    21, 0, 21, 0, 2, 0, 13, 20, 16, 0, 7, 17, 10, 18, 1, 
    16, 6, 25, 17, 7, 11, 20, 14, 21, 0, 19, 26, 6, 13, 10, 
    15, 10, 17, 32, 0, 3, 11, 16, 22, 0, 24, 19, 7, 6, 15, 
    11, 9, 6, 15, 0, 0, 27, 14, 25, 0, 24, 23, 4, 7, 20, 
    15, 0, 28, 3, 12, 5, 19, 15, 3, 5, 17, 28, 8, 13, 15, 
    16, 4, 30, 0, 16, 8, 0, 5, 7, 22, 22, 9, 0, 1, 20, 
    0, 2, 26, 0, 17, 1, 0, 8, 21, 9, 4, 0, 0, 1, 10, 
    0, 0, 8, 0, 29, 30, 5, 7, 14, 5, 2, 0, 0, 0, 2, 
    3, 0, 0, 7, 45, 3, 1, 2, 3, 1, 0, 0, 0, 0, 0, 
    7, 0, 0, 34, 19, 0, 4, 1, 0, 0, 0, 2, 3, 0, 3, 
    6, 0, 0, 8, 9, 4, 5, 4, 0, 0, 3, 0, 0, 0, 10, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 8, 6, 0, 
    13, 26, 0, 0, 0, 24, 11, 10, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 48, 9, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 17, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 19, 25, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 22, 7, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 20, 7, 0, 0, 0, 0, 10, 10, 
    46, 20, 0, 0, 31, 52, 28, 26, 13, 0, 0, 0, 0, 0, 0, 
    0, 33, 10, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 34, 32, 5, 0, 0, 0, 0, 0, 0, 5, 0, 0, 15, 
    0, 0, 1, 36, 8, 14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    27, 26, 30, 26, 27, 26, 28, 31, 29, 23, 25, 30, 27, 22, 21, 
    29, 27, 31, 25, 32, 11, 15, 24, 24, 22, 0, 0, 17, 31, 21, 
    8, 50, 30, 28, 30, 8, 13, 9, 17, 9, 0, 0, 0, 18, 26, 
    0, 28, 22, 33, 15, 32, 0, 0, 0, 26, 0, 0, 0, 0, 38, 
    0, 0, 9, 66, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 19, 
    0, 0, 9, 22, 20, 24, 0, 0, 0, 55, 0, 0, 1, 0, 0, 
    4, 0, 27, 0, 15, 26, 0, 0, 0, 25, 0, 0, 0, 1, 0, 
    0, 0, 2, 0, 25, 7, 0, 0, 0, 11, 0, 0, 8, 0, 11, 
    0, 0, 0, 10, 1, 13, 0, 0, 17, 0, 2, 0, 9, 13, 16, 
    0, 0, 0, 4, 0, 20, 28, 0, 0, 11, 0, 7, 12, 20, 21, 
    0, 0, 0, 37, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    29, 33, 29, 29, 29, 29, 31, 34, 30, 23, 23, 26, 26, 27, 27, 
    28, 33, 28, 30, 26, 25, 20, 30, 24, 14, 1, 10, 20, 24, 25, 
    29, 29, 31, 33, 29, 35, 34, 21, 4, 0, 0, 0, 0, 11, 27, 
    6, 3, 27, 29, 30, 13, 3, 0, 0, 0, 12, 5, 11, 9, 14, 
    0, 0, 19, 0, 0, 0, 9, 8, 11, 0, 0, 0, 2, 2, 5, 
    0, 4, 24, 25, 36, 10, 13, 0, 8, 0, 1, 11, 0, 0, 0, 
    0, 8, 25, 34, 8, 3, 2, 3, 6, 0, 7, 5, 1, 0, 0, 
    0, 1, 0, 14, 0, 0, 11, 13, 14, 1, 12, 11, 0, 4, 18, 
    0, 0, 0, 4, 1, 15, 17, 8, 0, 12, 17, 22, 13, 17, 16, 
    4, 0, 7, 0, 0, 0, 0, 0, 0, 15, 14, 3, 0, 8, 19, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 15, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 14, 21, 11, 12, 1, 0, 
    10, 0, 0, 0, 0, 0, 11, 6, 8, 21, 14, 13, 5, 0, 0, 
    21, 29, 0, 0, 27, 19, 22, 6, 8, 2, 21, 10, 7, 3, 0, 
    25, 37, 0, 0, 37, 20, 22, 12, 7, 16, 28, 9, 13, 8, 0, 
    17, 46, 5, 0, 18, 14, 44, 15, 17, 32, 26, 9, 8, 11, 7, 
    26, 40, 16, 5, 9, 46, 25, 21, 7, 20, 19, 11, 13, 14, 0, 
    37, 48, 18, 25, 3, 19, 11, 12, 13, 10, 19, 5, 1, 0, 0, 
    36, 43, 28, 30, 30, 2, 10, 31, 15, 15, 9, 3, 11, 3, 0, 
    48, 40, 31, 30, 37, 32, 45, 50, 29, 11, 13, 20, 32, 35, 29, 
    63, 46, 35, 58, 67, 30, 35, 33, 31, 30, 34, 36, 37, 41, 39, 
    44, 49, 32, 68, 29, 32, 34, 31, 30, 32, 37, 40, 45, 44, 43, 
    45, 41, 51, 60, 27, 34, 32, 33, 34, 37, 41, 45, 41, 45, 56, 
    44, 42, 40, 47, 30, 34, 37, 32, 35, 37, 39, 36, 41, 54, 43, 
    
    -- channel=61
    46, 47, 47, 49, 48, 46, 48, 54, 50, 39, 32, 31, 38, 45, 46, 
    46, 50, 50, 50, 49, 27, 50, 36, 35, 15, 11, 11, 15, 29, 40, 
    24, 28, 48, 52, 49, 36, 32, 28, 16, 0, 12, 13, 13, 13, 24, 
    36, 0, 43, 48, 36, 31, 19, 18, 4, 0, 16, 11, 14, 10, 11, 
    36, 0, 45, 41, 20, 22, 23, 16, 6, 0, 19, 24, 7, 16, 5, 
    22, 0, 45, 23, 0, 27, 18, 28, 15, 0, 17, 24, 7, 13, 14, 
    28, 0, 28, 47, 4, 0, 12, 16, 26, 0, 25, 16, 4, 4, 17, 
    13, 9, 21, 28, 23, 0, 19, 7, 24, 0, 16, 19, 3, 5, 32, 
    8, 0, 15, 0, 10, 15, 23, 4, 10, 15, 10, 19, 3, 19, 31, 
    1, 0, 18, 0, 21, 8, 8, 10, 7, 11, 14, 11, 1, 14, 38, 
    0, 0, 19, 0, 15, 10, 0, 0, 10, 3, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    34, 41, 38, 37, 35, 39, 41, 41, 36, 34, 33, 34, 33, 32, 27, 
    34, 42, 39, 40, 36, 43, 38, 44, 37, 18, 12, 13, 20, 28, 29, 
    37, 33, 39, 40, 37, 44, 34, 12, 4, 10, 14, 6, 8, 9, 30, 
    14, 5, 38, 39, 42, 21, 23, 6, 4, 13, 25, 15, 7, 1, 16, 
    14, 20, 36, 24, 48, 31, 34, 14, 6, 0, 22, 14, 4, 0, 2, 
    15, 34, 41, 36, 55, 43, 41, 14, 6, 8, 35, 15, 6, 2, 0, 
    12, 41, 35, 37, 25, 33, 48, 25, 15, 17, 30, 10, 2, 5, 6, 
    26, 33, 12, 28, 12, 45, 33, 26, 14, 20, 29, 11, 5, 15, 14, 
    33, 34, 18, 27, 19, 24, 21, 15, 9, 21, 26, 12, 1, 13, 28, 
    36, 30, 26, 12, 26, 9, 13, 27, 10, 27, 12, 0, 4, 27, 33, 
    34, 34, 26, 12, 32, 11, 27, 40, 20, 0, 0, 0, 0, 4, 5, 
    4, 28, 23, 41, 55, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 59, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    2, 0, 4, 0, 0, 4, 4, 0, 0, 0, 0, 2, 1, 0, 0, 
    4, 6, 6, 0, 6, 21, 0, 0, 0, 4, 0, 0, 7, 6, 0, 
    0, 14, 5, 0, 8, 11, 0, 0, 3, 42, 0, 0, 0, 12, 14, 
    0, 66, 3, 7, 0, 5, 0, 0, 0, 52, 0, 0, 0, 0, 42, 
    0, 49, 0, 35, 2, 5, 0, 0, 0, 59, 0, 0, 1, 0, 27, 
    0, 13, 0, 15, 36, 0, 0, 0, 0, 129, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 55, 36, 0, 0, 0, 111, 0, 0, 5, 11, 0, 
    0, 0, 0, 0, 35, 59, 0, 0, 0, 74, 0, 0, 15, 8, 0, 
    0, 2, 0, 19, 0, 0, 0, 0, 14, 0, 12, 0, 14, 13, 17, 
    0, 1, 0, 46, 0, 0, 15, 0, 2, 0, 0, 0, 32, 37, 0, 
    45, 0, 0, 108, 0, 0, 46, 0, 0, 0, 3, 15, 15, 6, 0, 
    48, 13, 0, 97, 0, 0, 0, 0, 0, 0, 0, 3, 1, 3, 0, 
    0, 47, 40, 5, 0, 0, 0, 0, 0, 2, 5, 7, 1, 0, 6, 
    0, 2, 90, 0, 0, 2, 0, 0, 1, 3, 1, 0, 0, 20, 0, 
    0, 0, 9, 0, 0, 7, 0, 0, 6, 1, 0, 0, 27, 0, 0, 
    
    
    others => 0);
end ifmap_package;
