library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    146, 118, 122, 126, 125, 121, 126, 124, 125, 123, 123, 123, 123, 125, 125, 127, 129, 126, 124, 125, 123, 120, 122, 122, 128, 124, 124, 123, 126, 126, 126, 165, 
    93, 103, 101, 113, 115, 108, 111, 112, 116, 112, 106, 104, 108, 113, 115, 121, 126, 118, 107, 102, 103, 98, 103, 102, 111, 113, 114, 113, 120, 122, 121, 213, 
    99, 111, 103, 115, 112, 110, 112, 112, 116, 116, 107, 107, 105, 112, 122, 121, 120, 110, 99, 101, 104, 97, 91, 92, 93, 97, 116, 117, 121, 123, 121, 214, 
    103, 119, 107, 117, 110, 106, 111, 113, 111, 106, 89, 120, 104, 101, 109, 105, 92, 107, 102, 104, 93, 96, 88, 84, 89, 81, 97, 110, 116, 118, 120, 218, 
    96, 108, 101, 111, 114, 105, 112, 115, 112, 97, 15, 91, 120, 99, 83, 97, 107, 107, 82, 67, 58, 74, 85, 86, 86, 84, 67, 86, 108, 120, 117, 222, 
    83, 90, 74, 107, 123, 111, 112, 121, 114, 102, 9, 68, 144, 129, 103, 104, 131, 78, 29, 40, 44, 49, 69, 80, 82, 94, 87, 67, 83, 119, 116, 220, 
    78, 120, 68, 82, 118, 116, 112, 119, 118, 110, 87, 90, 109, 129, 125, 85, 90, 57, 5, 31, 60, 57, 65, 62, 80, 105, 111, 70, 52, 103, 121, 222, 
    85, 138, 91, 54, 86, 114, 114, 112, 117, 116, 103, 96, 75, 92, 99, 63, 73, 77, 5, 0, 78, 98, 62, 53, 87, 109, 108, 97, 46, 78, 123, 225, 
    89, 128, 55, 57, 80, 105, 110, 102, 105, 137, 94, 48, 41, 70, 98, 69, 67, 81, 48, 0, 59, 107, 89, 70, 79, 104, 106, 112, 64, 46, 109, 231, 
    61, 108, 11, 31, 106, 103, 101, 41, 43, 88, 82, 0, 40, 72, 105, 86, 67, 87, 77, 21, 38, 70, 105, 84, 67, 83, 94, 122, 103, 38, 71, 231, 
    50, 34, 6, 26, 120, 109, 117, 0, 0, 27, 92, 23, 56, 86, 75, 98, 76, 112, 56, 2, 40, 31, 91, 85, 63, 78, 85, 108, 130, 76, 48, 202, 
    74, 0, 0, 38, 120, 109, 135, 12, 0, 27, 81, 25, 41, 105, 64, 88, 93, 128, 17, 0, 33, 34, 96, 95, 56, 61, 90, 91, 117, 96, 78, 175, 
    87, 4, 0, 29, 93, 112, 134, 126, 0, 10, 78, 23, 2, 97, 91, 64, 72, 143, 0, 0, 38, 70, 98, 92, 63, 47, 78, 85, 98, 89, 111, 177, 
    97, 2, 0, 58, 78, 93, 123, 157, 0, 26, 71, 25, 0, 50, 95, 73, 53, 121, 0, 0, 49, 82, 103, 85, 74, 65, 62, 69, 82, 78, 115, 197, 
    93, 0, 0, 101, 100, 52, 103, 159, 40, 38, 9, 25, 0, 15, 70, 69, 72, 105, 0, 0, 59, 76, 84, 82, 67, 70, 45, 44, 80, 85, 106, 214, 
    72, 0, 0, 87, 125, 29, 77, 139, 68, 23, 0, 0, 56, 40, 43, 52, 82, 109, 0, 0, 51, 82, 78, 92, 60, 51, 48, 44, 92, 107, 104, 218, 
    45, 0, 0, 43, 133, 18, 41, 107, 97, 1, 0, 0, 80, 102, 60, 76, 66, 94, 27, 11, 24, 91, 99, 87, 60, 37, 55, 77, 104, 103, 101, 224, 
    20, 4, 0, 3, 126, 46, 0, 77, 132, 25, 0, 40, 84, 99, 74, 84, 47, 63, 71, 75, 33, 50, 97, 105, 87, 63, 61, 99, 92, 83, 99, 231, 
    0, 15, 0, 0, 96, 93, 0, 25, 99, 84, 76, 34, 82, 68, 51, 96, 45, 4, 95, 124, 53, 36, 104, 130, 85, 89, 57, 85, 88, 94, 109, 237, 
    0, 24, 0, 0, 61, 108, 0, 15, 50, 63, 132, 11, 58, 48, 15, 94, 90, 0, 46, 65, 82, 111, 101, 103, 59, 72, 61, 74, 95, 105, 111, 232, 
    0, 33, 2, 0, 42, 97, 13, 7, 81, 47, 110, 64, 43, 11, 0, 57, 118, 57, 44, 60, 95, 128, 114, 77, 41, 39, 51, 66, 95, 88, 93, 216, 
    0, 22, 13, 0, 41, 97, 0, 0, 48, 106, 51, 14, 0, 0, 0, 23, 77, 80, 99, 95, 90, 75, 76, 51, 33, 19, 23, 39, 67, 57, 55, 187, 
    0, 0, 19, 0, 48, 102, 0, 0, 0, 46, 45, 0, 0, 0, 0, 16, 61, 66, 94, 86, 57, 35, 21, 22, 29, 18, 12, 17, 33, 32, 29, 163, 
    0, 0, 0, 0, 31, 47, 0, 0, 0, 14, 69, 64, 26, 26, 32, 32, 53, 52, 44, 33, 28, 28, 20, 18, 19, 21, 10, 9, 24, 21, 21, 166, 
    0, 0, 0, 0, 34, 0, 0, 0, 4, 70, 95, 58, 41, 37, 37, 33, 29, 33, 35, 27, 21, 25, 23, 19, 10, 12, 15, 13, 16, 15, 18, 171, 
    11, 7, 0, 0, 34, 0, 0, 0, 71, 81, 61, 33, 26, 29, 33, 34, 36, 37, 36, 29, 20, 21, 18, 7, 0, 2, 10, 6, 13, 6, 0, 172, 
    2, 27, 6, 0, 0, 0, 0, 42, 102, 70, 23, 25, 32, 30, 33, 35, 36, 33, 27, 22, 15, 4, 4, 1, 3, 7, 11, 1, 0, 0, 0, 183, 
    0, 24, 22, 13, 0, 0, 0, 102, 83, 52, 23, 17, 40, 38, 28, 27, 27, 24, 22, 15, 14, 2, 0, 7, 19, 23, 10, 0, 0, 0, 0, 191, 
    1, 15, 15, 16, 6, 0, 0, 107, 74, 35, 27, 15, 26, 36, 35, 27, 28, 22, 19, 13, 15, 16, 5, 8, 19, 24, 0, 0, 0, 38, 9, 174, 
    3, 18, 7, 15, 18, 0, 0, 60, 82, 32, 22, 13, 13, 20, 35, 32, 26, 18, 16, 20, 17, 16, 22, 17, 9, 0, 0, 0, 21, 55, 6, 146, 
    0, 36, 7, 13, 16, 31, 18, 29, 59, 46, 27, 24, 19, 19, 23, 20, 15, 14, 12, 19, 24, 24, 29, 8, 0, 0, 0, 8, 28, 42, 37, 140, 
    0, 31, 14, 11, 14, 23, 35, 32, 45, 48, 31, 37, 34, 36, 32, 22, 14, 3, 0, 5, 29, 29, 26, 0, 0, 0, 0, 27, 51, 28, 44, 149, 
    
    -- channel=1
    33, 94, 95, 98, 98, 97, 97, 98, 96, 97, 93, 95, 98, 101, 103, 100, 96, 93, 92, 92, 90, 87, 84, 84, 82, 81, 77, 75, 69, 63, 57, 0, 
    48, 156, 157, 159, 161, 159, 163, 165, 163, 161, 160, 161, 163, 166, 167, 168, 166, 163, 155, 146, 130, 123, 116, 120, 127, 130, 132, 133, 127, 122, 116, 44, 
    48, 155, 157, 155, 162, 164, 169, 171, 168, 167, 171, 177, 189, 178, 168, 171, 167, 152, 138, 116, 118, 113, 107, 99, 92, 107, 109, 126, 132, 130, 121, 47, 
    50, 159, 164, 161, 161, 164, 167, 169, 166, 168, 201, 214, 238, 191, 165, 153, 134, 103, 91, 112, 127, 124, 113, 99, 96, 89, 108, 116, 124, 129, 125, 47, 
    49, 155, 156, 153, 161, 164, 167, 166, 166, 165, 194, 199, 193, 159, 122, 94, 66, 72, 96, 114, 136, 139, 131, 113, 92, 92, 82, 86, 107, 126, 132, 52, 
    37, 119, 121, 109, 142, 168, 168, 168, 168, 167, 170, 167, 185, 144, 109, 89, 75, 79, 90, 122, 161, 160, 136, 120, 114, 92, 68, 70, 86, 110, 129, 51, 
    29, 107, 92, 104, 143, 167, 166, 167, 169, 167, 156, 143, 150, 146, 126, 97, 78, 84, 102, 136, 170, 170, 142, 123, 107, 84, 64, 42, 65, 93, 122, 53, 
    39, 130, 106, 100, 166, 176, 169, 172, 180, 167, 163, 145, 166, 171, 144, 107, 81, 84, 92, 123, 148, 165, 144, 111, 91, 81, 62, 46, 44, 69, 110, 59, 
    59, 167, 159, 151, 185, 189, 170, 187, 216, 246, 239, 222, 187, 184, 149, 114, 87, 81, 73, 91, 141, 181, 153, 118, 102, 85, 74, 50, 40, 53, 84, 45, 
    64, 215, 178, 203, 221, 197, 156, 197, 232, 293, 276, 226, 194, 197, 165, 117, 98, 60, 71, 98, 147, 211, 180, 141, 100, 89, 94, 65, 39, 33, 60, 26, 
    61, 233, 202, 224, 244, 218, 155, 167, 200, 243, 279, 251, 217, 212, 187, 131, 101, 72, 78, 117, 187, 240, 181, 140, 102, 96, 97, 89, 59, 43, 39, 10, 
    56, 232, 184, 241, 256, 219, 160, 136, 152, 207, 247, 233, 217, 241, 219, 160, 134, 87, 119, 138, 213, 238, 175, 135, 100, 97, 102, 92, 73, 63, 48, 4, 
    52, 235, 187, 237, 246, 193, 163, 134, 136, 143, 211, 223, 263, 273, 261, 192, 155, 111, 135, 151, 224, 241, 166, 126, 86, 84, 91, 100, 99, 92, 72, 20, 
    56, 250, 198, 224, 224, 183, 160, 136, 133, 115, 197, 231, 268, 269, 248, 198, 168, 132, 144, 152, 228, 230, 167, 135, 105, 93, 108, 121, 118, 115, 97, 31, 
    67, 263, 214, 232, 216, 175, 156, 151, 143, 129, 220, 260, 298, 281, 228, 197, 155, 120, 145, 158, 212, 215, 171, 113, 87, 89, 107, 125, 125, 120, 109, 50, 
    81, 278, 229, 249, 222, 189, 153, 171, 151, 143, 177, 247, 249, 203, 181, 149, 143, 129, 140, 146, 209, 201, 164, 134, 107, 93, 106, 116, 116, 120, 127, 58, 
    94, 292, 251, 264, 229, 193, 150, 169, 177, 155, 161, 177, 194, 184, 144, 129, 137, 133, 148, 143, 143, 141, 154, 112, 60, 56, 78, 101, 125, 140, 142, 64, 
    103, 297, 266, 273, 244, 205, 159, 174, 189, 174, 127, 137, 139, 167, 160, 139, 147, 142, 149, 143, 153, 148, 115, 67, 53, 41, 77, 106, 139, 149, 147, 70, 
    105, 295, 275, 273, 257, 214, 166, 151, 192, 178, 129, 148, 112, 151, 166, 164, 166, 146, 136, 163, 141, 97, 77, 50, 42, 58, 107, 132, 161, 160, 158, 74, 
    99, 276, 284, 275, 260, 222, 182, 161, 196, 206, 122, 101, 102, 160, 208, 223, 195, 149, 125, 118, 91, 54, 35, 22, 30, 68, 111, 140, 163, 163, 151, 69, 
    90, 254, 291, 274, 255, 216, 185, 185, 247, 264, 228, 184, 174, 239, 262, 264, 242, 184, 120, 101, 61, 56, 45, 46, 66, 91, 131, 148, 153, 151, 140, 66, 
    80, 236, 296, 279, 252, 218, 217, 246, 337, 341, 270, 232, 185, 194, 214, 219, 194, 156, 100, 69, 65, 65, 67, 71, 70, 89, 106, 125, 136, 131, 115, 69, 
    50, 192, 258, 270, 260, 248, 270, 297, 371, 365, 281, 159, 132, 133, 141, 142, 127, 120, 101, 87, 70, 68, 74, 81, 85, 88, 97, 110, 108, 105, 99, 60, 
    11, 138, 201, 224, 243, 262, 276, 327, 374, 314, 210, 148, 108, 101, 105, 98, 96, 94, 77, 72, 74, 78, 79, 80, 90, 97, 105, 108, 107, 105, 98, 59, 
    0, 111, 145, 186, 202, 258, 305, 350, 335, 235, 147, 106, 85, 80, 76, 71, 67, 69, 68, 69, 75, 80, 86, 93, 101, 113, 114, 111, 109, 113, 119, 88, 
    0, 103, 101, 121, 164, 239, 303, 337, 285, 180, 116, 89, 86, 81, 75, 75, 75, 75, 75, 78, 80, 88, 98, 107, 111, 108, 103, 105, 111, 134, 152, 100, 
    0, 107, 92, 91, 123, 214, 269, 310, 259, 155, 97, 93, 84, 84, 78, 73, 75, 77, 80, 83, 85, 93, 97, 100, 102, 101, 97, 106, 130, 147, 136, 76, 
    0, 107, 91, 86, 94, 153, 223, 236, 229, 119, 92, 94, 97, 96, 86, 81, 73, 74, 77, 85, 87, 88, 95, 98, 96, 92, 100, 118, 127, 106, 100, 55, 
    1, 115, 92, 82, 87, 103, 146, 164, 152, 94, 77, 78, 88, 99, 94, 88, 84, 89, 95, 94, 91, 91, 86, 83, 91, 107, 128, 135, 125, 106, 94, 37, 
    4, 108, 92, 81, 85, 89, 96, 107, 117, 70, 63, 65, 72, 77, 79, 83, 87, 95, 103, 111, 112, 100, 86, 87, 105, 135, 157, 160, 139, 97, 66, 28, 
    4, 113, 95, 80, 83, 84, 84, 74, 75, 58, 49, 46, 56, 58, 63, 62, 64, 84, 108, 120, 116, 102, 89, 95, 109, 147, 168, 162, 126, 90, 65, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 11, 0, 0, 0, 0, 
    
    -- channel=2
    41, 13, 19, 13, 8, 16, 14, 12, 11, 13, 18, 19, 13, 10, 12, 10, 12, 17, 21, 18, 15, 16, 14, 16, 13, 12, 12, 12, 12, 12, 13, 0, 
    66, 23, 32, 23, 20, 30, 26, 23, 21, 26, 31, 29, 23, 23, 28, 29, 30, 33, 31, 26, 25, 26, 29, 32, 29, 29, 20, 20, 23, 23, 21, 0, 
    64, 21, 34, 28, 27, 31, 26, 23, 22, 27, 41, 29, 5, 16, 32, 35, 36, 27, 25, 33, 23, 16, 13, 25, 30, 32, 30, 25, 23, 22, 20, 0, 
    69, 29, 34, 27, 30, 33, 27, 21, 25, 34, 71, 24, 0, 3, 33, 27, 20, 24, 46, 34, 12, 0, 0, 1, 11, 28, 22, 28, 27, 21, 17, 0, 
    76, 32, 33, 30, 27, 32, 27, 21, 26, 36, 80, 13, 0, 0, 19, 21, 24, 31, 52, 32, 2, 0, 0, 0, 0, 0, 10, 35, 37, 20, 14, 0, 
    79, 14, 19, 49, 34, 27, 28, 24, 27, 33, 75, 22, 0, 0, 1, 13, 5, 25, 62, 36, 0, 0, 0, 0, 0, 0, 0, 22, 45, 24, 11, 0, 
    79, 0, 11, 58, 32, 18, 28, 30, 31, 33, 37, 34, 28, 0, 0, 7, 7, 10, 49, 40, 0, 0, 0, 0, 0, 0, 0, 12, 48, 36, 12, 0, 
    72, 0, 5, 65, 8, 6, 32, 37, 39, 20, 16, 47, 42, 0, 0, 0, 1, 0, 27, 46, 0, 0, 0, 0, 0, 0, 0, 0, 37, 55, 22, 0, 
    70, 0, 3, 27, 0, 0, 31, 62, 71, 0, 0, 16, 22, 0, 0, 0, 0, 0, 7, 67, 25, 0, 0, 0, 0, 0, 0, 0, 7, 56, 44, 0, 
    67, 0, 23, 0, 0, 0, 23, 91, 97, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 85, 43, 0, 0, 0, 2, 0, 0, 0, 0, 44, 54, 0, 
    66, 0, 18, 0, 0, 0, 4, 88, 111, 3, 0, 0, 0, 0, 0, 0, 0, 0, 26, 114, 16, 0, 0, 0, 3, 3, 0, 0, 0, 11, 45, 0, 
    46, 0, 36, 0, 0, 0, 0, 49, 123, 21, 0, 0, 21, 0, 0, 0, 0, 0, 42, 122, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 7, 0, 
    36, 0, 50, 0, 0, 0, 3, 0, 108, 50, 0, 23, 38, 0, 0, 0, 0, 0, 57, 108, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    34, 0, 48, 0, 0, 0, 12, 0, 78, 57, 10, 36, 25, 0, 0, 0, 0, 0, 58, 85, 0, 0, 0, 0, 0, 5, 8, 2, 0, 0, 0, 0, 
    45, 0, 33, 0, 0, 0, 21, 0, 50, 54, 62, 43, 0, 0, 0, 0, 0, 0, 46, 61, 0, 0, 0, 0, 0, 10, 13, 0, 0, 0, 0, 0, 
    63, 0, 16, 0, 0, 0, 25, 0, 1, 46, 97, 15, 0, 0, 0, 0, 0, 0, 39, 48, 0, 0, 0, 0, 0, 15, 7, 0, 0, 0, 7, 0, 
    82, 0, 0, 0, 0, 0, 19, 0, 0, 36, 67, 12, 0, 0, 0, 0, 0, 0, 18, 3, 19, 1, 0, 0, 0, 24, 16, 0, 0, 10, 13, 0, 
    96, 0, 0, 0, 0, 0, 17, 0, 0, 0, 12, 7, 0, 0, 4, 0, 0, 10, 2, 0, 26, 0, 0, 0, 2, 23, 15, 0, 0, 10, 8, 0, 
    109, 0, 0, 0, 0, 0, 8, 13, 0, 0, 0, 8, 16, 0, 37, 0, 0, 14, 0, 0, 3, 0, 0, 0, 28, 25, 22, 19, 7, 10, 12, 0, 
    128, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 31, 29, 36, 42, 0, 0, 0, 0, 0, 0, 0, 0, 10, 44, 24, 28, 30, 9, 14, 22, 0, 
    154, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 2, 26, 30, 16, 0, 0, 0, 0, 0, 0, 0, 3, 19, 27, 22, 23, 25, 13, 20, 25, 0, 
    180, 3, 0, 0, 0, 0, 14, 83, 0, 0, 0, 0, 7, 17, 0, 0, 0, 0, 0, 0, 1, 1, 0, 4, 1, 0, 3, 0, 0, 0, 0, 0, 
    175, 11, 0, 0, 0, 0, 34, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    141, 1, 0, 0, 0, 0, 58, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    100, 0, 0, 2, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    78, 0, 0, 7, 0, 42, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 72, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 0, 0, 0, 67, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 0, 0, 0, 23, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    163, 153, 154, 144, 139, 140, 144, 142, 145, 146, 144, 134, 138, 151, 155, 160, 158, 151, 147, 149, 143, 142, 142, 139, 137, 126, 123, 132, 139, 137, 132, 105, 
    165, 155, 154, 144, 140, 145, 144, 144, 145, 143, 126, 104, 125, 154, 155, 150, 144, 133, 143, 137, 134, 127, 139, 149, 144, 150, 139, 134, 137, 135, 129, 101, 
    163, 147, 144, 141, 137, 145, 145, 146, 147, 145, 118, 57, 80, 128, 144, 136, 143, 152, 124, 101, 70, 57, 66, 90, 122, 130, 158, 150, 138, 132, 132, 101, 
    156, 139, 141, 142, 147, 151, 156, 152, 154, 153, 142, 126, 88, 120, 149, 159, 150, 144, 112, 63, 35, 28, 25, 38, 42, 77, 118, 153, 147, 131, 130, 105, 
    153, 132, 176, 179, 158, 152, 153, 151, 150, 159, 175, 201, 188, 140, 134, 141, 123, 89, 75, 53, 43, 53, 62, 49, 47, 62, 89, 138, 153, 131, 119, 98, 
    125, 113, 147, 197, 178, 154, 152, 150, 143, 147, 156, 155, 133, 91, 58, 48, 51, 55, 77, 75, 46, 58, 82, 79, 74, 69, 81, 93, 140, 147, 128, 101, 
    74, 49, 68, 84, 139, 157, 155, 150, 138, 122, 138, 114, 80, 55, 41, 52, 62, 63, 81, 120, 92, 54, 66, 96, 95, 83, 67, 84, 117, 150, 137, 101, 
    60, 0, 16, 33, 70, 138, 152, 138, 77, 39, 24, 63, 46, 48, 53, 67, 81, 86, 99, 119, 123, 78, 50, 70, 91, 76, 54, 56, 93, 150, 157, 101, 
    74, 23, 0, 28, 78, 127, 145, 135, 48, 0, 0, 0, 38, 50, 61, 46, 71, 77, 99, 89, 64, 58, 40, 44, 58, 59, 59, 50, 59, 111, 167, 128, 
    84, 50, 48, 34, 87, 126, 138, 133, 153, 68, 48, 39, 49, 31, 48, 57, 46, 72, 77, 57, 25, 30, 51, 59, 70, 69, 54, 60, 50, 67, 115, 135, 
    77, 55, 74, 65, 92, 114, 121, 121, 165, 166, 113, 92, 58, 27, 29, 60, 49, 35, 60, 53, 44, 47, 83, 78, 83, 85, 76, 53, 40, 39, 71, 100, 
    78, 50, 59, 67, 119, 140, 130, 107, 101, 129, 125, 96, 88, 41, 21, 40, 50, 33, 32, 68, 70, 81, 83, 81, 76, 89, 96, 66, 46, 42, 60, 73, 
    73, 33, 41, 53, 105, 166, 153, 117, 99, 120, 104, 58, 56, 85, 57, 38, 48, 63, 60, 72, 74, 75, 61, 60, 71, 73, 79, 65, 42, 56, 80, 68, 
    68, 21, 46, 49, 54, 120, 147, 124, 98, 104, 95, 40, 26, 106, 110, 89, 69, 61, 77, 97, 84, 62, 69, 58, 57, 58, 50, 60, 66, 85, 100, 88, 
    66, 19, 42, 39, 20, 65, 111, 100, 79, 104, 72, 79, 66, 53, 110, 111, 107, 84, 79, 94, 106, 78, 63, 83, 89, 86, 78, 85, 106, 105, 109, 91, 
    63, 15, 35, 37, 14, 34, 96, 66, 79, 99, 138, 155, 178, 143, 110, 108, 99, 86, 78, 130, 146, 104, 62, 65, 72, 93, 104, 102, 111, 110, 111, 91, 
    72, 11, 30, 49, 33, 25, 74, 83, 52, 60, 116, 155, 134, 119, 88, 66, 72, 85, 84, 107, 137, 157, 128, 102, 115, 103, 114, 106, 93, 108, 121, 100, 
    98, 35, 35, 51, 43, 21, 49, 89, 75, 45, 50, 109, 96, 65, 44, 15, 28, 93, 99, 52, 35, 82, 130, 117, 77, 63, 75, 93, 99, 118, 133, 110, 
    123, 60, 48, 58, 50, 31, 37, 65, 54, 79, 62, 48, 104, 68, 44, 20, 2, 58, 135, 118, 104, 92, 95, 94, 60, 63, 73, 100, 120, 137, 138, 109, 
    133, 76, 52, 61, 56, 47, 46, 21, 0, 0, 62, 49, 30, 25, 15, 14, 1, 14, 79, 149, 148, 122, 74, 44, 54, 66, 105, 121, 125, 127, 129, 99, 
    113, 83, 48, 58, 58, 55, 53, 19, 0, 0, 0, 0, 0, 8, 42, 64, 46, 35, 45, 44, 52, 41, 21, 0, 0, 30, 74, 96, 104, 98, 93, 73, 
    91, 105, 62, 49, 43, 23, 3, 9, 22, 27, 28, 41, 109, 140, 154, 164, 135, 105, 88, 46, 9, 5, 15, 26, 25, 27, 36, 47, 45, 37, 31, 30, 
    74, 132, 137, 77, 46, 42, 8, 21, 52, 118, 127, 130, 113, 111, 116, 112, 96, 70, 56, 48, 38, 35, 32, 32, 30, 20, 18, 26, 29, 24, 20, 19, 
    32, 80, 135, 137, 94, 75, 67, 54, 94, 119, 90, 52, 27, 20, 21, 26, 28, 35, 39, 36, 35, 33, 27, 22, 10, 9, 9, 10, 12, 11, 0, 0, 
    9, 11, 57, 110, 125, 70, 52, 61, 105, 91, 67, 24, 22, 27, 29, 34, 36, 36, 30, 26, 21, 15, 10, 5, 13, 19, 28, 27, 13, 0, 0, 0, 
    21, 12, 28, 61, 95, 105, 66, 69, 77, 59, 30, 31, 23, 29, 35, 31, 26, 22, 19, 17, 13, 16, 17, 13, 22, 38, 48, 32, 11, 6, 25, 36, 
    24, 16, 16, 23, 47, 102, 148, 88, 68, 46, 25, 26, 26, 16, 20, 31, 30, 26, 19, 16, 20, 21, 35, 42, 35, 27, 15, 1, 13, 40, 73, 66, 
    11, 10, 16, 10, 24, 72, 161, 171, 80, 73, 53, 38, 30, 18, 11, 15, 21, 20, 20, 19, 20, 22, 26, 36, 32, 11, 0, 0, 12, 47, 63, 57, 
    14, 0, 14, 13, 13, 40, 92, 142, 102, 64, 67, 65, 63, 56, 41, 24, 13, 6, 2, 1, 8, 20, 27, 27, 16, 0, 0, 0, 0, 13, 13, 48, 
    29, 14, 11, 16, 16, 24, 38, 51, 58, 41, 42, 48, 59, 69, 75, 71, 55, 41, 24, 9, 5, 13, 20, 21, 12, 3, 0, 0, 13, 21, 24, 31, 
    108, 100, 87, 90, 96, 100, 101, 101, 98, 92, 89, 93, 91, 96, 101, 117, 129, 128, 125, 123, 113, 102, 98, 97, 114, 128, 139, 130, 105, 93, 90, 76, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 3, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 68, 12, 0, 0, 0, 0, 0, 10, 37, 52, 48, 26, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 80, 27, 0, 0, 0, 0, 2, 25, 67, 86, 85, 65, 38, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 38, 16, 11, 9, 1, 0, 34, 91, 104, 94, 75, 62, 52, 22, 0, 0, 0, 0, 0, 
    0, 40, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 39, 51, 24, 8, 15, 6, 35, 96, 114, 87, 61, 61, 60, 37, 0, 0, 0, 0, 0, 
    0, 92, 47, 0, 0, 0, 0, 0, 0, 0, 7, 0, 19, 64, 82, 48, 25, 34, 16, 19, 74, 116, 85, 49, 47, 50, 36, 10, 0, 0, 0, 2, 
    0, 141, 82, 23, 42, 8, 0, 0, 12, 85, 103, 64, 56, 105, 107, 67, 36, 41, 27, 0, 42, 115, 101, 63, 44, 37, 37, 22, 0, 0, 0, 0, 
    0, 180, 98, 88, 111, 37, 0, 0, 27, 159, 198, 125, 103, 143, 124, 76, 48, 33, 29, 0, 30, 121, 121, 92, 44, 32, 46, 37, 13, 0, 0, 0, 
    0, 184, 115, 133, 148, 66, 0, 0, 17, 160, 243, 181, 135, 161, 132, 85, 57, 45, 22, 0, 63, 150, 130, 107, 47, 36, 48, 51, 41, 0, 0, 0, 
    0, 187, 97, 156, 169, 76, 0, 0, 0, 112, 208, 157, 116, 169, 154, 95, 74, 63, 33, 0, 104, 176, 138, 106, 44, 34, 50, 51, 50, 32, 0, 0, 
    0, 195, 88, 160, 176, 69, 1, 4, 0, 35, 149, 112, 107, 172, 193, 115, 80, 87, 42, 0, 135, 192, 133, 90, 39, 28, 36, 49, 60, 51, 18, 0, 
    0, 197, 89, 177, 180, 61, 0, 4, 0, 4, 97, 91, 113, 173, 197, 133, 96, 102, 53, 18, 150, 183, 127, 89, 55, 37, 36, 48, 66, 59, 25, 1, 
    0, 200, 107, 200, 192, 67, 2, 20, 4, 0, 66, 103, 181, 204, 173, 132, 104, 94, 49, 29, 138, 165, 123, 81, 48, 35, 37, 50, 69, 54, 6, 0, 
    0, 214, 138, 205, 210, 108, 24, 54, 27, 4, 21, 107, 201, 180, 124, 90, 89, 85, 36, 14, 110, 139, 117, 92, 56, 31, 46, 54, 56, 29, 0, 0, 
    0, 233, 170, 203, 224, 151, 55, 74, 73, 22, 20, 92, 155, 147, 84, 63, 69, 61, 31, 21, 53, 74, 108, 84, 30, 10, 27, 42, 36, 7, 0, 8, 
    0, 244, 196, 204, 231, 184, 79, 90, 116, 65, 33, 77, 75, 92, 67, 59, 80, 53, 45, 52, 41, 45, 82, 60, 23, 0, 7, 12, 10, 0, 0, 8, 
    0, 233, 207, 202, 223, 202, 102, 76, 133, 111, 80, 65, 30, 71, 57, 90, 117, 56, 48, 80, 50, 38, 54, 33, 3, 0, 3, 0, 4, 0, 0, 8, 
    0, 200, 209, 196, 206, 209, 134, 88, 138, 148, 107, 45, 21, 71, 77, 145, 168, 81, 41, 52, 53, 52, 24, 1, 0, 5, 4, 0, 7, 2, 0, 15, 
    0, 164, 212, 188, 192, 204, 141, 87, 173, 207, 167, 103, 71, 110, 132, 190, 212, 143, 64, 52, 41, 45, 29, 17, 24, 38, 40, 37, 49, 41, 30, 59, 
    0, 145, 225, 194, 193, 204, 138, 87, 213, 284, 215, 154, 110, 120, 159, 190, 196, 162, 98, 60, 45, 41, 46, 54, 63, 77, 74, 81, 93, 88, 78, 103, 
    0, 129, 215, 201, 205, 213, 141, 110, 231, 300, 277, 169, 119, 128, 149, 152, 158, 148, 113, 88, 70, 69, 74, 90, 105, 111, 112, 116, 119, 119, 114, 139, 
    0, 114, 173, 178, 200, 206, 134, 156, 264, 294, 257, 177, 116, 114, 122, 112, 117, 116, 95, 87, 90, 97, 101, 106, 117, 123, 128, 125, 130, 132, 129, 156, 
    0, 124, 123, 139, 178, 182, 142, 206, 292, 273, 195, 130, 103, 103, 102, 92, 88, 93, 91, 88, 95, 104, 111, 116, 121, 132, 137, 135, 139, 143, 142, 178, 
    0, 145, 110, 98, 143, 148, 142, 243, 301, 225, 140, 113, 111, 111, 106, 98, 95, 95, 94, 95, 100, 110, 121, 125, 131, 136, 135, 136, 142, 153, 159, 201, 
    0, 161, 130, 106, 108, 115, 144, 273, 289, 174, 108, 114, 114, 116, 107, 99, 99, 99, 102, 105, 109, 119, 124, 131, 139, 141, 134, 132, 147, 166, 166, 197, 
    0, 163, 140, 126, 110, 87, 131, 249, 257, 129, 107, 111, 119, 123, 110, 105, 102, 102, 107, 114, 119, 124, 126, 133, 139, 136, 131, 134, 154, 167, 155, 164, 
    0, 167, 142, 133, 130, 97, 94, 187, 194, 104, 97, 98, 107, 121, 120, 114, 109, 111, 118, 123, 124, 128, 123, 121, 125, 131, 139, 157, 176, 176, 137, 128, 
    0, 169, 141, 133, 136, 121, 93, 121, 144, 90, 81, 83, 93, 102, 110, 111, 107, 112, 121, 132, 137, 133, 123, 116, 115, 130, 158, 190, 196, 169, 113, 114, 
    0, 172, 141, 127, 131, 124, 110, 93, 99, 88, 72, 71, 81, 83, 91, 87, 84, 98, 116, 133, 144, 135, 119, 111, 106, 131, 172, 204, 194, 156, 117, 119, 
    0, 66, 50, 39, 43, 38, 34, 24, 20, 20, 8, 8, 12, 11, 12, 7, 7, 16, 28, 44, 58, 50, 36, 26, 23, 40, 70, 98, 90, 56, 36, 48, 
    
    -- channel=5
    66, 97, 98, 97, 95, 97, 95, 97, 96, 96, 96, 93, 97, 102, 102, 104, 104, 100, 98, 94, 89, 86, 84, 86, 85, 83, 79, 79, 80, 78, 74, 30, 
    145, 165, 165, 158, 158, 167, 165, 165, 162, 165, 160, 154, 159, 170, 173, 171, 167, 160, 154, 147, 143, 136, 138, 141, 138, 143, 139, 137, 136, 132, 123, 40, 
    142, 165, 167, 158, 157, 164, 168, 166, 163, 164, 168, 162, 149, 159, 166, 162, 157, 150, 138, 142, 122, 110, 100, 108, 119, 123, 140, 143, 138, 134, 129, 44, 
    140, 161, 165, 155, 160, 167, 173, 168, 169, 172, 189, 184, 150, 156, 155, 150, 138, 129, 134, 111, 101, 91, 90, 85, 82, 105, 105, 130, 141, 138, 130, 48, 
    136, 149, 163, 167, 164, 170, 170, 169, 167, 177, 210, 193, 195, 164, 139, 129, 126, 95, 94, 109, 119, 107, 94, 87, 89, 77, 97, 117, 136, 139, 131, 43, 
    129, 132, 132, 170, 176, 170, 168, 167, 167, 176, 229, 190, 150, 136, 112, 83, 58, 70, 111, 140, 137, 122, 116, 110, 95, 79, 83, 88, 118, 134, 133, 44, 
    122, 89, 102, 123, 156, 170, 171, 168, 167, 166, 174, 159, 140, 110, 79, 76, 73, 90, 122, 152, 159, 135, 114, 115, 105, 82, 56, 80, 103, 125, 136, 44, 
    123, 53, 71, 129, 141, 164, 173, 169, 162, 155, 136, 147, 143, 121, 98, 94, 95, 99, 128, 152, 165, 142, 116, 108, 102, 82, 56, 47, 86, 118, 136, 45, 
    132, 89, 86, 127, 162, 161, 168, 178, 188, 147, 125, 118, 156, 141, 115, 101, 93, 80, 105, 157, 148, 127, 120, 100, 84, 74, 66, 49, 60, 92, 128, 56, 
    147, 110, 165, 156, 163, 168, 164, 184, 223, 188, 167, 185, 175, 144, 105, 99, 81, 80, 70, 135, 158, 136, 114, 92, 98, 92, 72, 52, 48, 79, 101, 42, 
    161, 143, 174, 201, 171, 165, 153, 198, 230, 268, 199, 196, 173, 151, 109, 98, 99, 52, 77, 153, 168, 163, 131, 108, 103, 102, 102, 64, 37, 54, 87, 18, 
    145, 163, 192, 198, 168, 176, 149, 185, 218, 209, 182, 193, 204, 165, 140, 103, 101, 62, 90, 183, 189, 191, 130, 106, 103, 103, 99, 88, 56, 52, 69, 15, 
    138, 159, 194, 184, 158, 182, 163, 132, 180, 178, 177, 199, 205, 189, 158, 131, 112, 70, 135, 206, 201, 168, 119, 94, 96, 105, 105, 102, 73, 71, 69, 20, 
    135, 159, 198, 177, 150, 147, 166, 127, 158, 157, 171, 202, 232, 199, 183, 166, 138, 76, 151, 208, 191, 156, 123, 93, 84, 97, 99, 104, 99, 93, 86, 34, 
    140, 179, 203, 158, 128, 131, 159, 128, 149, 144, 185, 227, 239, 183, 168, 149, 145, 110, 150, 193, 190, 157, 109, 104, 100, 100, 121, 125, 116, 115, 116, 35, 
    154, 187, 206, 169, 116, 124, 148, 131, 140, 142, 231, 225, 226, 212, 156, 158, 129, 103, 160, 199, 172, 163, 138, 91, 87, 99, 120, 132, 120, 124, 126, 43, 
    176, 193, 204, 190, 127, 131, 138, 156, 139, 160, 193, 236, 183, 150, 144, 127, 116, 118, 155, 151, 180, 171, 122, 88, 99, 104, 115, 127, 115, 124, 136, 53, 
    195, 208, 209, 208, 144, 136, 136, 146, 137, 159, 144, 155, 152, 115, 130, 113, 105, 121, 158, 152, 142, 108, 112, 98, 67, 88, 98, 112, 130, 145, 153, 56, 
    210, 220, 217, 219, 163, 126, 146, 149, 139, 156, 122, 98, 117, 128, 157, 129, 110, 128, 141, 122, 131, 121, 78, 50, 59, 72, 106, 125, 147, 158, 156, 51, 
    214, 232, 218, 218, 185, 129, 144, 156, 149, 105, 98, 142, 114, 158, 176, 139, 124, 131, 118, 135, 119, 97, 62, 36, 66, 77, 141, 161, 164, 160, 157, 55, 
    207, 229, 218, 219, 193, 131, 145, 182, 180, 155, 65, 106, 120, 149, 194, 180, 125, 122, 115, 92, 76, 45, 41, 44, 56, 82, 118, 139, 141, 135, 124, 42, 
    195, 217, 219, 215, 191, 139, 164, 223, 197, 189, 158, 113, 162, 208, 225, 205, 154, 120, 102, 81, 47, 39, 39, 61, 75, 88, 113, 129, 114, 112, 108, 26, 
    172, 203, 229, 221, 188, 144, 198, 275, 296, 227, 180, 198, 180, 181, 181, 162, 133, 109, 71, 58, 63, 76, 81, 83, 84, 90, 94, 99, 98, 94, 87, 11, 
    140, 170, 194, 226, 196, 172, 270, 307, 303, 232, 170, 117, 108, 100, 93, 94, 73, 69, 75, 77, 79, 82, 86, 88, 86, 87, 93, 98, 93, 89, 87, 11, 
    96, 128, 152, 181, 196, 218, 278, 298, 250, 170, 107, 74, 74, 71, 68, 74, 77, 75, 75, 78, 78, 80, 81, 83, 92, 91, 96, 97, 94, 95, 98, 5, 
    72, 92, 123, 153, 149, 231, 289, 280, 189, 124, 73, 82, 78, 76, 77, 76, 75, 73, 73, 74, 80, 83, 87, 90, 95, 103, 103, 103, 107, 109, 109, 16, 
    78, 83, 91, 115, 127, 213, 303, 246, 144, 97, 81, 82, 87, 76, 70, 73, 75, 75, 76, 81, 85, 86, 95, 107, 106, 98, 94, 106, 107, 115, 132, 33, 
    81, 82, 78, 80, 113, 198, 255, 216, 129, 103, 95, 93, 81, 80, 75, 69, 73, 78, 83, 85, 86, 96, 97, 94, 92, 90, 91, 100, 110, 122, 119, 16, 
    83, 79, 76, 77, 84, 160, 199, 146, 137, 92, 89, 98, 95, 91, 84, 80, 77, 78, 77, 84, 85, 83, 89, 90, 91, 90, 102, 112, 115, 78, 74, 0, 
    82, 92, 80, 77, 76, 100, 148, 95, 83, 82, 79, 84, 88, 94, 92, 90, 86, 92, 98, 95, 86, 80, 82, 85, 94, 113, 131, 118, 88, 61, 80, 0, 
    86, 87, 82, 75, 80, 77, 89, 85, 65, 63, 67, 73, 78, 79, 73, 83, 98, 106, 110, 108, 100, 92, 81, 87, 116, 144, 149, 131, 96, 70, 64, 0, 
    58, 93, 94, 85, 84, 85, 81, 80, 70, 63, 64, 61, 65, 65, 71, 73, 76, 91, 109, 115, 107, 96, 89, 103, 120, 151, 154, 133, 99, 80, 61, 14, 
    
    -- channel=6
    58, 50, 53, 60, 56, 51, 57, 56, 57, 53, 54, 55, 54, 56, 58, 59, 59, 56, 52, 53, 53, 50, 51, 50, 56, 54, 53, 52, 54, 54, 53, 93, 
    36, 52, 53, 60, 56, 56, 58, 58, 60, 58, 56, 54, 53, 57, 60, 60, 62, 58, 55, 50, 50, 45, 43, 45, 47, 52, 55, 52, 57, 59, 57, 110, 
    37, 56, 53, 60, 53, 55, 58, 60, 58, 58, 52, 61, 57, 52, 59, 60, 60, 63, 47, 46, 43, 41, 34, 32, 36, 33, 48, 53, 57, 60, 60, 112, 
    34, 57, 55, 58, 56, 53, 59, 60, 58, 53, 27, 82, 68, 50, 53, 59, 51, 48, 36, 42, 38, 43, 40, 36, 31, 29, 30, 43, 53, 59, 58, 115, 
    32, 52, 48, 54, 59, 55, 59, 61, 57, 53, 12, 60, 73, 57, 45, 42, 49, 29, 22, 29, 29, 34, 40, 38, 36, 41, 24, 25, 41, 59, 56, 115, 
    27, 57, 20, 37, 62, 61, 58, 62, 60, 56, 32, 30, 49, 61, 52, 28, 44, 27, 4, 19, 29, 25, 26, 25, 40, 39, 35, 15, 21, 53, 57, 115, 
    31, 67, 15, 12, 51, 61, 58, 60, 63, 57, 53, 37, 37, 61, 59, 34, 39, 30, 0, 6, 39, 33, 16, 21, 33, 39, 39, 25, 5, 34, 56, 116, 
    50, 66, 19, 24, 42, 55, 56, 55, 55, 71, 47, 37, 38, 54, 52, 28, 27, 33, 5, 0, 29, 50, 29, 19, 26, 42, 37, 35, 5, 13, 53, 118, 
    50, 65, 3, 32, 52, 51, 54, 38, 48, 86, 62, 21, 37, 42, 50, 27, 23, 28, 17, 0, 12, 43, 48, 30, 22, 35, 41, 44, 22, 0, 35, 122, 
    38, 35, 10, 19, 60, 51, 59, 0, 29, 67, 80, 14, 35, 39, 40, 43, 22, 38, 8, 0, 23, 27, 55, 40, 21, 34, 34, 47, 44, 4, 8, 110, 
    44, 0, 1, 19, 63, 53, 71, 0, 0, 30, 55, 16, 27, 54, 29, 45, 32, 50, 0, 0, 40, 23, 53, 36, 18, 28, 37, 38, 49, 27, 13, 83, 
    53, 0, 0, 19, 56, 54, 72, 45, 0, 5, 33, 1, 12, 65, 42, 31, 40, 64, 0, 0, 34, 31, 44, 35, 19, 14, 35, 33, 45, 34, 35, 73, 
    57, 0, 0, 28, 29, 46, 66, 80, 0, 2, 21, 3, 0, 57, 58, 33, 29, 67, 0, 0, 28, 40, 40, 33, 24, 13, 20, 30, 38, 32, 46, 83, 
    56, 0, 0, 45, 23, 23, 56, 87, 5, 4, 5, 24, 0, 29, 46, 41, 34, 47, 0, 0, 33, 35, 44, 37, 23, 21, 13, 24, 37, 31, 38, 100, 
    49, 0, 0, 47, 49, 4, 43, 82, 26, 10, 0, 24, 42, 8, 23, 30, 39, 45, 0, 0, 31, 39, 36, 38, 19, 23, 20, 20, 41, 34, 37, 111, 
    36, 0, 0, 35, 70, 0, 30, 66, 52, 0, 0, 0, 50, 33, 16, 20, 27, 44, 0, 1, 15, 42, 39, 37, 15, 8, 19, 21, 34, 34, 44, 112, 
    28, 7, 0, 17, 75, 6, 2, 53, 69, 0, 0, 0, 14, 39, 13, 28, 17, 27, 20, 14, 0, 30, 54, 37, 23, 6, 11, 28, 28, 36, 45, 117, 
    15, 14, 0, 3, 64, 36, 0, 24, 62, 37, 12, 0, 27, 30, 20, 47, 14, 6, 48, 42, 9, 18, 38, 38, 19, 20, 7, 34, 41, 47, 53, 128, 
    0, 18, 0, 0, 44, 57, 0, 0, 31, 51, 54, 0, 35, 17, 17, 64, 32, 0, 34, 50, 51, 29, 23, 39, 13, 33, 14, 30, 42, 45, 51, 122, 
    0, 21, 3, 0, 29, 58, 0, 0, 32, 20, 60, 5, 11, 3, 10, 53, 58, 2, 6, 26, 36, 41, 32, 20, 10, 13, 17, 32, 44, 42, 50, 121, 
    0, 23, 9, 0, 25, 49, 0, 0, 57, 47, 25, 25, 4, 2, 6, 33, 59, 36, 24, 17, 16, 25, 32, 17, 9, 0, 4, 16, 34, 29, 30, 110, 
    0, 14, 14, 3, 28, 45, 0, 0, 22, 74, 54, 13, 0, 0, 0, 12, 35, 28, 40, 33, 25, 15, 16, 17, 11, 0, 0, 12, 29, 27, 25, 95, 
    0, 0, 10, 5, 26, 40, 0, 0, 0, 41, 43, 4, 0, 0, 0, 0, 7, 8, 16, 22, 18, 12, 3, 1, 1, 1, 0, 0, 9, 8, 8, 70, 
    0, 0, 0, 0, 24, 5, 0, 0, 14, 29, 15, 8, 0, 0, 0, 0, 0, 5, 6, 4, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 
    0, 0, 0, 0, 17, 0, 0, 2, 40, 20, 23, 9, 5, 6, 4, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 
    1, 0, 0, 0, 0, 0, 0, 31, 41, 16, 8, 2, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 
    0, 0, 0, 0, 0, 0, 0, 54, 36, 21, 0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 
    0, 0, 0, 0, 0, 0, 0, 63, 26, 15, 3, 0, 4, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 
    0, 0, 0, 0, 0, 0, 0, 29, 23, 3, 0, 0, 0, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 45, 
    0, 4, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 6, 4, 0, 6, 43, 
    0, 5, 2, 0, 0, 1, 6, 8, 12, 13, 6, 8, 7, 9, 6, 0, 0, 0, 0, 0, 5, 5, 5, 0, 0, 0, 0, 6, 12, 3, 9, 36, 
    
    -- channel=7
    109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 23, 13, 12, 5, 6, 12, 12, 10, 0, 0, 0, 0, 0, 
    134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 40, 57, 29, 22, 5, 9, 14, 9, 0, 22, 18, 0, 0, 0, 
    141, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 19, 71, 81, 30, 7, 11, 17, 18, 1, 0, 21, 45, 17, 0, 0, 
    153, 0, 0, 52, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 23, 58, 93, 35, 0, 0, 23, 22, 0, 1, 19, 48, 46, 0, 0, 
    177, 0, 0, 75, 21, 0, 0, 0, 0, 0, 0, 0, 23, 2, 0, 0, 35, 24, 32, 79, 62, 0, 0, 15, 22, 12, 6, 13, 32, 65, 18, 0, 
    217, 0, 0, 86, 0, 0, 0, 0, 11, 0, 0, 0, 28, 0, 0, 0, 28, 21, 26, 70, 88, 4, 0, 0, 16, 26, 14, 10, 7, 51, 56, 0, 
    233, 0, 25, 67, 0, 0, 0, 0, 77, 0, 0, 0, 26, 0, 0, 0, 10, 20, 18, 89, 103, 4, 0, 0, 12, 35, 12, 7, 0, 26, 66, 0, 
    247, 0, 72, 52, 0, 0, 0, 0, 107, 61, 0, 0, 27, 0, 0, 0, 0, 7, 16, 131, 98, 0, 0, 0, 12, 46, 17, 8, 1, 12, 50, 8, 
    247, 0, 102, 54, 0, 0, 0, 0, 61, 110, 0, 0, 51, 0, 0, 0, 5, 0, 4, 159, 80, 0, 0, 0, 21, 44, 28, 11, 16, 11, 30, 0, 
    250, 0, 114, 44, 0, 0, 0, 0, 0, 115, 0, 4, 62, 12, 0, 0, 4, 0, 0, 165, 53, 0, 0, 0, 23, 37, 45, 32, 24, 12, 18, 0, 
    252, 0, 117, 26, 0, 0, 0, 0, 0, 90, 24, 41, 27, 5, 0, 0, 0, 0, 12, 153, 34, 0, 0, 0, 18, 36, 44, 47, 25, 1, 9, 0, 
    259, 0, 104, 13, 0, 0, 25, 0, 0, 64, 56, 93, 0, 0, 0, 0, 0, 0, 23, 129, 37, 0, 0, 0, 13, 47, 45, 44, 18, 0, 5, 0, 
    268, 0, 80, 19, 0, 0, 53, 0, 0, 29, 77, 77, 0, 0, 0, 12, 6, 1, 29, 95, 22, 0, 0, 0, 8, 52, 49, 30, 13, 0, 2, 0, 
    284, 0, 54, 30, 0, 0, 72, 21, 0, 0, 83, 51, 0, 0, 0, 22, 12, 29, 12, 20, 10, 41, 0, 0, 8, 50, 61, 36, 7, 0, 0, 0, 
    297, 0, 35, 39, 0, 0, 42, 71, 0, 0, 30, 25, 38, 3, 10, 25, 0, 44, 39, 0, 0, 42, 0, 0, 19, 58, 61, 50, 5, 0, 0, 0, 
    297, 0, 20, 37, 0, 0, 2, 87, 9, 0, 0, 0, 70, 4, 44, 31, 0, 32, 63, 0, 0, 2, 0, 11, 37, 71, 37, 37, 0, 0, 0, 0, 
    283, 18, 6, 27, 8, 0, 0, 99, 28, 0, 0, 0, 84, 36, 72, 22, 0, 0, 45, 1, 1, 0, 0, 39, 57, 76, 34, 20, 0, 0, 0, 0, 
    261, 65, 0, 16, 9, 0, 0, 124, 81, 0, 0, 12, 66, 55, 67, 8, 0, 0, 3, 2, 20, 31, 46, 54, 74, 65, 47, 26, 0, 0, 0, 0, 
    246, 118, 0, 10, 10, 0, 8, 146, 78, 0, 0, 0, 39, 58, 45, 12, 0, 0, 4, 6, 36, 56, 65, 66, 71, 65, 78, 62, 41, 29, 46, 5, 
    227, 149, 35, 25, 17, 0, 23, 144, 46, 0, 0, 0, 50, 69, 54, 50, 41, 28, 40, 38, 61, 71, 77, 80, 79, 81, 87, 86, 77, 66, 76, 26, 
    213, 132, 95, 78, 27, 0, 63, 109, 0, 0, 0, 9, 66, 75, 71, 73, 72, 64, 70, 75, 84, 84, 84, 89, 92, 95, 86, 86, 81, 75, 84, 32, 
    211, 102, 111, 121, 71, 21, 108, 63, 0, 0, 0, 50, 72, 72, 69, 73, 78, 77, 81, 85, 91, 93, 89, 95, 97, 93, 81, 80, 84, 88, 98, 31, 
    214, 74, 95, 117, 103, 78, 131, 19, 0, 0, 52, 76, 75, 73, 75, 78, 76, 77, 81, 86, 90, 95, 95, 91, 90, 83, 81, 88, 104, 100, 96, 20, 
    220, 70, 84, 100, 102, 135, 159, 0, 0, 0, 69, 82, 80, 66, 76, 81, 79, 79, 82, 87, 89, 89, 98, 97, 87, 80, 91, 109, 117, 93, 84, 21, 
    221, 76, 86, 93, 97, 129, 178, 22, 0, 34, 72, 82, 85, 67, 72, 76, 80, 85, 89, 87, 91, 90, 97, 97, 89, 89, 102, 115, 105, 82, 76, 46, 
    223, 68, 89, 97, 93, 106, 139, 79, 0, 56, 77, 90, 93, 76, 72, 71, 83, 86, 87, 86, 87, 86, 88, 95, 101, 107, 107, 109, 84, 64, 66, 69, 
    228, 63, 84, 102, 90, 93, 100, 93, 30, 64, 84, 97, 91, 87, 84, 77, 85, 87, 89, 85, 75, 74, 82, 92, 110, 120, 110, 75, 51, 55, 71, 62, 
    228, 68, 74, 98, 90, 87, 79, 79, 69, 64, 84, 97, 89, 91, 84, 87, 98, 97, 94, 87, 66, 63, 76, 88, 116, 118, 99, 53, 39, 57, 86, 40, 
    170, 76, 74, 89, 87, 85, 77, 75, 77, 70, 80, 87, 79, 85, 80, 84, 92, 92, 91, 87, 68, 64, 76, 79, 101, 101, 90, 64, 52, 68, 89, 45, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 46, 64, 55, 31, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 38, 60, 68, 62, 50, 33, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 24, 40, 42, 38, 34, 26, 29, 31, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 27, 16, 26, 23, 13, 6, 7, 16, 24, 25, 0, 0, 0, 0, 0, 
    37, 53, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 18, 30, 29, 9, 6, 13, 13, 5, 6, 11, 23, 25, 7, 0, 0, 0, 0, 
    66, 96, 83, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 18, 14, 27, 22, 14, 3, 13, 30, 19, 14, 16, 22, 30, 20, 0, 0, 0, 0, 
    79, 124, 114, 52, 0, 0, 0, 0, 0, 28, 36, 5, 15, 14, 16, 12, 23, 20, 19, 19, 32, 43, 30, 23, 21, 27, 32, 35, 14, 0, 0, 0, 
    89, 125, 133, 69, 0, 0, 0, 0, 0, 18, 28, 0, 10, 13, 9, 15, 22, 25, 28, 34, 57, 49, 40, 28, 25, 32, 34, 42, 37, 11, 0, 0, 
    94, 125, 131, 79, 0, 0, 0, 0, 0, 0, 2, 0, 10, 25, 16, 14, 27, 31, 33, 50, 73, 54, 43, 30, 28, 29, 38, 44, 47, 23, 0, 0, 
    93, 119, 122, 96, 0, 0, 0, 0, 0, 0, 0, 0, 22, 49, 37, 25, 28, 40, 39, 64, 76, 63, 46, 38, 40, 34, 42, 48, 43, 9, 0, 0, 
    93, 110, 117, 118, 34, 0, 0, 0, 0, 0, 1, 28, 50, 77, 50, 35, 26, 27, 29, 55, 68, 56, 47, 38, 42, 39, 40, 40, 16, 0, 0, 0, 
    99, 115, 122, 132, 77, 13, 0, 0, 0, 0, 0, 52, 64, 55, 35, 27, 22, 4, 0, 0, 29, 32, 41, 38, 39, 44, 36, 13, 0, 0, 0, 0, 
    109, 136, 140, 144, 113, 66, 25, 0, 0, 0, 0, 37, 48, 17, 12, 14, 21, 0, 0, 0, 0, 7, 21, 23, 20, 30, 23, 0, 0, 0, 0, 0, 
    118, 152, 161, 159, 141, 97, 82, 34, 0, 0, 0, 8, 0, 0, 0, 20, 38, 12, 0, 0, 0, 0, 10, 8, 11, 2, 0, 0, 0, 0, 0, 0, 
    109, 145, 163, 164, 152, 110, 92, 76, 49, 14, 0, 0, 0, 0, 9, 42, 52, 30, 0, 0, 0, 0, 10, 5, 18, 0, 0, 0, 0, 0, 0, 0, 
    88, 119, 141, 145, 141, 118, 106, 111, 92, 67, 25, 0, 11, 21, 37, 76, 64, 30, 7, 0, 1, 18, 18, 34, 43, 0, 0, 0, 0, 0, 0, 0, 
    77, 106, 120, 121, 122, 115, 114, 133, 132, 108, 88, 50, 72, 81, 92, 118, 98, 54, 26, 19, 41, 64, 76, 95, 108, 84, 22, 0, 0, 0, 0, 0, 
    97, 145, 134, 120, 119, 115, 117, 132, 168, 150, 129, 128, 132, 144, 150, 157, 144, 116, 86, 85, 107, 140, 161, 175, 195, 188, 168, 151, 138, 140, 149, 105, 
    141, 221, 179, 150, 138, 125, 115, 125, 165, 179, 171, 178, 182, 193, 189, 198, 201, 191, 184, 182, 200, 224, 238, 256, 273, 284, 292, 288, 281, 284, 291, 188, 
    192, 291, 239, 193, 157, 134, 109, 133, 157, 191, 213, 218, 221, 228, 222, 232, 245, 245, 246, 257, 272, 285, 289, 302, 316, 321, 326, 322, 321, 324, 332, 207, 
    236, 332, 285, 234, 179, 143, 117, 142, 167, 218, 232, 251, 254, 256, 251, 253, 261, 269, 274, 288, 301, 311, 318, 325, 332, 330, 328, 327, 335, 344, 353, 217, 
    264, 363, 311, 263, 214, 157, 145, 160, 197, 228, 255, 275, 276, 277, 269, 266, 266, 274, 283, 295, 312, 325, 335, 339, 340, 337, 335, 346, 363, 371, 372, 232, 
    274, 384, 343, 293, 250, 204, 189, 195, 215, 232, 266, 284, 282, 281, 275, 271, 272, 281, 291, 305, 323, 338, 351, 351, 352, 350, 357, 374, 389, 384, 374, 232, 
    274, 394, 371, 335, 287, 248, 237, 225, 226, 245, 272, 288, 288, 285, 279, 278, 279, 289, 301, 315, 332, 344, 356, 358, 357, 361, 377, 394, 403, 381, 361, 212, 
    271, 395, 384, 363, 328, 274, 264, 251, 237, 257, 277, 286, 293, 293, 286, 285, 285, 295, 307, 318, 333, 341, 346, 349, 352, 365, 384, 406, 410, 377, 343, 199, 
    265, 384, 377, 367, 348, 305, 271, 273, 251, 265, 278, 284, 290, 292, 288, 284, 284, 294, 307, 319, 326, 330, 330, 332, 338, 358, 381, 404, 398, 370, 327, 201, 
    260, 368, 356, 354, 345, 322, 288, 276, 268, 272, 276, 279, 283, 284, 279, 273, 272, 286, 302, 313, 316, 315, 310, 313, 321, 340, 364, 377, 377, 362, 329, 201, 
    177, 237, 224, 225, 223, 214, 197, 183, 182, 181, 181, 183, 183, 182, 177, 172, 172, 181, 193, 204, 205, 199, 196, 195, 202, 213, 230, 239, 240, 231, 221, 136, 
    
    -- channel=10
    89, 61, 67, 61, 56, 61, 61, 59, 55, 55, 60, 60, 62, 64, 59, 56, 51, 50, 55, 56, 54, 52, 52, 55, 52, 48, 43, 41, 37, 32, 28, 0, 
    148, 94, 102, 92, 88, 96, 98, 94, 92, 91, 95, 96, 97, 97, 91, 90, 86, 84, 81, 77, 70, 68, 74, 77, 81, 82, 78, 73, 68, 60, 53, 0, 
    145, 87, 99, 93, 90, 100, 101, 96, 92, 98, 124, 122, 100, 96, 92, 90, 90, 70, 72, 79, 81, 71, 63, 67, 62, 72, 80, 78, 73, 66, 59, 0, 
    147, 89, 97, 94, 90, 99, 99, 93, 92, 106, 184, 171, 111, 94, 96, 78, 55, 54, 78, 102, 109, 100, 91, 73, 73, 70, 76, 81, 81, 70, 62, 0, 
    145, 83, 96, 99, 96, 98, 98, 90, 91, 103, 171, 167, 93, 68, 57, 51, 43, 52, 103, 140, 146, 134, 105, 96, 85, 62, 57, 77, 93, 82, 68, 0, 
    145, 46, 59, 100, 105, 98, 96, 92, 90, 100, 155, 139, 90, 74, 55, 52, 44, 67, 146, 184, 168, 142, 126, 117, 100, 68, 38, 58, 96, 91, 71, 0, 
    148, 40, 41, 105, 118, 99, 92, 95, 92, 88, 95, 105, 116, 96, 58, 69, 81, 85, 150, 206, 182, 134, 117, 120, 103, 54, 29, 40, 86, 101, 80, 0, 
    171, 33, 69, 139, 133, 103, 97, 104, 115, 86, 83, 123, 157, 132, 78, 82, 93, 86, 117, 187, 184, 126, 100, 104, 90, 64, 37, 21, 58, 103, 93, 0, 
    221, 82, 129, 187, 143, 104, 100, 154, 205, 183, 132, 167, 187, 149, 93, 88, 90, 68, 86, 170, 191, 144, 110, 92, 87, 75, 59, 29, 24, 77, 100, 0, 
    235, 138, 207, 228, 144, 105, 90, 185, 282, 246, 176, 204, 207, 148, 110, 83, 86, 54, 68, 183, 220, 182, 119, 85, 100, 95, 74, 38, 12, 47, 86, 0, 
    248, 169, 251, 252, 155, 110, 89, 149, 295, 289, 206, 210, 227, 160, 119, 102, 84, 35, 88, 239, 244, 193, 128, 81, 99, 115, 95, 63, 21, 35, 64, 0, 
    232, 177, 276, 253, 158, 115, 90, 110, 243, 264, 184, 211, 261, 196, 139, 118, 113, 44, 123, 282, 257, 182, 120, 79, 101, 114, 99, 82, 53, 48, 49, 0, 
    227, 180, 291, 231, 138, 120, 102, 56, 167, 225, 193, 226, 300, 240, 156, 138, 132, 60, 156, 306, 249, 162, 104, 78, 88, 103, 112, 107, 86, 75, 55, 0, 
    231, 190, 302, 215, 111, 121, 121, 47, 113, 183, 206, 253, 289, 236, 172, 165, 144, 71, 174, 296, 229, 161, 121, 93, 97, 107, 125, 136, 111, 87, 70, 0, 
    252, 214, 305, 208, 97, 129, 141, 71, 109, 170, 262, 329, 276, 216, 170, 156, 136, 87, 173, 269, 223, 149, 109, 82, 90, 113, 137, 147, 110, 91, 86, 0, 
    280, 230, 303, 236, 113, 135, 163, 107, 86, 167, 257, 292, 222, 157, 156, 147, 120, 90, 177, 235, 201, 165, 131, 87, 89, 118, 129, 125, 102, 92, 95, 0, 
    316, 245, 296, 269, 142, 125, 190, 152, 106, 148, 221, 235, 166, 122, 136, 123, 119, 129, 146, 139, 160, 161, 98, 57, 63, 95, 117, 113, 102, 105, 103, 0, 
    346, 261, 297, 292, 180, 125, 191, 200, 132, 130, 142, 157, 150, 129, 150, 126, 112, 152, 163, 128, 126, 128, 80, 33, 48, 76, 113, 117, 111, 113, 100, 0, 
    358, 270, 291, 296, 213, 123, 178, 205, 163, 155, 96, 119, 137, 142, 200, 160, 100, 158, 160, 112, 112, 93, 42, 22, 61, 87, 127, 136, 122, 111, 94, 0, 
    351, 280, 281, 291, 237, 139, 175, 245, 185, 130, 76, 107, 156, 193, 254, 202, 117, 127, 131, 96, 72, 34, 15, 30, 68, 100, 134, 141, 111, 98, 90, 0, 
    333, 291, 273, 283, 238, 132, 178, 304, 296, 200, 137, 168, 216, 260, 304, 249, 152, 134, 110, 77, 52, 43, 56, 74, 109, 129, 143, 144, 119, 106, 102, 0, 
    315, 314, 275, 281, 239, 150, 234, 375, 359, 268, 186, 181, 219, 258, 265, 225, 150, 109, 91, 70, 70, 85, 93, 113, 126, 141, 158, 157, 134, 126, 124, 0, 
    265, 308, 282, 289, 253, 192, 300, 432, 411, 265, 167, 162, 186, 197, 188, 177, 144, 121, 100, 88, 104, 123, 134, 140, 144, 153, 161, 164, 155, 147, 145, 2, 
    212, 247, 267, 293, 243, 236, 363, 436, 353, 236, 139, 130, 151, 151, 146, 145, 128, 120, 118, 123, 132, 136, 143, 151, 160, 165, 169, 172, 162, 157, 162, 10, 
    180, 198, 229, 273, 246, 285, 406, 398, 256, 142, 106, 123, 131, 128, 122, 124, 126, 125, 125, 132, 143, 147, 151, 164, 176, 178, 176, 175, 172, 183, 199, 22, 
    167, 157, 185, 223, 229, 322, 426, 338, 174, 104, 127, 142, 138, 132, 130, 130, 128, 129, 131, 138, 150, 160, 170, 175, 177, 174, 166, 178, 198, 212, 218, 28, 
    176, 151, 157, 180, 202, 341, 425, 279, 126, 116, 139, 151, 143, 129, 128, 131, 132, 134, 139, 150, 154, 160, 174, 181, 174, 161, 168, 198, 216, 210, 207, 19, 
    177, 156, 151, 155, 180, 291, 381, 220, 110, 130, 147, 158, 152, 141, 135, 131, 130, 139, 147, 153, 159, 164, 171, 169, 161, 162, 184, 203, 205, 173, 172, 10, 
    183, 157, 158, 154, 160, 220, 277, 179, 102, 120, 132, 152, 158, 151, 144, 142, 148, 154, 156, 160, 157, 153, 154, 159, 171, 190, 212, 222, 194, 134, 139, 12, 
    186, 155, 158, 159, 153, 167, 199, 151, 102, 112, 123, 135, 139, 141, 139, 142, 152, 165, 177, 176, 161, 151, 146, 159, 192, 233, 249, 215, 160, 122, 124, 9, 
    189, 155, 153, 155, 153, 143, 142, 131, 106, 97, 112, 121, 126, 123, 115, 125, 146, 166, 183, 182, 162, 149, 141, 164, 210, 252, 249, 197, 146, 125, 121, 1, 
    89, 51, 50, 54, 54, 50, 40, 37, 29, 21, 29, 31, 30, 32, 32, 39, 51, 63, 76, 74, 55, 46, 47, 61, 89, 112, 106, 72, 39, 39, 34, 0, 
    
    -- channel=11
    37, 42, 41, 44, 42, 38, 41, 40, 42, 41, 42, 45, 40, 38, 42, 43, 44, 43, 42, 44, 45, 46, 46, 44, 45, 43, 45, 45, 46, 48, 49, 83, 
    2, 19, 20, 29, 25, 20, 22, 22, 24, 20, 18, 24, 24, 20, 24, 22, 23, 23, 27, 35, 42, 44, 41, 37, 36, 31, 31, 28, 29, 31, 34, 87, 
    4, 20, 17, 25, 20, 18, 19, 21, 23, 20, 7, 9, 16, 18, 23, 22, 24, 36, 39, 34, 31, 32, 35, 39, 42, 42, 39, 30, 28, 30, 32, 86, 
    1, 20, 16, 24, 23, 20, 23, 25, 23, 17, 0, 5, 17, 15, 24, 36, 49, 59, 34, 24, 19, 25, 19, 20, 26, 24, 31, 34, 31, 32, 34, 89, 
    1, 31, 26, 26, 25, 20, 23, 25, 22, 17, 0, 55, 57, 40, 49, 61, 54, 34, 17, 17, 17, 26, 31, 29, 22, 35, 33, 33, 29, 30, 28, 88, 
    5, 53, 47, 37, 27, 19, 20, 23, 20, 16, 0, 33, 50, 39, 33, 28, 38, 22, 2, 4, 14, 29, 36, 27, 33, 45, 39, 29, 25, 33, 31, 89, 
    2, 60, 23, 11, 21, 22, 22, 22, 22, 23, 24, 28, 22, 32, 38, 22, 28, 22, 0, 5, 21, 28, 29, 31, 44, 53, 56, 34, 16, 30, 32, 88, 
    2, 62, 15, 0, 2, 17, 18, 17, 17, 27, 26, 9, 2, 26, 43, 34, 38, 37, 14, 9, 35, 38, 28, 34, 43, 48, 48, 48, 22, 21, 30, 89, 
    13, 45, 0, 0, 6, 12, 18, 0, 0, 0, 0, 0, 4, 30, 44, 31, 33, 48, 35, 0, 13, 36, 30, 24, 29, 41, 43, 47, 32, 20, 34, 94, 
    21, 43, 0, 0, 27, 15, 24, 0, 0, 16, 28, 0, 10, 28, 37, 33, 33, 49, 31, 0, 0, 9, 36, 36, 24, 31, 39, 54, 49, 18, 26, 100, 
    22, 15, 0, 5, 30, 12, 27, 0, 0, 31, 41, 0, 8, 24, 26, 40, 28, 58, 11, 0, 0, 8, 48, 45, 29, 33, 32, 43, 53, 28, 19, 87, 
    39, 5, 0, 14, 38, 17, 30, 5, 0, 24, 43, 8, 0, 26, 17, 27, 26, 53, 0, 0, 15, 22, 52, 43, 27, 30, 41, 39, 48, 34, 31, 71, 
    46, 0, 0, 24, 46, 28, 28, 41, 0, 18, 19, 0, 0, 22, 25, 17, 25, 64, 0, 0, 16, 34, 48, 43, 35, 30, 33, 29, 38, 31, 40, 67, 
    44, 0, 0, 37, 34, 21, 23, 49, 0, 23, 0, 0, 0, 38, 45, 20, 20, 60, 0, 0, 23, 33, 34, 29, 26, 20, 12, 19, 33, 33, 40, 76, 
    35, 0, 0, 41, 39, 5, 12, 43, 1, 4, 0, 0, 0, 15, 33, 35, 41, 47, 0, 0, 24, 31, 47, 53, 37, 30, 15, 19, 41, 34, 25, 82, 
    22, 0, 0, 23, 51, 0, 7, 32, 23, 8, 0, 12, 63, 36, 32, 29, 38, 49, 0, 0, 20, 33, 26, 34, 26, 26, 29, 32, 45, 27, 20, 86, 
    6, 0, 0, 8, 62, 12, 7, 19, 26, 0, 5, 17, 52, 54, 26, 31, 30, 27, 0, 35, 38, 45, 56, 61, 46, 35, 34, 31, 24, 17, 22, 91, 
    0, 0, 0, 0, 52, 23, 0, 22, 34, 0, 26, 23, 23, 25, 2, 24, 23, 15, 14, 9, 0, 36, 70, 61, 44, 31, 17, 20, 9, 12, 21, 92, 
    0, 6, 0, 0, 36, 42, 0, 18, 37, 20, 30, 3, 34, 20, 0, 26, 25, 5, 31, 31, 23, 36, 55, 60, 27, 25, 0, 8, 16, 19, 26, 97, 
    0, 8, 0, 0, 22, 48, 0, 0, 11, 38, 72, 8, 24, 0, 0, 27, 35, 3, 33, 55, 75, 72, 57, 51, 30, 40, 10, 15, 29, 31, 34, 100, 
    0, 9, 0, 0, 20, 58, 4, 0, 0, 0, 1, 0, 0, 0, 0, 9, 39, 16, 14, 37, 52, 51, 35, 14, 12, 13, 11, 26, 39, 35, 41, 109, 
    0, 5, 1, 0, 19, 43, 0, 0, 0, 14, 0, 7, 10, 11, 24, 43, 70, 65, 54, 35, 29, 24, 29, 26, 24, 21, 16, 16, 28, 25, 26, 97, 
    0, 15, 12, 0, 13, 21, 0, 0, 0, 45, 80, 47, 34, 40, 43, 47, 60, 48, 45, 43, 38, 28, 24, 28, 31, 25, 22, 23, 29, 26, 28, 102, 
    1, 13, 24, 7, 26, 17, 0, 0, 0, 57, 67, 41, 21, 21, 23, 20, 34, 37, 32, 31, 32, 31, 29, 26, 23, 24, 20, 20, 26, 29, 30, 105, 
    22, 2, 0, 7, 32, 0, 0, 0, 48, 71, 60, 36, 29, 31, 33, 31, 34, 35, 32, 28, 27, 27, 24, 21, 16, 21, 22, 22, 24, 18, 7, 101, 
    43, 27, 6, 2, 28, 0, 0, 10, 70, 53, 42, 28, 30, 34, 33, 30, 31, 31, 29, 27, 25, 23, 19, 17, 24, 29, 32, 28, 20, 7, 9, 120, 
    43, 37, 24, 10, 7, 0, 0, 42, 61, 41, 30, 29, 32, 31, 33, 33, 31, 29, 29, 25, 25, 27, 28, 27, 28, 30, 27, 11, 10, 23, 31, 129, 
    41, 35, 30, 24, 9, 0, 0, 77, 60, 42, 31, 21, 30, 27, 26, 30, 34, 32, 30, 26, 29, 25, 23, 30, 34, 28, 11, 9, 26, 47, 33, 117, 
    35, 31, 30, 29, 24, 0, 0, 89, 60, 45, 42, 32, 32, 32, 31, 24, 21, 18, 22, 24, 27, 31, 30, 29, 23, 12, 2, 12, 22, 43, 21, 110, 
    44, 34, 26, 30, 28, 19, 0, 43, 53, 37, 31, 32, 38, 41, 43, 33, 27, 23, 17, 17, 22, 29, 31, 21, 8, 0, 1, 18, 40, 50, 24, 102, 
    40, 37, 25, 31, 30, 34, 29, 30, 45, 42, 32, 33, 30, 33, 42, 41, 36, 29, 23, 28, 34, 30, 31, 19, 6, 0, 17, 38, 49, 42, 39, 93, 
    82, 93, 82, 81, 81, 82, 82, 79, 83, 79, 72, 76, 75, 76, 70, 63, 66, 72, 77, 89, 95, 89, 86, 73, 73, 79, 97, 110, 102, 82, 85, 110, 
    
    -- channel=12
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 
    13, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 0, 0, 
    1, 0, 6, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 0, 0, 0, 
    0, 0, 0, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=13
    3, 105, 109, 113, 110, 105, 103, 108, 100, 98, 98, 106, 112, 108, 106, 103, 95, 92, 93, 95, 97, 94, 90, 91, 86, 86, 78, 75, 65, 58, 50, 0, 
    83, 204, 209, 214, 215, 208, 211, 213, 208, 203, 206, 217, 219, 211, 205, 201, 193, 192, 188, 188, 176, 171, 167, 167, 174, 178, 175, 169, 154, 143, 132, 17, 
    77, 190, 198, 206, 215, 213, 218, 218, 212, 211, 239, 253, 250, 223, 200, 199, 199, 184, 189, 179, 184, 174, 158, 149, 139, 155, 157, 163, 156, 149, 140, 22, 
    75, 188, 196, 202, 208, 213, 216, 217, 212, 221, 306, 324, 333, 252, 208, 196, 179, 164, 171, 193, 228, 226, 209, 170, 159, 143, 148, 153, 159, 156, 149, 24, 
    75, 191, 201, 201, 206, 211, 214, 212, 209, 215, 297, 348, 342, 238, 175, 160, 136, 134, 172, 241, 302, 307, 273, 235, 191, 156, 137, 131, 153, 166, 165, 31, 
    82, 166, 173, 162, 186, 208, 211, 208, 205, 210, 275, 315, 308, 230, 178, 149, 111, 130, 208, 303, 365, 358, 322, 283, 243, 201, 134, 111, 135, 160, 171, 36, 
    95, 178, 150, 134, 175, 206, 205, 206, 206, 203, 208, 230, 250, 234, 200, 168, 150, 172, 240, 332, 389, 371, 314, 276, 256, 199, 131, 89, 115, 149, 172, 43, 
    132, 220, 178, 157, 219, 223, 208, 215, 237, 217, 222, 229, 279, 304, 267, 220, 196, 198, 224, 310, 365, 358, 295, 251, 227, 190, 137, 84, 87, 125, 159, 49, 
    205, 328, 284, 272, 299, 252, 210, 267, 339, 380, 358, 347, 359, 379, 310, 249, 208, 188, 192, 262, 331, 368, 313, 250, 214, 185, 158, 104, 70, 92, 132, 41, 
    243, 436, 393, 415, 379, 286, 205, 314, 435, 545, 510, 471, 435, 421, 341, 249, 218, 160, 165, 239, 337, 423, 347, 276, 227, 202, 193, 134, 76, 66, 99, 20, 
    266, 496, 466, 506, 436, 321, 214, 292, 475, 611, 608, 541, 491, 449, 373, 280, 230, 150, 175, 277, 407, 488, 379, 298, 231, 228, 224, 185, 112, 79, 77, 2, 
    257, 510, 482, 534, 464, 334, 223, 248, 409, 517, 548, 515, 508, 495, 431, 322, 274, 181, 232, 335, 491, 516, 384, 288, 228, 232, 230, 212, 160, 127, 91, 0, 
    258, 515, 485, 525, 464, 316, 231, 192, 300, 382, 478, 474, 549, 558, 496, 375, 316, 229, 288, 396, 529, 503, 358, 262, 208, 215, 227, 233, 215, 191, 133, 11, 
    263, 526, 500, 527, 437, 291, 232, 180, 242, 300, 420, 466, 569, 576, 518, 418, 357, 273, 322, 415, 522, 485, 355, 273, 230, 218, 238, 263, 260, 232, 173, 26, 
    283, 554, 534, 538, 415, 300, 240, 206, 237, 278, 449, 556, 629, 601, 486, 412, 357, 282, 322, 414, 504, 454, 347, 260, 221, 218, 255, 289, 277, 247, 188, 44, 
    314, 589, 568, 572, 439, 354, 274, 264, 227, 289, 415, 559, 595, 504, 413, 363, 323, 265, 314, 379, 467, 440, 367, 278, 231, 228, 259, 277, 257, 223, 189, 58, 
    353, 631, 603, 609, 486, 393, 335, 329, 294, 298, 371, 497, 480, 396, 336, 290, 291, 275, 279, 296, 359, 349, 319, 243, 175, 182, 224, 241, 232, 210, 204, 67, 
    386, 665, 637, 643, 539, 427, 375, 380, 354, 312, 299, 354, 329, 328, 318, 283, 298, 288, 298, 301, 289, 284, 273, 184, 137, 133, 189, 213, 229, 227, 223, 73, 
    397, 671, 655, 653, 575, 444, 392, 380, 403, 364, 278, 289, 246, 317, 351, 349, 335, 314, 298, 298, 263, 242, 186, 109, 111, 126, 197, 220, 251, 245, 224, 71, 
    381, 641, 654, 646, 593, 473, 420, 423, 433, 397, 270, 246, 256, 359, 434, 464, 401, 319, 276, 264, 232, 170, 98, 70, 97, 153, 211, 234, 250, 234, 207, 64, 
    350, 593, 647, 630, 583, 472, 431, 477, 562, 541, 409, 342, 365, 463, 559, 579, 483, 374, 270, 226, 171, 133, 112, 121, 167, 220, 250, 263, 256, 237, 216, 76, 
    322, 571, 651, 626, 579, 485, 483, 571, 714, 697, 540, 449, 434, 502, 569, 560, 472, 368, 256, 189, 154, 156, 169, 199, 231, 266, 292, 309, 299, 288, 270, 128, 
    273, 539, 626, 630, 595, 526, 561, 687, 852, 778, 624, 472, 422, 444, 458, 445, 400, 346, 269, 223, 212, 231, 256, 282, 300, 314, 329, 342, 339, 331, 319, 173, 
    222, 461, 545, 588, 577, 575, 636, 775, 848, 746, 555, 397, 339, 334, 333, 324, 307, 291, 267, 263, 273, 285, 298, 310, 330, 343, 357, 364, 358, 351, 348, 190, 
    188, 396, 440, 513, 539, 604, 691, 805, 771, 598, 394, 309, 283, 278, 272, 266, 267, 270, 269, 273, 289, 303, 313, 330, 350, 369, 375, 374, 371, 381, 392, 226, 
    182, 359, 359, 407, 461, 577, 715, 786, 677, 459, 330, 309, 303, 298, 287, 280, 275, 275, 275, 283, 300, 321, 341, 357, 370, 377, 369, 377, 396, 424, 444, 270, 
    199, 369, 335, 343, 384, 552, 710, 743, 586, 379, 312, 321, 312, 303, 286, 279, 280, 284, 291, 306, 317, 337, 356, 373, 379, 368, 364, 386, 420, 449, 460, 262, 
    201, 376, 338, 323, 345, 477, 643, 624, 514, 337, 318, 329, 326, 319, 298, 288, 284, 293, 306, 322, 335, 348, 359, 364, 361, 354, 367, 394, 433, 420, 405, 202, 
    206, 387, 350, 331, 335, 392, 495, 481, 408, 299, 292, 308, 325, 331, 318, 310, 306, 316, 329, 339, 341, 339, 337, 339, 351, 372, 410, 450, 449, 376, 331, 151, 
    212, 388, 354, 338, 337, 339, 374, 358, 315, 263, 260, 273, 294, 306, 307, 308, 313, 334, 358, 369, 362, 347, 328, 330, 360, 424, 483, 495, 436, 345, 281, 139, 
    218, 386, 352, 334, 335, 316, 305, 285, 258, 234, 228, 237, 259, 261, 263, 269, 289, 328, 367, 385, 379, 352, 319, 332, 378, 464, 518, 503, 426, 338, 275, 138, 
    103, 205, 182, 171, 173, 167, 150, 135, 119, 106, 100, 101, 106, 106, 109, 114, 130, 161, 196, 216, 207, 182, 162, 172, 208, 267, 299, 283, 223, 172, 136, 55, 
    
    -- channel=14
    0, 18, 17, 16, 21, 26, 23, 25, 25, 25, 21, 18, 21, 24, 27, 27, 29, 30, 27, 21, 16, 14, 11, 14, 15, 19, 18, 18, 18, 19, 21, 0, 
    107, 174, 174, 166, 167, 173, 175, 175, 175, 182, 174, 165, 166, 176, 188, 192, 190, 184, 168, 152, 137, 129, 129, 133, 135, 140, 143, 149, 152, 151, 144, 64, 
    110, 178, 180, 173, 175, 176, 181, 179, 179, 177, 179, 176, 172, 179, 188, 184, 175, 155, 143, 144, 134, 126, 113, 110, 112, 115, 128, 146, 152, 151, 147, 68, 
    111, 179, 181, 170, 170, 176, 179, 178, 180, 179, 190, 164, 160, 172, 167, 150, 127, 115, 132, 110, 93, 81, 89, 97, 99, 120, 119, 130, 142, 146, 142, 65, 
    101, 156, 160, 167, 172, 183, 182, 183, 183, 182, 169, 106, 132, 139, 122, 109, 119, 125, 94, 67, 60, 52, 43, 47, 67, 63, 90, 114, 131, 141, 148, 67, 
    84, 124, 127, 150, 171, 183, 187, 186, 187, 189, 202, 198, 164, 141, 138, 133, 91, 71, 70, 75, 69, 56, 51, 60, 42, 51, 77, 96, 110, 121, 134, 61, 
    79, 103, 143, 154, 158, 175, 185, 183, 181, 180, 170, 170, 152, 109, 81, 69, 51, 56, 73, 72, 73, 79, 77, 59, 49, 50, 41, 69, 99, 113, 131, 63, 
    57, 67, 89, 129, 150, 175, 190, 187, 182, 166, 158, 155, 126, 86, 63, 51, 46, 51, 70, 78, 74, 81, 78, 66, 67, 55, 51, 42, 76, 108, 126, 61, 
    33, 70, 75, 73, 130, 169, 180, 192, 197, 168, 163, 125, 93, 81, 71, 70, 61, 46, 59, 113, 101, 81, 80, 84, 72, 52, 44, 44, 63, 92, 108, 54, 
    35, 55, 69, 82, 113, 161, 165, 175, 128, 81, 56, 96, 91, 90, 73, 60, 54, 51, 66, 97, 99, 98, 67, 56, 64, 58, 44, 30, 41, 85, 104, 38, 
    45, 90, 56, 99, 127, 165, 159, 161, 111, 105, 88, 108, 96, 89, 76, 52, 68, 37, 72, 92, 74, 89, 59, 63, 60, 52, 60, 49, 35, 53, 89, 36, 
    31, 89, 85, 98, 114, 152, 148, 150, 186, 125, 93, 104, 111, 87, 94, 79, 64, 47, 83, 77, 69, 96, 76, 74, 65, 62, 48, 48, 33, 37, 59, 36, 
    30, 98, 94, 83, 109, 145, 152, 124, 147, 110, 122, 148, 131, 100, 97, 89, 64, 31, 83, 87, 103, 98, 81, 62, 53, 62, 65, 62, 44, 43, 56, 31, 
    35, 94, 74, 77, 129, 141, 151, 126, 130, 110, 124, 116, 122, 88, 88, 90, 80, 48, 80, 92, 94, 95, 85, 70, 64, 74, 76, 61, 53, 55, 69, 29, 
    37, 94, 79, 74, 94, 128, 142, 130, 143, 130, 136, 127, 134, 134, 109, 71, 65, 73, 92, 91, 98, 92, 50, 36, 46, 45, 57, 63, 58, 80, 107, 37, 
    45, 89, 88, 82, 61, 106, 114, 121, 108, 102, 114, 67, 56, 104, 88, 92, 88, 66, 93, 113, 106, 91, 98, 81, 67, 56, 54, 65, 79, 109, 117, 50, 
    52, 90, 88, 77, 45, 77, 85, 107, 107, 140, 99, 128, 127, 89, 100, 87, 84, 90, 97, 72, 100, 88, 51, 34, 41, 50, 63, 88, 113, 119, 126, 62, 
    52, 89, 88, 87, 60, 68, 86, 72, 93, 107, 99, 122, 123, 111, 113, 80, 82, 84, 91, 153, 168, 86, 59, 70, 59, 67, 83, 95, 116, 127, 146, 69, 
    67, 93, 90, 95, 72, 50, 77, 68, 70, 83, 97, 104, 59, 81, 89, 64, 74, 83, 75, 81, 66, 81, 83, 48, 57, 59, 91, 106, 123, 146, 157, 69, 
    82, 106, 100, 99, 84, 55, 78, 94, 89, 50, 25, 79, 70, 112, 100, 62, 68, 91, 69, 54, 38, 51, 46, 29, 26, 33, 80, 118, 142, 154, 153, 69, 
    98, 104, 105, 106, 85, 50, 64, 84, 87, 135, 112, 98, 116, 99, 87, 85, 61, 73, 94, 91, 88, 59, 43, 47, 33, 61, 73, 96, 111, 117, 108, 44, 
    98, 89, 106, 105, 89, 81, 114, 102, 53, 43, 60, 24, 15, 20, 45, 44, 23, 17, 22, 54, 47, 24, 0, 0, 0, 19, 47, 81, 80, 77, 77, 25, 
    58, 54, 83, 95, 90, 86, 110, 103, 124, 58, 4, 40, 48, 55, 70, 62, 54, 53, 29, 2, 0, 0, 0, 0, 0, 0, 7, 9, 8, 10, 2, 0, 
    39, 50, 55, 72, 63, 67, 102, 120, 123, 95, 105, 72, 62, 62, 59, 55, 35, 14, 5, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    16, 43, 65, 58, 65, 125, 128, 125, 96, 93, 52, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 18, 47, 55, 105, 117, 107, 97, 76, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 46, 71, 98, 94, 91, 35, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 61, 71, 61, 57, 13, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 34, 76, 33, 48, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 56, 56, 23, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    44, 68, 69, 67, 68, 72, 70, 70, 70, 70, 72, 70, 69, 73, 77, 78, 79, 77, 72, 66, 61, 60, 60, 63, 64, 67, 68, 69, 71, 70, 67, 50, 
    109, 84, 91, 88, 86, 88, 89, 87, 86, 89, 88, 83, 84, 92, 98, 99, 97, 91, 80, 70, 63, 61, 64, 68, 71, 72, 76, 82, 85, 82, 77, 50, 
    110, 87, 97, 96, 93, 90, 90, 86, 90, 85, 84, 76, 74, 87, 95, 94, 89, 76, 62, 55, 38, 34, 38, 47, 60, 60, 68, 74, 81, 79, 76, 52, 
    111, 87, 95, 96, 94, 95, 91, 89, 90, 89, 79, 53, 46, 73, 81, 77, 72, 58, 55, 25, 10, 0, 6, 23, 27, 47, 51, 61, 71, 75, 74, 51, 
    107, 77, 77, 86, 87, 95, 93, 92, 92, 92, 89, 51, 37, 52, 65, 57, 52, 50, 21, 8, 0, 0, 0, 0, 14, 11, 41, 55, 63, 66, 72, 50, 
    95, 58, 58, 73, 80, 88, 97, 93, 94, 91, 79, 86, 22, 26, 37, 39, 19, 15, 18, 2, 0, 0, 0, 0, 0, 0, 16, 41, 58, 64, 69, 51, 
    80, 18, 39, 62, 68, 84, 98, 97, 91, 87, 73, 69, 40, 18, 8, 10, 11, 3, 14, 0, 0, 0, 0, 0, 0, 0, 0, 28, 57, 64, 63, 49, 
    52, 0, 0, 52, 63, 77, 92, 92, 83, 70, 60, 48, 23, 3, 0, 0, 4, 0, 6, 14, 0, 0, 0, 0, 4, 0, 1, 9, 49, 69, 60, 41, 
    30, 0, 0, 8, 43, 67, 84, 78, 60, 16, 18, 11, 6, 0, 0, 0, 1, 0, 0, 29, 8, 0, 0, 2, 2, 0, 0, 8, 31, 66, 62, 35, 
    38, 0, 0, 0, 3, 51, 79, 74, 26, 0, 0, 3, 0, 0, 0, 0, 0, 2, 10, 15, 10, 0, 0, 0, 2, 1, 0, 0, 11, 54, 70, 30, 
    29, 0, 0, 0, 0, 35, 70, 72, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 63, 41, 
    27, 0, 0, 0, 0, 28, 73, 48, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 0, 0, 0, 0, 0, 2, 0, 0, 0, 5, 33, 45, 
    28, 0, 0, 0, 0, 25, 72, 53, 54, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 21, 32, 
    31, 0, 0, 0, 0, 19, 61, 58, 40, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 23, 
    32, 0, 0, 0, 0, 12, 46, 42, 31, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 25, 
    34, 0, 0, 0, 0, 0, 23, 18, 11, 33, 13, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 8, 30, 50, 43, 
    31, 0, 0, 0, 0, 0, 7, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 1, 17, 14, 0, 0, 0, 1, 12, 5, 5, 26, 38, 59, 44, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 2, 0, 0, 0, 0, 0, 0, 0, 26, 17, 0, 0, 0, 1, 17, 27, 32, 48, 63, 75, 42, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 3, 0, 0, 0, 0, 6, 0, 0, 18, 10, 0, 15, 13, 30, 53, 55, 71, 72, 43, 
    47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 0, 0, 0, 0, 0, 12, 0, 0, 0, 1, 9, 7, 13, 25, 54, 54, 57, 56, 34, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    107, 40, 42, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 42, 40, 41, 41, 42, 42, 41, 42, 41, 41, 41, 41, 42, 187, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 299, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 300, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 300, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 300, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 301, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 302, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 301, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 302, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 303, 
    26, 24, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 23, 14, 0, 0, 0, 0, 0, 302, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 11, 13, 0, 17, 31, 0, 0, 0, 0, 0, 302, 
    0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 302, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 11, 113, 63, 40, 40, 40, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 298, 
    0, 43, 35, 0, 0, 0, 0, 0, 0, 30, 130, 92, 48, 31, 8, 0, 0, 0, 0, 0, 0, 0, 6, 9, 0, 0, 7, 25, 1, 0, 0, 281, 
    10, 42, 48, 5, 0, 8, 0, 0, 0, 22, 58, 40, 0, 0, 0, 0, 0, 0, 12, 30, 47, 44, 45, 44, 33, 16, 17, 19, 0, 0, 0, 261, 
    41, 0, 0, 29, 62, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 29, 21, 28, 20, 33, 29, 14, 5, 3, 0, 0, 0, 0, 0, 0, 260, 
    63, 0, 0, 4, 43, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 8, 243, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 11, 26, 23, 19, 15, 8, 225, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 8, 0, 0, 36, 21, 0, 2, 25, 41, 33, 21, 20, 13, 7, 8, 10, 226, 
    0, 0, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 3, 0, 0, 22, 18, 12, 21, 31, 32, 23, 17, 22, 22, 17, 15, 6, 224, 
    49, 59, 57, 62, 50, 45, 41, 39, 31, 26, 21, 12, 6, 7, 8, 8, 14, 23, 29, 34, 39, 40, 41, 39, 36, 36, 42, 31, 13, 9, 8, 230, 
    119, 104, 70, 85, 104, 96, 90, 89, 86, 83, 79, 63, 59, 63, 48, 41, 39, 52, 58, 59, 58, 56, 55, 53, 43, 26, 21, 24, 20, 19, 10, 238, 
    108, 124, 70, 47, 99, 114, 112, 113, 116, 113, 113, 87, 58, 109, 97, 74, 68, 75, 78, 72, 66, 60, 46, 22, 6, 6, 27, 45, 34, 18, 0, 245, 
    111, 121, 98, 39, 62, 106, 120, 127, 129, 124, 123, 97, 0, 31, 97, 79, 70, 68, 61, 53, 40, 24, 11, 12, 30, 50, 61, 47, 17, 0, 0, 252, 
    141, 117, 113, 86, 76, 104, 122, 130, 134, 128, 123, 116, 0, 0, 43, 71, 59, 52, 49, 46, 43, 44, 56, 82, 90, 61, 30, 21, 6, 0, 0, 259, 
    148, 137, 114, 118, 109, 111, 123, 128, 128, 125, 122, 124, 65, 0, 38, 89, 83, 80, 82, 89, 100, 111, 100, 74, 49, 28, 21, 17, 0, 0, 0, 262, 
    130, 158, 120, 122, 119, 116, 122, 126, 125, 124, 123, 123, 107, 41, 68, 112, 107, 109, 115, 120, 112, 89, 54, 27, 28, 38, 30, 10, 0, 0, 0, 264, 
    108, 164, 136, 123, 122, 120, 122, 124, 124, 124, 123, 122, 116, 59, 61, 119, 130, 129, 112, 90, 64, 43, 31, 33, 40, 43, 27, 6, 0, 0, 0, 265, 
    108, 157, 145, 126, 123, 122, 123, 124, 125, 125, 124, 122, 122, 85, 75, 125, 133, 104, 64, 41, 36, 39, 44, 46, 36, 29, 22, 5, 0, 0, 0, 265, 
    115, 142, 135, 126, 121, 121, 123, 124, 123, 122, 122, 117, 118, 103, 89, 93, 79, 59, 47, 39, 43, 50, 50, 43, 31, 21, 15, 2, 0, 0, 0, 267, 
    81, 119, 111, 109, 108, 106, 104, 103, 100, 98, 97, 93, 89, 79, 59, 48, 39, 39, 44, 34, 38, 42, 33, 23, 14, 6, 0, 0, 0, 0, 0, 256, 
    
    -- channel=17
    138, 279, 277, 277, 277, 277, 277, 277, 277, 278, 278, 279, 279, 279, 278, 278, 276, 276, 276, 278, 278, 277, 278, 279, 279, 278, 278, 277, 278, 278, 278, 155, 
    153, 392, 389, 389, 389, 389, 389, 389, 389, 390, 390, 390, 390, 391, 391, 391, 389, 388, 390, 389, 389, 386, 390, 390, 390, 390, 390, 389, 390, 390, 391, 253, 
    153, 395, 392, 392, 392, 392, 392, 391, 391, 391, 391, 391, 391, 392, 392, 392, 390, 388, 386, 373, 368, 351, 372, 375, 388, 392, 391, 391, 391, 392, 392, 255, 
    153, 394, 391, 392, 392, 392, 392, 391, 391, 390, 391, 391, 391, 391, 391, 393, 392, 388, 379, 348, 339, 329, 362, 380, 388, 392, 391, 391, 392, 393, 393, 255, 
    154, 396, 392, 392, 392, 392, 392, 392, 391, 391, 392, 392, 391, 391, 390, 387, 376, 356, 338, 314, 313, 314, 349, 367, 385, 392, 392, 393, 393, 394, 395, 256, 
    150, 386, 384, 387, 388, 391, 393, 394, 393, 393, 394, 391, 389, 386, 383, 373, 348, 322, 304, 289, 283, 271, 302, 335, 372, 394, 393, 393, 394, 395, 396, 257, 
    144, 380, 385, 388, 389, 392, 395, 396, 395, 395, 396, 382, 379, 367, 375, 364, 336, 318, 307, 296, 281, 274, 295, 336, 370, 397, 396, 395, 396, 397, 398, 258, 
    146, 388, 388, 391, 393, 396, 397, 396, 395, 395, 395, 375, 373, 361, 373, 368, 354, 335, 327, 328, 319, 320, 331, 359, 385, 398, 396, 396, 398, 399, 399, 259, 
    97, 271, 279, 298, 327, 362, 393, 393, 392, 393, 394, 378, 377, 363, 380, 381, 370, 365, 363, 364, 358, 355, 345, 334, 330, 334, 334, 349, 372, 398, 401, 260, 
    50, 227, 228, 253, 301, 345, 387, 385, 385, 390, 392, 386, 389, 376, 387, 390, 385, 380, 379, 374, 353, 324, 298, 283, 271, 265, 270, 303, 350, 394, 401, 261, 
    82, 273, 271, 292, 328, 356, 372, 364, 364, 370, 376, 376, 373, 366, 375, 382, 387, 387, 385, 370, 345, 322, 312, 305, 289, 270, 268, 293, 355, 393, 401, 262, 
    114, 295, 295, 311, 326, 338, 346, 332, 322, 330, 324, 287, 244, 248, 260, 274, 287, 314, 339, 364, 367, 357, 345, 335, 319, 300, 303, 319, 357, 387, 396, 262, 
    77, 243, 241, 253, 271, 293, 316, 323, 338, 337, 280, 209, 148, 152, 161, 180, 217, 283, 348, 386, 388, 373, 358, 350, 335, 329, 333, 321, 331, 345, 367, 248, 
    22, 157, 160, 179, 212, 269, 289, 306, 332, 323, 266, 193, 132, 142, 172, 224, 281, 326, 347, 354, 339, 314, 289, 273, 262, 264, 263, 251, 263, 284, 316, 226, 
    0, 86, 114, 158, 196, 204, 216, 257, 295, 305, 289, 253, 218, 237, 264, 277, 265, 256, 258, 260, 241, 223, 207, 201, 202, 213, 226, 239, 252, 279, 309, 221, 
    0, 43, 118, 196, 216, 192, 207, 237, 291, 324, 341, 333, 319, 325, 318, 301, 272, 257, 255, 254, 245, 240, 229, 229, 229, 238, 255, 274, 283, 288, 288, 188, 
    0, 59, 185, 281, 288, 281, 279, 299, 338, 360, 372, 367, 369, 364, 365, 351, 325, 307, 292, 296, 289, 282, 276, 270, 265, 262, 260, 256, 245, 240, 237, 158, 
    0, 117, 238, 301, 326, 306, 307, 314, 328, 336, 348, 348, 351, 340, 332, 306, 276, 260, 256, 245, 234, 241, 243, 225, 211, 199, 194, 200, 209, 218, 224, 143, 
    44, 180, 232, 274, 283, 274, 275, 277, 280, 281, 284, 282, 281, 262, 253, 236, 232, 228, 214, 209, 204, 207, 201, 185, 174, 170, 176, 182, 185, 188, 191, 118, 
    31, 110, 154, 175, 178, 184, 193, 195, 197, 202, 211, 220, 224, 215, 214, 201, 200, 195, 185, 171, 152, 145, 143, 133, 125, 122, 127, 132, 139, 156, 182, 120, 
    0, 34, 46, 46, 52, 51, 52, 55, 64, 74, 84, 96, 107, 117, 122, 118, 119, 120, 120, 106, 87, 81, 83, 81, 80, 87, 101, 119, 141, 163, 183, 117, 
    0, 0, 0, 0, 11, 4, 0, 0, 0, 0, 0, 0, 11, 22, 28, 31, 41, 48, 47, 39, 35, 38, 43, 50, 64, 93, 123, 144, 153, 160, 185, 121, 
    0, 0, 0, 0, 2, 13, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 0, 0, 0, 0, 7, 24, 48, 78, 112, 140, 146, 140, 142, 167, 206, 137, 
    0, 0, 0, 0, 1, 12, 0, 0, 0, 0, 0, 0, 0, 17, 86, 101, 78, 68, 69, 71, 82, 99, 117, 133, 133, 117, 112, 135, 168, 194, 231, 157, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 113, 147, 139, 133, 129, 125, 121, 113, 98, 83, 85, 108, 142, 167, 184, 213, 256, 171, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 88, 126, 116, 107, 97, 84, 71, 57, 58, 81, 116, 144, 157, 172, 204, 240, 274, 183, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 70, 71, 57, 43, 31, 33, 51, 82, 114, 137, 149, 163, 187, 220, 250, 284, 191, 
    0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 13, 58, 94, 120, 136, 149, 166, 184, 201, 226, 258, 289, 194, 
    0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 75, 107, 131, 148, 156, 167, 181, 196, 214, 237, 269, 298, 199, 
    0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 61, 88, 110, 132, 151, 161, 168, 178, 190, 205, 224, 249, 276, 300, 201, 
    0, 75, 31, 9, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 33, 58, 84, 99, 121, 142, 152, 159, 166, 175, 186, 197, 215, 234, 254, 278, 299, 200, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 19, 23, 27, 31, 32, 35, 40, 46, 55, 63, 73, 82, 30, 
    
    -- channel=18
    94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    161, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    125, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    116, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 
    116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    112, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    87, 0, 4, 17, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    69, 43, 58, 0, 0, 0, 22, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    77, 124, 95, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    111, 152, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    146, 88, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    131, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 21, 17, 0, 0, 0, 0, 1, 4, 5, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 33, 38, 5, 0, 0, 0, 3, 12, 17, 31, 43, 14, 0, 0, 0, 0, 0, 0, 0, 1, 3, 6, 0, 0, 0, 0, 0, 1, 3, 0, 
    23, 0, 36, 53, 14, 0, 0, 0, 0, 10, 20, 36, 84, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 0, 
    27, 0, 26, 55, 33, 2, 0, 0, 0, 13, 21, 34, 107, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 9, 12, 5, 0, 
    19, 0, 15, 37, 39, 26, 17, 11, 10, 17, 24, 27, 96, 120, 31, 0, 0, 2, 2, 0, 1, 9, 20, 20, 11, 10, 12, 9, 11, 5, 0, 0, 
    18, 0, 1, 25, 30, 32, 27, 24, 23, 24, 26, 25, 56, 108, 78, 44, 45, 45, 41, 39, 37, 33, 36, 34, 21, 11, 6, 6, 9, 0, 0, 0, 
    25, 0, 0, 22, 26, 29, 26, 24, 25, 25, 26, 27, 34, 77, 86, 68, 67, 75, 79, 71, 55, 42, 34, 24, 9, 0, 0, 3, 7, 0, 0, 0, 
    27, 0, 0, 17, 23, 25, 21, 20, 23, 24, 25, 27, 28, 58, 76, 65, 74, 80, 72, 56, 42, 26, 9, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    26, 0, 0, 10, 17, 18, 15, 16, 19, 21, 21, 23, 21, 38, 56, 52, 54, 51, 46, 38, 26, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 2, 9, 10, 10, 10, 12, 14, 14, 15, 11, 19, 32, 32, 33, 29, 20, 17, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 11, 17, 20, 21, 21, 20, 21, 23, 23, 24, 25, 29, 37, 38, 38, 34, 28, 29, 22, 14, 14, 12, 12, 12, 12, 10, 10, 7, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 48, 48, 49, 49, 49, 49, 49, 49, 49, 50, 50, 50, 49, 49, 48, 49, 49, 50, 49, 49, 46, 49, 50, 50, 49, 49, 49, 49, 49, 49, 29, 
    90, 52, 53, 53, 53, 53, 53, 53, 54, 54, 54, 55, 55, 55, 54, 55, 57, 57, 57, 60, 76, 69, 69, 61, 55, 54, 54, 54, 54, 54, 53, 33, 
    90, 51, 51, 51, 51, 51, 51, 51, 52, 52, 52, 52, 52, 52, 52, 53, 53, 55, 60, 73, 93, 100, 75, 68, 54, 50, 52, 52, 51, 52, 51, 31, 
    90, 52, 52, 52, 52, 52, 52, 52, 52, 51, 51, 50, 51, 53, 52, 56, 65, 70, 71, 74, 71, 79, 60, 49, 50, 50, 51, 51, 50, 50, 50, 30, 
    95, 55, 53, 54, 52, 51, 52, 52, 51, 50, 49, 49, 54, 56, 54, 63, 86, 105, 100, 81, 74, 84, 93, 74, 55, 53, 53, 53, 52, 52, 51, 30, 
    102, 63, 58, 57, 57, 55, 53, 51, 48, 47, 49, 52, 70, 67, 60, 62, 61, 64, 63, 57, 60, 83, 105, 104, 71, 55, 55, 54, 53, 53, 52, 31, 
    85, 55, 47, 47, 53, 57, 56, 53, 49, 48, 49, 55, 70, 77, 61, 44, 32, 12, 0, 0, 0, 0, 8, 39, 64, 58, 54, 54, 54, 54, 52, 32, 
    137, 110, 113, 107, 88, 63, 59, 56, 54, 53, 54, 53, 47, 60, 54, 37, 17, 14, 5, 0, 0, 0, 0, 26, 71, 96, 95, 84, 63, 57, 54, 32, 
    158, 196, 196, 191, 159, 99, 66, 61, 55, 55, 58, 51, 36, 40, 49, 46, 29, 25, 29, 30, 47, 70, 97, 121, 138, 154, 161, 143, 94, 62, 56, 33, 
    26, 12, 17, 29, 56, 80, 75, 76, 71, 63, 66, 65, 55, 51, 57, 56, 51, 46, 47, 57, 78, 99, 99, 90, 72, 73, 93, 91, 86, 64, 57, 35, 
    6, 0, 0, 0, 0, 26, 73, 102, 101, 85, 102, 143, 148, 144, 137, 127, 115, 101, 70, 49, 29, 14, 0, 0, 0, 0, 0, 6, 38, 61, 57, 33, 
    117, 92, 94, 88, 82, 71, 73, 71, 76, 80, 108, 180, 226, 228, 226, 217, 193, 146, 98, 50, 16, 1, 0, 8, 10, 0, 0, 18, 59, 80, 72, 39, 
    150, 172, 185, 191, 159, 140, 100, 37, 14, 27, 36, 45, 75, 82, 69, 51, 40, 35, 46, 56, 70, 85, 100, 110, 120, 113, 99, 105, 125, 129, 105, 63, 
    105, 109, 91, 76, 94, 118, 127, 106, 79, 63, 14, 0, 0, 0, 0, 0, 0, 4, 73, 122, 146, 165, 176, 169, 168, 173, 161, 133, 110, 103, 100, 68, 
    92, 85, 11, 0, 27, 79, 111, 113, 107, 78, 15, 0, 0, 0, 0, 19, 89, 126, 132, 120, 100, 86, 74, 57, 44, 39, 32, 13, 1, 14, 56, 54, 
    85, 65, 6, 0, 0, 0, 0, 4, 12, 14, 4, 1, 11, 19, 33, 36, 42, 39, 11, 0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 49, 81, 77, 
    24, 0, 3, 4, 0, 0, 0, 0, 0, 16, 40, 61, 76, 89, 80, 48, 11, 0, 6, 22, 27, 17, 18, 35, 58, 77, 95, 119, 129, 117, 100, 76, 
    0, 0, 25, 82, 84, 74, 75, 85, 94, 101, 109, 108, 104, 116, 132, 141, 125, 108, 107, 129, 144, 144, 138, 141, 143, 143, 132, 112, 92, 72, 59, 44, 
    38, 44, 94, 120, 118, 121, 123, 120, 113, 107, 107, 101, 88, 76, 70, 69, 69, 74, 62, 49, 56, 72, 79, 70, 54, 45, 47, 50, 50, 52, 54, 43, 
    146, 185, 184, 158, 145, 134, 126, 124, 121, 113, 101, 91, 74, 53, 34, 26, 29, 40, 46, 41, 42, 51, 55, 51, 47, 47, 55, 60, 59, 57, 53, 43, 
    100, 146, 154, 133, 125, 134, 142, 151, 161, 168, 170, 167, 151, 136, 128, 124, 118, 108, 102, 98, 92, 87, 79, 70, 59, 46, 34, 29, 37, 47, 56, 42, 
    54, 45, 62, 55, 17, 16, 38, 65, 88, 106, 119, 122, 106, 75, 86, 103, 109, 103, 89, 78, 69, 58, 46, 24, 0, 0, 0, 19, 36, 52, 55, 33, 
    85, 76, 74, 86, 62, 14, 6, 21, 43, 58, 66, 64, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 34, 51, 58, 53, 44, 27, 
    80, 99, 99, 112, 133, 113, 84, 73, 69, 70, 72, 72, 70, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 61, 89, 86, 64, 48, 45, 48, 30, 
    49, 54, 80, 92, 110, 122, 110, 98, 88, 80, 75, 75, 93, 129, 108, 22, 0, 0, 0, 0, 34, 72, 105, 114, 93, 66, 53, 52, 53, 54, 58, 42, 
    54, 35, 64, 77, 82, 86, 85, 81, 79, 77, 75, 76, 83, 104, 117, 79, 57, 69, 91, 114, 125, 117, 91, 61, 42, 43, 59, 67, 64, 58, 60, 43, 
    70, 47, 57, 75, 76, 78, 78, 78, 77, 76, 75, 76, 76, 76, 70, 37, 36, 67, 87, 85, 65, 43, 28, 35, 55, 70, 75, 74, 72, 71, 65, 42, 
    87, 70, 62, 72, 76, 76, 77, 77, 76, 75, 75, 76, 76, 82, 96, 92, 84, 90, 76, 48, 24, 23, 43, 65, 77, 74, 65, 66, 69, 70, 68, 44, 
    100, 86, 73, 63, 67, 69, 70, 71, 69, 67, 66, 66, 67, 76, 96, 97, 66, 39, 25, 29, 41, 61, 78, 85, 82, 76, 68, 63, 64, 60, 61, 43, 
    96, 82, 70, 57, 55, 56, 55, 51, 48, 45, 42, 40, 40, 43, 43, 37, 21, 17, 36, 62, 78, 85, 89, 85, 81, 78, 78, 74, 72, 72, 68, 45, 
    144, 119, 107, 97, 90, 87, 85, 80, 76, 75, 75, 75, 77, 83, 90, 99, 109, 127, 144, 155, 164, 164, 163, 163, 163, 168, 172, 180, 188, 198, 204, 172, 
    
    -- channel=20
    0, 171, 168, 168, 168, 168, 168, 168, 168, 168, 168, 169, 169, 169, 170, 170, 170, 168, 167, 167, 170, 172, 170, 168, 167, 168, 169, 168, 168, 168, 169, 189, 
    0, 282, 277, 278, 278, 278, 278, 278, 278, 277, 278, 278, 278, 278, 279, 280, 278, 275, 275, 277, 279, 280, 281, 277, 276, 277, 278, 278, 277, 278, 279, 328, 
    0, 283, 279, 279, 279, 279, 279, 279, 279, 278, 279, 279, 279, 279, 279, 280, 277, 273, 275, 275, 272, 259, 271, 269, 276, 279, 279, 279, 278, 279, 280, 330, 
    0, 283, 279, 279, 279, 279, 279, 279, 279, 278, 278, 279, 279, 278, 278, 279, 276, 275, 277, 277, 256, 233, 257, 264, 276, 280, 279, 279, 279, 279, 280, 330, 
    0, 283, 280, 280, 280, 279, 279, 280, 279, 278, 279, 280, 280, 279, 278, 277, 271, 265, 264, 266, 237, 208, 239, 255, 275, 281, 279, 279, 279, 280, 281, 331, 
    0, 278, 276, 278, 277, 279, 279, 280, 281, 280, 281, 281, 281, 275, 276, 278, 266, 250, 243, 242, 217, 187, 209, 234, 265, 281, 278, 278, 279, 281, 283, 332, 
    0, 272, 277, 278, 276, 278, 280, 280, 282, 283, 283, 282, 278, 258, 270, 282, 266, 241, 233, 233, 218, 199, 196, 213, 252, 281, 279, 279, 280, 281, 283, 334, 
    0, 274, 281, 282, 278, 279, 280, 280, 282, 284, 283, 287, 274, 239, 264, 280, 268, 244, 241, 250, 242, 231, 217, 219, 254, 282, 280, 279, 281, 282, 284, 334, 
    0, 214, 222, 228, 236, 255, 277, 279, 280, 282, 281, 290, 272, 231, 262, 280, 271, 258, 265, 272, 266, 262, 249, 235, 240, 251, 246, 249, 262, 279, 284, 335, 
    0, 178, 175, 177, 186, 226, 272, 273, 275, 278, 277, 286, 275, 247, 266, 280, 279, 270, 278, 282, 272, 261, 244, 230, 220, 210, 199, 197, 229, 273, 283, 335, 
    0, 188, 181, 181, 177, 221, 266, 257, 258, 264, 266, 271, 266, 258, 268, 275, 279, 279, 283, 286, 276, 256, 241, 230, 220, 210, 184, 160, 212, 270, 281, 334, 
    0, 219, 215, 221, 216, 239, 260, 239, 225, 237, 247, 227, 195, 199, 206, 214, 221, 234, 251, 281, 282, 256, 245, 239, 237, 240, 208, 180, 225, 268, 279, 336, 
    0, 212, 205, 214, 225, 238, 249, 233, 218, 243, 257, 200, 128, 129, 133, 141, 158, 184, 226, 276, 283, 266, 264, 261, 255, 263, 240, 221, 243, 249, 261, 330, 
    0, 158, 152, 152, 166, 203, 217, 212, 217, 254, 277, 199, 103, 101, 111, 133, 159, 182, 219, 260, 262, 250, 241, 229, 210, 210, 210, 211, 213, 203, 220, 310, 
    0, 96, 101, 98, 124, 149, 144, 163, 207, 251, 273, 219, 151, 146, 155, 173, 176, 181, 207, 226, 218, 201, 186, 174, 158, 156, 171, 188, 186, 176, 198, 293, 
    0, 36, 58, 109, 156, 142, 113, 131, 191, 231, 254, 240, 213, 207, 219, 236, 220, 208, 211, 211, 205, 193, 172, 165, 159, 157, 165, 184, 192, 186, 194, 268, 
    0, 0, 47, 186, 233, 188, 152, 170, 210, 233, 255, 257, 253, 248, 278, 285, 249, 221, 210, 216, 217, 215, 203, 197, 195, 189, 185, 190, 196, 194, 190, 241, 
    0, 0, 88, 232, 265, 218, 208, 220, 238, 250, 264, 269, 259, 249, 268, 259, 231, 207, 206, 207, 199, 210, 216, 209, 197, 182, 178, 178, 182, 187, 181, 213, 
    0, 59, 161, 244, 247, 235, 241, 247, 254, 257, 257, 255, 243, 233, 237, 219, 213, 210, 216, 209, 186, 194, 205, 198, 179, 164, 163, 157, 151, 151, 152, 188, 
    0, 94, 174, 195, 192, 199, 212, 215, 217, 219, 221, 224, 227, 231, 228, 201, 188, 191, 205, 188, 159, 159, 165, 155, 138, 126, 125, 122, 122, 129, 140, 182, 
    0, 71, 94, 97, 106, 113, 120, 122, 124, 128, 133, 141, 157, 177, 181, 165, 156, 157, 165, 154, 135, 130, 127, 119, 111, 110, 113, 115, 117, 123, 129, 173, 
    0, 16, 2, 17, 43, 51, 47, 40, 35, 34, 40, 49, 70, 97, 111, 109, 110, 115, 119, 111, 101, 95, 90, 90, 94, 103, 112, 117, 113, 109, 119, 168, 
    0, 0, 0, 0, 7, 29, 15, 0, 0, 0, 0, 0, 0, 35, 68, 59, 54, 62, 68, 65, 62, 62, 68, 81, 99, 113, 119, 117, 105, 103, 116, 172, 
    0, 0, 0, 0, 0, 22, 12, 0, 0, 0, 0, 0, 0, 10, 93, 100, 78, 76, 80, 78, 80, 84, 90, 100, 106, 105, 105, 109, 107, 106, 118, 188, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 152, 131, 122, 117, 110, 103, 97, 92, 90, 91, 90, 94, 99, 98, 108, 133, 210, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 162, 152, 137, 126, 114, 101, 85, 74, 73, 75, 72, 71, 85, 102, 122, 151, 229, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 122, 136, 115, 99, 82, 66, 54, 45, 42, 50, 62, 75, 90, 107, 132, 166, 239, 
    0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 82, 54, 38, 27, 24, 22, 28, 42, 62, 81, 89, 95, 109, 140, 173, 245, 
    0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 40, 14, 5, 7, 17, 30, 50, 66, 78, 87, 94, 103, 119, 147, 178, 251, 
    0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 5, 32, 59, 73, 76, 78, 86, 99, 112, 129, 153, 182, 254, 
    0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 20, 32, 51, 72, 76, 75, 79, 88, 104, 120, 135, 158, 186, 255, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 1, 6, 13, 20, 29, 39, 51, 68, 139, 
    
    -- channel=21
    113, 173, 172, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 172, 173, 174, 174, 171, 172, 173, 174, 174, 173, 173, 173, 173, 173, 173, 85, 
    271, 295, 295, 295, 295, 295, 295, 295, 295, 295, 296, 296, 296, 296, 296, 295, 294, 295, 295, 295, 293, 294, 294, 297, 297, 295, 295, 295, 296, 296, 295, 84, 
    273, 296, 295, 295, 295, 295, 295, 295, 295, 296, 296, 296, 296, 296, 297, 296, 295, 295, 294, 288, 287, 298, 295, 301, 298, 295, 295, 295, 296, 297, 296, 84, 
    272, 296, 296, 296, 296, 296, 296, 295, 295, 295, 295, 295, 295, 296, 296, 295, 296, 292, 285, 268, 275, 276, 287, 285, 293, 295, 295, 295, 296, 296, 296, 84, 
    273, 296, 295, 296, 296, 296, 296, 295, 295, 296, 295, 295, 295, 296, 296, 291, 289, 288, 280, 243, 254, 253, 280, 293, 295, 296, 296, 296, 297, 297, 297, 85, 
    270, 297, 296, 295, 297, 298, 298, 296, 295, 295, 296, 295, 292, 298, 296, 285, 274, 263, 249, 217, 227, 251, 278, 302, 303, 297, 298, 298, 299, 299, 298, 85, 
    268, 295, 291, 292, 295, 298, 299, 298, 296, 297, 297, 290, 286, 301, 291, 268, 252, 236, 219, 206, 211, 224, 246, 273, 295, 300, 299, 299, 300, 300, 300, 85, 
    265, 285, 290, 294, 297, 298, 300, 299, 298, 298, 299, 281, 280, 289, 286, 264, 236, 238, 234, 219, 211, 215, 240, 272, 285, 301, 302, 302, 302, 303, 302, 85, 
    232, 293, 295, 304, 318, 318, 302, 299, 298, 298, 301, 270, 278, 284, 284, 273, 265, 262, 258, 256, 248, 249, 262, 293, 298, 297, 302, 313, 317, 306, 303, 87, 
    208, 213, 217, 233, 269, 294, 297, 298, 298, 297, 300, 275, 281, 290, 294, 284, 284, 289, 284, 281, 273, 278, 278, 271, 260, 248, 255, 284, 304, 307, 304, 88, 
    165, 155, 161, 188, 238, 260, 288, 290, 292, 298, 299, 285, 291, 298, 300, 298, 295, 298, 294, 284, 270, 250, 227, 204, 190, 175, 196, 255, 278, 304, 306, 88, 
    172, 213, 213, 235, 279, 282, 273, 267, 283, 286, 264, 261, 280, 284, 286, 291, 297, 306, 312, 278, 252, 228, 218, 217, 206, 190, 209, 253, 287, 302, 307, 89, 
    199, 249, 253, 263, 279, 284, 262, 257, 256, 241, 209, 187, 181, 187, 197, 213, 235, 264, 273, 268, 268, 272, 268, 267, 258, 238, 254, 268, 290, 302, 306, 92, 
    162, 183, 189, 206, 225, 218, 226, 254, 269, 242, 159, 116, 92, 106, 126, 142, 161, 215, 259, 283, 284, 283, 274, 270, 265, 256, 270, 267, 261, 274, 293, 85, 
    93, 106, 126, 147, 153, 191, 229, 253, 279, 251, 166, 128, 113, 125, 140, 170, 225, 271, 280, 266, 247, 232, 212, 204, 204, 207, 207, 196, 199, 228, 251, 67, 
    48, 82, 135, 160, 152, 171, 190, 224, 246, 235, 203, 193, 204, 230, 250, 253, 249, 232, 212, 188, 165, 147, 136, 133, 141, 157, 165, 171, 183, 220, 240, 75, 
    30, 103, 170, 185, 184, 156, 179, 204, 229, 242, 259, 267, 282, 301, 277, 242, 201, 180, 178, 170, 163, 166, 166, 170, 176, 190, 202, 217, 228, 243, 241, 66, 
    31, 137, 207, 229, 215, 219, 237, 250, 270, 284, 294, 288, 293, 285, 257, 235, 227, 232, 216, 226, 236, 234, 228, 223, 220, 224, 231, 227, 210, 194, 185, 39, 
    88, 169, 241, 239, 232, 242, 254, 256, 255, 254, 253, 246, 252, 242, 234, 218, 209, 211, 205, 196, 192, 192, 190, 174, 166, 155, 147, 146, 146, 152, 167, 42, 
    127, 204, 213, 195, 198, 196, 192, 191, 192, 192, 190, 186, 186, 168, 157, 150, 155, 149, 133, 126, 132, 132, 123, 107, 104, 109, 115, 129, 145, 157, 162, 36, 
    111, 125, 118, 119, 118, 119, 121, 125, 129, 134, 141, 145, 146, 132, 125, 130, 141, 136, 115, 109, 109, 104, 96, 91, 93, 104, 114, 121, 128, 139, 161, 40, 
    47, 30, 36, 47, 41, 32, 36, 43, 54, 62, 72, 82, 87, 84, 86, 92, 96, 95, 84, 76, 70, 66, 68, 72, 78, 87, 95, 103, 121, 148, 171, 45, 
    0, 8, 10, 23, 32, 8, 0, 0, 0, 0, 3, 12, 24, 29, 12, 18, 26, 30, 30, 25, 29, 38, 47, 59, 70, 81, 98, 123, 148, 160, 177, 47, 
    1, 5, 24, 40, 41, 36, 16, 0, 0, 0, 0, 0, 14, 40, 31, 4, 5, 2, 2, 7, 17, 34, 51, 71, 95, 127, 147, 142, 140, 163, 200, 55, 
    8, 0, 4, 40, 41, 36, 22, 6, 0, 0, 0, 0, 45, 69, 99, 90, 69, 59, 57, 62, 74, 86, 108, 134, 146, 135, 116, 125, 158, 189, 220, 67, 
    10, 0, 0, 6, 17, 6, 0, 0, 0, 0, 0, 0, 57, 110, 107, 107, 103, 104, 106, 108, 112, 119, 118, 104, 93, 101, 128, 158, 185, 208, 236, 70, 
    28, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 76, 73, 55, 49, 53, 58, 65, 66, 60, 60, 74, 104, 140, 161, 175, 199, 225, 245, 72, 
    51, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 31, 10, 1, 10, 21, 27, 34, 53, 87, 124, 149, 159, 165, 182, 209, 230, 248, 73, 
    65, 25, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 25, 4, 1, 0, 9, 33, 76, 117, 143, 155, 157, 161, 173, 190, 215, 233, 247, 72, 
    70, 37, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 3, 0, 18, 65, 107, 135, 150, 158, 160, 163, 171, 185, 202, 220, 240, 253, 74, 
    71, 55, 35, 24, 18, 15, 14, 10, 7, 5, 7, 11, 13, 28, 44, 44, 56, 93, 126, 147, 152, 152, 156, 161, 171, 183, 192, 208, 227, 244, 255, 76, 
    40, 70, 54, 45, 40, 35, 33, 33, 34, 34, 35, 40, 47, 56, 75, 93, 108, 116, 128, 143, 142, 139, 142, 151, 162, 171, 184, 196, 213, 227, 236, 92, 
    
    -- channel=22
    57, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 55, 55, 55, 54, 55, 54, 55, 54, 54, 55, 54, 55, 54, 54, 54, 54, 55, 188, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 171, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 7, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 7, 13, 10, 2, 5, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 6, 16, 10, 5, 13, 9, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 22, 0, 0, 0, 15, 6, 0, 6, 2, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 172, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 5, 0, 0, 4, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 173, 
    17, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 5, 2, 12, 11, 0, 0, 0, 0, 0, 172, 
    10, 10, 13, 9, 0, 0, 4, 0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 14, 13, 12, 18, 12, 22, 30, 0, 0, 0, 0, 0, 172, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 18, 37, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 3, 7, 0, 0, 15, 1, 0, 0, 0, 0, 169, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 29, 65, 26, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 51, 45, 23, 11, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 144, 
    0, 0, 0, 32, 14, 0, 0, 0, 0, 3, 19, 26, 12, 6, 16, 2, 0, 0, 0, 1, 12, 9, 6, 9, 10, 2, 2, 8, 9, 0, 0, 134, 
    0, 0, 0, 35, 31, 20, 2, 0, 0, 0, 0, 7, 0, 0, 15, 21, 16, 3, 13, 11, 19, 21, 17, 15, 11, 8, 1, 0, 3, 0, 0, 121, 
    0, 0, 0, 4, 18, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 111, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 
    16, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 117, 
    40, 33, 6, 9, 38, 34, 25, 20, 17, 12, 9, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 8, 8, 7, 7, 1, 0, 0, 130, 
    27, 36, 17, 0, 26, 44, 42, 39, 36, 30, 29, 16, 0, 31, 49, 30, 21, 20, 19, 19, 17, 16, 15, 11, 7, 3, 4, 7, 3, 1, 0, 140, 
    36, 32, 27, 3, 3, 25, 33, 36, 37, 34, 33, 27, 0, 0, 56, 53, 43, 39, 37, 30, 24, 16, 9, 6, 1, 0, 6, 10, 3, 0, 0, 144, 
    58, 44, 32, 24, 12, 19, 29, 32, 34, 34, 33, 33, 0, 0, 10, 30, 22, 21, 18, 13, 9, 5, 0, 4, 13, 14, 12, 8, 2, 0, 0, 144, 
    61, 63, 34, 32, 27, 26, 32, 35, 34, 34, 33, 34, 17, 0, 0, 22, 12, 6, 1, 5, 8, 13, 17, 19, 22, 19, 12, 6, 0, 0, 0, 145, 
    52, 72, 39, 34, 32, 30, 33, 35, 35, 34, 33, 33, 27, 0, 3, 32, 21, 15, 17, 27, 30, 29, 26, 21, 17, 17, 12, 5, 0, 0, 0, 147, 
    45, 64, 47, 36, 35, 34, 34, 36, 36, 35, 34, 33, 31, 0, 0, 27, 30, 32, 32, 33, 31, 28, 23, 18, 16, 18, 14, 5, 0, 0, 0, 146, 
    43, 54, 51, 42, 40, 39, 38, 38, 38, 37, 37, 35, 34, 18, 8, 31, 44, 42, 32, 22, 21, 22, 18, 18, 16, 14, 12, 6, 0, 0, 0, 146, 
    41, 51, 50, 47, 44, 43, 42, 42, 41, 40, 41, 40, 39, 34, 28, 35, 36, 31, 24, 16, 21, 21, 20, 19, 15, 11, 8, 5, 0, 0, 0, 146, 
    15, 38, 35, 34, 34, 33, 32, 31, 31, 30, 30, 29, 27, 22, 15, 11, 7, 5, 8, 8, 10, 12, 8, 4, 0, 0, 0, 0, 0, 0, 0, 84, 
    
    -- channel=23
    253, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    346, 1, 5, 5, 5, 5, 5, 5, 5, 5, 6, 5, 5, 5, 5, 4, 3, 4, 6, 3, 6, 9, 6, 5, 4, 5, 4, 5, 6, 6, 4, 0, 
    347, 1, 6, 6, 6, 6, 6, 5, 5, 6, 6, 6, 6, 6, 7, 3, 2, 3, 4, 0, 0, 25, 13, 19, 9, 5, 5, 6, 6, 7, 5, 0, 
    347, 1, 6, 5, 5, 5, 5, 5, 4, 6, 6, 5, 5, 6, 6, 4, 4, 2, 0, 0, 0, 55, 25, 29, 12, 4, 6, 6, 6, 7, 5, 0, 
    347, 1, 6, 5, 5, 5, 5, 5, 4, 7, 6, 4, 4, 6, 7, 0, 0, 1, 2, 0, 0, 62, 40, 34, 15, 4, 5, 5, 6, 6, 5, 0, 
    343, 3, 7, 5, 8, 7, 5, 5, 4, 6, 6, 1, 0, 9, 10, 0, 0, 7, 18, 11, 12, 51, 57, 57, 31, 4, 4, 5, 6, 7, 5, 0, 
    339, 14, 11, 6, 10, 10, 5, 4, 5, 5, 5, 0, 0, 24, 15, 0, 0, 14, 27, 22, 24, 41, 57, 75, 53, 6, 5, 7, 7, 7, 6, 0, 
    339, 22, 16, 9, 13, 11, 6, 4, 5, 4, 5, 0, 0, 39, 22, 0, 0, 19, 26, 13, 21, 27, 41, 55, 49, 9, 7, 9, 9, 8, 6, 0, 
    301, 31, 32, 36, 49, 38, 9, 4, 5, 5, 6, 0, 0, 38, 19, 0, 0, 17, 20, 5, 16, 9, 12, 19, 24, 13, 21, 35, 32, 13, 7, 0, 
    263, 51, 58, 64, 92, 79, 9, 6, 8, 6, 7, 0, 0, 23, 13, 3, 0, 13, 15, 0, 1, 4, 10, 18, 23, 25, 40, 74, 75, 21, 7, 0, 
    261, 35, 50, 50, 75, 71, 1, 6, 15, 11, 7, 2, 4, 17, 16, 12, 12, 13, 12, 0, 0, 15, 21, 25, 27, 14, 36, 93, 88, 25, 8, 0, 
    287, 13, 31, 26, 38, 30, 0, 0, 32, 24, 0, 0, 28, 35, 35, 33, 35, 43, 48, 17, 0, 12, 15, 12, 19, 0, 12, 76, 54, 24, 15, 0, 
    284, 28, 42, 41, 46, 37, 12, 6, 42, 25, 0, 0, 59, 67, 67, 76, 90, 94, 85, 25, 0, 8, 7, 0, 16, 6, 3, 36, 19, 32, 33, 0, 
    238, 56, 57, 83, 91, 60, 41, 38, 44, 10, 0, 0, 57, 78, 92, 91, 82, 76, 60, 9, 0, 0, 5, 2, 21, 28, 25, 24, 21, 57, 66, 0, 
    183, 82, 82, 89, 79, 46, 64, 79, 54, 18, 0, 0, 39, 55, 55, 32, 25, 34, 25, 7, 6, 13, 29, 32, 44, 54, 56, 44, 42, 68, 79, 0, 
    134, 112, 140, 86, 14, 14, 69, 89, 59, 41, 8, 2, 17, 33, 25, 0, 4, 28, 31, 31, 29, 25, 38, 44, 45, 49, 57, 48, 36, 37, 51, 0, 
    114, 152, 194, 73, 0, 2, 46, 55, 35, 35, 16, 6, 7, 31, 11, 0, 0, 20, 37, 29, 31, 22, 25, 27, 26, 29, 32, 30, 27, 27, 38, 0, 
    130, 173, 172, 37, 0, 11, 22, 25, 20, 25, 19, 9, 3, 26, 0, 0, 8, 20, 25, 18, 44, 41, 25, 20, 23, 41, 43, 44, 50, 44, 41, 0, 
    176, 154, 95, 30, 24, 41, 38, 38, 37, 36, 37, 30, 23, 38, 18, 38, 45, 55, 38, 29, 64, 69, 47, 43, 47, 64, 60, 54, 57, 54, 52, 0, 
    204, 114, 58, 53, 62, 67, 63, 63, 64, 64, 65, 60, 56, 53, 37, 52, 58, 65, 41, 34, 60, 63, 52, 49, 53, 64, 62, 58, 64, 65, 58, 0, 
    172, 79, 74, 77, 75, 76, 76, 79, 79, 80, 77, 78, 77, 68, 56, 58, 62, 62, 49, 47, 57, 60, 60, 60, 66, 74, 75, 69, 69, 66, 57, 0, 
    121, 51, 87, 99, 76, 68, 73, 81, 83, 85, 85, 91, 96, 90, 84, 85, 84, 76, 65, 66, 71, 75, 76, 80, 86, 88, 79, 57, 53, 59, 58, 0, 
    98, 25, 62, 101, 78, 39, 40, 51, 56, 64, 71, 84, 112, 106, 74, 83, 92, 90, 80, 84, 89, 91, 93, 96, 89, 67, 47, 36, 42, 55, 57, 0, 
    88, 27, 50, 89, 91, 32, 17, 23, 30, 41, 54, 64, 116, 154, 62, 37, 62, 73, 73, 78, 79, 78, 70, 55, 41, 36, 40, 37, 43, 56, 57, 0, 
    80, 24, 48, 73, 90, 51, 24, 22, 28, 39, 51, 57, 98, 181, 87, 0, 6, 20, 23, 22, 19, 16, 18, 23, 29, 38, 45, 43, 48, 58, 56, 0, 
    90, 0, 33, 59, 70, 60, 41, 34, 36, 44, 51, 53, 82, 161, 117, 0, 0, 0, 0, 0, 0, 0, 18, 36, 37, 38, 45, 47, 51, 58, 51, 0, 
    116, 0, 9, 52, 54, 57, 49, 42, 44, 48, 51, 51, 63, 109, 112, 1, 0, 0, 0, 0, 5, 23, 37, 47, 44, 36, 38, 45, 54, 58, 45, 0, 
    136, 0, 0, 49, 50, 54, 53, 48, 48, 50, 51, 51, 53, 71, 87, 0, 0, 0, 1, 30, 39, 43, 44, 42, 37, 30, 32, 45, 55, 56, 45, 0, 
    144, 0, 0, 42, 48, 51, 52, 50, 50, 50, 50, 52, 51, 58, 77, 26, 0, 21, 47, 58, 49, 39, 30, 29, 31, 34, 34, 42, 52, 53, 45, 0, 
    146, 0, 2, 33, 41, 46, 47, 48, 48, 49, 50, 51, 53, 56, 76, 61, 33, 43, 48, 49, 38, 23, 17, 26, 33, 37, 38, 40, 48, 49, 41, 0, 
    146, 0, 13, 25, 32, 36, 40, 42, 42, 43, 44, 46, 48, 50, 61, 58, 42, 38, 28, 25, 26, 16, 20, 31, 35, 38, 38, 40, 44, 47, 40, 0, 
    109, 2, 22, 28, 30, 33, 35, 38, 38, 38, 39, 38, 37, 37, 41, 43, 37, 34, 28, 26, 31, 26, 31, 37, 37, 39, 40, 43, 45, 47, 44, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 2, 0, 0, 0, 0, 0, 0, 4, 8, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 6, 2, 0, 0, 0, 0, 4, 9, 11, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 9, 0, 0, 0, 4, 11, 15, 13, 13, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 6, 11, 7, 6, 10, 13, 14, 13, 13, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 13, 11, 10, 12, 14, 14, 14, 13, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 11, 11, 12, 12, 12, 13, 13, 13, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 6, 8, 8, 8, 9, 9, 9, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    
    -- channel=25
    75, 116, 115, 115, 115, 115, 115, 115, 115, 116, 116, 116, 116, 116, 116, 114, 114, 114, 116, 119, 120, 120, 117, 114, 113, 114, 116, 115, 116, 116, 116, 58, 
    118, 162, 162, 162, 162, 162, 162, 162, 162, 162, 162, 162, 162, 163, 162, 159, 157, 156, 160, 166, 172, 171, 166, 162, 160, 161, 162, 162, 162, 163, 163, 117, 
    119, 163, 163, 163, 163, 163, 163, 163, 163, 162, 163, 163, 163, 163, 162, 157, 154, 155, 161, 166, 175, 170, 170, 163, 162, 162, 162, 162, 163, 163, 163, 118, 
    119, 163, 163, 163, 163, 163, 163, 162, 162, 162, 162, 162, 162, 162, 162, 159, 158, 162, 171, 172, 176, 172, 170, 166, 163, 162, 163, 163, 163, 164, 163, 118, 
    118, 163, 162, 162, 162, 163, 163, 163, 163, 162, 162, 163, 163, 165, 164, 164, 166, 174, 183, 186, 177, 179, 172, 169, 165, 163, 162, 163, 163, 164, 164, 118, 
    117, 160, 159, 160, 160, 161, 162, 162, 162, 162, 162, 164, 165, 169, 168, 171, 178, 191, 201, 201, 186, 182, 178, 174, 167, 164, 161, 162, 164, 165, 164, 119, 
    121, 167, 166, 165, 164, 162, 162, 161, 161, 161, 162, 159, 165, 166, 169, 179, 188, 203, 214, 214, 202, 192, 186, 184, 175, 170, 165, 166, 168, 168, 166, 119, 
    135, 192, 190, 184, 178, 169, 163, 160, 160, 161, 162, 156, 158, 157, 165, 176, 188, 203, 214, 221, 216, 209, 199, 198, 194, 185, 178, 178, 176, 173, 168, 121, 
    138, 195, 192, 189, 184, 172, 164, 158, 159, 162, 163, 159, 150, 152, 162, 168, 179, 194, 206, 217, 222, 221, 214, 204, 199, 188, 182, 185, 180, 178, 171, 122, 
    134, 189, 184, 183, 184, 171, 162, 154, 156, 162, 166, 169, 156, 160, 165, 173, 177, 187, 200, 207, 216, 214, 211, 200, 190, 178, 175, 182, 181, 182, 174, 123, 
    132, 196, 189, 184, 181, 173, 156, 146, 150, 159, 167, 175, 171, 176, 178, 183, 186, 193, 201, 206, 214, 213, 208, 202, 191, 178, 174, 176, 185, 185, 176, 125, 
    146, 209, 204, 197, 185, 178, 151, 140, 146, 154, 159, 169, 168, 174, 175, 178, 181, 192, 199, 210, 213, 212, 207, 204, 200, 189, 182, 179, 192, 190, 182, 129, 
    151, 204, 200, 195, 191, 179, 161, 155, 162, 170, 164, 167, 165, 170, 167, 167, 174, 187, 197, 207, 204, 205, 203, 199, 200, 194, 181, 186, 190, 190, 188, 134, 
    142, 188, 181, 182, 182, 178, 175, 169, 180, 196, 188, 171, 172, 177, 176, 176, 180, 180, 186, 187, 182, 181, 177, 169, 168, 168, 165, 172, 174, 182, 189, 139, 
    125, 172, 169, 169, 162, 155, 149, 156, 179, 201, 202, 184, 188, 191, 189, 182, 173, 164, 165, 162, 159, 158, 156, 148, 145, 151, 160, 167, 170, 184, 195, 143, 
    95, 149, 158, 155, 156, 126, 108, 124, 155, 180, 191, 187, 191, 193, 191, 185, 174, 168, 169, 172, 174, 173, 172, 168, 166, 171, 179, 186, 189, 192, 202, 142, 
    68, 125, 152, 175, 164, 128, 114, 127, 150, 173, 183, 185, 190, 197, 205, 199, 190, 196, 203, 212, 216, 215, 212, 210, 209, 205, 205, 205, 203, 197, 199, 136, 
    75, 127, 177, 207, 189, 174, 167, 172, 183, 199, 202, 199, 201, 207, 219, 212, 213, 218, 225, 234, 240, 240, 238, 231, 225, 216, 210, 206, 201, 196, 188, 127, 
    103, 176, 225, 235, 232, 237, 237, 238, 241, 244, 242, 237, 231, 235, 238, 235, 238, 234, 238, 240, 245, 249, 246, 236, 226, 218, 210, 200, 191, 184, 178, 119, 
    116, 205, 227, 235, 244, 258, 265, 266, 267, 266, 267, 269, 269, 272, 263, 254, 247, 249, 245, 235, 237, 242, 236, 226, 219, 212, 204, 191, 180, 174, 170, 112, 
    103, 168, 174, 186, 199, 213, 221, 223, 224, 225, 229, 243, 258, 268, 258, 250, 243, 245, 240, 229, 226, 224, 217, 211, 210, 209, 201, 185, 168, 157, 152, 102, 
    63, 100, 107, 121, 133, 142, 143, 140, 139, 137, 144, 167, 197, 221, 226, 224, 224, 222, 218, 213, 209, 205, 200, 195, 196, 196, 182, 161, 142, 130, 129, 89, 
    34, 48, 54, 78, 87, 89, 81, 72, 65, 58, 61, 87, 131, 168, 191, 197, 198, 199, 197, 192, 190, 188, 187, 184, 176, 163, 141, 122, 110, 104, 114, 79, 
    18, 20, 21, 49, 58, 52, 41, 32, 24, 17, 16, 34, 89, 135, 167, 178, 178, 179, 178, 170, 161, 152, 147, 139, 121, 103, 89, 87, 88, 94, 111, 83, 
    0, 4, 3, 14, 23, 13, 6, 4, 3, 0, 0, 6, 42, 90, 103, 101, 93, 92, 88, 81, 69, 58, 52, 50, 48, 51, 57, 69, 85, 101, 121, 93, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 50, 75, 98, 116, 138, 105, 
    6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 38, 62, 83, 107, 130, 151, 112, 
    19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 37, 56, 72, 88, 113, 137, 157, 116, 
    23, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 40, 52, 64, 78, 96, 118, 140, 160, 118, 
    21, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 39, 53, 61, 72, 86, 102, 124, 143, 161, 119, 
    18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 44, 58, 68, 77, 93, 107, 128, 146, 162, 118, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 20, 28, 34, 40, 50, 60, 72, 84, 95, 84, 
    
    -- channel=26
    296, 263, 263, 263, 263, 263, 263, 263, 263, 264, 265, 265, 265, 265, 265, 263, 262, 263, 264, 264, 264, 264, 265, 265, 265, 264, 263, 263, 264, 265, 264, 30, 
    457, 387, 388, 388, 388, 388, 388, 388, 388, 389, 389, 389, 389, 390, 389, 387, 386, 388, 388, 386, 389, 389, 389, 388, 388, 388, 388, 388, 389, 390, 388, 36, 
    460, 389, 390, 390, 390, 390, 390, 389, 389, 390, 390, 390, 390, 391, 390, 387, 385, 385, 383, 357, 366, 372, 381, 390, 390, 389, 389, 389, 391, 391, 390, 37, 
    459, 389, 390, 390, 390, 390, 390, 389, 388, 389, 389, 389, 388, 390, 390, 390, 389, 381, 368, 325, 339, 368, 380, 392, 391, 389, 389, 390, 391, 392, 391, 37, 
    460, 390, 391, 391, 391, 391, 390, 389, 389, 391, 391, 390, 388, 391, 388, 374, 362, 352, 337, 298, 315, 358, 379, 396, 393, 390, 390, 391, 392, 393, 393, 38, 
    452, 385, 386, 387, 390, 392, 392, 390, 390, 392, 393, 386, 381, 390, 385, 355, 329, 319, 308, 275, 284, 319, 357, 393, 396, 392, 391, 391, 393, 394, 395, 38, 
    446, 387, 386, 387, 392, 394, 394, 393, 392, 393, 395, 367, 367, 388, 377, 340, 317, 317, 310, 292, 289, 304, 340, 393, 403, 395, 393, 394, 396, 397, 396, 38, 
    447, 395, 393, 393, 397, 396, 394, 393, 393, 393, 396, 352, 352, 387, 381, 340, 324, 340, 337, 327, 322, 333, 364, 404, 410, 397, 396, 397, 399, 399, 398, 39, 
    357, 310, 316, 341, 384, 397, 393, 391, 391, 393, 394, 350, 352, 390, 384, 361, 357, 371, 368, 362, 360, 352, 352, 361, 355, 344, 356, 387, 401, 401, 399, 39, 
    298, 256, 262, 295, 371, 395, 385, 387, 389, 390, 393, 365, 368, 394, 391, 379, 378, 391, 386, 366, 347, 327, 311, 300, 289, 278, 301, 369, 404, 403, 400, 40, 
    305, 279, 290, 320, 382, 390, 364, 366, 374, 379, 377, 365, 369, 383, 387, 388, 390, 396, 391, 361, 337, 323, 307, 300, 282, 252, 291, 374, 412, 405, 401, 41, 
    339, 306, 320, 342, 380, 371, 325, 324, 354, 345, 285, 266, 276, 288, 298, 312, 328, 366, 389, 367, 343, 339, 330, 329, 316, 284, 318, 386, 405, 403, 402, 42, 
    320, 273, 287, 301, 330, 338, 321, 332, 363, 329, 209, 167, 186, 196, 209, 241, 294, 364, 399, 382, 366, 370, 355, 348, 346, 324, 338, 357, 359, 379, 393, 41, 
    240, 199, 209, 257, 288, 295, 306, 336, 368, 313, 173, 127, 159, 192, 237, 279, 321, 370, 384, 356, 329, 317, 295, 282, 286, 286, 293, 285, 289, 341, 373, 37, 
    148, 147, 187, 228, 232, 237, 278, 324, 347, 307, 221, 201, 235, 266, 282, 285, 300, 318, 305, 276, 249, 234, 225, 221, 233, 251, 260, 258, 275, 333, 360, 35, 
    71, 146, 243, 252, 213, 203, 264, 315, 339, 334, 309, 304, 324, 353, 341, 304, 286, 281, 270, 261, 243, 232, 231, 234, 242, 262, 282, 290, 293, 316, 326, 27, 
    54, 215, 341, 317, 249, 257, 309, 339, 359, 372, 373, 362, 378, 397, 367, 317, 290, 296, 296, 293, 288, 282, 282, 278, 276, 280, 282, 281, 273, 277, 280, 15, 
    109, 286, 384, 324, 286, 309, 332, 344, 357, 370, 371, 355, 358, 350, 310, 278, 279, 285, 271, 268, 283, 282, 269, 249, 240, 244, 246, 249, 248, 244, 242, 10, 
    203, 324, 342, 300, 297, 309, 316, 318, 317, 317, 316, 301, 302, 290, 267, 259, 263, 269, 247, 237, 254, 252, 233, 211, 206, 210, 206, 206, 211, 216, 229, 10, 
    213, 249, 229, 227, 239, 245, 245, 249, 254, 260, 265, 263, 265, 248, 234, 234, 240, 235, 201, 188, 200, 192, 173, 158, 157, 165, 167, 176, 196, 214, 227, 10, 
    129, 109, 106, 113, 118, 121, 126, 132, 141, 150, 161, 174, 183, 176, 171, 177, 186, 180, 155, 143, 142, 137, 131, 129, 136, 151, 163, 176, 192, 208, 226, 10, 
    41, 22, 50, 67, 59, 47, 43, 44, 49, 55, 63, 82, 96, 100, 102, 110, 117, 112, 101, 95, 93, 96, 103, 115, 137, 163, 174, 174, 187, 207, 233, 11, 
    0, 0, 8, 55, 55, 29, 7, 0, 0, 0, 0, 14, 66, 73, 60, 59, 62, 60, 57, 62, 75, 93, 117, 148, 171, 178, 169, 168, 187, 213, 249, 17, 
    0, 0, 0, 40, 52, 22, 0, 0, 0, 0, 0, 0, 77, 147, 126, 108, 107, 104, 104, 111, 125, 145, 158, 159, 153, 158, 166, 171, 195, 233, 277, 25, 
    0, 0, 0, 7, 28, 5, 0, 0, 0, 0, 0, 0, 64, 180, 177, 150, 143, 143, 141, 138, 132, 125, 124, 131, 140, 151, 163, 182, 218, 258, 300, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 161, 169, 123, 109, 107, 100, 90, 82, 84, 98, 116, 130, 151, 180, 208, 243, 281, 313, 29, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 127, 82, 56, 44, 35, 38, 51, 69, 96, 128, 152, 171, 191, 217, 260, 295, 318, 30, 
    67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 67, 15, 0, 0, 10, 42, 73, 105, 135, 161, 175, 181, 196, 228, 268, 299, 321, 30, 
    77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 3, 0, 11, 51, 93, 127, 150, 162, 170, 180, 193, 211, 240, 276, 306, 325, 30, 
    80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 35, 32, 61, 102, 141, 158, 161, 164, 172, 187, 205, 224, 249, 283, 312, 327, 30, 
    86, 12, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 36, 66, 75, 91, 119, 139, 157, 162, 159, 166, 180, 198, 215, 233, 256, 285, 311, 325, 28, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 21, 30, 36, 41, 49, 51, 47, 52, 61, 70, 79, 90, 101, 116, 130, 134, 0, 
    
    -- channel=27
    16, 4, 5, 5, 5, 5, 5, 5, 5, 4, 5, 5, 5, 5, 5, 6, 5, 5, 4, 4, 6, 5, 4, 4, 4, 5, 5, 5, 4, 5, 5, 126, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 155, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 
    9, 33, 33, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 5, 0, 0, 0, 0, 157, 
    0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 18, 17, 14, 14, 4, 0, 0, 0, 0, 157, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 40, 46, 41, 38, 31, 24, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 157, 
    17, 34, 33, 31, 20, 8, 0, 0, 0, 0, 40, 27, 32, 31, 30, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 162, 
    14, 32, 25, 9, 0, 7, 7, 0, 0, 9, 51, 13, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 34, 31, 28, 34, 30, 28, 15, 0, 0, 162, 
    27, 29, 0, 0, 1, 13, 0, 0, 1, 18, 32, 0, 0, 0, 0, 0, 0, 6, 21, 32, 36, 33, 33, 23, 11, 4, 4, 1, 0, 0, 0, 149, 
    46, 20, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 150, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 24, 19, 13, 144, 
    0, 0, 0, 12, 11, 0, 0, 0, 0, 0, 0, 1, 0, 5, 28, 38, 28, 12, 27, 31, 30, 31, 34, 42, 42, 41, 35, 25, 20, 14, 8, 130, 
    0, 0, 0, 15, 16, 16, 15, 14, 15, 16, 18, 23, 12, 24, 24, 25, 20, 21, 27, 14, 8, 22, 28, 31, 20, 15, 15, 11, 11, 13, 10, 122, 
    16, 30, 38, 36, 28, 26, 25, 23, 20, 16, 12, 11, 8, 16, 7, 1, 0, 11, 26, 18, 14, 23, 30, 32, 26, 24, 28, 25, 18, 9, 4, 120, 
    40, 62, 67, 64, 64, 65, 64, 62, 59, 59, 55, 51, 51, 55, 52, 45, 38, 41, 50, 50, 48, 47, 45, 42, 38, 33, 25, 14, 7, 6, 3, 121, 
    40, 39, 35, 34, 36, 44, 50, 54, 54, 57, 59, 56, 58, 62, 64, 61, 59, 60, 60, 56, 52, 50, 44, 36, 26, 12, 5, 5, 6, 5, 0, 117, 
    67, 52, 37, 36, 36, 32, 36, 45, 49, 52, 52, 43, 28, 25, 28, 35, 42, 51, 49, 44, 37, 27, 15, 1, 0, 0, 14, 22, 10, 0, 0, 119, 
    70, 70, 51, 41, 61, 64, 62, 61, 63, 63, 62, 52, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 34, 30, 15, 2, 0, 0, 124, 
    53, 60, 58, 40, 55, 73, 76, 76, 73, 66, 63, 54, 7, 27, 46, 21, 10, 6, 6, 10, 16, 30, 45, 50, 36, 16, 11, 8, 0, 0, 0, 133, 
    55, 57, 61, 52, 48, 60, 68, 70, 70, 66, 63, 61, 15, 3, 52, 61, 57, 56, 58, 61, 64, 59, 43, 27, 14, 6, 5, 2, 0, 0, 0, 137, 
    57, 65, 61, 61, 55, 58, 65, 67, 67, 64, 63, 63, 43, 2, 19, 39, 44, 51, 58, 61, 50, 31, 12, 6, 10, 11, 7, 0, 0, 0, 0, 137, 
    54, 77, 62, 62, 59, 59, 63, 64, 64, 63, 62, 62, 57, 20, 20, 52, 66, 67, 52, 32, 14, 5, 5, 7, 11, 11, 4, 0, 0, 0, 0, 139, 
    57, 80, 63, 58, 57, 57, 60, 62, 62, 61, 61, 60, 58, 28, 25, 53, 49, 33, 17, 9, 4, 6, 11, 13, 12, 8, 1, 0, 0, 0, 0, 140, 
    55, 66, 57, 49, 49, 51, 52, 53, 52, 52, 51, 49, 47, 22, 7, 21, 21, 13, 6, 5, 11, 18, 18, 14, 9, 6, 3, 0, 0, 0, 0, 140, 
    48, 49, 44, 42, 42, 42, 40, 38, 37, 36, 35, 32, 31, 16, 2, 9, 16, 12, 7, 5, 16, 22, 17, 12, 5, 1, 0, 0, 0, 0, 0, 142, 
    85, 92, 85, 84, 82, 81, 80, 80, 80, 80, 81, 81, 82, 81, 79, 82, 87, 93, 95, 89, 94, 97, 95, 95, 94, 96, 97, 99, 98, 102, 109, 201, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 14, 18, 4, 0, 0, 0, 5, 10, 11, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 14, 23, 21, 0, 0, 0, 9, 20, 27, 29, 27, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 17, 24, 30, 15, 0, 0, 5, 18, 29, 32, 31, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 19, 30, 35, 32, 17, 10, 13, 22, 30, 35, 33, 37, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 4, 30, 37, 37, 32, 26, 26, 31, 35, 36, 35, 40, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 36, 37, 35, 32, 32, 35, 36, 37, 36, 42, 59, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 34, 34, 34, 34, 35, 36, 36, 36, 35, 40, 55, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 28, 29, 29, 31, 33, 33, 32, 31, 30, 32, 40, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 16, 19, 20, 21, 22, 22, 21, 20, 19, 18, 21, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 9, 19, 21, 23, 24, 25, 25, 25, 25, 24, 24, 24, 24, 21, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    276, 548, 544, 545, 545, 545, 545, 545, 545, 546, 547, 548, 548, 548, 548, 546, 545, 545, 545, 546, 546, 548, 546, 545, 545, 546, 546, 545, 546, 547, 547, 311, 
    516, 876, 871, 872, 872, 872, 872, 872, 872, 872, 873, 874, 874, 875, 875, 873, 871, 870, 871, 871, 874, 872, 874, 871, 872, 872, 872, 872, 873, 874, 874, 516, 
    520, 881, 876, 876, 876, 876, 876, 875, 875, 875, 875, 876, 876, 877, 877, 874, 870, 866, 865, 842, 846, 828, 855, 859, 872, 876, 875, 874, 876, 877, 878, 518, 
    518, 880, 875, 876, 876, 876, 876, 875, 874, 874, 874, 874, 874, 875, 875, 875, 872, 864, 852, 802, 793, 779, 827, 851, 870, 876, 875, 875, 876, 878, 878, 519, 
    520, 882, 877, 878, 878, 878, 878, 876, 875, 875, 877, 877, 875, 876, 873, 862, 844, 823, 799, 744, 725, 732, 798, 843, 870, 878, 877, 877, 879, 881, 882, 521, 
    512, 870, 867, 872, 874, 877, 879, 878, 878, 879, 881, 876, 871, 871, 865, 843, 803, 761, 728, 680, 659, 672, 741, 810, 857, 880, 878, 879, 881, 883, 885, 524, 
    504, 858, 864, 869, 871, 877, 881, 881, 882, 883, 886, 859, 857, 847, 850, 825, 770, 729, 703, 679, 657, 656, 700, 780, 844, 883, 880, 881, 884, 887, 888, 525, 
    501, 862, 871, 875, 876, 880, 882, 883, 884, 886, 888, 845, 834, 819, 845, 819, 776, 752, 742, 737, 713, 710, 737, 803, 858, 886, 883, 884, 888, 889, 891, 527, 
    414, 720, 735, 764, 811, 848, 878, 880, 881, 883, 885, 840, 822, 813, 846, 837, 820, 815, 816, 817, 801, 791, 784, 794, 801, 801, 806, 835, 864, 889, 894, 528, 
    337, 589, 593, 634, 724, 799, 864, 867, 870, 877, 880, 852, 838, 838, 861, 861, 855, 860, 864, 851, 825, 790, 752, 719, 690, 667, 678, 744, 817, 884, 894, 529, 
    312, 580, 582, 628, 715, 792, 836, 828, 836, 849, 853, 843, 836, 842, 858, 867, 872, 880, 879, 852, 813, 758, 712, 681, 642, 602, 616, 686, 804, 881, 894, 530, 
    366, 668, 673, 710, 767, 803, 784, 761, 770, 776, 745, 704, 662, 675, 693, 717, 742, 793, 830, 839, 808, 763, 735, 724, 700, 665, 669, 721, 824, 876, 889, 530, 
    376, 653, 660, 688, 731, 750, 742, 738, 753, 749, 653, 539, 445, 456, 479, 522, 595, 703, 798, 852, 844, 829, 810, 801, 783, 755, 750, 764, 803, 826, 854, 518, 
    277, 483, 491, 541, 591, 650, 680, 706, 759, 747, 602, 437, 335, 363, 418, 495, 590, 698, 787, 823, 802, 773, 733, 704, 682, 675, 683, 679, 683, 720, 776, 485, 
    150, 311, 357, 413, 471, 531, 572, 650, 741, 739, 635, 520, 468, 496, 536, 586, 631, 676, 703, 691, 647, 605, 564, 539, 532, 552, 573, 584, 598, 659, 723, 458, 
    48, 226, 347, 452, 504, 471, 500, 594, 700, 734, 720, 687, 682, 713, 733, 730, 686, 651, 630, 607, 568, 537, 507, 497, 502, 526, 558, 591, 615, 653, 688, 418, 
    9, 233, 449, 627, 623, 553, 575, 645, 726, 776, 809, 808, 827, 841, 839, 779, 692, 652, 630, 632, 621, 609, 599, 595, 594, 596, 608, 623, 624, 631, 633, 364, 
    49, 303, 582, 721, 703, 664, 688, 724, 768, 805, 828, 819, 818, 798, 774, 707, 663, 643, 632, 637, 635, 641, 640, 613, 589, 574, 574, 576, 571, 565, 556, 313, 
    157, 460, 656, 710, 702, 701, 718, 727, 736, 741, 740, 721, 711, 688, 669, 630, 620, 617, 605, 586, 572, 580, 572, 534, 503, 483, 473, 467, 466, 476, 494, 279, 
    204, 462, 542, 553, 562, 576, 588, 592, 598, 605, 614, 614, 615, 596, 570, 538, 535, 534, 506, 468, 450, 448, 430, 396, 373, 367, 371, 383, 409, 442, 476, 271, 
    133, 278, 292, 298, 312, 322, 334, 343, 355, 370, 391, 415, 438, 444, 436, 424, 428, 427, 405, 376, 354, 339, 325, 312, 311, 327, 346, 367, 393, 428, 465, 266, 
    8, 84, 90, 118, 144, 143, 133, 128, 134, 146, 166, 197, 233, 263, 275, 281, 290, 290, 281, 261, 244, 237, 237, 249, 275, 316, 348, 368, 391, 420, 466, 266, 
    0, 0, 0, 33, 75, 80, 42, 6, 0, 0, 0, 6, 77, 126, 158, 147, 145, 148, 148, 145, 154, 177, 212, 261, 310, 353, 373, 381, 392, 423, 484, 279, 
    0, 0, 0, 7, 62, 79, 39, 0, 0, 0, 0, 0, 26, 143, 234, 234, 206, 197, 198, 205, 226, 258, 295, 327, 348, 363, 371, 378, 401, 448, 524, 314, 
    0, 0, 0, 0, 14, 40, 16, 0, 0, 0, 0, 0, 5, 185, 332, 374, 343, 326, 319, 318, 313, 310, 314, 324, 332, 337, 346, 375, 425, 489, 575, 351, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152, 312, 384, 368, 350, 335, 312, 288, 269, 262, 265, 276, 302, 346, 402, 467, 540, 620, 376, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 174, 257, 264, 240, 214, 188, 172, 169, 188, 228, 282, 336, 381, 429, 499, 575, 648, 390, 
    24, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 92, 89, 61, 62, 83, 122, 169, 229, 294, 346, 377, 406, 449, 518, 594, 660, 398, 
    43, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 27, 23, 61, 128, 205, 269, 320, 352, 374, 396, 428, 476, 539, 610, 671, 405, 
    46, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 52, 84, 147, 226, 293, 339, 359, 367, 384, 414, 453, 500, 560, 625, 681, 411, 
    47, 106, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 50, 93, 147, 202, 253, 298, 330, 352, 360, 373, 401, 434, 475, 520, 575, 634, 684, 410, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 68, 97, 117, 135, 149, 158, 163, 175, 194, 215, 242, 271, 306, 342, 372, 221, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    94, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 136, 134, 133, 135, 138, 139, 138, 137, 137, 138, 138, 137, 27, 
    98, 142, 141, 141, 141, 141, 141, 141, 141, 141, 142, 142, 142, 142, 142, 142, 142, 141, 137, 123, 125, 122, 131, 138, 141, 142, 141, 141, 141, 141, 141, 29, 
    96, 140, 140, 140, 140, 140, 140, 139, 140, 140, 140, 140, 140, 140, 140, 143, 145, 141, 133, 119, 144, 136, 149, 139, 138, 140, 140, 141, 141, 141, 141, 28, 
    99, 142, 141, 141, 141, 141, 141, 140, 140, 141, 140, 140, 140, 140, 139, 132, 122, 115, 114, 110, 127, 119, 122, 131, 136, 140, 141, 140, 140, 141, 141, 28, 
    91, 136, 136, 137, 139, 141, 142, 142, 141, 140, 140, 137, 136, 139, 136, 131, 132, 128, 117, 98, 85, 93, 107, 125, 136, 140, 141, 141, 141, 141, 141, 28, 
    100, 143, 140, 142, 141, 141, 142, 142, 140, 140, 140, 129, 135, 141, 133, 128, 134, 132, 117, 106, 110, 126, 140, 140, 135, 142, 144, 144, 143, 143, 143, 28, 
    104, 134, 133, 138, 141, 143, 143, 142, 139, 139, 141, 129, 151, 141, 138, 131, 113, 102, 97, 97, 96, 107, 125, 141, 135, 141, 143, 142, 143, 143, 143, 29, 
    33, 69, 75, 91, 121, 139, 143, 142, 141, 140, 141, 130, 147, 140, 138, 125, 123, 112, 98, 96, 83, 72, 67, 85, 102, 105, 111, 128, 141, 144, 144, 30, 
    121, 148, 147, 148, 151, 135, 139, 141, 141, 141, 143, 136, 135, 137, 140, 130, 124, 122, 118, 105, 88, 86, 99, 113, 124, 126, 133, 144, 139, 143, 145, 30, 
    93, 122, 125, 142, 149, 126, 136, 135, 131, 134, 136, 128, 120, 126, 132, 136, 132, 131, 130, 124, 140, 152, 153, 146, 132, 119, 135, 149, 138, 143, 147, 31, 
    1, 29, 27, 44, 79, 117, 127, 126, 133, 124, 97, 83, 78, 78, 80, 84, 90, 109, 125, 129, 133, 116, 95, 86, 71, 73, 100, 102, 126, 139, 144, 31, 
    29, 51, 49, 50, 70, 104, 124, 158, 158, 124, 112, 136, 123, 118, 119, 127, 144, 162, 142, 124, 107, 97, 88, 85, 80, 73, 75, 78, 108, 126, 131, 25, 
    72, 90, 98, 117, 125, 104, 97, 99, 98, 93, 84, 96, 85, 101, 130, 146, 138, 117, 102, 101, 92, 87, 80, 85, 85, 71, 70, 92, 110, 121, 126, 25, 
    38, 49, 83, 99, 66, 82, 102, 88, 97, 102, 80, 58, 54, 57, 29, 0, 6, 39, 78, 96, 104, 113, 116, 122, 129, 136, 137, 133, 132, 141, 129, 31, 
    2, 23, 49, 43, 70, 114, 122, 129, 147, 135, 101, 62, 51, 49, 51, 83, 115, 133, 140, 140, 133, 129, 121, 107, 103, 110, 107, 94, 82, 85, 87, 18, 
    28, 76, 56, 51, 111, 110, 114, 122, 129, 115, 104, 93, 101, 112, 124, 145, 135, 120, 99, 80, 59, 52, 46, 40, 40, 39, 33, 30, 35, 58, 91, 25, 
    41, 50, 35, 64, 56, 42, 48, 56, 68, 84, 99, 108, 124, 105, 83, 48, 33, 36, 13, 13, 19, 15, 13, 16, 23, 31, 56, 86, 99, 101, 95, 17, 
    25, 3, 61, 83, 69, 60, 67, 75, 79, 83, 85, 87, 93, 91, 103, 95, 87, 71, 81, 101, 95, 80, 82, 85, 94, 96, 92, 84, 71, 58, 60, 8, 
    0, 0, 46, 51, 57, 64, 64, 62, 64, 69, 75, 76, 72, 71, 73, 72, 69, 57, 48, 40, 36, 41, 40, 31, 23, 20, 17, 22, 36, 52, 64, 3, 
    27, 40, 29, 17, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 22, 41, 50, 52, 60, 3, 
    48, 51, 50, 46, 41, 28, 22, 19, 21, 22, 20, 17, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 30, 36, 35, 39, 54, 74, 16, 
    0, 0, 3, 0, 3, 8, 6, 4, 7, 13, 16, 20, 27, 24, 17, 10, 4, 0, 0, 0, 0, 5, 15, 26, 27, 16, 6, 19, 53, 74, 90, 13, 
    0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 23, 22, 16, 13, 14, 16, 11, 0, 0, 0, 33, 66, 74, 83, 99, 14, 
    24, 15, 15, 31, 23, 7, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 83, 81, 66, 76, 92, 102, 18, 
    4, 14, 7, 13, 28, 24, 14, 9, 3, 0, 0, 0, 26, 51, 6, 0, 0, 0, 0, 0, 0, 22, 63, 89, 88, 70, 64, 78, 95, 102, 113, 26, 
    4, 12, 6, 0, 4, 4, 0, 0, 0, 0, 0, 0, 14, 59, 55, 40, 38, 33, 35, 47, 69, 83, 81, 64, 52, 62, 83, 93, 98, 106, 118, 28, 
    17, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 24, 12, 0, 0, 2, 33, 58, 64, 57, 52, 58, 76, 92, 97, 99, 105, 112, 119, 26, 
    20, 26, 19, 7, 5, 5, 3, 0, 0, 0, 0, 0, 4, 19, 12, 0, 30, 55, 60, 48, 45, 54, 70, 85, 94, 95, 97, 104, 114, 122, 122, 27, 
    35, 51, 30, 23, 19, 17, 16, 14, 12, 11, 11, 13, 17, 34, 51, 53, 51, 44, 44, 55, 67, 79, 93, 98, 96, 94, 96, 104, 110, 117, 120, 28, 
    44, 63, 48, 40, 34, 33, 34, 32, 29, 28, 28, 30, 32, 43, 55, 48, 38, 48, 71, 88, 91, 95, 100, 100, 100, 105, 107, 108, 112, 116, 119, 28, 
    0, 11, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 17, 20, 19, 15, 12, 10, 9, 9, 9, 11, 11, 7, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 13, 26, 12, 0, 0, 3, 9, 15, 21, 21, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 16, 30, 35, 9, 2, 11, 23, 29, 37, 39, 39, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    53, 27, 31, 41, 42, 23, 24, 28, 34, 40, 45, 43, 52, 26, 0, 0, 0, 0, 1, 4, 6, 6, 4, 3, 5, 0, 0, 0, 0, 0, 0, 0, 
    37, 29, 40, 43, 59, 51, 42, 42, 41, 43, 49, 47, 48, 87, 51, 44, 65, 66, 63, 57, 48, 41, 34, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 8, 37, 50, 55, 60, 54, 50, 48, 48, 51, 51, 52, 103, 133, 133, 142, 130, 109, 83, 65, 46, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 29, 50, 52, 54, 52, 49, 49, 50, 52, 50, 58, 104, 158, 165, 162, 144, 115, 79, 47, 25, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 19, 47, 48, 48, 46, 45, 48, 50, 50, 48, 54, 89, 135, 134, 120, 94, 63, 39, 22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 11, 40, 42, 41, 40, 41, 44, 45, 45, 43, 44, 60, 92, 88, 60, 41, 30, 27, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 13, 28, 32, 32, 31, 32, 32, 34, 32, 29, 30, 35, 50, 44, 28, 25, 21, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 7, 28, 34, 36, 36, 36, 37, 37, 38, 37, 33, 33, 35, 38, 38, 36, 32, 28, 25, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    94, 52, 46, 24, 38, 36, 30, 30, 31, 33, 37, 29, 37, 36, 34, 47, 28, 36, 34, 35, 37, 33, 37, 37, 42, 34, 34, 41, 38, 34, 39, 189, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 303, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 306, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 307, 
    0, 3, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 305, 
    0, 6, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 303, 
    0, 10, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 3, 0, 0, 0, 0, 89, 3, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 303, 
    0, 14, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 6, 0, 0, 18, 81, 54, 5, 21, 0, 0, 0, 0, 0, 0, 0, 0, 299, 
    0, 21, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 48, 63, 61, 55, 46, 42, 75, 35, 0, 0, 0, 4, 18, 0, 6, 281, 
    0, 33, 50, 13, 8, 30, 6, 0, 7, 16, 6, 0, 14, 5, 0, 41, 57, 42, 29, 33, 26, 27, 70, 38, 23, 0, 4, 56, 42, 0, 20, 248, 
    9, 48, 60, 45, 48, 47, 26, 24, 33, 41, 24, 23, 32, 12, 7, 38, 44, 30, 31, 47, 44, 31, 61, 14, 35, 3, 0, 112, 59, 25, 35, 209, 
    29, 48, 57, 15, 31, 50, 51, 37, 29, 47, 37, 16, 11, 4, 10, 29, 34, 28, 36, 49, 54, 0, 2, 14, 56, 43, 0, 83, 98, 37, 51, 191, 
    19, 27, 45, 0, 18, 58, 60, 14, 0, 17, 37, 4, 0, 10, 26, 29, 33, 31, 24, 36, 36, 0, 0, 0, 38, 104, 0, 5, 138, 45, 47, 190, 
    3, 15, 56, 31, 35, 53, 40, 4, 0, 2, 28, 26, 4, 15, 32, 32, 32, 26, 10, 21, 7, 0, 0, 0, 4, 84, 47, 0, 131, 84, 38, 187, 
    12, 27, 55, 46, 56, 56, 25, 10, 2, 0, 0, 6, 0, 0, 8, 0, 0, 3, 0, 0, 0, 0, 0, 6, 10, 34, 98, 23, 94, 124, 57, 171, 
    14, 15, 35, 32, 16, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 1, 8, 11, 12, 22, 16, 103, 107, 79, 104, 67, 164, 
    0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 69, 36, 18, 8, 0, 15, 8, 71, 84, 22, 48, 75, 190, 
    0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 13, 0, 23, 64, 26, 0, 5, 0, 9, 10, 35, 19, 0, 18, 73, 238, 
    0, 0, 25, 39, 20, 0, 0, 0, 0, 0, 0, 0, 5, 9, 6, 5, 7, 0, 0, 29, 8, 0, 9, 11, 9, 10, 16, 17, 24, 25, 18, 246, 
    20, 41, 19, 0, 0, 0, 0, 0, 1, 8, 2, 0, 0, 0, 0, 0, 1, 0, 0, 10, 5, 0, 0, 11, 7, 17, 37, 51, 63, 45, 0, 217, 
    17, 20, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 10, 27, 0, 2, 8, 1, 0, 0, 22, 38, 49, 65, 73, 74, 62, 16, 178, 
    0, 2, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 4, 36, 47, 57, 66, 0, 0, 0, 4, 16, 30, 52, 63, 62, 67, 74, 62, 71, 85, 163, 
    0, 0, 0, 0, 0, 0, 0, 17, 16, 14, 0, 0, 8, 62, 84, 59, 51, 0, 0, 16, 38, 48, 55, 59, 56, 70, 79, 70, 66, 94, 117, 153, 
    0, 0, 1, 0, 5, 43, 44, 45, 44, 42, 0, 0, 0, 38, 59, 42, 40, 26, 30, 47, 49, 49, 55, 73, 75, 80, 79, 77, 89, 105, 106, 144, 
    0, 0, 10, 3, 6, 61, 63, 35, 23, 17, 0, 0, 15, 46, 56, 55, 55, 46, 42, 46, 56, 64, 74, 76, 77, 77, 78, 89, 98, 98, 98, 144, 
    0, 0, 5, 2, 5, 39, 47, 28, 27, 32, 34, 49, 62, 64, 54, 45, 44, 42, 50, 68, 79, 80, 72, 54, 73, 93, 90, 87, 93, 94, 92, 145, 
    0, 7, 25, 36, 43, 52, 56, 56, 62, 68, 66, 59, 52, 47, 47, 54, 66, 72, 74, 75, 71, 72, 78, 68, 81, 97, 93, 86, 89, 89, 87, 142, 
    44, 61, 67, 71, 74, 74, 69, 60, 61, 59, 59, 61, 64, 64, 67, 78, 80, 67, 69, 64, 72, 85, 86, 81, 88, 93, 88, 86, 87, 87, 92, 142, 
    78, 90, 86, 79, 77, 79, 74, 65, 68, 74, 76, 78, 78, 74, 72, 80, 63, 34, 74, 89, 84, 86, 85, 87, 91, 89, 86, 86, 83, 93, 104, 142, 
    82, 97, 92, 88, 84, 85, 85, 82, 80, 80, 79, 72, 69, 67, 72, 85, 64, 33, 88, 102, 85, 84, 89, 92, 89, 86, 83, 85, 85, 111, 123, 139, 
    84, 97, 93, 88, 85, 84, 82, 79, 75, 70, 72, 71, 73, 75, 80, 95, 72, 40, 96, 101, 85, 90, 93, 90, 88, 87, 83, 82, 99, 127, 134, 132, 
    73, 84, 82, 78, 76, 76, 74, 73, 74, 75, 79, 83, 87, 94, 101, 114, 86, 39, 85, 101, 90, 89, 87, 88, 88, 89, 77, 86, 123, 136, 125, 128, 
    
    -- channel=33
    94, 205, 188, 188, 202, 234, 247, 251, 256, 261, 261, 265, 267, 278, 283, 276, 276, 272, 282, 287, 289, 288, 285, 288, 286, 284, 283, 286, 285, 282, 285, 166, 
    105, 295, 276, 269, 283, 331, 348, 353, 357, 365, 368, 369, 372, 384, 393, 386, 391, 379, 394, 400, 393, 389, 384, 402, 400, 402, 398, 401, 403, 399, 397, 269, 
    108, 303, 282, 277, 287, 336, 352, 358, 363, 370, 372, 369, 368, 378, 393, 385, 394, 382, 391, 380, 361, 345, 358, 398, 402, 405, 399, 402, 403, 398, 396, 269, 
    112, 308, 288, 281, 286, 338, 353, 360, 360, 366, 375, 365, 363, 367, 383, 374, 388, 380, 380, 358, 330, 324, 347, 394, 398, 403, 396, 398, 400, 395, 396, 268, 
    116, 313, 287, 281, 283, 338, 350, 360, 363, 368, 376, 361, 360, 353, 365, 348, 357, 363, 358, 332, 296, 269, 321, 390, 394, 398, 388, 385, 394, 390, 389, 262, 
    116, 312, 280, 275, 270, 333, 346, 361, 362, 365, 371, 355, 357, 345, 343, 313, 319, 338, 332, 298, 271, 251, 285, 341, 357, 377, 377, 371, 381, 378, 380, 254, 
    117, 313, 276, 271, 268, 332, 345, 354, 359, 359, 363, 349, 354, 341, 336, 309, 304, 277, 241, 197, 163, 142, 163, 206, 238, 290, 344, 357, 363, 357, 356, 239, 
    102, 277, 247, 248, 243, 286, 296, 305, 323, 328, 333, 327, 331, 326, 324, 290, 256, 211, 179, 169, 159, 136, 138, 159, 179, 231, 277, 295, 300, 301, 302, 205, 
    61, 208, 193, 189, 178, 201, 213, 230, 245, 254, 261, 262, 265, 267, 268, 250, 225, 184, 161, 140, 128, 119, 109, 115, 129, 200, 236, 247, 234, 221, 222, 144, 
    17, 136, 134, 132, 129, 155, 167, 163, 180, 187, 195, 193, 198, 208, 213, 205, 187, 152, 139, 125, 116, 114, 115, 150, 150, 167, 197, 213, 223, 177, 167, 105, 
    0, 97, 106, 125, 134, 148, 135, 125, 135, 154, 166, 164, 174, 191, 191, 182, 168, 153, 142, 138, 132, 144, 169, 214, 215, 219, 226, 203, 212, 157, 125, 76, 
    0, 97, 116, 130, 123, 129, 122, 120, 150, 175, 180, 178, 173, 170, 165, 156, 144, 134, 139, 143, 147, 170, 209, 258, 263, 241, 237, 218, 211, 161, 106, 61, 
    10, 111, 116, 119, 112, 119, 109, 121, 137, 159, 175, 172, 170, 170, 170, 163, 155, 157, 163, 166, 180, 208, 238, 284, 293, 263, 237, 212, 186, 153, 90, 41, 
    13, 112, 118, 121, 104, 108, 113, 121, 151, 191, 207, 209, 207, 210, 209, 206, 204, 212, 214, 214, 224, 238, 253, 279, 283, 274, 232, 187, 135, 103, 63, 32, 
    21, 142, 145, 149, 144, 153, 170, 188, 208, 223, 236, 246, 246, 244, 243, 244, 239, 238, 239, 223, 214, 205, 226, 250, 260, 261, 223, 176, 116, 104, 82, 37, 
    32, 162, 166, 176, 187, 192, 199, 212, 227, 244, 253, 261, 266, 269, 262, 250, 240, 236, 231, 208, 193, 185, 216, 245, 249, 254, 224, 200, 172, 174, 168, 80, 
    36, 172, 182, 185, 172, 177, 201, 234, 253, 262, 266, 266, 260, 252, 242, 230, 222, 227, 233, 225, 214, 207, 225, 239, 241, 245, 226, 225, 216, 198, 184, 100, 
    31, 164, 146, 138, 150, 179, 216, 236, 245, 245, 235, 230, 229, 233, 239, 242, 241, 242, 239, 235, 233, 221, 232, 241, 240, 240, 231, 227, 207, 195, 207, 116, 
    15, 127, 125, 155, 192, 207, 213, 223, 218, 214, 217, 229, 240, 248, 252, 251, 241, 236, 236, 246, 245, 239, 244, 245, 239, 227, 206, 181, 156, 149, 160, 95, 
    23, 159, 167, 176, 184, 193, 200, 205, 210, 219, 238, 242, 242, 239, 230, 213, 194, 195, 203, 237, 248, 243, 242, 230, 208, 178, 152, 135, 115, 102, 112, 60, 
    37, 170, 169, 179, 197, 209, 216, 209, 208, 209, 217, 224, 231, 220, 195, 151, 123, 146, 175, 221, 237, 220, 201, 178, 157, 141, 126, 101, 84, 76, 62, 11, 
    31, 160, 190, 199, 202, 200, 191, 175, 161, 155, 172, 191, 219, 210, 174, 135, 117, 138, 159, 186, 182, 165, 152, 140, 130, 104, 79, 68, 61, 44, 19, 0, 
    19, 150, 180, 188, 188, 174, 154, 123, 114, 115, 143, 175, 209, 207, 180, 142, 116, 115, 114, 134, 144, 136, 125, 103, 78, 60, 56, 47, 34, 15, 5, 0, 
    14, 130, 167, 183, 185, 169, 149, 123, 118, 127, 146, 162, 171, 156, 131, 105, 95, 105, 111, 122, 114, 96, 75, 66, 65, 57, 41, 23, 12, 6, 0, 0, 
    13, 125, 159, 174, 171, 158, 141, 117, 105, 101, 100, 93, 100, 105, 107, 107, 106, 103, 93, 82, 69, 61, 61, 63, 50, 33, 20, 7, 2, 0, 0, 0, 
    0, 94, 108, 113, 105, 97, 89, 72, 68, 73, 79, 86, 91, 89, 84, 79, 71, 63, 55, 55, 61, 55, 41, 33, 27, 22, 9, 0, 0, 0, 0, 0, 
    0, 39, 44, 49, 49, 51, 51, 52, 58, 66, 66, 61, 56, 50, 48, 49, 49, 52, 59, 66, 48, 29, 21, 19, 13, 10, 2, 0, 0, 0, 0, 0, 
    0, 11, 10, 14, 16, 19, 21, 24, 28, 31, 31, 31, 32, 37, 43, 44, 44, 52, 56, 52, 32, 17, 15, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 5, 8, 13, 21, 27, 33, 36, 36, 34, 29, 29, 40, 47, 50, 22, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 10, 13, 18, 24, 26, 26, 24, 24, 23, 15, 13, 23, 34, 45, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 5, 7, 9, 11, 13, 16, 17, 15, 11, 3, 0, 0, 0, 0, 12, 29, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    137, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    137, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    135, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 
    126, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 12, 0, 0, 0, 0, 0, 0, 
    115, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 50, 28, 0, 0, 0, 13, 0, 0, 
    102, 0, 0, 0, 10, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 0, 7, 0, 0, 
    91, 0, 0, 1, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    92, 3, 0, 0, 0, 0, 0, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 14, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    97, 0, 0, 0, 0, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    98, 0, 0, 0, 0, 0, 0, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    97, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    121, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    119, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    111, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 
    57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 0, 0, 0, 
    47, 0, 2, 9, 8, 2, 3, 7, 4, 0, 0, 0, 0, 0, 0, 0, 4, 32, 0, 0, 0, 0, 0, 1, 1, 3, 5, 4, 4, 0, 0, 0, 
    47, 3, 6, 12, 11, 5, 3, 5, 3, 0, 0, 0, 0, 0, 0, 0, 10, 42, 0, 0, 0, 1, 0, 3, 5, 5, 7, 7, 0, 0, 0, 2, 
    50, 5, 7, 9, 7, 3, 3, 4, 2, 0, 0, 0, 0, 0, 0, 0, 20, 55, 0, 0, 0, 3, 3, 6, 6, 5, 10, 5, 0, 0, 6, 14, 
    36, 11, 11, 12, 11, 9, 9, 9, 9, 7, 5, 4, 4, 3, 2, 1, 25, 47, 3, 0, 4, 9, 11, 11, 10, 9, 15, 9, 0, 0, 19, 20, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 12, 14, 26, 30, 21, 20, 29, 30, 25, 29, 36, 43, 41, 42, 38, 40, 47, 46, 45, 49, 61, 57, 51, 42, 43, 45, 41, 41, 47, 40, 20, 
    57, 31, 30, 36, 41, 36, 33, 37, 43, 41, 41, 49, 55, 54, 57, 50, 46, 52, 52, 62, 96, 99, 77, 56, 48, 47, 50, 46, 45, 50, 52, 28, 
    61, 33, 37, 46, 49, 48, 43, 44, 51, 48, 48, 53, 58, 58, 62, 58, 48, 54, 56, 72, 101, 113, 88, 58, 49, 50, 56, 54, 52, 51, 55, 32, 
    65, 35, 38, 53, 59, 55, 53, 54, 62, 61, 56, 56, 60, 60, 71, 84, 69, 68, 61, 70, 92, 78, 65, 62, 57, 57, 67, 66, 60, 55, 53, 36, 
    75, 46, 46, 61, 68, 63, 60, 55, 60, 66, 63, 60, 60, 63, 78, 104, 102, 92, 87, 70, 85, 108, 99, 91, 77, 66, 78, 79, 69, 66, 63, 44, 
    79, 51, 52, 58, 69, 60, 65, 58, 62, 70, 69, 62, 63, 69, 62, 70, 99, 119, 147, 126, 87, 128, 181, 202, 177, 108, 80, 81, 79, 84, 78, 53, 
    97, 64, 55, 54, 72, 70, 83, 77, 77, 83, 76, 70, 72, 79, 57, 46, 70, 121, 153, 157, 130, 125, 164, 211, 230, 195, 126, 104, 105, 117, 112, 82, 
    139, 120, 101, 94, 124, 143, 142, 143, 133, 133, 122, 113, 111, 111, 102, 93, 83, 74, 49, 27, 16, 13, 20, 28, 55, 123, 144, 146, 158, 161, 168, 125, 
    143, 144, 131, 129, 137, 151, 156, 161, 166, 161, 159, 155, 150, 137, 128, 115, 89, 57, 42, 41, 45, 56, 43, 25, 28, 41, 79, 73, 113, 138, 161, 130, 
    102, 103, 92, 86, 68, 62, 79, 106, 103, 93, 102, 111, 97, 81, 80, 81, 70, 63, 60, 60, 60, 58, 26, 0, 23, 64, 98, 44, 13, 64, 84, 82, 
    62, 42, 38, 43, 37, 27, 45, 49, 40, 21, 15, 36, 35, 23, 29, 42, 46, 44, 47, 38, 28, 13, 0, 0, 0, 0, 68, 102, 30, 52, 67, 57, 
    39, 24, 29, 49, 76, 76, 52, 39, 34, 23, 11, 10, 30, 37, 35, 42, 49, 51, 51, 41, 28, 23, 38, 52, 43, 14, 26, 101, 71, 52, 88, 62, 
    42, 37, 47, 55, 66, 68, 62, 48, 52, 61, 48, 21, 9, 12, 6, 0, 0, 0, 0, 5, 9, 25, 51, 75, 86, 69, 45, 88, 127, 70, 86, 85, 
    37, 28, 29, 25, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 61, 80, 80, 77, 71, 59, 76, 126, 93, 57, 63, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 9, 15, 39, 48, 49, 68, 102, 119, 109, 98, 76, 65, 52, 27, 11, 0, 0, 16, 
    41, 9, 14, 21, 25, 36, 23, 9, 13, 20, 26, 34, 45, 56, 65, 68, 71, 78, 68, 62, 60, 66, 62, 67, 66, 63, 50, 10, 0, 0, 0, 0, 
    45, 39, 56, 72, 75, 66, 63, 35, 24, 34, 48, 60, 69, 77, 79, 70, 53, 50, 41, 13, 0, 9, 27, 41, 57, 60, 56, 51, 72, 98, 82, 23, 
    56, 60, 73, 54, 24, 7, 19, 47, 56, 62, 68, 65, 54, 41, 32, 26, 27, 37, 51, 42, 29, 34, 43, 42, 48, 59, 71, 88, 112, 133, 121, 72, 
    43, 22, 14, 0, 0, 0, 15, 43, 61, 48, 37, 25, 21, 24, 37, 56, 79, 88, 73, 61, 52, 50, 55, 59, 73, 96, 106, 117, 125, 117, 121, 116, 
    23, 0, 0, 7, 36, 47, 45, 33, 34, 31, 27, 37, 48, 63, 98, 126, 137, 137, 106, 67, 60, 65, 79, 99, 111, 118, 118, 108, 91, 82, 103, 123, 
    69, 31, 20, 24, 29, 32, 43, 51, 57, 79, 92, 79, 64, 65, 80, 101, 98, 89, 98, 94, 92, 105, 114, 116, 114, 101, 95, 91, 83, 86, 92, 96, 
    77, 69, 41, 36, 38, 49, 81, 103, 104, 104, 105, 88, 58, 40, 23, 17, 21, 37, 78, 112, 121, 115, 107, 102, 99, 97, 95, 90, 96, 98, 92, 76, 
    58, 63, 58, 54, 50, 52, 63, 76, 66, 50, 42, 60, 73, 72, 57, 46, 52, 69, 84, 93, 92, 96, 97, 94, 86, 82, 78, 79, 81, 84, 74, 65, 
    53, 49, 48, 44, 45, 38, 18, 15, 23, 30, 50, 79, 110, 121, 113, 99, 85, 74, 71, 78, 89, 96, 99, 86, 62, 55, 68, 74, 69, 65, 62, 59, 
    67, 69, 74, 76, 86, 88, 76, 66, 77, 96, 111, 120, 110, 88, 68, 65, 74, 85, 94, 96, 93, 83, 73, 72, 79, 76, 72, 71, 70, 64, 58, 57, 
    93, 111, 131, 134, 134, 132, 124, 112, 99, 91, 80, 72, 72, 75, 80, 91, 101, 93, 76, 75, 71, 71, 74, 78, 84, 80, 71, 65, 64, 61, 58, 64, 
    87, 104, 111, 112, 104, 94, 86, 81, 78, 78, 84, 89, 92, 91, 91, 92, 86, 60, 37, 47, 73, 77, 71, 72, 71, 71, 66, 63, 62, 58, 68, 75, 
    70, 66, 68, 72, 76, 79, 80, 84, 91, 93, 91, 88, 80, 71, 64, 67, 70, 68, 61, 68, 74, 70, 68, 66, 68, 66, 63, 61, 60, 67, 82, 88, 
    77, 71, 69, 70, 70, 72, 72, 71, 70, 66, 60, 57, 60, 66, 73, 80, 86, 87, 79, 73, 69, 69, 65, 67, 65, 66, 67, 63, 63, 83, 90, 92, 
    72, 69, 62, 60, 58, 57, 56, 55, 56, 61, 68, 74, 81, 87, 93, 99, 101, 98, 82, 68, 67, 65, 64, 61, 63, 67, 68, 65, 76, 87, 89, 80, 
    93, 89, 89, 90, 92, 95, 98, 100, 103, 107, 109, 110, 111, 112, 112, 112, 110, 119, 124, 103, 94, 92, 89, 90, 90, 91, 91, 97, 94, 91, 87, 80, 
    
    -- channel=36
    0, 164, 154, 127, 128, 164, 176, 177, 179, 183, 185, 179, 170, 177, 179, 182, 177, 165, 177, 183, 186, 182, 174, 175, 180, 179, 171, 179, 185, 175, 174, 204, 
    0, 268, 256, 211, 205, 262, 283, 283, 282, 290, 297, 285, 274, 285, 287, 294, 291, 270, 284, 292, 298, 288, 271, 283, 294, 295, 280, 293, 303, 286, 283, 353, 
    0, 265, 255, 209, 198, 255, 280, 278, 270, 281, 292, 277, 266, 278, 284, 288, 293, 271, 279, 285, 286, 252, 242, 277, 295, 296, 278, 294, 305, 282, 280, 354, 
    0, 261, 250, 204, 191, 246, 271, 273, 256, 267, 284, 268, 257, 268, 274, 274, 288, 269, 273, 288, 272, 214, 218, 273, 292, 295, 274, 289, 302, 278, 279, 351, 
    0, 258, 244, 199, 181, 236, 258, 264, 245, 256, 276, 260, 249, 260, 264, 250, 267, 255, 260, 286, 246, 160, 195, 270, 288, 291, 266, 275, 289, 271, 277, 344, 
    0, 251, 240, 193, 167, 225, 244, 256, 235, 245, 265, 250, 241, 253, 255, 220, 230, 226, 242, 277, 219, 133, 176, 237, 257, 276, 255, 257, 270, 257, 272, 331, 
    0, 247, 238, 189, 161, 222, 239, 248, 231, 240, 253, 239, 234, 246, 248, 210, 211, 193, 191, 213, 155, 83, 114, 147, 163, 210, 230, 239, 253, 238, 246, 305, 
    0, 226, 219, 174, 147, 204, 216, 218, 217, 227, 230, 221, 223, 231, 227, 207, 205, 181, 162, 161, 140, 101, 106, 102, 84, 133, 180, 204, 216, 194, 196, 268, 
    0, 180, 177, 141, 118, 161, 164, 163, 175, 185, 184, 180, 191, 194, 187, 199, 208, 173, 146, 124, 114, 103, 102, 82, 47, 92, 140, 176, 178, 135, 137, 211, 
    0, 120, 123, 105, 91, 119, 119, 109, 127, 135, 137, 136, 150, 155, 156, 178, 181, 144, 125, 119, 113, 106, 108, 100, 84, 95, 108, 154, 165, 103, 104, 157, 
    0, 78, 89, 84, 83, 108, 100, 84, 88, 108, 119, 111, 124, 142, 154, 167, 156, 131, 119, 118, 115, 104, 108, 127, 140, 141, 107, 138, 169, 105, 87, 119, 
    0, 69, 90, 80, 76, 114, 110, 83, 89, 126, 142, 126, 125, 145, 161, 157, 136, 115, 108, 113, 117, 99, 105, 161, 188, 179, 113, 120, 184, 128, 75, 106, 
    0, 82, 105, 89, 80, 117, 106, 83, 89, 131, 157, 148, 143, 160, 174, 161, 140, 127, 120, 126, 133, 116, 126, 183, 211, 218, 151, 107, 169, 140, 56, 89, 
    0, 100, 119, 104, 88, 105, 98, 91, 114, 151, 175, 184, 177, 184, 192, 181, 166, 163, 158, 160, 159, 142, 155, 185, 195, 216, 185, 117, 127, 114, 33, 69, 
    0, 129, 134, 127, 120, 130, 133, 141, 161, 177, 192, 205, 207, 208, 213, 206, 195, 197, 193, 183, 164, 138, 151, 168, 177, 189, 193, 151, 95, 84, 41, 59, 
    0, 151, 149, 152, 152, 163, 173, 182, 197, 212, 219, 223, 226, 229, 230, 221, 206, 204, 203, 192, 159, 123, 133, 152, 169, 179, 190, 181, 106, 91, 102, 95, 
    0, 166, 166, 171, 161, 162, 187, 215, 231, 238, 239, 235, 228, 221, 214, 207, 191, 183, 193, 198, 160, 118, 130, 147, 165, 177, 182, 179, 124, 117, 142, 139, 
    0, 168, 159, 154, 152, 153, 180, 212, 227, 231, 225, 217, 208, 201, 194, 191, 183, 171, 177, 192, 169, 136, 152, 165, 173, 177, 175, 167, 136, 134, 155, 169, 
    0, 155, 144, 146, 157, 165, 178, 199, 210, 209, 203, 201, 198, 195, 190, 184, 181, 170, 168, 191, 186, 169, 180, 185, 181, 172, 161, 146, 124, 108, 98, 149, 
    0, 167, 145, 143, 159, 178, 192, 195, 195, 190, 190, 189, 188, 189, 188, 178, 168, 154, 145, 177, 189, 183, 185, 184, 172, 148, 133, 119, 99, 73, 55, 110, 
    0, 165, 151, 162, 184, 196, 203, 198, 181, 171, 177, 181, 186, 190, 184, 153, 125, 104, 106, 159, 182, 175, 167, 159, 142, 118, 103, 85, 64, 50, 40, 60, 
    0, 154, 178, 187, 188, 185, 183, 177, 156, 146, 156, 160, 178, 193, 179, 131, 97, 72, 77, 135, 152, 143, 135, 124, 108, 81, 64, 51, 37, 34, 32, 24, 
    0, 126, 168, 178, 176, 176, 167, 140, 124, 119, 120, 127, 164, 191, 178, 122, 86, 66, 65, 105, 119, 109, 100, 86, 66, 50, 45, 31, 22, 20, 15, 0, 
    0, 97, 150, 165, 167, 177, 165, 120, 104, 109, 104, 110, 145, 160, 143, 105, 84, 79, 78, 90, 86, 72, 59, 56, 50, 43, 33, 18, 13, 7, 0, 0, 
    0, 92, 136, 154, 155, 165, 152, 107, 90, 90, 84, 85, 106, 114, 107, 91, 81, 76, 70, 66, 59, 48, 41, 38, 32, 34, 24, 9, 4, 0, 0, 0, 
    0, 78, 105, 119, 115, 118, 111, 85, 74, 74, 70, 73, 77, 73, 67, 58, 53, 51, 48, 48, 47, 37, 25, 16, 20, 32, 16, 0, 0, 0, 0, 0, 
    0, 46, 61, 69, 65, 64, 61, 55, 53, 51, 44, 38, 36, 36, 39, 39, 37, 37, 39, 45, 33, 21, 18, 12, 11, 15, 3, 0, 0, 0, 0, 0, 
    0, 18, 19, 17, 13, 14, 13, 11, 14, 18, 18, 18, 20, 23, 29, 30, 22, 15, 30, 47, 29, 15, 13, 7, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 13, 13, 15, 17, 17, 5, 0, 31, 60, 23, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 5, 4, 7, 12, 12, 0, 0, 25, 56, 13, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 5, 40, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    80, 119, 109, 115, 129, 142, 147, 151, 156, 158, 156, 161, 167, 171, 173, 168, 169, 169, 176, 179, 176, 177, 180, 182, 175, 174, 177, 175, 173, 176, 177, 87, 
    209, 212, 195, 220, 245, 259, 263, 266, 275, 278, 270, 281, 287, 296, 301, 288, 290, 296, 303, 303, 297, 302, 311, 308, 299, 297, 305, 302, 294, 299, 306, 86, 
    219, 220, 199, 226, 254, 268, 270, 274, 281, 284, 275, 281, 290, 295, 300, 291, 291, 295, 304, 296, 278, 299, 310, 311, 298, 300, 309, 303, 294, 305, 308, 88, 
    222, 224, 201, 228, 259, 272, 269, 272, 288, 289, 277, 279, 286, 285, 297, 291, 292, 295, 300, 274, 251, 267, 285, 308, 300, 300, 310, 304, 293, 307, 304, 86, 
    225, 228, 205, 229, 258, 276, 274, 276, 290, 288, 278, 276, 284, 277, 287, 281, 291, 298, 293, 230, 213, 272, 292, 306, 299, 298, 308, 303, 293, 304, 304, 86, 
    228, 232, 201, 226, 255, 276, 273, 273, 292, 288, 278, 274, 285, 266, 268, 266, 271, 286, 272, 219, 200, 234, 276, 309, 305, 299, 302, 295, 292, 301, 300, 85, 
    228, 229, 190, 220, 243, 266, 262, 271, 288, 283, 275, 270, 281, 260, 255, 243, 224, 249, 230, 179, 192, 217, 238, 266, 286, 303, 301, 284, 283, 293, 295, 84, 
    214, 227, 188, 214, 230, 257, 259, 271, 279, 274, 272, 267, 274, 253, 245, 231, 215, 204, 182, 122, 111, 139, 139, 156, 189, 220, 272, 272, 269, 281, 280, 80, 
    188, 202, 172, 197, 211, 222, 231, 233, 248, 247, 250, 251, 250, 245, 249, 218, 181, 135, 111, 99, 94, 97, 85, 120, 169, 182, 218, 216, 207, 237, 231, 71, 
    143, 150, 134, 152, 165, 151, 159, 176, 185, 189, 193, 202, 196, 200, 203, 174, 145, 129, 123, 120, 116, 116, 108, 112, 128, 186, 206, 189, 141, 166, 164, 39, 
    99, 102, 101, 108, 113, 107, 115, 124, 142, 137, 138, 149, 148, 150, 151, 141, 129, 122, 125, 118, 109, 114, 124, 155, 146, 152, 172, 175, 146, 122, 130, 21, 
    80, 91, 85, 108, 125, 120, 109, 117, 124, 122, 128, 124, 134, 145, 140, 127, 123, 129, 127, 121, 113, 144, 167, 193, 188, 170, 202, 167, 155, 111, 118, 22, 
    85, 99, 104, 132, 124, 108, 103, 114, 142, 153, 150, 154, 153, 147, 135, 124, 120, 122, 127, 130, 133, 181, 217, 231, 215, 177, 212, 179, 142, 112, 97, 27, 
    96, 114, 103, 112, 108, 93, 92, 128, 150, 150, 144, 149, 152, 139, 129, 128, 131, 133, 144, 142, 156, 197, 224, 240, 229, 179, 179, 177, 106, 116, 94, 13, 
    104, 108, 100, 101, 96, 96, 99, 112, 132, 158, 163, 162, 169, 172, 164, 162, 168, 179, 182, 175, 185, 215, 224, 230, 220, 198, 151, 149, 89, 73, 76, 3, 
    105, 120, 122, 127, 122, 125, 150, 165, 179, 188, 198, 204, 206, 206, 199, 203, 201, 203, 201, 182, 179, 190, 197, 200, 203, 200, 145, 118, 109, 82, 73, 2, 
    118, 144, 141, 144, 166, 178, 193, 197, 196, 200, 204, 209, 213, 217, 211, 203, 202, 196, 183, 149, 146, 154, 176, 193, 194, 196, 160, 133, 149, 153, 154, 44, 
    122, 131, 147, 158, 160, 166, 168, 190, 198, 198, 202, 206, 207, 202, 195, 180, 177, 178, 177, 158, 160, 178, 190, 198, 190, 192, 173, 171, 197, 193, 161, 47, 
    114, 130, 129, 121, 119, 147, 175, 183, 191, 195, 190, 183, 178, 177, 181, 182, 185, 202, 200, 185, 190, 197, 195, 196, 188, 183, 173, 173, 167, 161, 169, 44, 
    109, 100, 94, 117, 157, 176, 187, 179, 171, 173, 168, 176, 186, 192, 195, 198, 189, 201, 214, 200, 196, 197, 193, 185, 181, 176, 164, 137, 116, 121, 135, 21, 
    103, 125, 150, 166, 173, 170, 161, 158, 157, 169, 192, 204, 206, 193, 170, 163, 155, 167, 190, 197, 190, 188, 185, 173, 165, 141, 112, 98, 90, 83, 100, 16, 
    125, 163, 160, 160, 160, 162, 157, 154, 169, 172, 185, 198, 193, 165, 134, 105, 92, 129, 157, 177, 186, 176, 162, 136, 110, 104, 95, 83, 78, 68, 62, 0, 
    125, 148, 160, 164, 165, 156, 144, 136, 137, 134, 146, 164, 176, 146, 110, 90, 86, 129, 160, 161, 148, 131, 112, 99, 99, 90, 73, 67, 65, 51, 25, 0, 
    116, 145, 156, 157, 157, 134, 111, 95, 93, 95, 126, 147, 159, 144, 125, 124, 121, 127, 125, 114, 105, 102, 106, 94, 76, 53, 50, 53, 44, 27, 17, 0, 
    106, 138, 144, 146, 146, 118, 102, 94, 99, 109, 135, 157, 152, 128, 108, 99, 95, 97, 99, 102, 102, 95, 75, 63, 63, 56, 48, 38, 31, 24, 19, 0, 
    94, 127, 136, 143, 142, 121, 109, 112, 115, 117, 115, 101, 87, 78, 80, 91, 95, 95, 96, 90, 70, 58, 59, 71, 62, 46, 37, 30, 26, 24, 21, 0, 
    75, 104, 103, 104, 99, 89, 81, 78, 75, 72, 73, 76, 80, 84, 87, 89, 85, 79, 66, 50, 57, 60, 54, 55, 45, 34, 28, 28, 29, 27, 24, 0, 
    49, 52, 48, 47, 48, 51, 52, 56, 62, 70, 74, 77, 78, 73, 65, 59, 57, 65, 68, 63, 57, 48, 38, 35, 34, 28, 28, 28, 29, 30, 20, 0, 
    26, 28, 27, 32, 38, 42, 47, 55, 58, 59, 57, 52, 50, 52, 54, 51, 60, 85, 77, 56, 45, 35, 31, 32, 27, 27, 29, 30, 32, 25, 13, 0, 
    24, 27, 26, 29, 34, 36, 38, 40, 43, 43, 45, 51, 56, 59, 55, 47, 55, 84, 68, 43, 34, 30, 28, 22, 23, 26, 29, 32, 31, 11, 5, 0, 
    24, 23, 26, 28, 32, 35, 38, 41, 47, 52, 53, 54, 51, 49, 43, 32, 41, 68, 56, 38, 31, 26, 20, 20, 22, 24, 29, 31, 18, 1, 0, 0, 
    10, 28, 31, 35, 38, 40, 41, 43, 45, 47, 45, 42, 38, 31, 23, 10, 14, 36, 33, 37, 27, 21, 21, 20, 21, 21, 26, 26, 14, 0, 0, 0, 
    
    -- channel=38
    45, 60, 52, 23, 38, 48, 48, 47, 49, 52, 56, 45, 52, 53, 52, 64, 46, 50, 51, 55, 59, 53, 54, 55, 62, 51, 50, 60, 57, 49, 55, 195, 
    0, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 1, 0, 0, 0, 5, 0, 0, 3, 1, 0, 0, 174, 
    0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 4, 0, 0, 0, 0, 6, 0, 0, 3, 3, 0, 0, 173, 
    0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 2, 0, 5, 0, 0, 0, 21, 0, 0, 0, 0, 7, 0, 0, 3, 2, 0, 0, 173, 
    0, 11, 16, 0, 0, 0, 3, 0, 0, 4, 5, 0, 0, 10, 0, 0, 0, 0, 10, 35, 0, 0, 0, 0, 8, 0, 0, 5, 0, 0, 0, 170, 
    0, 11, 24, 0, 0, 0, 5, 1, 0, 7, 6, 2, 0, 19, 0, 0, 0, 0, 12, 49, 0, 0, 0, 0, 4, 6, 0, 6, 0, 0, 4, 167, 
    0, 14, 29, 0, 0, 0, 3, 2, 0, 10, 6, 4, 0, 21, 11, 5, 0, 0, 0, 28, 3, 0, 0, 0, 0, 4, 0, 8, 4, 0, 8, 165, 
    0, 13, 27, 0, 0, 0, 0, 0, 0, 9, 5, 2, 2, 9, 9, 27, 14, 7, 0, 9, 10, 0, 3, 0, 0, 0, 0, 7, 9, 0, 6, 150, 
    0, 3, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 22, 22, 16, 16, 19, 14, 14, 30, 6, 0, 0, 0, 7, 3, 0, 0, 124, 
    0, 0, 7, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 11, 8, 12, 7, 0, 16, 3, 21, 0, 0, 45, 10, 0, 0, 103, 
    0, 5, 12, 0, 15, 20, 11, 0, 0, 15, 3, 0, 3, 1, 2, 9, 11, 5, 5, 12, 13, 0, 10, 16, 24, 9, 0, 65, 42, 14, 9, 91, 
    0, 10, 20, 0, 13, 26, 16, 0, 3, 19, 20, 4, 2, 8, 6, 6, 8, 3, 4, 15, 15, 0, 0, 15, 41, 54, 0, 26, 73, 9, 14, 84, 
    0, 7, 19, 0, 2, 11, 9, 0, 0, 2, 19, 9, 0, 2, 5, 3, 2, 4, 2, 13, 7, 0, 0, 0, 20, 60, 9, 0, 81, 16, 4, 81, 
    0, 0, 13, 7, 9, 6, 0, 0, 0, 0, 1, 7, 0, 0, 8, 5, 10, 12, 7, 11, 1, 0, 0, 0, 5, 29, 48, 0, 46, 38, 3, 72, 
    2, 0, 13, 11, 11, 18, 3, 0, 0, 0, 0, 1, 2, 2, 8, 0, 3, 9, 10, 12, 0, 0, 0, 5, 11, 11, 57, 24, 12, 43, 20, 69, 
    4, 0, 6, 13, 1, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 0, 0, 0, 1, 12, 9, 46, 45, 18, 51, 43, 82, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 8, 27, 5, 0, 6, 0, 10, 8, 27, 28, 15, 35, 50, 114, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 6, 27, 15, 5, 12, 8, 8, 7, 15, 13, 1, 2, 16, 129, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 10, 0, 0, 12, 9, 1, 7, 13, 7, 10, 11, 10, 9, 0, 0, 119, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 5, 4, 1, 2, 12, 7, 7, 12, 15, 14, 9, 0, 83, 
    0, 5, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 8, 1, 0, 0, 0, 0, 5, 2, 4, 2, 7, 11, 12, 17, 18, 15, 24, 10, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 18, 6, 11, 0, 0, 0, 2, 3, 6, 11, 14, 19, 20, 17, 19, 26, 26, 48, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 1, 24, 31, 19, 16, 0, 0, 0, 5, 9, 12, 18, 14, 19, 20, 18, 19, 23, 29, 51, 
    0, 0, 0, 0, 0, 19, 8, 0, 2, 3, 0, 0, 0, 9, 15, 13, 12, 7, 4, 9, 13, 12, 14, 18, 21, 22, 19, 22, 22, 26, 28, 49, 
    0, 0, 0, 0, 0, 18, 20, 8, 7, 4, 0, 0, 0, 3, 5, 5, 10, 11, 11, 13, 17, 16, 17, 13, 25, 26, 20, 20, 24, 25, 26, 51, 
    0, 0, 0, 0, 0, 2, 8, 4, 3, 3, 0, 1, 5, 10, 11, 11, 13, 10, 8, 16, 18, 21, 21, 10, 19, 25, 22, 20, 23, 24, 26, 52, 
    0, 0, 0, 0, 0, 1, 2, 2, 6, 11, 14, 14, 13, 11, 10, 13, 15, 10, 18, 20, 19, 20, 19, 17, 18, 23, 23, 21, 23, 23, 26, 47, 
    7, 10, 7, 7, 9, 14, 12, 9, 11, 14, 14, 14, 14, 13, 14, 19, 14, 8, 30, 25, 17, 20, 22, 21, 21, 22, 22, 22, 22, 27, 28, 41, 
    19, 23, 20, 17, 16, 18, 17, 14, 13, 15, 17, 16, 17, 18, 19, 24, 12, 0, 29, 29, 19, 23, 22, 22, 22, 21, 21, 22, 22, 34, 28, 38, 
    18, 26, 23, 22, 21, 21, 21, 20, 19, 19, 21, 20, 19, 18, 19, 25, 11, 0, 30, 29, 21, 22, 22, 22, 21, 21, 19, 20, 29, 35, 31, 37, 
    20, 25, 24, 23, 23, 23, 22, 22, 22, 20, 21, 21, 21, 22, 21, 26, 11, 0, 29, 30, 22, 21, 22, 23, 22, 22, 17, 24, 34, 33, 34, 39, 
    17, 23, 23, 22, 21, 20, 19, 18, 18, 19, 19, 20, 21, 23, 23, 25, 18, 3, 17, 27, 22, 22, 21, 23, 24, 23, 18, 23, 32, 35, 34, 37, 
    
    -- channel=39
    238, 11, 0, 25, 64, 30, 12, 11, 10, 6, 0, 0, 6, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    318, 33, 9, 47, 104, 64, 37, 33, 43, 35, 18, 17, 35, 20, 17, 10, 0, 28, 20, 16, 0, 0, 22, 14, 4, 0, 22, 15, 0, 8, 25, 0, 
    319, 29, 5, 40, 99, 59, 33, 22, 39, 33, 7, 11, 32, 20, 14, 17, 0, 22, 18, 0, 0, 13, 53, 19, 4, 0, 22, 14, 0, 6, 30, 0, 
    319, 22, 0, 34, 93, 53, 29, 10, 34, 31, 0, 5, 25, 19, 8, 28, 0, 17, 16, 0, 0, 36, 81, 24, 6, 0, 19, 13, 0, 7, 26, 0, 
    319, 16, 0, 26, 93, 46, 29, 4, 27, 29, 0, 0, 21, 17, 0, 31, 2, 21, 22, 0, 0, 76, 96, 26, 11, 0, 15, 15, 0, 12, 20, 0, 
    315, 10, 0, 15, 96, 40, 30, 0, 21, 21, 0, 2, 18, 11, 0, 24, 20, 23, 35, 0, 0, 88, 90, 36, 33, 0, 7, 17, 0, 18, 18, 0, 
    311, 1, 0, 8, 99, 30, 20, 0, 14, 8, 0, 5, 11, 6, 0, 8, 2, 1, 16, 0, 0, 73, 72, 48, 86, 51, 19, 17, 0, 13, 21, 0, 
    293, 1, 0, 4, 85, 19, 10, 12, 11, 0, 0, 7, 5, 0, 0, 0, 0, 1, 24, 27, 31, 67, 62, 45, 98, 101, 50, 22, 0, 7, 30, 0, 
    256, 18, 3, 12, 66, 31, 21, 38, 25, 9, 2, 16, 10, 1, 15, 12, 0, 5, 28, 39, 39, 48, 41, 40, 90, 85, 67, 16, 0, 13, 46, 0, 
    208, 45, 30, 36, 67, 45, 38, 55, 44, 33, 25, 34, 32, 28, 43, 23, 0, 31, 47, 45, 40, 61, 61, 40, 64, 37, 80, 20, 0, 22, 49, 0, 
    174, 68, 53, 55, 73, 38, 26, 50, 64, 53, 30, 50, 57, 51, 52, 37, 29, 46, 54, 48, 42, 66, 94, 59, 33, 0, 55, 56, 0, 3, 38, 0, 
    170, 82, 52, 47, 80, 32, 21, 55, 82, 63, 25, 38, 62, 59, 45, 36, 42, 49, 55, 50, 42, 65, 103, 51, 6, 0, 0, 86, 0, 0, 45, 0, 
    178, 81, 49, 39, 72, 38, 35, 63, 86, 68, 41, 35, 57, 65, 47, 45, 54, 55, 61, 61, 48, 71, 91, 36, 8, 0, 0, 55, 0, 0, 51, 11, 
    190, 74, 49, 39, 61, 42, 59, 86, 91, 75, 61, 47, 54, 59, 46, 48, 57, 52, 51, 52, 41, 61, 59, 23, 15, 0, 0, 0, 18, 0, 46, 23, 
    206, 64, 56, 44, 60, 58, 62, 75, 74, 65, 58, 49, 49, 51, 43, 37, 52, 43, 32, 21, 19, 49, 44, 25, 16, 1, 0, 0, 19, 12, 32, 12, 
    220, 56, 66, 50, 50, 62, 55, 61, 62, 57, 52, 49, 50, 46, 41, 32, 43, 48, 33, 8, 8, 59, 50, 36, 23, 8, 0, 0, 23, 45, 0, 0, 
    235, 64, 65, 46, 46, 75, 85, 67, 60, 57, 51, 46, 45, 45, 43, 38, 41, 59, 46, 9, 3, 57, 48, 31, 27, 15, 13, 0, 19, 34, 0, 0, 
    232, 56, 58, 58, 69, 84, 95, 75, 56, 48, 49, 50, 53, 53, 49, 47, 37, 44, 49, 14, 5, 45, 38, 20, 27, 21, 19, 4, 23, 24, 10, 0, 
    221, 52, 77, 84, 78, 78, 70, 65, 54, 53, 63, 61, 57, 51, 43, 37, 31, 31, 50, 30, 17, 36, 33, 19, 16, 15, 11, 8, 13, 21, 53, 0, 
    228, 47, 70, 85, 74, 69, 56, 52, 58, 63, 61, 54, 48, 42, 31, 25, 24, 39, 72, 46, 28, 32, 29, 15, 2, 16, 17, 13, 22, 36, 55, 17, 
    230, 56, 71, 79, 70, 65, 58, 44, 47, 65, 56, 53, 48, 32, 9, 22, 37, 64, 110, 61, 24, 24, 21, 19, 16, 23, 24, 25, 37, 43, 38, 14, 
    235, 94, 72, 62, 61, 56, 47, 42, 46, 64, 66, 78, 58, 28, 0, 24, 53, 68, 106, 58, 25, 31, 31, 28, 24, 30, 32, 36, 45, 42, 25, 13, 
    216, 117, 73, 59, 61, 45, 28, 49, 62, 69, 78, 104, 70, 26, 0, 15, 42, 52, 81, 57, 39, 39, 33, 31, 35, 46, 39, 42, 50, 40, 30, 25, 
    199, 118, 77, 62, 64, 45, 16, 53, 72, 71, 74, 89, 55, 23, 13, 33, 49, 53, 61, 47, 36, 36, 44, 50, 46, 44, 38, 48, 46, 41, 43, 32, 
    193, 104, 77, 57, 58, 42, 16, 44, 60, 54, 61, 70, 57, 48, 47, 53, 53, 47, 48, 44, 43, 45, 48, 51, 55, 37, 35, 50, 48, 46, 50, 35, 
    181, 87, 74, 53, 55, 47, 38, 54, 63, 60, 62, 62, 56, 55, 53, 53, 49, 48, 57, 56, 45, 45, 47, 52, 60, 38, 40, 55, 55, 53, 54, 35, 
    157, 76, 75, 64, 67, 63, 63, 69, 67, 58, 53, 52, 52, 55, 58, 56, 53, 61, 64, 47, 42, 50, 48, 51, 56, 44, 49, 58, 58, 56, 54, 31, 
    129, 64, 64, 65, 68, 64, 62, 66, 66, 58, 56, 57, 59, 60, 61, 55, 51, 69, 70, 28, 36, 53, 50, 50, 52, 51, 56, 59, 58, 54, 43, 27, 
    110, 52, 52, 60, 63, 61, 60, 64, 67, 64, 61, 60, 59, 58, 57, 50, 49, 79, 74, 14, 35, 57, 50, 50, 53, 56, 59, 60, 57, 46, 26, 31, 
    104, 53, 51, 59, 61, 60, 58, 60, 60, 60, 58, 56, 58, 56, 54, 46, 48, 84, 76, 12, 39, 59, 50, 52, 55, 57, 60, 63, 53, 32, 22, 41, 
    104, 57, 53, 58, 57, 57, 56, 57, 57, 56, 56, 53, 52, 50, 48, 44, 49, 89, 84, 19, 44, 56, 53, 55, 54, 57, 62, 63, 43, 21, 32, 47, 
    86, 57, 55, 57, 57, 57, 57, 58, 56, 55, 54, 53, 53, 52, 50, 49, 53, 79, 79, 38, 49, 56, 56, 57, 56, 57, 58, 63, 44, 30, 45, 51, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 12, 11, 15, 
    
    -- channel=41
    139, 212, 198, 199, 203, 210, 208, 203, 196, 189, 177, 169, 158, 152, 149, 142, 143, 142, 145, 144, 140, 136, 133, 134, 134, 136, 137, 136, 134, 132, 131, 69, 
    211, 292, 269, 264, 274, 283, 276, 269, 261, 251, 237, 221, 211, 204, 202, 197, 193, 194, 198, 195, 186, 178, 173, 179, 182, 186, 188, 189, 184, 180, 181, 132, 
    197, 272, 249, 239, 248, 256, 248, 240, 231, 223, 211, 197, 193, 189, 192, 189, 186, 187, 189, 181, 171, 159, 156, 169, 174, 177, 180, 182, 175, 172, 174, 128, 
    182, 250, 227, 215, 220, 227, 219, 208, 200, 194, 185, 175, 173, 172, 178, 179, 176, 179, 184, 177, 166, 152, 155, 166, 169, 168, 170, 172, 168, 163, 167, 123, 
    168, 229, 206, 194, 195, 199, 191, 180, 172, 169, 164, 157, 158, 158, 160, 165, 161, 168, 176, 174, 161, 149, 162, 170, 166, 158, 157, 157, 158, 156, 161, 119, 
    150, 204, 183, 171, 170, 171, 163, 152, 142, 144, 144, 143, 147, 146, 139, 144, 143, 153, 166, 166, 155, 150, 162, 164, 158, 146, 139, 135, 139, 143, 147, 110, 
    130, 176, 159, 144, 143, 137, 130, 119, 109, 113, 117, 123, 128, 132, 126, 127, 135, 136, 153, 152, 132, 136, 138, 132, 135, 127, 122, 115, 110, 113, 106, 83, 
    110, 146, 135, 115, 115, 102, 97, 86, 78, 81, 86, 96, 101, 114, 116, 122, 139, 145, 157, 163, 152, 151, 135, 114, 112, 112, 104, 94, 78, 71, 56, 51, 
    93, 123, 115, 95, 96, 86, 79, 71, 62, 61, 61, 73, 82, 100, 113, 140, 158, 173, 176, 180, 180, 171, 147, 116, 92, 103, 92, 78, 58, 42, 36, 39, 
    84, 114, 110, 100, 102, 99, 89, 84, 77, 69, 69, 80, 96, 116, 138, 165, 176, 184, 188, 191, 188, 181, 160, 126, 97, 89, 82, 64, 62, 50, 69, 54, 
    88, 130, 128, 129, 129, 129, 116, 110, 110, 107, 112, 122, 143, 167, 189, 201, 193, 187, 183, 183, 177, 175, 155, 129, 113, 81, 80, 60, 69, 78, 102, 71, 
    106, 160, 153, 151, 152, 153, 143, 141, 151, 164, 167, 177, 197, 218, 231, 225, 204, 189, 182, 179, 174, 162, 148, 134, 115, 73, 63, 67, 65, 94, 114, 82, 
    123, 183, 171, 160, 160, 163, 159, 160, 180, 200, 204, 212, 232, 248, 248, 235, 219, 204, 201, 195, 184, 156, 140, 129, 114, 84, 45, 66, 60, 81, 108, 80, 
    133, 199, 184, 164, 162, 169, 174, 188, 208, 223, 233, 240, 252, 261, 258, 249, 239, 232, 226, 214, 187, 151, 126, 107, 99, 91, 51, 55, 61, 59, 92, 74, 
    148, 218, 201, 188, 190, 197, 213, 230, 240, 247, 256, 263, 270, 274, 271, 264, 257, 248, 229, 203, 166, 128, 105, 87, 83, 91, 78, 58, 66, 55, 76, 62, 
    164, 238, 225, 216, 221, 234, 248, 263, 272, 275, 277, 281, 285, 284, 278, 262, 254, 239, 213, 177, 139, 108, 90, 84, 87, 99, 106, 88, 77, 73, 78, 57, 
    180, 256, 245, 233, 231, 250, 267, 284, 292, 293, 292, 289, 287, 277, 265, 243, 226, 214, 194, 165, 130, 108, 95, 100, 107, 117, 125, 110, 85, 85, 82, 53, 
    183, 257, 244, 235, 233, 246, 269, 284, 291, 291, 287, 280, 273, 260, 245, 226, 205, 194, 183, 166, 141, 127, 122, 125, 131, 133, 131, 112, 89, 91, 91, 57, 
    173, 251, 244, 242, 248, 254, 268, 274, 278, 278, 273, 266, 256, 243, 228, 214, 197, 187, 183, 175, 160, 150, 147, 142, 144, 136, 125, 107, 88, 82, 92, 68, 
    178, 255, 252, 256, 264, 271, 266, 263, 265, 263, 261, 252, 241, 228, 215, 201, 188, 181, 178, 179, 170, 162, 157, 148, 139, 128, 116, 103, 90, 83, 87, 74, 
    186, 267, 268, 277, 280, 278, 268, 254, 249, 246, 247, 243, 235, 218, 201, 180, 165, 166, 170, 176, 171, 162, 153, 144, 131, 123, 113, 102, 94, 83, 77, 64, 
    192, 279, 284, 284, 278, 266, 256, 241, 228, 227, 231, 231, 229, 213, 190, 167, 151, 150, 161, 167, 160, 154, 147, 139, 129, 117, 111, 104, 90, 80, 68, 41, 
    179, 266, 274, 274, 267, 253, 237, 220, 209, 208, 212, 218, 220, 212, 186, 162, 150, 142, 149, 154, 150, 146, 141, 130, 122, 113, 109, 99, 87, 76, 60, 30, 
    154, 242, 252, 256, 256, 244, 225, 208, 203, 204, 202, 205, 202, 193, 173, 158, 151, 145, 145, 143, 137, 136, 134, 128, 118, 108, 102, 93, 83, 68, 56, 30, 
    143, 225, 233, 238, 239, 234, 213, 198, 192, 190, 181, 177, 171, 165, 159, 154, 149, 144, 138, 132, 127, 126, 125, 121, 109, 100, 95, 89, 80, 71, 63, 35, 
    131, 202, 208, 207, 204, 200, 186, 178, 171, 164, 155, 149, 143, 143, 141, 140, 137, 133, 131, 126, 120, 112, 109, 106, 103, 96, 89, 85, 82, 80, 73, 43, 
    109, 162, 166, 162, 158, 154, 152, 151, 143, 135, 126, 122, 121, 127, 128, 125, 124, 128, 126, 121, 110, 101, 97, 92, 93, 90, 85, 83, 84, 84, 74, 44, 
    78, 112, 113, 112, 113, 115, 116, 117, 116, 113, 111, 110, 113, 119, 118, 111, 110, 119, 119, 118, 104, 94, 87, 85, 85, 85, 84, 83, 81, 75, 63, 34, 
    52, 76, 74, 78, 84, 89, 92, 94, 100, 103, 106, 107, 109, 114, 108, 96, 93, 107, 119, 114, 96, 85, 81, 80, 80, 83, 84, 82, 75, 60, 42, 17, 
    41, 62, 62, 67, 75, 82, 85, 88, 94, 100, 102, 104, 105, 109, 100, 83, 75, 94, 111, 107, 87, 79, 76, 76, 78, 81, 84, 82, 65, 45, 18, 0, 
    42, 66, 67, 73, 79, 84, 85, 86, 89, 92, 93, 92, 91, 90, 78, 58, 52, 76, 99, 97, 80, 75, 71, 72, 77, 80, 82, 76, 55, 29, 0, 0, 
    27, 43, 43, 47, 50, 53, 53, 53, 53, 53, 52, 50, 48, 47, 38, 25, 19, 37, 61, 57, 47, 43, 42, 43, 46, 49, 49, 44, 30, 6, 0, 0, 
    
    -- channel=42
    241, 203, 178, 211, 248, 254, 254, 258, 264, 265, 255, 262, 272, 273, 276, 259, 260, 272, 279, 282, 274, 271, 276, 279, 267, 267, 280, 274, 264, 275, 282, 35, 
    383, 309, 271, 323, 379, 384, 376, 381, 395, 393, 377, 385, 399, 399, 406, 383, 383, 402, 409, 407, 384, 388, 403, 410, 393, 394, 415, 406, 386, 406, 415, 43, 
    389, 311, 271, 322, 378, 386, 375, 377, 396, 392, 371, 377, 395, 391, 405, 387, 382, 399, 404, 366, 331, 367, 404, 413, 394, 393, 418, 405, 382, 407, 417, 40, 
    392, 311, 268, 318, 373, 384, 367, 365, 392, 387, 363, 366, 385, 374, 392, 386, 376, 393, 390, 329, 291, 357, 405, 412, 393, 389, 413, 399, 380, 405, 412, 38, 
    394, 309, 260, 312, 365, 377, 365, 359, 387, 381, 355, 354, 377, 356, 359, 365, 356, 387, 370, 257, 244, 356, 407, 412, 390, 377, 401, 389, 375, 400, 402, 35, 
    391, 304, 243, 297, 354, 368, 359, 352, 380, 371, 346, 349, 372, 336, 316, 331, 330, 359, 347, 232, 222, 324, 363, 384, 381, 362, 383, 375, 367, 392, 388, 31, 
    388, 296, 232, 289, 351, 355, 348, 346, 368, 354, 338, 343, 359, 328, 309, 304, 282, 270, 237, 152, 154, 225, 232, 261, 322, 341, 366, 357, 341, 370, 365, 22, 
    355, 268, 213, 262, 315, 304, 309, 320, 334, 322, 317, 329, 332, 307, 295, 274, 231, 211, 196, 154, 153, 187, 170, 183, 247, 291, 317, 306, 279, 319, 319, 8, 
    286, 214, 178, 208, 241, 230, 240, 260, 267, 260, 263, 276, 271, 267, 279, 244, 189, 166, 157, 150, 143, 142, 120, 159, 222, 269, 278, 237, 202, 238, 246, 0, 
    205, 160, 140, 165, 189, 174, 185, 201, 207, 201, 206, 218, 217, 227, 239, 200, 164, 163, 165, 153, 141, 159, 152, 165, 183, 220, 275, 211, 161, 182, 190, 0, 
    149, 138, 132, 160, 173, 152, 139, 158, 184, 178, 176, 196, 207, 217, 216, 191, 171, 175, 177, 162, 149, 191, 229, 254, 220, 185, 262, 216, 137, 143, 147, 0, 
    145, 150, 131, 158, 177, 143, 131, 166, 207, 206, 185, 193, 209, 211, 195, 172, 164, 169, 175, 167, 164, 226, 283, 293, 254, 190, 252, 247, 128, 115, 133, 0, 
    158, 163, 141, 158, 160, 133, 127, 164, 208, 215, 201, 202, 219, 218, 198, 188, 185, 185, 196, 194, 202, 270, 315, 307, 276, 200, 209, 246, 126, 81, 118, 0, 
    172, 170, 142, 145, 146, 127, 147, 198, 231, 242, 238, 236, 247, 244, 228, 231, 236, 236, 241, 236, 243, 287, 303, 298, 282, 225, 172, 175, 102, 59, 98, 0, 
    195, 185, 170, 170, 181, 188, 210, 236, 257, 274, 276, 273, 279, 282, 267, 264, 273, 269, 258, 229, 228, 255, 267, 271, 266, 246, 167, 125, 103, 77, 92, 0, 
    211, 201, 211, 209, 218, 233, 249, 272, 287, 295, 300, 304, 306, 302, 289, 276, 276, 272, 252, 202, 199, 232, 248, 260, 254, 251, 185, 141, 178, 168, 125, 0, 
    233, 226, 225, 211, 219, 256, 284, 298, 306, 309, 306, 300, 293, 285, 272, 256, 258, 273, 255, 202, 200, 235, 248, 257, 249, 247, 210, 179, 211, 212, 170, 0, 
    228, 198, 196, 197, 218, 254, 286, 296, 291, 283, 277, 274, 273, 271, 268, 259, 251, 264, 261, 221, 223, 255, 259, 254, 251, 247, 225, 211, 226, 211, 192, 0, 
    201, 177, 196, 215, 236, 263, 276, 274, 264, 264, 268, 271, 272, 272, 269, 263, 252, 263, 271, 252, 250, 265, 263, 252, 242, 224, 200, 180, 159, 158, 200, 2, 
    216, 184, 204, 230, 250, 260, 257, 252, 257, 263, 269, 271, 272, 264, 249, 230, 208, 235, 268, 264, 260, 263, 255, 227, 200, 184, 159, 129, 115, 120, 148, 0, 
    222, 210, 239, 256, 260, 260, 250, 234, 239, 254, 264, 271, 270, 234, 188, 163, 148, 202, 262, 259, 244, 230, 212, 186, 164, 143, 115, 98, 96, 88, 88, 0, 
    238, 242, 247, 247, 246, 238, 220, 201, 205, 212, 235, 260, 259, 210, 152, 135, 135, 188, 234, 219, 199, 186, 172, 143, 119, 103, 87, 77, 75, 58, 29, 0, 
    220, 238, 236, 235, 234, 201, 171, 159, 164, 170, 209, 252, 254, 201, 143, 130, 129, 161, 192, 178, 163, 147, 123, 100, 92, 81, 66, 58, 55, 30, 2, 0, 
    199, 230, 227, 229, 230, 186, 147, 149, 160, 168, 201, 225, 205, 159, 127, 130, 135, 148, 154, 139, 118, 104, 98, 92, 81, 62, 49, 45, 31, 13, 4, 0, 
    186, 216, 215, 213, 210, 169, 135, 139, 143, 139, 154, 165, 154, 139, 129, 130, 126, 120, 114, 104, 95, 87, 75, 74, 70, 47, 34, 30, 21, 14, 12, 0, 
    154, 168, 165, 157, 152, 126, 109, 117, 121, 124, 126, 122, 114, 108, 106, 107, 98, 91, 95, 88, 73, 61, 58, 68, 59, 33, 25, 26, 23, 20, 16, 0, 
    105, 105, 102, 98, 97, 90, 88, 95, 95, 90, 87, 85, 84, 85, 87, 84, 80, 90, 87, 70, 58, 53, 47, 48, 40, 23, 21, 26, 25, 25, 16, 0, 
    63, 51, 48, 49, 52, 52, 54, 62, 66, 64, 64, 67, 71, 74, 73, 63, 64, 92, 89, 58, 47, 43, 35, 32, 26, 22, 25, 26, 29, 22, 3, 0, 
    33, 19, 18, 26, 32, 34, 39, 48, 55, 58, 59, 60, 60, 61, 59, 48, 59, 104, 85, 38, 33, 32, 27, 22, 20, 22, 26, 28, 29, 4, 0, 0, 
    25, 14, 16, 23, 30, 34, 38, 44, 48, 51, 51, 54, 56, 55, 48, 31, 43, 94, 72, 26, 25, 28, 20, 17, 18, 20, 25, 31, 16, 0, 0, 0, 
    27, 21, 24, 29, 32, 35, 37, 40, 44, 48, 46, 42, 36, 26, 13, 0, 11, 69, 55, 18, 20, 18, 15, 15, 15, 16, 27, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    24, 18, 18, 0, 3, 4, 3, 4, 3, 3, 7, 0, 1, 1, 0, 11, 0, 3, 2, 1, 4, 3, 3, 1, 8, 2, 0, 6, 7, 0, 0, 127, 
    0, 5, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 161, 
    0, 4, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 161, 
    0, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 161, 
    0, 2, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 160, 
    0, 4, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 
    0, 3, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 14, 53, 94, 46, 22, 45, 38, 30, 11, 0, 0, 0, 0, 0, 153, 
    0, 21, 35, 0, 0, 5, 7, 0, 0, 2, 0, 0, 0, 5, 0, 14, 22, 24, 17, 27, 18, 0, 6, 0, 0, 13, 6, 15, 18, 0, 10, 158, 
    10, 40, 47, 15, 21, 35, 22, 22, 24, 27, 21, 18, 24, 19, 13, 36, 37, 32, 24, 25, 26, 28, 41, 0, 0, 0, 0, 23, 34, 9, 33, 155, 
    15, 38, 44, 23, 14, 21, 15, 17, 21, 24, 22, 22, 27, 16, 18, 41, 43, 33, 30, 34, 35, 29, 27, 3, 20, 0, 0, 11, 10, 4, 21, 125, 
    15, 27, 26, 5, 7, 18, 20, 17, 7, 12, 9, 5, 4, 1, 11, 23, 21, 17, 17, 21, 21, 0, 0, 0, 0, 0, 0, 38, 21, 21, 22, 109, 
    13, 14, 25, 10, 24, 37, 29, 2, 0, 5, 3, 0, 7, 16, 24, 29, 30, 24, 21, 25, 22, 0, 0, 0, 2, 9, 0, 27, 49, 32, 29, 104, 
    12, 21, 34, 11, 30, 46, 34, 15, 15, 26, 28, 12, 7, 16, 20, 15, 12, 9, 6, 13, 4, 0, 0, 0, 15, 40, 0, 3, 71, 37, 37, 109, 
    17, 23, 35, 20, 25, 28, 20, 1, 0, 0, 5, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 29, 12, 87, 55, 31, 104, 
    11, 9, 15, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 18, 16, 9, 8, 2, 3, 9, 45, 23, 39, 40, 21, 89, 
    17, 9, 10, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 7, 14, 21, 34, 17, 5, 0, 0, 5, 2, 39, 22, 0, 0, 4, 81, 
    16, 6, 11, 23, 21, 12, 6, 0, 0, 0, 0, 1, 7, 12, 17, 19, 6, 0, 6, 17, 0, 0, 0, 0, 6, 5, 27, 21, 1, 24, 30, 96, 
    13, 26, 34, 30, 11, 0, 0, 0, 3, 9, 14, 15, 10, 5, 0, 0, 0, 0, 6, 18, 0, 0, 0, 0, 4, 2, 13, 16, 12, 24, 34, 127, 
    31, 29, 13, 0, 0, 0, 0, 6, 16, 12, 5, 0, 0, 0, 0, 0, 7, 0, 0, 12, 3, 0, 2, 4, 7, 15, 29, 35, 39, 32, 17, 132, 
    13, 2, 0, 3, 6, 11, 8, 7, 3, 0, 0, 0, 1, 9, 18, 27, 38, 19, 6, 6, 2, 0, 5, 22, 31, 38, 41, 43, 43, 28, 18, 133, 
    21, 14, 0, 0, 1, 2, 9, 10, 5, 11, 9, 6, 6, 22, 40, 48, 46, 11, 3, 7, 10, 19, 28, 41, 37, 34, 43, 45, 36, 39, 39, 105, 
    15, 12, 6, 5, 6, 12, 24, 35, 27, 31, 22, 11, 7, 27, 30, 22, 18, 0, 0, 27, 34, 36, 35, 37, 42, 46, 49, 45, 44, 58, 60, 85, 
    0, 12, 17, 14, 15, 30, 38, 41, 33, 27, 5, 2, 8, 30, 32, 22, 28, 13, 17, 29, 30, 31, 39, 50, 47, 48, 47, 46, 50, 57, 60, 80, 
    1, 6, 13, 10, 11, 31, 24, 14, 10, 9, 0, 4, 32, 56, 60, 46, 36, 23, 20, 27, 38, 47, 48, 43, 36, 44, 48, 50, 51, 53, 54, 77, 
    8, 5, 14, 14, 20, 41, 35, 25, 30, 38, 37, 39, 41, 39, 33, 27, 30, 33, 40, 47, 48, 42, 41, 40, 46, 53, 51, 52, 53, 52, 51, 76, 
    26, 28, 42, 46, 49, 61, 60, 50, 45, 38, 30, 29, 30, 34, 36, 38, 45, 48, 45, 42, 42, 46, 48, 40, 50, 58, 51, 49, 50, 50, 49, 78, 
    41, 44, 52, 51, 47, 47, 44, 38, 37, 36, 38, 40, 43, 45, 48, 47, 44, 31, 29, 40, 46, 50, 48, 44, 51, 54, 51, 48, 48, 47, 51, 80, 
    41, 44, 44, 44, 45, 45, 44, 43, 47, 49, 50, 49, 44, 38, 39, 43, 37, 27, 42, 48, 48, 48, 48, 49, 51, 51, 47, 47, 46, 49, 59, 79, 
    49, 52, 50, 47, 48, 49, 47, 43, 43, 42, 38, 37, 38, 40, 45, 49, 38, 25, 53, 58, 48, 49, 52, 51, 51, 49, 47, 47, 47, 60, 67, 76, 
    49, 53, 49, 46, 44, 43, 41, 39, 38, 40, 42, 42, 43, 45, 50, 55, 42, 27, 56, 57, 48, 51, 50, 51, 50, 49, 48, 47, 54, 70, 67, 69, 
    44, 47, 44, 43, 45, 45, 45, 45, 45, 45, 47, 49, 53, 57, 62, 67, 51, 34, 61, 59, 51, 51, 51, 51, 51, 51, 46, 49, 66, 71, 65, 65, 
    67, 73, 73, 73, 74, 74, 73, 74, 74, 74, 75, 75, 74, 73, 70, 68, 57, 52, 81, 81, 72, 71, 71, 73, 72, 71, 67, 73, 80, 71, 65, 68, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 9, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 4, 12, 
    10, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 4, 1, 10, 19, 
    14, 3, 5, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 3, 3, 3, 7, 18, 26, 
    15, 4, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 8, 0, 0, 0, 0, 3, 1, 2, 3, 5, 6, 3, 4, 17, 25, 31, 
    22, 16, 15, 14, 12, 11, 10, 9, 9, 8, 8, 8, 9, 10, 15, 19, 21, 16, 3, 4, 13, 14, 14, 13, 14, 15, 17, 14, 16, 25, 32, 34, 
    
    -- channel=45
    225, 441, 406, 408, 440, 497, 519, 527, 536, 543, 539, 543, 542, 557, 565, 551, 551, 543, 566, 576, 575, 571, 566, 570, 564, 563, 562, 565, 565, 562, 566, 334, 
    439, 727, 673, 678, 731, 814, 838, 848, 860, 870, 866, 863, 867, 886, 901, 880, 880, 873, 900, 909, 895, 890, 882, 906, 900, 900, 902, 908, 900, 899, 904, 553, 
    446, 736, 678, 681, 731, 818, 839, 845, 856, 867, 861, 851, 859, 872, 897, 878, 882, 872, 892, 868, 832, 818, 837, 900, 900, 903, 906, 910, 900, 900, 905, 555, 
    446, 735, 673, 676, 720, 810, 825, 830, 842, 851, 848, 831, 839, 842, 876, 860, 872, 867, 871, 823, 760, 744, 800, 892, 895, 898, 899, 901, 895, 892, 899, 549, 
    446, 735, 665, 668, 702, 797, 812, 819, 830, 837, 837, 812, 821, 812, 832, 814, 825, 844, 831, 746, 668, 665, 775, 887, 887, 883, 880, 877, 878, 878, 887, 538, 
    442, 728, 645, 649, 673, 778, 793, 805, 815, 820, 820, 795, 809, 782, 775, 744, 748, 782, 779, 691, 608, 603, 713, 822, 838, 847, 848, 838, 849, 858, 868, 522, 
    436, 716, 628, 632, 656, 758, 777, 788, 800, 800, 798, 778, 792, 767, 746, 693, 674, 653, 614, 517, 441, 446, 507, 586, 658, 728, 790, 795, 801, 814, 817, 490, 
    399, 662, 583, 583, 609, 685, 709, 720, 744, 746, 745, 741, 751, 732, 705, 652, 610, 545, 491, 420, 380, 378, 374, 404, 464, 570, 669, 698, 693, 708, 704, 427, 
    323, 542, 488, 483, 502, 543, 560, 579, 611, 619, 623, 633, 641, 640, 637, 605, 544, 450, 389, 350, 332, 314, 286, 309, 353, 488, 566, 581, 550, 538, 542, 322, 
    217, 388, 367, 371, 384, 402, 416, 431, 463, 469, 481, 494, 507, 523, 533, 513, 462, 402, 381, 363, 344, 344, 330, 343, 355, 436, 502, 498, 470, 411, 417, 225, 
    133, 285, 293, 316, 328, 345, 330, 332, 359, 379, 399, 408, 430, 462, 477, 463, 423, 396, 387, 371, 349, 372, 403, 474, 477, 457, 499, 465, 444, 360, 332, 166, 
    118, 274, 287, 317, 333, 347, 326, 322, 367, 415, 420, 412, 427, 453, 457, 426, 390, 372, 370, 363, 359, 407, 482, 578, 575, 502, 519, 491, 449, 368, 295, 150, 
    137, 310, 323, 336, 331, 338, 308, 321, 385, 444, 457, 455, 466, 477, 469, 439, 411, 397, 405, 409, 427, 487, 573, 655, 649, 561, 512, 496, 416, 347, 257, 125, 
    161, 345, 338, 327, 312, 307, 311, 360, 432, 493, 516, 522, 525, 527, 514, 500, 487, 491, 498, 498, 512, 552, 605, 651, 647, 593, 496, 445, 338, 270, 211, 96, 
    192, 388, 374, 368, 366, 377, 408, 449, 503, 549, 577, 591, 598, 604, 593, 585, 581, 584, 576, 541, 528, 531, 566, 592, 600, 588, 488, 405, 293, 225, 205, 87, 
    218, 433, 435, 440, 455, 479, 514, 556, 596, 627, 646, 662, 669, 670, 657, 637, 625, 616, 596, 533, 493, 476, 513, 553, 568, 575, 499, 422, 357, 323, 314, 141, 
    251, 480, 485, 485, 492, 532, 582, 635, 665, 680, 684, 680, 670, 656, 634, 603, 587, 588, 576, 521, 471, 457, 498, 542, 554, 564, 519, 467, 439, 441, 427, 207, 
    249, 464, 458, 454, 465, 508, 576, 630, 653, 654, 642, 630, 620, 610, 597, 578, 560, 564, 563, 532, 506, 506, 538, 559, 561, 562, 532, 510, 501, 491, 472, 242, 
    220, 425, 419, 431, 470, 519, 570, 600, 607, 605, 596, 595, 594, 592, 587, 579, 565, 572, 576, 575, 568, 568, 578, 575, 562, 534, 498, 458, 410, 387, 410, 225, 
    231, 423, 415, 449, 507, 548, 566, 569, 569, 567, 577, 584, 589, 588, 577, 553, 518, 522, 540, 577, 587, 583, 580, 553, 513, 466, 415, 359, 309, 281, 303, 171, 
    236, 453, 478, 521, 556, 569, 564, 544, 535, 540, 569, 586, 594, 564, 513, 445, 388, 417, 475, 547, 566, 543, 518, 478, 428, 370, 316, 267, 230, 204, 210, 91, 
    259, 486, 527, 542, 542, 535, 520, 491, 476, 477, 513, 539, 564, 527, 447, 356, 304, 347, 415, 483, 487, 457, 426, 375, 322, 271, 231, 198, 173, 154, 120, 9, 
    229, 452, 511, 525, 522, 491, 454, 400, 381, 380, 424, 477, 534, 507, 419, 331, 286, 313, 360, 398, 392, 359, 320, 273, 238, 202, 176, 148, 132, 101, 54, 0, 
    191, 414, 481, 503, 505, 464, 405, 343, 329, 344, 385, 436, 470, 437, 371, 321, 301, 312, 320, 319, 294, 266, 239, 216, 191, 162, 136, 110, 87, 55, 24, 0, 
    175, 390, 446, 470, 469, 430, 369, 318, 307, 311, 331, 354, 366, 348, 321, 299, 284, 274, 263, 250, 232, 209, 183, 171, 154, 135, 106, 77, 57, 38, 24, 0, 
    144, 331, 365, 380, 370, 341, 305, 280, 276, 278, 279, 274, 263, 249, 241, 236, 226, 219, 215, 202, 183, 155, 138, 140, 131, 112, 79, 57, 49, 41, 33, 0, 
    89, 227, 243, 247, 237, 226, 215, 211, 208, 203, 192, 186, 184, 188, 192, 190, 184, 185, 178, 170, 147, 125, 113, 106, 96, 77, 55, 47, 47, 46, 38, 0, 
    28, 119, 115, 112, 112, 112, 114, 122, 133, 140, 142, 144, 148, 154, 156, 146, 140, 158, 169, 167, 129, 100, 86, 77, 64, 53, 47, 46, 51, 44, 29, 0, 
    0, 46, 40, 41, 52, 62, 71, 84, 99, 112, 117, 120, 120, 123, 123, 112, 115, 158, 175, 160, 101, 70, 68, 55, 46, 43, 44, 49, 52, 30, 0, 0, 
    0, 28, 28, 31, 44, 55, 64, 72, 82, 92, 97, 103, 108, 112, 108, 87, 88, 133, 151, 136, 75, 56, 51, 41, 36, 36, 42, 50, 41, 7, 0, 0, 
    0, 33, 37, 41, 51, 59, 66, 73, 82, 91, 95, 94, 87, 74, 55, 24, 22, 74, 104, 104, 58, 39, 37, 31, 30, 29, 39, 39, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 7, 9, 7, 3, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 56, 54, 74, 77, 85, 89, 95, 100, 100, 102, 114, 116, 122, 129, 122, 130, 131, 134, 128, 121, 134, 140, 140, 136, 138, 138, 134, 135, 138, 133, 22, 
    60, 71, 66, 84, 88, 97, 101, 112, 116, 114, 117, 121, 127, 130, 138, 129, 135, 134, 135, 122, 117, 140, 140, 147, 138, 140, 141, 136, 135, 143, 137, 28, 
    65, 83, 75, 91, 97, 110, 108, 112, 123, 123, 124, 127, 132, 125, 138, 128, 133, 135, 133, 125, 147, 153, 134, 142, 137, 142, 144, 137, 138, 147, 140, 29, 
    67, 86, 79, 100, 102, 119, 119, 129, 139, 132, 133, 131, 134, 123, 134, 121, 124, 137, 127, 98, 103, 121, 128, 144, 138, 142, 145, 141, 143, 141, 138, 29, 
    70, 92, 79, 104, 102, 124, 124, 131, 141, 136, 138, 133, 139, 122, 131, 132, 130, 136, 113, 106, 125, 101, 99, 126, 131, 141, 150, 143, 144, 144, 140, 33, 
    78, 102, 85, 114, 109, 129, 126, 133, 142, 141, 144, 136, 137, 127, 145, 141, 115, 100, 73, 42, 48, 60, 73, 91, 102, 123, 149, 144, 140, 144, 141, 35, 
    58, 85, 75, 93, 83, 95, 109, 118, 127, 130, 134, 128, 129, 125, 114, 86, 96, 112, 138, 119, 92, 116, 136, 155, 149, 112, 113, 114, 119, 139, 130, 33, 
    58, 80, 66, 72, 76, 89, 107, 99, 105, 111, 112, 108, 105, 112, 107, 90, 89, 72, 48, 24, 16, 11, 6, 59, 104, 131, 130, 120, 117, 132, 113, 41, 
    67, 79, 68, 78, 103, 107, 104, 107, 114, 115, 112, 111, 109, 111, 101, 81, 60, 37, 22, 17, 19, 26, 39, 40, 15, 73, 110, 121, 126, 120, 117, 51, 
    52, 59, 63, 75, 69, 59, 62, 74, 90, 87, 93, 99, 98, 86, 75, 71, 62, 49, 50, 52, 52, 69, 68, 82, 96, 98, 98, 61, 78, 68, 75, 18, 
    33, 38, 28, 32, 22, 25, 41, 66, 59, 51, 60, 55, 39, 28, 30, 28, 22, 31, 38, 35, 36, 56, 43, 50, 69, 81, 133, 82, 61, 63, 49, 8, 
    20, 11, 15, 44, 37, 29, 31, 19, 12, 21, 21, 35, 41, 36, 38, 41, 49, 53, 54, 51, 57, 71, 82, 96, 83, 69, 107, 105, 54, 67, 36, 1, 
    11, 20, 28, 37, 44, 45, 32, 45, 69, 72, 58, 55, 59, 51, 43, 45, 50, 53, 61, 57, 63, 74, 95, 120, 120, 94, 74, 94, 38, 52, 52, 8, 
    26, 38, 38, 41, 48, 48, 52, 46, 40, 47, 50, 42, 34, 36, 32, 29, 21, 26, 30, 28, 41, 63, 91, 108, 111, 107, 72, 95, 94, 60, 54, 13, 
    9, 17, 19, 25, 17, 0, 0, 5, 19, 28, 37, 45, 49, 48, 42, 45, 50, 50, 54, 61, 89, 105, 116, 110, 105, 102, 73, 83, 107, 71, 55, 11, 
    13, 26, 20, 6, 11, 25, 32, 44, 49, 53, 54, 54, 54, 57, 59, 62, 79, 88, 89, 88, 104, 99, 95, 101, 95, 91, 74, 55, 28, 7, 36, 7, 
    20, 4, 7, 35, 61, 71, 51, 44, 41, 39, 42, 52, 68, 83, 93, 92, 85, 78, 65, 58, 58, 65, 77, 91, 91, 93, 81, 66, 73, 89, 74, 0, 
    2, 24, 56, 65, 50, 37, 45, 41, 42, 58, 72, 79, 79, 76, 71, 65, 57, 74, 79, 69, 69, 75, 80, 81, 82, 72, 61, 65, 76, 84, 88, 6, 
    38, 48, 26, 0, 0, 13, 36, 53, 66, 72, 63, 54, 50, 46, 44, 46, 47, 67, 80, 82, 82, 83, 77, 64, 61, 62, 73, 73, 72, 78, 69, 0, 
    1, 0, 6, 28, 47, 55, 47, 45, 43, 30, 40, 53, 66, 61, 53, 57, 67, 85, 79, 77, 73, 63, 58, 62, 79, 83, 65, 56, 55, 36, 40, 31, 
    17, 24, 30, 36, 36, 31, 24, 17, 25, 32, 51, 67, 73, 65, 77, 82, 74, 83, 65, 54, 61, 66, 76, 77, 59, 44, 42, 42, 28, 15, 31, 21, 
    46, 27, 27, 31, 33, 26, 32, 38, 44, 54, 71, 63, 59, 52, 42, 28, 13, 24, 50, 74, 81, 75, 58, 38, 40, 42, 40, 32, 25, 31, 22, 0, 
    33, 36, 44, 47, 47, 42, 56, 56, 48, 45, 50, 39, 30, 18, 6, 10, 28, 49, 65, 62, 46, 35, 39, 51, 49, 30, 21, 20, 25, 20, 10, 0, 
    24, 36, 38, 37, 31, 18, 15, 6, 0, 0, 0, 24, 52, 65, 65, 57, 46, 35, 25, 23, 34, 52, 48, 32, 10, 9, 15, 13, 10, 7, 7, 0, 
    10, 13, 9, 13, 15, 10, 0, 2, 19, 40, 61, 67, 56, 37, 24, 19, 18, 23, 35, 45, 44, 27, 17, 23, 15, 13, 14, 11, 7, 7, 5, 0, 
    11, 22, 29, 38, 43, 45, 43, 42, 41, 36, 29, 23, 17, 15, 20, 29, 41, 54, 47, 24, 16, 16, 21, 21, 19, 16, 8, 7, 8, 7, 0, 0, 
    25, 30, 34, 30, 26, 23, 19, 14, 9, 12, 17, 24, 34, 40, 40, 36, 34, 26, 5, 12, 21, 20, 14, 9, 13, 10, 8, 8, 9, 4, 0, 0, 
    5, 6, 7, 9, 13, 14, 16, 22, 28, 35, 40, 38, 30, 20, 16, 13, 20, 25, 13, 19, 21, 9, 4, 8, 7, 7, 6, 6, 8, 0, 4, 1, 
    8, 10, 12, 15, 19, 23, 24, 25, 25, 20, 14, 12, 13, 15, 17, 14, 21, 34, 24, 22, 11, 4, 8, 4, 4, 5, 6, 8, 3, 0, 14, 6, 
    15, 15, 15, 12, 11, 9, 8, 8, 9, 12, 14, 14, 13, 12, 11, 7, 14, 26, 15, 11, 5, 6, 2, 1, 3, 4, 10, 6, 0, 8, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 7, 13, 13, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 
    32, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 3, 16, 27, 
    36, 5, 5, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 1, 0, 0, 1, 2, 10, 25, 36, 
    36, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 10, 0, 0, 0, 8, 4, 5, 4, 1, 2, 3, 5, 23, 29, 43, 
    42, 25, 22, 22, 20, 19, 18, 17, 15, 14, 15, 14, 16, 16, 21, 28, 30, 31, 22, 5, 20, 24, 25, 24, 23, 23, 23, 21, 29, 31, 40, 48, 
    
    -- channel=48
    95, 58, 46, 56, 57, 48, 56, 56, 52, 53, 54, 54, 52, 55, 52, 57, 57, 52, 53, 52, 53, 54, 53, 55, 56, 57, 56, 55, 51, 47, 65, 170, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 268, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 272, 
    0, 0, 0, 0, 0, 0, 31, 33, 5, 1, 0, 0, 7, 7, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 272, 
    0, 0, 0, 0, 0, 0, 58, 64, 16, 24, 27, 27, 42, 39, 32, 23, 31, 31, 22, 28, 25, 23, 44, 0, 0, 0, 0, 0, 0, 0, 8, 273, 
    0, 0, 0, 0, 0, 0, 41, 23, 17, 45, 33, 19, 33, 31, 29, 17, 21, 20, 10, 18, 15, 9, 21, 0, 0, 0, 0, 0, 0, 0, 6, 273, 
    0, 0, 0, 0, 0, 0, 52, 16, 15, 35, 13, 4, 38, 29, 18, 0, 2, 0, 0, 11, 2, 9, 0, 4, 0, 0, 0, 0, 0, 0, 6, 274, 
    0, 0, 0, 0, 0, 28, 83, 42, 8, 23, 22, 15, 46, 34, 22, 13, 23, 11, 17, 43, 15, 31, 5, 38, 17, 0, 0, 0, 0, 0, 5, 270, 
    0, 0, 0, 0, 0, 26, 38, 19, 0, 0, 12, 0, 8, 11, 8, 6, 11, 4, 5, 27, 5, 8, 0, 16, 22, 0, 0, 0, 0, 0, 4, 267, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 266, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 2, 0, 2, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 266, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 267, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 269, 
    0, 0, 6, 25, 52, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 269, 
    0, 0, 0, 13, 33, 75, 74, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 265, 
    0, 0, 0, 0, 0, 26, 81, 101, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 262, 
    0, 0, 0, 0, 0, 0, 0, 75, 123, 53, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 262, 
    0, 0, 0, 0, 0, 0, 0, 6, 125, 109, 46, 55, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 263, 
    0, 0, 0, 0, 0, 0, 0, 0, 87, 125, 61, 72, 71, 58, 34, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 263, 
    0, 0, 0, 0, 0, 0, 0, 0, 79, 144, 85, 70, 75, 71, 72, 72, 58, 43, 30, 27, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 263, 
    0, 0, 0, 0, 0, 0, 0, 13, 100, 167, 131, 70, 57, 65, 59, 81, 95, 88, 85, 82, 79, 30, 7, 7, 0, 3, 0, 0, 0, 0, 4, 264, 
    0, 0, 0, 0, 0, 0, 0, 58, 100, 98, 125, 107, 63, 87, 55, 34, 54, 67, 98, 72, 85, 86, 81, 73, 14, 0, 0, 0, 0, 0, 1, 261, 
    0, 0, 0, 0, 0, 0, 0, 21, 23, 0, 38, 102, 64, 50, 6, 0, 0, 17, 87, 35, 0, 29, 65, 50, 0, 0, 0, 0, 0, 0, 0, 255, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 9, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 250, 
    0, 0, 13, 17, 21, 23, 25, 27, 29, 24, 30, 31, 28, 22, 10, 6, 14, 6, 0, 0, 4, 0, 0, 0, 0, 2, 0, 0, 0, 0, 8, 234, 
    31, 25, 34, 39, 40, 38, 38, 41, 42, 38, 43, 44, 41, 33, 21, 6, 19, 27, 21, 21, 21, 23, 17, 13, 13, 13, 14, 22, 22, 18, 34, 218, 
    23, 23, 31, 30, 34, 36, 38, 42, 45, 48, 50, 49, 50, 47, 49, 42, 47, 62, 58, 55, 58, 63, 61, 58, 57, 57, 59, 70, 75, 67, 63, 202, 
    61, 56, 62, 65, 66, 74, 77, 74, 80, 84, 84, 81, 82, 80, 79, 79, 79, 89, 91, 89, 88, 86, 86, 87, 86, 85, 86, 91, 93, 63, 40, 179, 
    97, 78, 82, 83, 81, 86, 87, 82, 88, 92, 92, 88, 87, 86, 87, 86, 84, 87, 93, 95, 92, 88, 87, 89, 90, 88, 87, 82, 56, 16, 32, 195, 
    97, 81, 87, 85, 82, 90, 87, 83, 90, 93, 93, 89, 88, 89, 88, 86, 89, 92, 95, 91, 90, 86, 90, 90, 89, 86, 71, 38, 15, 41, 89, 206, 
    101, 83, 88, 88, 83, 86, 86, 85, 90, 90, 79, 79, 78, 84, 81, 74, 82, 83, 84, 81, 88, 84, 90, 92, 82, 59, 22, 18, 62, 106, 103, 184, 
    77, 85, 82, 82, 79, 78, 80, 81, 83, 82, 61, 64, 73, 77, 75, 67, 71, 71, 72, 74, 90, 87, 82, 75, 43, 18, 30, 77, 109, 94, 79, 174, 
    
    -- channel=49
    74, 181, 206, 210, 204, 192, 174, 173, 179, 183, 187, 189, 192, 186, 185, 181, 182, 185, 183, 185, 186, 189, 193, 191, 192, 199, 211, 227, 234, 235, 228, 122, 
    80, 251, 285, 294, 296, 288, 275, 267, 264, 266, 282, 292, 298, 295, 293, 291, 291, 294, 294, 296, 300, 300, 299, 296, 298, 306, 317, 326, 327, 331, 328, 213, 
    79, 251, 287, 300, 309, 307, 280, 250, 220, 222, 260, 272, 272, 268, 261, 263, 269, 279, 274, 278, 282, 279, 276, 279, 282, 308, 319, 326, 333, 338, 333, 218, 
    77, 249, 283, 298, 310, 318, 292, 249, 213, 215, 221, 212, 215, 214, 218, 219, 222, 229, 227, 230, 235, 231, 230, 247, 255, 300, 326, 330, 332, 334, 329, 215, 
    75, 248, 281, 295, 304, 312, 296, 263, 224, 225, 226, 219, 227, 231, 222, 225, 232, 247, 248, 250, 257, 250, 255, 267, 275, 315, 334, 336, 338, 339, 335, 218, 
    73, 248, 278, 290, 301, 304, 281, 236, 201, 229, 231, 223, 226, 221, 207, 218, 234, 248, 248, 257, 252, 245, 260, 253, 257, 281, 310, 332, 332, 337, 332, 215, 
    74, 248, 277, 288, 300, 296, 258, 202, 194, 222, 221, 218, 218, 221, 203, 210, 217, 227, 232, 227, 228, 220, 238, 233, 245, 251, 284, 326, 333, 335, 327, 211, 
    77, 252, 276, 286, 298, 291, 265, 228, 217, 230, 231, 235, 240, 242, 233, 236, 233, 241, 246, 243, 240, 234, 251, 251, 262, 263, 287, 319, 324, 326, 322, 210, 
    83, 260, 279, 282, 295, 296, 290, 262, 242, 233, 240, 239, 238, 243, 243, 246, 243, 251, 254, 247, 240, 235, 250, 264, 285, 282, 296, 324, 326, 325, 320, 209, 
    91, 271, 291, 286, 297, 302, 296, 275, 263, 248, 250, 250, 244, 256, 259, 261, 262, 261, 259, 255, 260, 254, 269, 289, 303, 308, 313, 324, 321, 322, 318, 208, 
    99, 287, 305, 298, 304, 305, 296, 293, 292, 281, 280, 278, 282, 285, 287, 290, 287, 289, 291, 291, 289, 289, 291, 299, 307, 317, 318, 318, 316, 322, 319, 210, 
    104, 296, 312, 294, 271, 259, 261, 283, 308, 302, 301, 299, 297, 301, 304, 306, 306, 302, 299, 299, 302, 302, 304, 303, 309, 322, 325, 327, 329, 333, 326, 213, 
    108, 303, 310, 277, 241, 212, 202, 206, 235, 271, 301, 314, 313, 313, 317, 322, 323, 322, 321, 321, 320, 320, 320, 323, 324, 325, 326, 327, 326, 327, 321, 208, 
    111, 309, 321, 303, 286, 254, 208, 177, 177, 199, 236, 275, 306, 321, 327, 330, 331, 330, 328, 324, 318, 316, 317, 318, 317, 316, 318, 319, 319, 322, 317, 206, 
    112, 312, 335, 326, 312, 289, 253, 205, 173, 156, 177, 223, 269, 308, 328, 332, 330, 329, 326, 322, 320, 318, 318, 321, 322, 321, 321, 320, 317, 319, 314, 204, 
    114, 316, 342, 338, 342, 340, 326, 274, 203, 147, 113, 143, 195, 237, 280, 314, 330, 331, 327, 323, 320, 319, 319, 319, 319, 319, 319, 319, 317, 318, 313, 204, 
    115, 318, 349, 346, 349, 350, 348, 331, 261, 178, 108, 87, 122, 160, 198, 232, 266, 295, 312, 320, 321, 319, 318, 322, 321, 320, 320, 320, 318, 319, 313, 204, 
    116, 320, 352, 347, 351, 351, 348, 343, 296, 214, 117, 74, 87, 97, 124, 156, 179, 200, 224, 246, 269, 288, 309, 323, 323, 321, 319, 319, 317, 318, 312, 201, 
    117, 321, 353, 348, 351, 352, 351, 346, 294, 211, 102, 44, 58, 66, 78, 93, 114, 133, 143, 144, 148, 169, 205, 250, 282, 303, 317, 325, 324, 322, 313, 202, 
    117, 322, 352, 345, 347, 349, 351, 330, 269, 172, 83, 36, 37, 52, 67, 73, 79, 84, 88, 89, 89, 100, 124, 157, 179, 200, 232, 261, 285, 305, 309, 200, 
    115, 315, 346, 340, 342, 344, 343, 312, 259, 200, 133, 86, 58, 29, 51, 82, 129, 161, 137, 100, 67, 86, 101, 103, 130, 175, 237, 274, 281, 292, 296, 195, 
    113, 310, 342, 337, 340, 343, 342, 324, 310, 287, 245, 192, 154, 136, 159, 198, 234, 247, 218, 200, 188, 187, 178, 177, 192, 222, 255, 275, 291, 303, 302, 196, 
    106, 295, 324, 322, 321, 320, 317, 312, 303, 279, 263, 250, 223, 202, 211, 222, 246, 264, 251, 238, 225, 235, 235, 225, 225, 229, 248, 259, 258, 267, 272, 177, 
    60, 204, 215, 214, 209, 206, 200, 196, 191, 189, 185, 184, 170, 151, 157, 168, 187, 208, 210, 205, 189, 195, 205, 208, 203, 201, 210, 216, 219, 222, 221, 139, 
    33, 177, 188, 185, 184, 184, 181, 179, 176, 176, 172, 169, 165, 164, 166, 172, 169, 168, 164, 161, 165, 163, 160, 161, 165, 166, 162, 157, 153, 149, 153, 92, 
    25, 137, 131, 134, 130, 127, 119, 112, 107, 104, 99, 96, 91, 87, 84, 88, 94, 96, 91, 85, 82, 80, 79, 79, 80, 83, 84, 81, 75, 72, 84, 47, 
    0, 90, 78, 78, 76, 76, 73, 75, 75, 75, 70, 66, 60, 61, 62, 64, 67, 70, 68, 61, 57, 57, 58, 59, 61, 61, 60, 59, 58, 63, 96, 77, 
    0, 81, 66, 68, 67, 66, 64, 63, 64, 64, 58, 52, 51, 51, 50, 53, 55, 57, 54, 45, 42, 41, 41, 40, 39, 37, 39, 45, 62, 98, 136, 79, 
    0, 58, 35, 41, 39, 38, 41, 41, 41, 41, 35, 33, 33, 37, 41, 43, 46, 47, 45, 43, 40, 41, 41, 42, 40, 40, 48, 75, 116, 134, 115, 48, 
    0, 58, 38, 43, 43, 43, 45, 45, 45, 46, 47, 52, 62, 62, 61, 64, 67, 70, 68, 65, 59, 54, 46, 45, 46, 56, 90, 129, 135, 101, 89, 43, 
    0, 58, 34, 39, 37, 38, 40, 40, 40, 42, 47, 50, 54, 56, 57, 59, 59, 62, 60, 59, 52, 49, 44, 49, 67, 101, 129, 117, 87, 79, 73, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 11, 9, 0, 0, 0, 
    
    -- channel=50
    92, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    147, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    145, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 
    143, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 16, 0, 0, 7, 19, 9, 0, 6, 0, 0, 0, 0, 12, 28, 0, 0, 0, 0, 0, 0, 0, 
    141, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 8, 0, 0, 10, 18, 4, 0, 2, 0, 0, 0, 0, 3, 15, 0, 0, 0, 0, 0, 0, 0, 
    141, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    140, 0, 0, 0, 0, 0, 0, 10, 30, 0, 0, 0, 0, 0, 5, 8, 0, 1, 0, 0, 4, 0, 3, 0, 0, 31, 2, 0, 0, 0, 0, 0, 
    140, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    152, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    157, 0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    160, 0, 0, 0, 0, 0, 0, 0, 0, 17, 22, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 30, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    165, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 28, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    165, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 32, 26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    166, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 18, 22, 25, 19, 10, 1, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    166, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 17, 10, 9, 9, 13, 10, 0, 7, 30, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 17, 30, 43, 16, 0, 0, 0, 17, 21, 9, 10, 42, 42, 0, 0, 0, 0, 0, 0, 
    163, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 38, 4, 0, 0, 0, 0, 0, 0, 0, 30, 32, 0, 0, 0, 0, 0, 0, 
    158, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 
    130, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    117, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 23, 21, 0, 
    61, 4, 3, 1, 2, 0, 0, 4, 1, 0, 2, 6, 5, 5, 6, 6, 6, 0, 0, 1, 5, 7, 6, 3, 5, 7, 7, 10, 22, 29, 0, 0, 
    44, 2, 6, 3, 11, 4, 3, 10, 4, 0, 3, 9, 9, 5, 5, 9, 8, 1, 0, 3, 7, 8, 5, 2, 4, 9, 20, 27, 12, 0, 0, 0, 
    44, 2, 5, 3, 8, 3, 5, 9, 3, 3, 11, 13, 2, 0, 3, 9, 4, 0, 0, 0, 0, 0, 3, 3, 10, 26, 28, 2, 0, 0, 0, 0, 
    43, 2, 7, 3, 9, 6, 4, 4, 4, 4, 14, 13, 3, 0, 2, 7, 3, 1, 0, 1, 0, 0, 5, 10, 24, 23, 0, 0, 0, 0, 0, 0, 
    35, 18, 20, 18, 20, 18, 17, 18, 18, 20, 30, 25, 16, 15, 17, 22, 20, 18, 17, 16, 8, 13, 20, 24, 34, 29, 3, 0, 0, 1, 19, 0, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 35, 26, 22, 12, 15, 36, 43, 43, 40, 36, 38, 38, 42, 42, 46, 39, 35, 41, 42, 43, 42, 42, 45, 43, 36, 28, 23, 23, 28, 37, 37, 
    75, 32, 29, 28, 16, 0, 0, 30, 35, 19, 16, 16, 11, 13, 10, 9, 5, 5, 2, 0, 2, 7, 7, 14, 0, 0, 13, 22, 31, 36, 42, 41, 
    71, 30, 34, 36, 29, 20, 13, 38, 42, 52, 60, 59, 66, 63, 66, 60, 54, 55, 60, 54, 56, 60, 54, 68, 41, 16, 32, 36, 38, 35, 38, 37, 
    69, 33, 37, 36, 35, 32, 23, 12, 0, 11, 38, 37, 44, 47, 37, 38, 30, 37, 42, 38, 41, 43, 44, 45, 40, 31, 32, 32, 33, 31, 36, 37, 
    70, 39, 39, 33, 34, 30, 39, 34, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 31, 26, 30, 32, 32, 35, 36, 
    64, 34, 39, 33, 29, 31, 44, 50, 52, 42, 26, 33, 29, 36, 30, 32, 38, 40, 41, 40, 50, 45, 45, 37, 64, 79, 51, 41, 43, 42, 42, 40, 
    58, 25, 34, 30, 26, 27, 12, 3, 8, 22, 15, 20, 24, 14, 12, 14, 16, 22, 31, 34, 35, 41, 32, 27, 23, 39, 44, 41, 42, 39, 43, 43, 
    53, 17, 30, 28, 29, 23, 0, 0, 0, 6, 13, 13, 23, 24, 17, 9, 0, 0, 2, 7, 3, 12, 15, 7, 0, 0, 10, 34, 36, 31, 39, 41, 
    55, 10, 24, 28, 29, 28, 20, 20, 34, 45, 46, 55, 50, 51, 47, 40, 42, 44, 48, 48, 52, 51, 54, 46, 24, 7, 19, 30, 30, 30, 37, 39, 
    61, 16, 18, 20, 20, 32, 30, 18, 11, 14, 12, 9, 8, 0, 0, 0, 0, 10, 15, 14, 11, 14, 10, 18, 32, 31, 33, 35, 36, 35, 37, 37, 
    70, 25, 22, 31, 46, 65, 57, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 22, 34, 34, 33, 32, 29, 32, 34, 
    77, 34, 35, 53, 88, 110, 130, 112, 60, 28, 16, 17, 18, 19, 19, 18, 18, 19, 20, 22, 25, 24, 22, 24, 28, 30, 29, 27, 25, 24, 31, 36, 
    80, 34, 24, 10, 19, 41, 90, 164, 178, 133, 76, 36, 24, 24, 22, 21, 20, 20, 18, 19, 23, 26, 27, 27, 28, 31, 34, 37, 40, 40, 44, 45, 
    82, 35, 15, 0, 0, 0, 0, 0, 100, 157, 155, 111, 54, 24, 18, 21, 25, 30, 32, 32, 34, 36, 37, 38, 38, 37, 36, 38, 38, 37, 40, 40, 
    81, 39, 30, 23, 25, 11, 0, 0, 0, 50, 119, 144, 137, 95, 53, 33, 30, 33, 36, 35, 31, 31, 30, 28, 26, 25, 25, 26, 27, 28, 32, 35, 
    79, 36, 32, 25, 26, 31, 27, 4, 0, 0, 73, 118, 158, 182, 160, 109, 65, 41, 30, 29, 31, 32, 28, 29, 29, 31, 31, 30, 29, 27, 29, 31, 
    79, 39, 41, 35, 33, 35, 38, 35, 9, 0, 40, 79, 99, 135, 174, 194, 176, 137, 98, 65, 51, 38, 25, 20, 23, 28, 31, 34, 34, 31, 30, 32, 
    82, 42, 46, 44, 42, 42, 39, 36, 34, 38, 63, 87, 82, 79, 89, 118, 162, 195, 204, 191, 163, 133, 94, 61, 45, 35, 29, 28, 30, 27, 28, 32, 
    86, 43, 43, 42, 41, 39, 37, 41, 71, 71, 83, 112, 102, 87, 76, 64, 68, 92, 127, 165, 195, 215, 215, 196, 166, 126, 90, 59, 37, 24, 22, 25, 
    92, 47, 42, 41, 42, 41, 39, 56, 68, 46, 3, 24, 81, 85, 86, 63, 20, 6, 20, 44, 39, 60, 126, 181, 201, 171, 134, 112, 83, 54, 37, 31, 
    95, 47, 38, 37, 37, 39, 41, 33, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 0, 0, 27, 44, 47, 38, 
    97, 49, 39, 44, 46, 50, 52, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 8, 24, 37, 37, 
    140, 116, 109, 115, 122, 130, 135, 137, 141, 144, 142, 122, 89, 64, 62, 67, 86, 102, 91, 64, 50, 62, 64, 47, 35, 46, 69, 79, 81, 82, 79, 66, 
    137, 143, 153, 148, 148, 149, 149, 150, 151, 152, 155, 152, 150, 145, 137, 129, 109, 96, 101, 104, 104, 102, 104, 105, 99, 87, 73, 68, 77, 91, 103, 94, 
    82, 44, 39, 34, 26, 25, 30, 32, 33, 35, 36, 34, 30, 29, 34, 46, 62, 67, 73, 80, 82, 85, 88, 94, 97, 98, 98, 97, 99, 113, 119, 106, 
    117, 97, 99, 94, 91, 91, 99, 109, 113, 118, 122, 124, 120, 120, 121, 120, 125, 127, 127, 133, 138, 135, 131, 130, 134, 138, 140, 138, 138, 129, 113, 98, 
    118, 115, 126, 128, 126, 123, 121, 119, 120, 120, 117, 110, 107, 105, 103, 105, 104, 102, 98, 95, 96, 96, 93, 89, 87, 87, 88, 90, 81, 59, 65, 69, 
    95, 69, 73, 77, 76, 75, 78, 80, 82, 83, 81, 74, 71, 75, 81, 83, 83, 85, 86, 84, 80, 80, 82, 83, 80, 78, 75, 60, 48, 65, 96, 103, 
    96, 75, 80, 80, 80, 80, 79, 81, 84, 85, 78, 63, 61, 62, 66, 70, 68, 68, 67, 66, 67, 73, 78, 80, 84, 75, 57, 50, 79, 115, 138, 125, 
    92, 70, 77, 77, 70, 68, 67, 71, 74, 75, 70, 59, 51, 56, 61, 66, 65, 58, 54, 52, 58, 68, 81, 87, 82, 67, 68, 94, 120, 133, 118, 88, 
    138, 112, 121, 123, 120, 116, 114, 115, 118, 119, 123, 133, 135, 134, 133, 137, 142, 140, 137, 135, 130, 122, 124, 125, 127, 137, 154, 169, 167, 140, 127, 118, 
    
    -- channel=52
    0, 102, 138, 150, 160, 145, 119, 113, 114, 120, 128, 130, 128, 125, 125, 120, 121, 121, 119, 122, 123, 124, 126, 124, 124, 125, 129, 140, 150, 152, 153, 154, 
    0, 180, 232, 248, 268, 256, 228, 214, 205, 207, 226, 237, 234, 232, 231, 223, 226, 228, 226, 228, 229, 233, 235, 231, 231, 229, 235, 249, 255, 252, 259, 277, 
    0, 188, 239, 252, 276, 275, 252, 224, 188, 187, 215, 231, 232, 229, 227, 215, 222, 233, 223, 227, 233, 229, 234, 224, 218, 241, 252, 264, 268, 262, 268, 288, 
    0, 189, 233, 244, 263, 275, 280, 241, 181, 186, 206, 203, 205, 204, 206, 200, 207, 215, 206, 210, 220, 212, 212, 201, 199, 245, 264, 266, 266, 263, 269, 289, 
    0, 190, 230, 240, 259, 276, 295, 253, 188, 202, 201, 193, 210, 208, 191, 187, 207, 218, 211, 217, 225, 213, 222, 202, 202, 258, 272, 269, 268, 268, 275, 293, 
    0, 188, 225, 236, 255, 277, 297, 226, 179, 220, 209, 194, 209, 203, 188, 187, 207, 218, 213, 226, 221, 208, 223, 202, 197, 225, 246, 264, 267, 267, 276, 294, 
    0, 189, 224, 235, 258, 280, 277, 198, 167, 209, 206, 198, 207, 202, 192, 193, 206, 210, 214, 222, 211, 199, 207, 211, 216, 198, 226, 263, 265, 264, 276, 295, 
    0, 198, 227, 236, 256, 277, 267, 203, 184, 203, 212, 210, 217, 209, 200, 205, 213, 215, 220, 229, 211, 203, 207, 227, 230, 189, 215, 259, 265, 261, 273, 292, 
    0, 210, 233, 234, 260, 277, 266, 233, 216, 206, 217, 207, 208, 208, 206, 214, 218, 222, 224, 226, 209, 198, 196, 220, 241, 218, 230, 260, 265, 263, 270, 288, 
    0, 222, 243, 236, 256, 257, 254, 255, 239, 212, 213, 211, 210, 213, 215, 220, 222, 226, 225, 221, 216, 205, 209, 221, 245, 258, 257, 262, 262, 262, 269, 287, 
    0, 230, 252, 239, 255, 252, 253, 264, 250, 228, 230, 226, 228, 229, 232, 240, 242, 244, 240, 235, 228, 225, 226, 227, 245, 265, 263, 260, 260, 261, 268, 287, 
    0, 229, 257, 242, 245, 228, 220, 242, 257, 247, 248, 246, 244, 249, 254, 259, 261, 257, 250, 246, 243, 241, 245, 247, 253, 263, 263, 263, 262, 262, 271, 289, 
    0, 228, 263, 248, 230, 189, 158, 170, 208, 235, 254, 263, 265, 266, 269, 275, 276, 274, 269, 267, 264, 262, 263, 264, 263, 263, 262, 263, 262, 261, 270, 289, 
    0, 227, 274, 269, 247, 204, 152, 123, 133, 163, 204, 238, 258, 267, 272, 276, 277, 274, 271, 269, 264, 260, 262, 263, 262, 261, 261, 264, 264, 262, 271, 288, 
    0, 227, 276, 275, 260, 237, 207, 151, 109, 100, 130, 179, 221, 252, 271, 276, 275, 271, 269, 269, 264, 259, 260, 264, 265, 264, 264, 264, 262, 261, 270, 286, 
    0, 228, 274, 274, 279, 271, 264, 231, 171, 107, 69, 94, 143, 189, 231, 260, 272, 273, 271, 267, 261, 257, 259, 261, 261, 261, 263, 263, 261, 260, 270, 287, 
    0, 229, 274, 271, 278, 272, 271, 276, 253, 172, 74, 45, 70, 103, 147, 188, 223, 247, 260, 264, 264, 260, 261, 265, 265, 264, 265, 264, 262, 261, 272, 290, 
    0, 229, 272, 266, 276, 273, 270, 273, 283, 232, 97, 33, 41, 42, 66, 101, 134, 163, 190, 215, 234, 244, 259, 272, 269, 266, 264, 261, 260, 260, 271, 290, 
    0, 228, 270, 262, 273, 272, 272, 271, 279, 248, 102, 17, 26, 26, 34, 47, 62, 81, 101, 124, 141, 153, 184, 219, 236, 247, 257, 262, 263, 263, 274, 291, 
    0, 227, 272, 261, 269, 271, 275, 270, 274, 223, 90, 11, 9, 18, 32, 38, 40, 41, 47, 60, 65, 63, 85, 121, 141, 162, 193, 218, 239, 254, 272, 292, 
    0, 223, 275, 265, 267, 270, 273, 277, 267, 204, 114, 55, 23, 7, 20, 33, 66, 92, 86, 64, 32, 32, 43, 54, 64, 95, 157, 199, 218, 237, 259, 288, 
    0, 220, 277, 269, 267, 268, 274, 286, 273, 217, 188, 164, 107, 76, 77, 81, 125, 170, 174, 138, 100, 111, 116, 105, 82, 99, 160, 197, 216, 232, 251, 282, 
    0, 211, 267, 262, 257, 255, 256, 262, 251, 219, 220, 232, 185, 142, 139, 132, 171, 222, 234, 198, 157, 180, 195, 179, 153, 156, 200, 225, 226, 227, 239, 271, 
    0, 158, 202, 201, 193, 189, 184, 181, 179, 176, 177, 185, 167, 146, 150, 158, 183, 211, 216, 208, 190, 195, 205, 209, 205, 208, 218, 227, 229, 222, 224, 246, 
    0, 131, 167, 170, 166, 164, 158, 155, 152, 146, 144, 145, 141, 143, 146, 155, 168, 177, 172, 170, 174, 173, 171, 174, 183, 188, 186, 186, 184, 171, 169, 186, 
    0, 100, 117, 125, 124, 121, 112, 103, 94, 87, 84, 84, 83, 83, 84, 88, 100, 108, 101, 93, 93, 93, 91, 90, 93, 96, 99, 104, 101, 85, 79, 105, 
    0, 66, 71, 76, 80, 81, 76, 68, 59, 55, 51, 49, 48, 49, 50, 50, 49, 53, 48, 40, 37, 36, 36, 35, 37, 37, 38, 39, 33, 19, 24, 70, 
    0, 44, 36, 41, 41, 43, 39, 26, 21, 20, 15, 14, 16, 14, 11, 11, 9, 11, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 63, 
    0, 21, 3, 9, 6, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 28, 55, 
    0, 20, 3, 8, 6, 9, 6, 1, 2, 2, 1, 5, 15, 15, 9, 4, 6, 14, 12, 8, 5, 2, 0, 0, 0, 0, 0, 14, 31, 35, 33, 35, 
    0, 16, 0, 0, 0, 5, 6, 2, 0, 0, 0, 0, 11, 14, 8, 2, 5, 12, 12, 11, 11, 7, 0, 0, 0, 0, 6, 31, 41, 32, 10, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    73, 114, 122, 121, 117, 110, 113, 118, 117, 118, 122, 125, 125, 125, 123, 125, 124, 121, 123, 125, 128, 129, 126, 127, 128, 130, 136, 135, 136, 140, 140, 69, 
    190, 212, 226, 226, 212, 204, 191, 189, 198, 207, 210, 212, 215, 207, 206, 204, 206, 209, 208, 209, 210, 210, 211, 210, 212, 219, 228, 240, 249, 253, 235, 70, 
    190, 213, 225, 229, 211, 204, 192, 171, 188, 202, 201, 202, 208, 199, 202, 209, 206, 206, 211, 211, 212, 214, 212, 213, 227, 233, 243, 247, 248, 253, 236, 68, 
    187, 214, 227, 235, 232, 222, 196, 167, 163, 164, 179, 192, 195, 195, 185, 189, 192, 195, 198, 202, 199, 200, 203, 205, 226, 247, 249, 248, 247, 255, 239, 69, 
    184, 212, 227, 233, 235, 227, 180, 150, 155, 154, 157, 153, 141, 139, 149, 157, 162, 160, 164, 168, 163, 164, 163, 190, 202, 227, 245, 248, 245, 251, 233, 64, 
    183, 208, 226, 231, 234, 222, 161, 159, 166, 154, 146, 143, 142, 137, 142, 150, 151, 157, 168, 156, 166, 168, 156, 196, 213, 238, 256, 255, 255, 256, 237, 67, 
    181, 206, 222, 226, 228, 208, 157, 158, 148, 156, 162, 167, 172, 157, 151, 164, 170, 181, 186, 183, 182, 190, 194, 198, 201, 220, 241, 248, 250, 253, 235, 65, 
    181, 203, 219, 223, 226, 200, 152, 140, 142, 158, 161, 160, 152, 159, 153, 157, 156, 169, 168, 156, 162, 161, 178, 162, 176, 194, 219, 244, 249, 252, 231, 62, 
    186, 202, 217, 223, 220, 195, 166, 152, 161, 170, 163, 173, 168, 180, 177, 172, 166, 171, 170, 158, 167, 166, 195, 185, 186, 210, 229, 239, 238, 245, 229, 62, 
    194, 210, 219, 221, 219, 218, 215, 199, 190, 189, 191, 190, 192, 190, 193, 194, 191, 197, 203, 196, 193, 197, 206, 215, 219, 228, 238, 243, 242, 246, 229, 63, 
    207, 216, 228, 226, 224, 227, 225, 205, 196, 188, 191, 189, 183, 190, 195, 196, 197, 193, 191, 190, 196, 195, 206, 226, 234, 239, 241, 246, 244, 246, 228, 63, 
    219, 228, 233, 223, 223, 227, 231, 222, 215, 213, 209, 212, 215, 218, 220, 220, 215, 214, 217, 218, 222, 224, 226, 237, 241, 239, 238, 240, 239, 243, 228, 63, 
    225, 237, 231, 215, 199, 195, 197, 220, 248, 249, 241, 233, 232, 236, 238, 237, 235, 234, 233, 233, 233, 236, 238, 236, 238, 241, 242, 244, 247, 252, 233, 66, 
    227, 244, 227, 201, 169, 153, 157, 157, 180, 214, 241, 250, 242, 238, 239, 239, 240, 241, 239, 237, 238, 240, 239, 241, 243, 244, 245, 245, 245, 249, 230, 62, 
    230, 249, 231, 206, 197, 180, 161, 142, 128, 152, 186, 219, 245, 250, 246, 245, 245, 247, 246, 242, 240, 241, 241, 239, 238, 238, 237, 237, 237, 240, 222, 60, 
    232, 253, 257, 247, 241, 219, 183, 159, 129, 113, 147, 181, 213, 250, 265, 258, 247, 242, 239, 236, 238, 238, 238, 237, 238, 238, 238, 237, 237, 239, 221, 59, 
    233, 257, 263, 255, 257, 258, 241, 196, 147, 107, 103, 143, 170, 192, 220, 249, 258, 253, 246, 236, 233, 237, 239, 236, 238, 239, 239, 239, 239, 241, 221, 58, 
    236, 258, 267, 263, 263, 264, 263, 239, 159, 102, 90, 95, 118, 147, 166, 182, 207, 230, 243, 245, 242, 243, 240, 237, 238, 238, 239, 240, 240, 241, 222, 58, 
    238, 260, 268, 265, 264, 265, 260, 254, 176, 98, 87, 83, 89, 98, 115, 135, 148, 162, 175, 184, 203, 226, 248, 257, 253, 249, 244, 239, 236, 238, 219, 55, 
    239, 257, 265, 261, 261, 263, 258, 249, 171, 104, 68, 52, 71, 76, 80, 88, 99, 113, 120, 112, 117, 143, 172, 198, 223, 242, 249, 253, 250, 245, 220, 56, 
    239, 255, 260, 259, 259, 260, 260, 229, 158, 85, 53, 29, 30, 61, 79, 99, 101, 79, 59, 57, 83, 93, 99, 124, 159, 188, 194, 199, 217, 236, 222, 55, 
    238, 252, 251, 254, 257, 258, 255, 212, 161, 115, 86, 78, 65, 49, 68, 92, 121, 139, 115, 90, 72, 91, 94, 80, 105, 137, 181, 210, 212, 222, 214, 50, 
    231, 249, 249, 249, 253, 255, 249, 218, 204, 217, 193, 148, 137, 118, 143, 188, 204, 196, 159, 164, 164, 155, 145, 144, 172, 197, 204, 211, 221, 230, 218, 54, 
    203, 232, 238, 235, 237, 237, 236, 234, 230, 234, 218, 189, 185, 191, 201, 222, 220, 202, 178, 181, 199, 199, 185, 184, 197, 204, 196, 189, 185, 195, 193, 48, 
    175, 169, 155, 156, 149, 146, 144, 140, 137, 137, 134, 134, 131, 128, 130, 132, 139, 143, 146, 148, 145, 146, 152, 156, 151, 148, 147, 148, 145, 154, 155, 31, 
    118, 126, 122, 115, 111, 111, 112, 114, 116, 117, 115, 111, 107, 109, 117, 126, 123, 122, 120, 119, 121, 121, 123, 124, 126, 128, 127, 124, 120, 120, 130, 30, 
    112, 123, 123, 122, 118, 117, 115, 112, 114, 112, 108, 103, 104, 104, 100, 104, 104, 100, 97, 92, 91, 88, 87, 88, 86, 87, 87, 82, 81, 93, 108, 18, 
    94, 87, 82, 82, 81, 75, 74, 78, 78, 76, 74, 68, 64, 65, 69, 71, 74, 70, 68, 67, 64, 63, 63, 63, 64, 64, 64, 68, 83, 100, 107, 44, 
    65, 68, 66, 64, 65, 65, 63, 67, 68, 67, 62, 60, 62, 63, 65, 70, 72, 70, 67, 63, 64, 65, 67, 64, 60, 60, 73, 91, 103, 126, 149, 66, 
    66, 64, 61, 62, 58, 57, 60, 63, 63, 62, 62, 61, 54, 58, 62, 68, 70, 66, 63, 62, 59, 60, 67, 70, 72, 86, 100, 111, 133, 152, 127, 28, 
    61, 61, 61, 63, 61, 58, 60, 61, 63, 62, 67, 73, 80, 78, 79, 84, 84, 83, 80, 81, 77, 72, 70, 78, 94, 108, 124, 147, 147, 102, 80, 22, 
    37, 67, 57, 61, 58, 57, 57, 58, 57, 60, 71, 73, 73, 72, 73, 79, 77, 77, 76, 75, 66, 64, 61, 65, 87, 124, 150, 123, 76, 63, 66, 21, 
    
    -- channel=54
    32, 40, 38, 49, 56, 43, 43, 45, 42, 43, 44, 46, 44, 49, 44, 45, 48, 43, 44, 44, 44, 47, 45, 46, 45, 42, 43, 47, 47, 44, 63, 157, 
    0, 0, 0, 0, 12, 9, 6, 9, 0, 0, 0, 5, 2, 8, 3, 0, 7, 5, 3, 2, 0, 5, 3, 3, 2, 0, 0, 1, 1, 0, 18, 148, 
    0, 0, 0, 0, 0, 9, 25, 16, 0, 3, 1, 7, 12, 9, 11, 3, 8, 10, 6, 7, 8, 8, 8, 0, 0, 0, 0, 0, 0, 0, 13, 144, 
    0, 0, 0, 0, 0, 0, 29, 12, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 0, 0, 0, 0, 0, 0, 15, 146, 
    0, 0, 0, 0, 0, 0, 29, 18, 12, 18, 2, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 12, 145, 
    0, 0, 0, 0, 0, 3, 31, 0, 12, 24, 20, 18, 31, 28, 18, 10, 22, 20, 22, 31, 18, 22, 25, 19, 0, 0, 0, 0, 0, 0, 13, 146, 
    0, 0, 0, 0, 0, 17, 25, 0, 0, 6, 11, 4, 13, 8, 5, 4, 6, 0, 5, 13, 0, 8, 0, 10, 0, 0, 0, 0, 0, 0, 10, 143, 
    0, 0, 0, 0, 0, 4, 5, 14, 0, 0, 1, 0, 4, 3, 5, 2, 0, 0, 0, 3, 0, 0, 0, 9, 6, 0, 0, 0, 0, 0, 8, 141, 
    0, 0, 0, 0, 0, 0, 11, 27, 15, 9, 7, 7, 10, 9, 11, 8, 11, 12, 13, 17, 12, 13, 2, 6, 20, 2, 0, 0, 0, 0, 10, 140, 
    0, 0, 0, 0, 0, 0, 3, 11, 0, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 10, 139, 
    0, 3, 0, 0, 0, 0, 0, 5, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 10, 140, 
    0, 0, 0, 0, 0, 0, 0, 5, 6, 2, 3, 3, 1, 0, 0, 0, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 11, 142, 
    0, 0, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 141, 
    0, 0, 10, 16, 21, 32, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 139, 
    0, 0, 0, 9, 17, 44, 57, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 137, 
    0, 0, 0, 0, 0, 12, 38, 71, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 138, 
    0, 0, 0, 0, 0, 0, 1, 34, 85, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 138, 
    0, 0, 0, 0, 0, 0, 0, 3, 70, 66, 11, 18, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 136, 
    0, 0, 0, 0, 0, 0, 0, 0, 57, 62, 15, 19, 20, 19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 136, 
    0, 0, 0, 0, 0, 0, 0, 14, 45, 59, 29, 9, 14, 18, 17, 23, 21, 15, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 138, 
    0, 0, 0, 0, 0, 0, 0, 28, 34, 51, 62, 30, 7, 17, 3, 11, 35, 41, 45, 23, 28, 15, 0, 0, 0, 0, 0, 0, 0, 0, 4, 138, 
    0, 0, 0, 0, 0, 0, 0, 25, 34, 35, 65, 70, 28, 29, 8, 0, 25, 45, 62, 24, 26, 44, 45, 30, 0, 0, 6, 0, 0, 0, 4, 133, 
    0, 0, 0, 0, 0, 0, 0, 4, 15, 9, 25, 51, 41, 32, 20, 0, 0, 12, 37, 29, 10, 16, 33, 33, 12, 0, 0, 0, 0, 0, 4, 128, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 
    12, 10, 9, 12, 14, 14, 14, 15, 17, 18, 17, 19, 16, 11, 9, 0, 2, 6, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 
    10, 4, 5, 5, 5, 8, 7, 4, 8, 9, 9, 8, 8, 8, 7, 6, 5, 12, 11, 8, 7, 8, 8, 8, 6, 5, 6, 8, 5, 0, 3, 91, 
    24, 11, 9, 10, 10, 13, 15, 14, 20, 22, 22, 19, 18, 17, 18, 17, 17, 23, 26, 26, 24, 23, 24, 27, 27, 26, 24, 21, 16, 20, 33, 96, 
    38, 27, 25, 25, 26, 27, 25, 25, 29, 31, 31, 28, 30, 29, 28, 28, 30, 31, 32, 32, 32, 31, 31, 30, 31, 26, 17, 15, 26, 31, 26, 83, 
    36, 26, 25, 26, 25, 28, 27, 27, 27, 29, 27, 29, 29, 30, 28, 27, 33, 32, 33, 31, 33, 29, 30, 28, 21, 16, 18, 27, 30, 29, 23, 79, 
    40, 29, 27, 28, 28, 28, 30, 28, 30, 30, 23, 28, 28, 30, 29, 25, 30, 30, 31, 31, 36, 29, 28, 27, 18, 21, 28, 30, 27, 27, 28, 78, 
    17, 23, 19, 20, 18, 17, 18, 18, 18, 19, 12, 11, 15, 17, 18, 15, 15, 16, 15, 17, 23, 22, 20, 18, 12, 13, 18, 18, 20, 20, 17, 55, 
    
    -- channel=55
    191, 35, 17, 14, 0, 0, 6, 7, 8, 10, 6, 0, 0, 0, 0, 2, 0, 0, 2, 0, 2, 0, 0, 0, 0, 4, 9, 5, 0, 0, 0, 0, 
    259, 69, 53, 51, 22, 6, 25, 26, 25, 39, 41, 32, 22, 25, 16, 29, 31, 22, 28, 27, 29, 28, 21, 24, 26, 31, 36, 27, 18, 20, 11, 0, 
    262, 75, 58, 55, 36, 19, 10, 0, 11, 46, 31, 27, 14, 10, 11, 21, 26, 13, 15, 18, 17, 16, 12, 17, 32, 33, 33, 26, 20, 21, 12, 0, 
    266, 73, 57, 56, 43, 24, 0, 0, 0, 28, 0, 13, 8, 0, 5, 9, 11, 0, 3, 9, 4, 3, 2, 4, 53, 43, 23, 25, 24, 21, 12, 0, 
    266, 73, 56, 53, 47, 37, 0, 0, 7, 8, 0, 10, 5, 0, 1, 11, 10, 0, 4, 9, 0, 5, 6, 4, 60, 43, 22, 25, 24, 22, 14, 0, 
    264, 72, 57, 51, 46, 39, 0, 0, 30, 0, 0, 16, 5, 0, 1, 13, 18, 7, 15, 8, 0, 16, 6, 11, 38, 39, 33, 24, 22, 24, 14, 0, 
    264, 68, 56, 54, 45, 22, 0, 0, 30, 6, 4, 13, 4, 0, 5, 13, 14, 4, 18, 0, 0, 18, 2, 16, 0, 36, 59, 31, 24, 27, 17, 0, 
    268, 62, 52, 55, 41, 8, 0, 0, 7, 10, 11, 6, 8, 0, 13, 13, 7, 6, 13, 0, 0, 15, 6, 28, 0, 29, 60, 32, 24, 28, 21, 0, 
    276, 54, 45, 55, 40, 21, 7, 9, 2, 22, 23, 24, 25, 17, 25, 23, 25, 22, 17, 10, 10, 25, 26, 42, 15, 26, 44, 36, 29, 29, 22, 0, 
    286, 50, 33, 54, 42, 37, 33, 17, 10, 39, 32, 37, 40, 37, 42, 37, 36, 32, 32, 28, 30, 39, 35, 51, 50, 28, 30, 30, 28, 29, 22, 0, 
    293, 51, 25, 49, 33, 32, 41, 25, 15, 36, 31, 32, 36, 36, 36, 32, 31, 29, 28, 30, 29, 35, 34, 44, 50, 30, 27, 26, 29, 32, 23, 0, 
    297, 51, 15, 29, 19, 25, 60, 55, 23, 27, 26, 28, 32, 31, 31, 26, 23, 21, 24, 26, 26, 28, 27, 32, 38, 33, 30, 29, 30, 30, 21, 0, 
    298, 49, 12, 7, 8, 10, 48, 81, 63, 53, 39, 30, 31, 34, 35, 31, 28, 28, 29, 26, 27, 31, 31, 28, 28, 29, 28, 26, 24, 26, 17, 0, 
    299, 51, 18, 9, 4, 0, 0, 43, 72, 82, 75, 54, 39, 35, 32, 29, 26, 25, 24, 20, 23, 28, 28, 25, 27, 28, 28, 28, 27, 29, 19, 0, 
    300, 56, 17, 13, 4, 0, 0, 0, 14, 64, 93, 91, 70, 47, 30, 23, 22, 22, 23, 19, 21, 28, 29, 27, 28, 29, 27, 27, 28, 32, 21, 0, 
    301, 61, 25, 30, 20, 8, 0, 0, 0, 0, 70, 94, 89, 79, 58, 35, 23, 19, 20, 20, 21, 26, 27, 26, 27, 29, 26, 27, 29, 32, 23, 0, 
    303, 61, 22, 29, 22, 19, 10, 0, 0, 0, 16, 76, 72, 81, 80, 68, 52, 38, 28, 21, 20, 27, 29, 24, 27, 29, 27, 28, 29, 30, 24, 0, 
    305, 59, 19, 27, 18, 17, 16, 8, 0, 0, 0, 53, 43, 63, 72, 71, 67, 60, 54, 42, 35, 44, 41, 25, 24, 25, 25, 27, 29, 29, 23, 0, 
    304, 58, 15, 25, 17, 17, 16, 10, 0, 0, 0, 51, 35, 46, 51, 55, 57, 58, 56, 52, 50, 75, 80, 52, 39, 34, 29, 25, 26, 28, 21, 0, 
    302, 55, 11, 21, 17, 19, 17, 0, 0, 0, 0, 42, 53, 52, 42, 39, 34, 39, 46, 45, 52, 82, 95, 67, 59, 62, 54, 47, 41, 33, 20, 0, 
    299, 58, 15, 20, 19, 23, 16, 0, 0, 0, 0, 0, 29, 55, 54, 80, 60, 17, 0, 3, 50, 54, 56, 55, 82, 111, 75, 51, 53, 44, 26, 0, 
    295, 60, 21, 23, 21, 22, 20, 1, 0, 0, 0, 0, 0, 47, 45, 79, 69, 11, 0, 0, 44, 36, 11, 11, 48, 91, 60, 35, 41, 37, 27, 0, 
    287, 60, 24, 22, 18, 18, 17, 4, 0, 8, 7, 0, 0, 18, 23, 50, 50, 11, 0, 0, 32, 25, 5, 0, 24, 51, 35, 25, 32, 32, 26, 0, 
    246, 54, 36, 27, 26, 26, 28, 29, 30, 34, 34, 15, 17, 34, 43, 58, 53, 36, 31, 30, 42, 42, 38, 35, 40, 44, 45, 46, 46, 45, 40, 0, 
    220, 53, 56, 45, 44, 44, 47, 47, 46, 49, 53, 47, 52, 56, 59, 66, 62, 49, 54, 60, 56, 54, 59, 63, 59, 54, 55, 53, 52, 55, 53, 0, 
    188, 32, 47, 37, 35, 31, 33, 33, 33, 34, 32, 31, 35, 39, 47, 51, 54, 41, 40, 49, 50, 50, 50, 55, 56, 56, 55, 52, 45, 51, 60, 6, 
    170, 24, 52, 44, 42, 41, 39, 41, 44, 39, 38, 43, 46, 47, 50, 49, 52, 44, 38, 43, 47, 48, 48, 49, 48, 49, 50, 45, 41, 60, 78, 14, 
    149, 16, 54, 44, 45, 44, 38, 42, 42, 31, 32, 37, 41, 42, 42, 42, 42, 38, 30, 32, 36, 40, 41, 39, 36, 38, 38, 43, 57, 71, 62, 0, 
    132, 2, 43, 32, 36, 36, 32, 38, 37, 27, 30, 35, 40, 36, 35, 37, 37, 33, 30, 32, 36, 37, 38, 37, 35, 36, 48, 65, 65, 48, 31, 0, 
    132, 5, 46, 36, 40, 39, 35, 39, 36, 34, 41, 46, 40, 33, 33, 39, 39, 29, 30, 31, 30, 27, 33, 29, 35, 54, 69, 62, 41, 23, 15, 0, 
    129, 1, 41, 34, 40, 39, 35, 35, 34, 32, 36, 45, 33, 27, 26, 31, 33, 25, 28, 27, 25, 19, 31, 36, 51, 68, 59, 40, 18, 12, 23, 1, 
    101, 17, 42, 37, 41, 41, 40, 38, 38, 37, 41, 50, 40, 37, 37, 39, 41, 37, 39, 37, 34, 28, 38, 41, 51, 67, 55, 26, 19, 30, 38, 28, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=57
    75, 122, 152, 158, 148, 140, 124, 117, 117, 117, 116, 113, 112, 109, 109, 108, 107, 108, 109, 110, 111, 111, 110, 109, 108, 110, 114, 117, 123, 129, 103, 52, 
    119, 191, 231, 242, 232, 208, 180, 160, 160, 172, 179, 181, 174, 169, 168, 168, 167, 167, 168, 169, 171, 170, 169, 168, 169, 173, 177, 179, 183, 190, 155, 105, 
    136, 216, 261, 266, 257, 221, 149, 103, 83, 107, 141, 144, 139, 133, 129, 136, 135, 137, 140, 138, 144, 146, 135, 156, 169, 185, 202, 196, 194, 199, 167, 115, 
    141, 220, 261, 261, 264, 232, 126, 57, 0, 18, 44, 35, 40, 32, 30, 34, 34, 35, 42, 45, 53, 57, 41, 83, 126, 177, 208, 194, 191, 196, 165, 114, 
    149, 219, 259, 263, 269, 235, 131, 58, 0, 2, 8, 0, 1, 0, 0, 0, 4, 14, 21, 28, 36, 34, 25, 59, 120, 184, 208, 199, 198, 202, 168, 112, 
    146, 212, 253, 261, 269, 220, 111, 54, 12, 37, 28, 21, 12, 0, 0, 10, 28, 50, 48, 54, 57, 48, 62, 62, 108, 164, 190, 203, 204, 205, 170, 113, 
    146, 213, 254, 259, 254, 180, 50, 0, 0, 29, 32, 46, 25, 5, 0, 12, 32, 51, 43, 40, 34, 34, 62, 47, 72, 114, 160, 202, 209, 212, 177, 117, 
    149, 214, 255, 258, 246, 178, 55, 0, 0, 48, 57, 64, 52, 42, 31, 36, 44, 50, 49, 34, 19, 31, 54, 54, 62, 95, 160, 205, 216, 220, 186, 123, 
    152, 217, 255, 256, 251, 213, 139, 98, 101, 118, 124, 119, 122, 125, 120, 115, 114, 116, 114, 100, 80, 91, 112, 126, 123, 142, 191, 216, 222, 226, 193, 127, 
    155, 217, 253, 253, 255, 245, 223, 203, 189, 182, 183, 183, 185, 188, 186, 181, 183, 188, 187, 178, 164, 166, 179, 194, 196, 201, 217, 225, 226, 230, 196, 129, 
    155, 215, 249, 247, 254, 253, 246, 234, 219, 213, 210, 209, 208, 208, 207, 205, 205, 209, 211, 206, 198, 196, 200, 213, 225, 223, 222, 219, 222, 229, 195, 128, 
    147, 209, 239, 233, 229, 224, 227, 229, 228, 227, 226, 222, 220, 219, 219, 219, 218, 218, 217, 219, 214, 211, 213, 218, 227, 225, 221, 216, 219, 225, 190, 125, 
    139, 201, 229, 216, 200, 176, 172, 186, 204, 221, 231, 234, 232, 231, 232, 232, 231, 229, 228, 227, 226, 223, 223, 223, 224, 224, 222, 218, 218, 221, 184, 121, 
    134, 197, 235, 217, 192, 149, 119, 124, 142, 173, 199, 215, 221, 224, 226, 226, 225, 222, 220, 217, 216, 216, 219, 219, 220, 221, 221, 217, 217, 221, 184, 122, 
    134, 199, 240, 226, 206, 170, 124, 95, 94, 119, 154, 183, 201, 211, 216, 218, 214, 211, 209, 207, 205, 206, 211, 216, 220, 220, 220, 218, 220, 227, 193, 127, 
    136, 199, 238, 228, 222, 203, 170, 124, 91, 88, 102, 128, 153, 175, 191, 202, 207, 207, 207, 206, 204, 205, 209, 214, 218, 220, 222, 221, 225, 234, 201, 132, 
    137, 197, 230, 219, 217, 209, 192, 169, 122, 88, 72, 70, 88, 114, 140, 161, 178, 190, 199, 203, 206, 210, 213, 216, 218, 221, 224, 223, 227, 236, 204, 135, 
    136, 187, 215, 204, 205, 201, 191, 187, 152, 98, 59, 39, 38, 52, 76, 99, 119, 138, 156, 172, 190, 204, 212, 216, 217, 219, 221, 219, 222, 231, 202, 134, 
    130, 176, 201, 190, 194, 195, 192, 185, 157, 103, 49, 28, 23, 25, 32, 43, 56, 71, 90, 112, 135, 157, 174, 184, 191, 199, 209, 211, 216, 225, 197, 131, 
    123, 171, 195, 185, 191, 195, 195, 176, 148, 90, 38, 28, 23, 22, 23, 21, 24, 33, 46, 63, 78, 97, 109, 116, 127, 144, 167, 183, 199, 215, 194, 128, 
    119, 172, 196, 190, 193, 198, 196, 171, 140, 90, 49, 40, 37, 27, 30, 37, 46, 54, 51, 54, 53, 57, 60, 62, 80, 107, 137, 160, 178, 198, 187, 124, 
    117, 177, 204, 196, 194, 199, 195, 181, 149, 123, 109, 91, 85, 75, 73, 87, 102, 111, 102, 97, 94, 92, 87, 83, 93, 118, 141, 158, 173, 190, 183, 124, 
    113, 177, 202, 193, 187, 188, 187, 182, 163, 157, 163, 153, 135, 131, 126, 138, 161, 172, 168, 149, 155, 162, 157, 150, 149, 169, 185, 191, 192, 199, 190, 128, 
    94, 148, 170, 163, 153, 152, 152, 150, 149, 150, 155, 155, 149, 150, 154, 164, 182, 195, 202, 194, 195, 199, 203, 204, 205, 214, 220, 224, 219, 217, 198, 134, 
    78, 125, 150, 146, 141, 143, 141, 138, 137, 135, 137, 139, 143, 148, 155, 166, 176, 183, 188, 189, 190, 189, 192, 198, 203, 206, 206, 203, 196, 192, 167, 114, 
    62, 98, 125, 124, 122, 122, 117, 110, 103, 98, 100, 101, 104, 109, 114, 122, 128, 127, 124, 122, 122, 122, 123, 126, 127, 129, 131, 124, 114, 116, 100, 71, 
    41, 64, 85, 85, 86, 88, 84, 75, 66, 59, 55, 56, 61, 63, 66, 66, 65, 60, 54, 52, 51, 52, 52, 53, 54, 54, 54, 49, 46, 66, 67, 58, 
    21, 30, 46, 43, 42, 42, 38, 29, 21, 16, 18, 24, 28, 27, 24, 22, 21, 19, 16, 14, 13, 13, 14, 15, 16, 17, 20, 25, 41, 70, 75, 70, 
    2, 5, 19, 19, 17, 18, 15, 9, 6, 3, 6, 12, 15, 13, 7, 6, 7, 10, 11, 10, 8, 9, 10, 9, 8, 16, 37, 59, 78, 95, 80, 57, 
    1, 3, 18, 22, 21, 22, 18, 15, 13, 11, 16, 20, 23, 19, 14, 11, 12, 16, 16, 15, 14, 12, 8, 5, 13, 35, 70, 93, 99, 88, 46, 22, 
    0, 0, 9, 13, 14, 17, 15, 11, 6, 3, 8, 12, 15, 12, 6, 5, 7, 9, 10, 10, 9, 5, 2, 9, 34, 64, 91, 99, 83, 49, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 24, 48, 63, 57, 31, 5, 0, 0, 
    
    -- channel=58
    202, 199, 218, 219, 188, 176, 178, 178, 183, 189, 193, 191, 190, 183, 182, 186, 183, 184, 185, 187, 192, 191, 189, 189, 192, 206, 222, 228, 229, 233, 207, 13, 
    321, 305, 330, 335, 305, 285, 284, 277, 282, 297, 309, 312, 311, 303, 297, 304, 304, 304, 307, 308, 313, 310, 306, 304, 309, 323, 337, 342, 342, 350, 312, 14, 
    325, 316, 341, 347, 327, 306, 266, 233, 246, 276, 287, 286, 282, 271, 271, 286, 287, 287, 290, 291, 297, 291, 283, 303, 316, 337, 353, 352, 350, 357, 318, 16, 
    323, 312, 336, 344, 339, 322, 261, 218, 222, 237, 235, 234, 233, 224, 228, 240, 241, 236, 244, 246, 245, 247, 236, 273, 320, 341, 348, 349, 347, 354, 317, 15, 
    322, 311, 333, 339, 341, 334, 259, 220, 234, 232, 225, 235, 231, 222, 226, 244, 251, 249, 261, 261, 255, 261, 255, 287, 338, 350, 350, 355, 354, 359, 321, 16, 
    319, 307, 329, 334, 340, 319, 236, 220, 234, 225, 224, 236, 217, 207, 217, 240, 245, 254, 260, 254, 254, 256, 254, 267, 308, 332, 339, 350, 354, 360, 321, 15, 
    319, 304, 327, 331, 332, 286, 207, 205, 228, 224, 223, 240, 219, 209, 219, 235, 237, 240, 249, 230, 234, 241, 254, 247, 259, 309, 340, 349, 348, 355, 318, 16, 
    323, 301, 325, 329, 323, 281, 223, 219, 239, 246, 245, 252, 246, 241, 245, 251, 250, 259, 263, 238, 245, 253, 271, 269, 259, 304, 340, 345, 346, 353, 317, 17, 
    335, 301, 321, 328, 326, 305, 276, 250, 248, 256, 257, 258, 255, 254, 259, 264, 267, 268, 263, 245, 248, 257, 280, 293, 291, 321, 346, 347, 344, 351, 315, 17, 
    354, 308, 323, 329, 328, 325, 315, 281, 269, 275, 270, 274, 274, 278, 286, 286, 284, 283, 282, 272, 277, 283, 297, 326, 333, 335, 342, 345, 342, 349, 314, 18, 
    370, 318, 331, 336, 326, 329, 329, 305, 297, 300, 299, 299, 300, 308, 313, 314, 313, 309, 305, 303, 305, 307, 316, 341, 348, 340, 339, 342, 343, 351, 315, 18, 
    380, 329, 321, 308, 284, 287, 320, 324, 319, 319, 315, 318, 322, 327, 331, 328, 322, 318, 319, 319, 321, 323, 326, 341, 348, 345, 346, 348, 348, 355, 319, 18, 
    385, 336, 311, 275, 238, 215, 240, 280, 309, 332, 337, 337, 339, 345, 349, 348, 346, 345, 342, 339, 339, 344, 345, 343, 344, 346, 344, 344, 345, 353, 315, 17, 
    388, 345, 329, 298, 265, 222, 197, 203, 229, 273, 314, 335, 345, 351, 354, 353, 350, 349, 345, 338, 337, 340, 340, 338, 339, 341, 342, 342, 342, 349, 312, 15, 
    392, 351, 337, 314, 299, 263, 218, 181, 175, 206, 255, 304, 339, 354, 355, 352, 348, 347, 344, 337, 336, 341, 342, 340, 342, 342, 340, 339, 339, 346, 308, 15, 
    396, 359, 364, 357, 349, 319, 275, 213, 139, 135, 184, 229, 274, 319, 344, 351, 349, 344, 340, 335, 336, 339, 339, 338, 340, 341, 339, 339, 340, 346, 310, 17, 
    399, 363, 369, 365, 364, 360, 339, 283, 164, 92, 122, 163, 194, 228, 266, 300, 324, 336, 340, 335, 333, 339, 341, 339, 342, 342, 340, 340, 341, 347, 311, 18, 
    403, 362, 367, 366, 363, 362, 358, 334, 204, 82, 87, 108, 125, 159, 186, 207, 231, 258, 283, 295, 311, 336, 345, 343, 342, 340, 338, 340, 339, 344, 310, 18, 
    404, 362, 365, 364, 363, 362, 358, 346, 214, 59, 51, 74, 78, 98, 123, 146, 162, 173, 180, 180, 200, 252, 294, 314, 329, 339, 342, 342, 341, 345, 311, 17, 
    403, 359, 358, 359, 361, 361, 359, 314, 187, 54, 27, 50, 66, 78, 87, 95, 104, 117, 124, 116, 123, 165, 195, 208, 234, 264, 290, 315, 330, 340, 311, 16, 
    398, 356, 353, 356, 357, 359, 352, 286, 180, 115, 81, 46, 52, 60, 93, 149, 165, 139, 85, 81, 108, 127, 133, 139, 201, 264, 283, 299, 315, 331, 307, 13, 
    393, 355, 353, 356, 357, 359, 354, 303, 245, 231, 196, 140, 137, 147, 174, 235, 258, 236, 176, 160, 185, 191, 171, 164, 216, 277, 298, 313, 324, 333, 307, 14, 
    377, 343, 342, 340, 337, 336, 328, 295, 277, 289, 260, 203, 195, 207, 233, 285, 295, 265, 222, 225, 253, 244, 223, 220, 257, 289, 283, 286, 297, 309, 288, 12, 
    290, 255, 253, 248, 240, 236, 233, 229, 226, 230, 216, 183, 180, 190, 214, 248, 254, 241, 223, 225, 240, 243, 237, 237, 250, 259, 259, 259, 257, 263, 246, 3, 
    248, 214, 217, 212, 206, 204, 203, 200, 197, 197, 194, 189, 189, 193, 199, 210, 209, 203, 207, 209, 205, 204, 209, 215, 211, 208, 208, 204, 201, 202, 189, 0, 
    183, 155, 163, 158, 151, 144, 139, 133, 129, 127, 122, 116, 116, 121, 131, 142, 142, 131, 127, 127, 127, 125, 125, 130, 133, 134, 134, 127, 118, 122, 135, 0, 
    143, 104, 117, 116, 113, 109, 105, 106, 105, 99, 93, 90, 92, 94, 95, 99, 102, 93, 86, 84, 83, 82, 85, 86, 86, 87, 87, 77, 76, 111, 141, 0, 
    115, 77, 92, 89, 86, 80, 74, 77, 74, 66, 62, 62, 62, 65, 65, 69, 70, 62, 54, 51, 50, 52, 52, 50, 49, 50, 50, 64, 100, 135, 139, 0, 
    77, 41, 53, 50, 52, 51, 49, 53, 50, 42, 39, 43, 48, 48, 49, 53, 55, 51, 45, 44, 46, 49, 50, 49, 46, 49, 76, 115, 136, 137, 118, 0, 
    80, 43, 57, 55, 55, 53, 53, 56, 53, 51, 62, 70, 69, 65, 66, 74, 74, 69, 65, 64, 55, 51, 51, 47, 57, 92, 134, 144, 132, 107, 77, 0, 
    75, 36, 48, 48, 51, 51, 49, 49, 48, 45, 57, 68, 67, 63, 61, 68, 69, 65, 66, 66, 56, 49, 51, 63, 98, 129, 138, 126, 90, 56, 53, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 8, 5, 5, 9, 10, 9, 9, 7, 0, 0, 0, 1, 25, 56, 56, 21, 0, 0, 0, 0, 
    
    -- channel=59
    17, 19, 10, 16, 26, 24, 26, 25, 24, 25, 25, 26, 26, 30, 29, 28, 27, 26, 28, 29, 27, 27, 27, 28, 26, 19, 10, 9, 10, 8, 23, 107, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 132, 
    0, 0, 0, 0, 0, 0, 7, 16, 4, 0, 0, 2, 4, 10, 7, 0, 1, 1, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 6, 134, 
    0, 0, 0, 0, 0, 0, 21, 6, 0, 18, 22, 23, 24, 21, 21, 14, 20, 20, 16, 21, 21, 17, 23, 0, 0, 0, 0, 0, 0, 0, 6, 134, 
    0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 135, 
    0, 0, 0, 0, 0, 1, 31, 0, 11, 9, 0, 0, 12, 8, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 6, 136, 
    0, 0, 0, 0, 0, 14, 28, 0, 12, 14, 8, 9, 15, 5, 7, 5, 14, 7, 15, 21, 10, 19, 2, 12, 2, 0, 0, 0, 0, 0, 8, 137, 
    0, 0, 0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 6, 136, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 134, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 133, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 132, 
    0, 0, 0, 4, 19, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 132, 
    0, 0, 0, 11, 23, 21, 21, 32, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 137, 
    0, 0, 0, 0, 0, 0, 0, 3, 24, 27, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 135, 
    0, 0, 0, 3, 2, 6, 0, 0, 0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 133, 
    0, 0, 0, 0, 0, 0, 12, 16, 12, 5, 5, 11, 17, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 132, 
    0, 0, 0, 0, 0, 0, 0, 18, 45, 27, 13, 10, 7, 18, 28, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 133, 
    0, 0, 0, 0, 0, 0, 0, 0, 51, 55, 23, 26, 17, 6, 8, 22, 35, 37, 30, 22, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 135, 
    0, 0, 0, 0, 0, 0, 0, 0, 53, 81, 48, 48, 42, 32, 20, 9, 8, 18, 35, 56, 54, 41, 30, 14, 0, 0, 0, 0, 0, 0, 5, 133, 
    0, 0, 0, 0, 0, 0, 0, 5, 65, 78, 45, 42, 39, 37, 36, 34, 27, 17, 14, 18, 18, 15, 30, 45, 45, 39, 28, 12, 0, 0, 6, 134, 
    0, 0, 0, 0, 0, 0, 0, 19, 40, 33, 17, 15, 30, 43, 28, 8, 0, 0, 25, 26, 9, 0, 2, 12, 0, 0, 0, 0, 0, 0, 9, 140, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 138, 
    0, 0, 0, 0, 0, 0, 1, 16, 19, 9, 27, 40, 10, 1, 0, 0, 0, 25, 39, 6, 0, 13, 22, 9, 0, 0, 9, 12, 9, 1, 14, 143, 
    0, 41, 44, 43, 48, 49, 48, 49, 50, 46, 56, 69, 65, 57, 46, 29, 27, 31, 40, 39, 30, 27, 33, 34, 27, 18, 16, 15, 19, 17, 31, 143, 
    0, 3, 8, 4, 5, 3, 1, 2, 1, 0, 3, 2, 0, 0, 0, 3, 13, 14, 11, 12, 14, 16, 15, 15, 20, 21, 21, 22, 23, 23, 35, 128, 
    12, 28, 26, 26, 30, 32, 35, 38, 38, 40, 41, 43, 45, 43, 40, 35, 41, 47, 45, 47, 49, 49, 46, 46, 47, 47, 49, 53, 50, 46, 41, 113, 
    31, 50, 49, 49, 51, 51, 48, 45, 45, 46, 47, 48, 45, 42, 41, 38, 39, 41, 39, 39, 40, 39, 37, 35, 35, 36, 37, 41, 38, 18, 10, 88, 
    23, 32, 31, 30, 33, 38, 37, 33, 36, 37, 36, 36, 37, 37, 37, 36, 36, 41, 43, 41, 39, 40, 41, 43, 41, 40, 39, 33, 11, 0, 20, 97, 
    41, 46, 43, 43, 43, 45, 43, 42, 46, 46, 46, 44, 41, 40, 40, 38, 39, 42, 43, 42, 40, 38, 38, 39, 40, 37, 26, 8, 6, 29, 52, 102, 
    37, 40, 39, 36, 37, 39, 37, 37, 39, 38, 31, 26, 28, 30, 29, 26, 28, 29, 29, 28, 34, 38, 39, 40, 37, 21, 2, 11, 39, 50, 46, 89, 
    39, 44, 44, 42, 42, 42, 42, 41, 42, 41, 37, 42, 43, 44, 42, 40, 45, 44, 44, 42, 46, 43, 41, 33, 12, 5, 24, 50, 54, 49, 44, 84, 
    76, 85, 79, 78, 79, 81, 82, 81, 81, 81, 73, 77, 82, 83, 81, 77, 80, 81, 82, 83, 88, 82, 79, 78, 75, 82, 89, 90, 88, 82, 79, 106, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 2, 10, 9, 7, 6, 6, 8, 8, 8, 8, 3, 0, 0, 2, 3, 1, 0, 0, 0, 0, 4, 7, 7, 5, 0, 0, 0, 0, 4, 12, 3, 
    
    -- channel=61
    158, 371, 424, 436, 423, 396, 367, 364, 372, 383, 396, 398, 400, 389, 388, 384, 382, 384, 382, 388, 394, 395, 397, 394, 395, 408, 427, 448, 464, 474, 451, 242, 
    331, 627, 707, 732, 721, 684, 643, 626, 634, 651, 678, 690, 693, 682, 676, 671, 672, 678, 679, 683, 689, 691, 691, 685, 688, 703, 728, 755, 768, 777, 741, 421, 
    338, 641, 723, 751, 746, 717, 649, 599, 584, 603, 657, 672, 666, 656, 646, 654, 660, 672, 670, 673, 681, 681, 672, 684, 698, 735, 767, 784, 788, 794, 756, 433, 
    341, 643, 715, 746, 759, 748, 670, 589, 530, 541, 583, 586, 589, 582, 577, 586, 598, 605, 606, 610, 618, 619, 601, 633, 676, 749, 783, 784, 784, 793, 757, 434, 
    344, 642, 707, 738, 758, 755, 676, 588, 525, 536, 543, 534, 537, 531, 523, 545, 564, 577, 584, 586, 596, 590, 581, 616, 674, 761, 792, 789, 793, 802, 764, 437, 
    339, 634, 697, 727, 751, 734, 650, 582, 534, 554, 536, 526, 525, 512, 503, 532, 554, 581, 583, 589, 594, 579, 591, 602, 657, 729, 766, 787, 791, 800, 766, 438, 
    338, 632, 693, 721, 739, 702, 612, 527, 515, 555, 552, 565, 552, 536, 520, 548, 572, 593, 600, 595, 593, 582, 616, 602, 630, 665, 725, 783, 788, 796, 761, 436, 
    345, 638, 693, 717, 732, 691, 596, 511, 515, 553, 563, 572, 558, 553, 541, 559, 570, 584, 590, 575, 568, 561, 597, 597, 608, 631, 704, 768, 777, 787, 753, 431, 
    361, 653, 698, 713, 730, 701, 643, 587, 574, 569, 577, 577, 574, 577, 573, 584, 588, 596, 595, 575, 562, 560, 600, 625, 644, 676, 726, 767, 773, 782, 748, 428, 
    383, 675, 713, 716, 733, 727, 714, 678, 646, 617, 616, 619, 616, 624, 632, 641, 645, 649, 647, 630, 625, 623, 649, 688, 720, 748, 760, 774, 774, 781, 745, 426, 
    402, 700, 735, 730, 739, 740, 733, 709, 682, 658, 658, 654, 655, 665, 675, 686, 689, 688, 680, 670, 666, 666, 681, 719, 753, 769, 768, 770, 769, 779, 745, 427, 
    412, 719, 740, 717, 690, 677, 689, 707, 725, 715, 708, 706, 710, 721, 731, 735, 731, 723, 717, 714, 714, 715, 723, 743, 761, 771, 772, 773, 774, 786, 754, 432, 
    418, 728, 738, 692, 620, 554, 551, 599, 671, 721, 750, 761, 763, 770, 778, 784, 784, 779, 773, 769, 765, 767, 770, 772, 772, 774, 774, 775, 777, 786, 751, 430, 
    420, 738, 760, 712, 636, 544, 482, 466, 503, 581, 664, 725, 761, 778, 789, 794, 793, 789, 782, 774, 767, 766, 768, 768, 767, 768, 771, 773, 774, 781, 745, 425, 
    424, 746, 777, 742, 698, 624, 534, 443, 405, 431, 514, 620, 707, 765, 792, 798, 793, 789, 784, 775, 767, 765, 769, 771, 771, 769, 769, 766, 764, 771, 736, 419, 
    428, 756, 810, 806, 797, 752, 680, 560, 423, 351, 358, 447, 562, 663, 738, 780, 792, 787, 778, 767, 760, 758, 761, 763, 765, 766, 766, 764, 762, 771, 737, 420, 
    432, 764, 818, 816, 820, 811, 786, 712, 544, 379, 286, 300, 387, 473, 565, 647, 708, 748, 765, 766, 762, 763, 764, 768, 770, 770, 770, 768, 766, 774, 740, 424, 
    436, 766, 820, 816, 823, 817, 810, 782, 631, 435, 273, 209, 251, 303, 375, 449, 516, 578, 633, 671, 707, 737, 761, 778, 777, 773, 769, 767, 765, 772, 740, 425, 
    437, 765, 817, 813, 821, 818, 812, 796, 655, 441, 243, 152, 171, 191, 235, 286, 336, 382, 421, 450, 487, 550, 626, 693, 731, 754, 766, 771, 768, 774, 742, 425, 
    434, 761, 810, 803, 811, 812, 812, 765, 628, 398, 196, 120, 127, 152, 182, 198, 218, 239, 259, 270, 287, 339, 407, 474, 531, 584, 644, 695, 730, 759, 740, 425, 
    426, 753, 804, 798, 804, 809, 805, 738, 598, 405, 247, 159, 126, 115, 168, 230, 287, 303, 249, 213, 188, 222, 262, 295, 372, 468, 573, 645, 687, 730, 722, 419, 
    418, 746, 803, 797, 801, 807, 804, 747, 645, 543, 457, 371, 303, 263, 302, 377, 462, 503, 442, 380, 341, 361, 354, 336, 371, 463, 574, 643, 685, 722, 712, 413, 
    400, 723, 779, 774, 770, 769, 759, 721, 676, 655, 621, 549, 473, 430, 458, 529, 603, 627, 570, 524, 515, 531, 516, 490, 510, 569, 620, 646, 662, 684, 673, 391, 
    310, 581, 616, 614, 600, 592, 583, 575, 568, 568, 552, 517, 480, 465, 491, 537, 578, 595, 572, 556, 558, 569, 570, 569, 577, 594, 605, 611, 613, 618, 599, 343, 
    247, 473, 499, 496, 484, 477, 467, 460, 453, 447, 442, 438, 432, 435, 445, 467, 480, 486, 487, 487, 488, 486, 492, 500, 506, 506, 501, 496, 493, 489, 476, 260, 
    164, 355, 367, 369, 361, 351, 337, 324, 313, 305, 298, 288, 282, 285, 297, 320, 334, 333, 323, 314, 313, 312, 312, 315, 323, 330, 332, 328, 314, 308, 313, 151, 
    121, 279, 279, 287, 287, 283, 272, 263, 253, 246, 234, 227, 225, 226, 228, 234, 238, 231, 217, 205, 199, 195, 195, 196, 198, 198, 199, 190, 182, 201, 232, 117, 
    78, 206, 195, 201, 198, 192, 182, 172, 164, 157, 144, 139, 136, 137, 137, 141, 143, 138, 127, 113, 105, 103, 104, 106, 106, 105, 106, 117, 146, 191, 242, 135, 
    30, 135, 113, 117, 115, 114, 111, 108, 108, 102, 92, 93, 97, 101, 102, 105, 109, 112, 104, 95, 91, 94, 97, 100, 98, 101, 124, 165, 208, 255, 269, 117, 
    32, 134, 113, 118, 116, 115, 113, 112, 112, 109, 114, 124, 137, 136, 132, 137, 142, 146, 138, 132, 120, 116, 105, 99, 106, 137, 189, 240, 277, 265, 213, 63, 
    26, 123, 98, 104, 105, 110, 110, 109, 105, 101, 111, 127, 145, 143, 137, 140, 144, 148, 146, 145, 133, 123, 108, 115, 146, 191, 245, 278, 249, 184, 136, 22, 
    0, 16, 4, 6, 8, 13, 14, 12, 8, 7, 20, 35, 46, 43, 38, 40, 43, 48, 48, 47, 35, 21, 10, 14, 42, 95, 138, 122, 67, 24, 11, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 83, 77, 73, 76, 90, 91, 87, 91, 95, 97, 99, 109, 107, 110, 108, 104, 110, 111, 114, 113, 108, 111, 111, 110, 109, 98, 95, 97, 101, 103, 21, 
    58, 79, 72, 72, 63, 60, 54, 42, 57, 58, 56, 55, 52, 50, 50, 58, 55, 54, 57, 58, 57, 59, 60, 63, 74, 77, 81, 93, 97, 103, 106, 21, 
    54, 78, 74, 80, 78, 75, 65, 79, 89, 58, 59, 66, 65, 78, 73, 68, 64, 67, 66, 67, 64, 69, 71, 79, 77, 86, 94, 100, 98, 102, 105, 21, 
    50, 76, 74, 80, 79, 80, 70, 67, 71, 80, 100, 103, 91, 89, 91, 94, 102, 105, 110, 110, 108, 109, 109, 120, 100, 92, 100, 103, 100, 102, 101, 16, 
    52, 78, 74, 79, 80, 73, 45, 34, 41, 46, 44, 36, 35, 42, 42, 43, 35, 38, 44, 34, 43, 43, 41, 45, 53, 77, 92, 95, 96, 98, 99, 16, 
    51, 77, 73, 77, 79, 67, 65, 73, 70, 64, 55, 62, 73, 73, 62, 61, 61, 66, 58, 60, 67, 63, 81, 71, 85, 96, 93, 99, 99, 100, 98, 14, 
    48, 74, 71, 75, 75, 77, 84, 66, 78, 77, 73, 81, 70, 74, 74, 76, 80, 88, 93, 87, 97, 91, 95, 82, 103, 104, 93, 97, 97, 101, 98, 15, 
    48, 72, 69, 73, 73, 73, 55, 31, 46, 48, 44, 44, 47, 56, 53, 47, 42, 44, 46, 40, 46, 46, 58, 65, 55, 65, 87, 95, 91, 94, 94, 15, 
    49, 75, 74, 76, 76, 74, 66, 65, 74, 74, 79, 77, 85, 87, 84, 82, 74, 72, 80, 85, 85, 89, 96, 93, 69, 73, 86, 91, 88, 91, 93, 15, 
    59, 78, 80, 81, 76, 77, 78, 77, 81, 78, 80, 84, 76, 75, 75, 74, 80, 85, 86, 81, 85, 82, 85, 89, 85, 87, 87, 91, 91, 94, 94, 15, 
    63, 87, 75, 63, 52, 64, 73, 67, 64, 65, 61, 58, 59, 60, 60, 61, 57, 55, 59, 62, 67, 70, 67, 74, 88, 91, 94, 98, 97, 97, 96, 14, 
    72, 98, 79, 83, 81, 82, 61, 38, 52, 70, 79, 79, 77, 78, 80, 81, 83, 85, 86, 88, 88, 88, 89, 91, 92, 92, 91, 89, 87, 89, 89, 11, 
    75, 102, 92, 106, 110, 110, 121, 108, 76, 57, 60, 75, 85, 88, 88, 87, 86, 86, 83, 82, 82, 83, 81, 81, 83, 86, 88, 90, 91, 94, 96, 17, 
    77, 102, 80, 54, 41, 50, 78, 107, 111, 100, 81, 69, 76, 84, 86, 87, 88, 89, 91, 92, 94, 95, 96, 97, 97, 96, 95, 94, 93, 93, 91, 13, 
    79, 106, 98, 97, 94, 81, 54, 41, 55, 67, 75, 73, 62, 67, 83, 95, 97, 97, 94, 91, 91, 91, 89, 87, 87, 86, 86, 88, 87, 88, 88, 12, 
    77, 107, 101, 101, 100, 105, 99, 67, 41, 53, 61, 78, 99, 89, 69, 66, 76, 88, 94, 93, 89, 89, 90, 90, 88, 88, 88, 88, 85, 87, 86, 7, 
    78, 109, 105, 106, 103, 107, 110, 105, 53, 35, 51, 50, 74, 102, 113, 97, 73, 58, 56, 61, 73, 85, 86, 89, 90, 90, 89, 91, 89, 88, 84, 6, 
    79, 113, 113, 115, 112, 113, 112, 108, 59, 29, 34, 28, 41, 49, 68, 98, 116, 113, 91, 60, 45, 39, 45, 64, 79, 90, 95, 97, 92, 90, 87, 8, 
    82, 112, 110, 110, 109, 109, 107, 88, 61, 59, 54, 44, 46, 42, 40, 41, 55, 81, 104, 114, 112, 105, 85, 66, 59, 56, 59, 70, 79, 83, 82, 6, 
    81, 111, 107, 109, 108, 107, 105, 91, 102, 83, 60, 53, 32, 27, 45, 68, 83, 75, 45, 44, 65, 89, 101, 119, 149, 154, 142, 117, 93, 85, 81, 4, 
    86, 112, 103, 103, 106, 108, 107, 109, 109, 71, 29, 43, 84, 87, 99, 79, 46, 48, 64, 87, 53, 47, 76, 97, 104, 77, 76, 98, 102, 99, 91, 12, 
    76, 101, 91, 89, 91, 93, 89, 68, 33, 23, 15, 0, 2, 0, 2, 21, 28, 25, 11, 14, 17, 9, 0, 0, 10, 29, 37, 34, 42, 60, 68, 2, 
    43, 63, 49, 49, 55, 58, 60, 59, 57, 61, 54, 31, 5, 1, 10, 34, 58, 63, 42, 18, 28, 40, 32, 18, 22, 45, 59, 59, 54, 53, 55, 0, 
    102, 136, 117, 120, 122, 125, 126, 125, 128, 129, 126, 128, 126, 121, 109, 90, 74, 69, 70, 72, 69, 64, 65, 64, 58, 48, 40, 35, 36, 42, 52, 5, 
    30, 47, 33, 24, 20, 17, 12, 14, 14, 13, 13, 8, 0, 0, 0, 11, 11, 10, 13, 10, 10, 13, 17, 16, 16, 16, 14, 14, 19, 26, 54, 15, 
    23, 46, 26, 21, 22, 24, 31, 40, 43, 48, 50, 48, 49, 51, 50, 53, 58, 62, 64, 65, 66, 65, 65, 67, 68, 67, 68, 67, 67, 83, 101, 33, 
    55, 86, 70, 70, 71, 65, 65, 70, 70, 72, 69, 66, 58, 54, 56, 57, 60, 56, 53, 55, 54, 52, 49, 46, 47, 49, 50, 59, 79, 82, 62, 14, 
    24, 48, 35, 35, 36, 36, 39, 40, 42, 45, 41, 39, 39, 43, 47, 51, 50, 50, 50, 48, 48, 50, 50, 49, 46, 44, 56, 74, 63, 38, 63, 42, 
    31, 55, 42, 46, 46, 44, 46, 48, 49, 51, 54, 54, 47, 47, 53, 58, 59, 62, 60, 58, 49, 47, 48, 50, 52, 68, 77, 56, 44, 79, 109, 43, 
    25, 47, 36, 36, 35, 34, 34, 37, 41, 41, 37, 26, 29, 33, 37, 39, 36, 36, 32, 34, 36, 46, 49, 60, 81, 77, 48, 50, 89, 91, 72, 22, 
    0, 14, 9, 11, 6, 1, 0, 3, 4, 6, 11, 12, 11, 10, 12, 18, 19, 16, 13, 11, 7, 9, 8, 8, 0, 0, 28, 56, 37, 15, 13, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 5, 21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 10, 24, 0, 0, 0, 0, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 6, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 13, 11, 9, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 16, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 4, 2, 1, 4, 2, 5, 2, 1, 6, 8, 9, 10, 10, 11, 12, 10, 5, 0, 0, 0, 0, 
    54, 7, 16, 13, 12, 11, 11, 13, 15, 15, 16, 16, 15, 16, 15, 16, 13, 12, 11, 11, 13, 14, 13, 14, 15, 13, 3, 0, 0, 0, 0, 0, 
    54, 7, 13, 11, 11, 10, 10, 12, 13, 10, 12, 11, 8, 8, 11, 11, 9, 8, 6, 9, 9, 11, 12, 12, 7, 0, 0, 0, 0, 0, 0, 0, 
    55, 9, 18, 13, 16, 17, 15, 17, 18, 19, 19, 12, 11, 10, 11, 13, 12, 9, 9, 9, 10, 14, 15, 9, 1, 0, 0, 0, 0, 0, 0, 12, 
    59, 24, 30, 28, 29, 28, 28, 29, 29, 29, 31, 32, 23, 22, 23, 26, 27, 22, 24, 23, 23, 23, 28, 25, 12, 0, 0, 0, 0, 10, 29, 31, 
    
    -- channel=64
    118, 118, 111, 111, 106, 108, 99, 98, 104, 122, 102, 103, 116, 108, 103, 94, 93, 95, 94, 89, 102, 106, 95, 72, 108, 131, 70, 102, 117, 100, 101, 144, 
    61, 102, 122, 105, 81, 78, 67, 75, 95, 140, 104, 63, 77, 90, 86, 58, 56, 57, 67, 63, 81, 109, 80, 9, 62, 165, 73, 73, 113, 89, 71, 167, 
    49, 84, 132, 85, 63, 79, 76, 74, 108, 140, 91, 53, 63, 98, 99, 52, 72, 89, 79, 60, 70, 116, 75, 0, 58, 191, 99, 76, 86, 67, 78, 165, 
    58, 70, 129, 63, 63, 80, 75, 72, 121, 133, 84, 64, 71, 106, 115, 48, 55, 99, 83, 46, 57, 123, 73, 0, 51, 191, 94, 41, 50, 76, 113, 177, 
    60, 55, 108, 60, 71, 81, 68, 67, 137, 129, 95, 86, 93, 95, 97, 46, 36, 77, 81, 53, 57, 131, 68, 0, 36, 150, 72, 27, 46, 99, 109, 188, 
    50, 53, 75, 90, 83, 79, 74, 63, 145, 130, 108, 93, 87, 67, 64, 53, 51, 72, 97, 79, 49, 122, 66, 0, 17, 112, 72, 50, 42, 80, 60, 187, 
    53, 99, 65, 94, 78, 69, 95, 74, 137, 120, 90, 68, 56, 58, 72, 80, 71, 60, 127, 116, 27, 81, 73, 0, 0, 100, 69, 56, 24, 72, 75, 185, 
    66, 130, 68, 74, 68, 61, 100, 107, 137, 90, 50, 48, 54, 77, 111, 130, 100, 33, 102, 135, 22, 55, 73, 0, 0, 89, 59, 47, 19, 114, 127, 168, 
    86, 107, 34, 43, 82, 86, 69, 111, 149, 60, 27, 55, 69, 107, 147, 129, 73, 49, 70, 95, 40, 45, 55, 5, 0, 68, 53, 42, 31, 148, 139, 155, 
    93, 85, 0, 17, 63, 128, 81, 69, 109, 48, 31, 59, 94, 147, 141, 65, 25, 76, 83, 44, 32, 49, 55, 14, 38, 57, 42, 40, 52, 170, 129, 148, 
    94, 86, 0, 8, 32, 109, 136, 77, 45, 40, 40, 55, 114, 153, 103, 31, 30, 69, 64, 41, 33, 80, 98, 9, 33, 53, 32, 42, 73, 188, 119, 137, 
    101, 92, 0, 3, 20, 60, 141, 126, 34, 35, 57, 59, 97, 80, 43, 41, 55, 58, 52, 61, 56, 97, 109, 0, 23, 59, 18, 41, 86, 187, 130, 139, 
    114, 108, 6, 9, 13, 27, 95, 107, 42, 50, 76, 63, 89, 53, 13, 40, 63, 68, 74, 70, 79, 78, 70, 0, 39, 84, 27, 31, 93, 183, 134, 154, 
    109, 103, 22, 24, 20, 1, 48, 54, 60, 63, 75, 68, 92, 86, 52, 47, 63, 64, 64, 57, 71, 61, 69, 26, 33, 79, 54, 19, 87, 159, 91, 167, 
    85, 85, 38, 35, 50, 0, 23, 49, 85, 83, 58, 55, 76, 68, 72, 78, 75, 65, 52, 52, 59, 36, 63, 56, 53, 52, 44, 30, 83, 120, 58, 193, 
    78, 85, 39, 41, 67, 14, 7, 46, 48, 106, 97, 24, 59, 62, 54, 57, 63, 80, 79, 65, 76, 28, 11, 38, 83, 68, 18, 45, 102, 125, 60, 208, 
    73, 88, 46, 27, 45, 23, 12, 38, 0, 54, 181, 60, 17, 52, 49, 40, 47, 57, 63, 51, 70, 60, 16, 0, 42, 91, 45, 36, 144, 143, 16, 194, 
    60, 64, 59, 19, 38, 22, 41, 45, 35, 0, 112, 113, 12, 16, 47, 56, 60, 40, 34, 49, 51, 64, 74, 9, 14, 60, 78, 36, 129, 144, 1, 193, 
    52, 31, 50, 29, 75, 36, 52, 45, 62, 16, 0, 88, 85, 20, 46, 40, 43, 59, 46, 47, 51, 33, 59, 51, 57, 62, 71, 71, 77, 124, 47, 196, 
    42, 17, 45, 50, 102, 67, 39, 49, 30, 82, 0, 0, 108, 50, 28, 36, 24, 32, 40, 51, 61, 45, 47, 59, 60, 119, 88, 82, 63, 53, 27, 210, 
    33, 38, 72, 80, 88, 86, 28, 62, 31, 63, 99, 0, 17, 61, 16, 31, 48, 23, 12, 61, 66, 38, 41, 66, 59, 112, 81, 74, 73, 15, 0, 224, 
    40, 91, 65, 67, 85, 87, 28, 65, 93, 7, 94, 78, 0, 8, 30, 26, 31, 48, 23, 43, 60, 53, 45, 74, 70, 81, 77, 56, 34, 24, 23, 224, 
    58, 123, 59, 50, 89, 91, 36, 29, 88, 45, 15, 85, 23, 0, 14, 45, 16, 43, 60, 50, 48, 62, 48, 63, 68, 81, 88, 31, 3, 40, 58, 220, 
    69, 79, 35, 47, 74, 101, 66, 7, 27, 84, 51, 21, 28, 19, 3, 44, 35, 31, 60, 62, 40, 56, 42, 55, 69, 85, 70, 25, 32, 49, 60, 216, 
    32, 0, 0, 32, 84, 101, 85, 34, 34, 60, 74, 30, 0, 36, 19, 34, 38, 28, 58, 59, 16, 59, 48, 55, 78, 93, 56, 21, 67, 43, 48, 214, 
    1, 0, 0, 9, 59, 85, 82, 59, 79, 66, 11, 22, 18, 21, 34, 43, 35, 21, 55, 64, 7, 31, 78, 74, 65, 96, 91, 16, 60, 39, 53, 214, 
    31, 59, 0, 0, 12, 52, 77, 75, 77, 86, 27, 2, 39, 42, 65, 93, 57, 8, 33, 44, 37, 35, 70, 71, 60, 93, 127, 29, 38, 57, 85, 214, 
    45, 114, 62, 0, 0, 30, 40, 70, 73, 75, 78, 55, 40, 54, 83, 116, 80, 0, 4, 34, 43, 54, 57, 51, 84, 123, 107, 34, 37, 98, 105, 190, 
    46, 129, 128, 67, 0, 3, 12, 21, 66, 82, 75, 72, 60, 61, 53, 67, 73, 17, 4, 49, 29, 40, 76, 71, 110, 141, 60, 49, 40, 62, 97, 194, 
    50, 122, 124, 143, 28, 0, 0, 3, 21, 59, 74, 62, 58, 69, 49, 59, 65, 44, 29, 44, 21, 30, 76, 104, 143, 112, 52, 95, 23, 0, 87, 236, 
    54, 120, 87, 150, 107, 20, 0, 0, 6, 9, 41, 58, 53, 66, 57, 82, 102, 66, 28, 52, 43, 68, 87, 75, 103, 80, 64, 67, 7, 0, 93, 237, 
    69, 137, 56, 92, 129, 101, 28, 0, 5, 0, 0, 4, 27, 41, 13, 14, 81, 108, 52, 80, 76, 54, 25, 0, 23, 41, 33, 2, 6, 4, 69, 230, 
    
    -- channel=65
    0, 34, 27, 2, 0, 14, 38, 37, 32, 6, 0, 0, 19, 42, 35, 37, 54, 83, 89, 88, 82, 69, 53, 70, 94, 86, 57, 17, 23, 26, 33, 7, 
    10, 89, 77, 52, 46, 61, 80, 78, 68, 38, 9, 7, 53, 72, 63, 66, 84, 114, 120, 116, 122, 118, 102, 113, 146, 146, 106, 33, 66, 90, 81, 36, 
    19, 114, 89, 83, 71, 90, 97, 88, 73, 40, 6, 7, 47, 58, 50, 63, 87, 121, 122, 119, 125, 116, 102, 116, 157, 161, 123, 61, 100, 112, 87, 29, 
    25, 133, 115, 123, 91, 104, 102, 93, 71, 40, 0, 0, 20, 38, 47, 73, 97, 117, 113, 111, 118, 107, 107, 121, 175, 191, 165, 105, 122, 130, 118, 50, 
    24, 130, 112, 111, 98, 103, 95, 89, 58, 35, 0, 0, 27, 59, 82, 94, 101, 120, 117, 100, 97, 87, 115, 141, 188, 218, 201, 137, 155, 164, 164, 82, 
    15, 103, 91, 85, 89, 104, 92, 81, 44, 29, 0, 26, 75, 108, 111, 105, 90, 89, 91, 90, 76, 84, 132, 157, 203, 243, 229, 175, 188, 182, 165, 55, 
    4, 74, 77, 75, 109, 106, 86, 73, 33, 24, 20, 79, 133, 143, 122, 80, 40, 62, 78, 79, 83, 91, 146, 173, 221, 245, 247, 198, 204, 171, 131, 27, 
    0, 79, 89, 101, 144, 134, 103, 69, 41, 49, 62, 127, 167, 155, 108, 47, 38, 74, 101, 98, 99, 127, 180, 206, 230, 248, 245, 206, 204, 152, 104, 0, 
    5, 92, 107, 126, 183, 157, 128, 82, 55, 81, 112, 169, 183, 135, 70, 43, 70, 110, 124, 142, 150, 166, 202, 215, 219, 241, 246, 211, 201, 136, 77, 0, 
    11, 103, 106, 140, 210, 198, 144, 92, 72, 89, 133, 180, 167, 124, 92, 85, 117, 148, 169, 175, 191, 196, 192, 192, 199, 237, 240, 211, 197, 123, 65, 0, 
    13, 108, 95, 135, 216, 223, 182, 118, 92, 117, 160, 176, 151, 139, 132, 153, 182, 201, 208, 197, 201, 189, 171, 197, 216, 244, 231, 209, 199, 125, 54, 0, 
    3, 87, 78, 117, 198, 220, 215, 179, 157, 163, 187, 181, 148, 142, 143, 154, 190, 205, 200, 196, 184, 176, 175, 201, 210, 237, 225, 200, 192, 131, 56, 0, 
    4, 102, 89, 113, 180, 212, 224, 234, 204, 183, 186, 176, 144, 143, 152, 173, 181, 175, 179, 181, 174, 176, 177, 197, 210, 227, 217, 209, 204, 145, 85, 0, 
    17, 122, 97, 120, 163, 194, 213, 243, 218, 186, 165, 154, 159, 172, 165, 171, 174, 171, 170, 160, 158, 174, 175, 200, 208, 215, 204, 212, 200, 156, 109, 9, 
    21, 125, 108, 122, 154, 180, 203, 234, 236, 204, 181, 156, 137, 168, 182, 183, 189, 188, 173, 167, 160, 174, 179, 211, 217, 209, 212, 201, 191, 139, 80, 2, 
    21, 129, 120, 138, 169, 194, 207, 225, 242, 213, 171, 164, 138, 171, 198, 209, 205, 193, 197, 208, 201, 201, 202, 213, 220, 225, 213, 195, 169, 118, 83, 29, 
    24, 139, 136, 162, 176, 193, 183, 205, 211, 223, 197, 188, 173, 183, 199, 207, 211, 219, 215, 204, 201, 196, 186, 213, 225, 220, 186, 189, 155, 118, 99, 17, 
    31, 157, 163, 183, 176, 176, 161, 182, 187, 197, 215, 211, 197, 187, 186, 209, 212, 220, 226, 230, 227, 228, 210, 204, 195, 196, 174, 129, 128, 118, 113, 47, 
    42, 177, 177, 185, 141, 146, 138, 158, 183, 177, 196, 202, 200, 212, 205, 225, 237, 229, 231, 234, 222, 206, 208, 213, 194, 165, 136, 116, 119, 125, 141, 93, 
    52, 183, 162, 151, 134, 136, 123, 134, 164, 155, 148, 177, 184, 201, 226, 237, 237, 246, 247, 235, 230, 219, 210, 211, 198, 157, 136, 120, 119, 140, 186, 113, 
    52, 170, 143, 133, 145, 135, 125, 129, 145, 163, 148, 155, 183, 208, 236, 259, 255, 243, 246, 228, 218, 208, 200, 193, 190, 161, 147, 122, 138, 169, 199, 131, 
    41, 148, 134, 134, 142, 139, 130, 129, 157, 168, 177, 166, 176, 214, 254, 259, 268, 253, 236, 225, 215, 197, 205, 205, 196, 172, 153, 152, 173, 191, 199, 129, 
    33, 163, 171, 192, 221, 181, 149, 148, 169, 178, 165, 180, 180, 211, 256, 260, 259, 245, 237, 218, 210, 210, 213, 201, 200, 177, 166, 169, 182, 202, 213, 135, 
    52, 216, 247, 265, 272, 243, 200, 181, 181, 185, 164, 173, 216, 215, 246, 251, 252, 241, 236, 226, 219, 209, 230, 209, 193, 179, 169, 158, 163, 211, 213, 136, 
    61, 211, 228, 270, 308, 297, 269, 225, 195, 187, 184, 182, 219, 243, 236, 226, 216, 210, 216, 225, 231, 227, 224, 199, 187, 175, 153, 136, 153, 207, 198, 125, 
    44, 171, 192, 235, 287, 316, 300, 278, 240, 206, 193, 193, 196, 207, 203, 170, 153, 159, 192, 226, 230, 226, 217, 204, 194, 162, 111, 112, 137, 192, 173, 93, 
    31, 133, 138, 152, 205, 267, 306, 298, 290, 261, 216, 195, 207, 202, 184, 158, 142, 158, 181, 225, 232, 221, 230, 208, 168, 131, 96, 91, 132, 176, 150, 94, 
    29, 118, 89, 67, 118, 189, 274, 313, 311, 294, 269, 230, 216, 216, 204, 189, 176, 179, 192, 207, 221, 227, 214, 201, 151, 97, 80, 94, 133, 162, 194, 134, 
    33, 119, 92, 38, 67, 124, 205, 282, 320, 321, 310, 289, 262, 242, 232, 208, 187, 171, 172, 194, 211, 217, 210, 173, 121, 100, 88, 81, 128, 187, 214, 135, 
    32, 118, 97, 38, 53, 67, 143, 214, 283, 319, 324, 317, 306, 281, 264, 241, 224, 195, 157, 146, 166, 146, 143, 151, 149, 154, 136, 132, 195, 226, 234, 163, 
    12, 88, 73, 59, 76, 49, 75, 149, 217, 281, 306, 314, 315, 310, 306, 293, 273, 228, 184, 138, 128, 125, 159, 200, 215, 219, 192, 204, 226, 244, 256, 170, 
    0, 0, 7, 0, 6, 0, 0, 27, 79, 102, 116, 123, 120, 107, 103, 100, 88, 56, 25, 14, 24, 24, 31, 45, 50, 57, 55, 59, 65, 79, 77, 24, 
    
    -- channel=66
    53, 0, 0, 0, 28, 20, 3, 1, 0, 0, 2, 46, 22, 0, 0, 14, 21, 0, 0, 0, 0, 0, 0, 42, 8, 0, 0, 22, 0, 13, 16, 0, 
    78, 0, 0, 0, 31, 10, 0, 0, 0, 0, 0, 60, 21, 0, 0, 21, 27, 0, 0, 4, 0, 0, 0, 64, 9, 0, 0, 38, 3, 4, 0, 0, 
    77, 0, 0, 0, 27, 0, 0, 0, 0, 0, 15, 55, 20, 0, 0, 36, 29, 0, 0, 8, 0, 0, 0, 75, 10, 0, 0, 40, 9, 0, 0, 0, 
    68, 0, 0, 0, 8, 0, 0, 0, 0, 0, 19, 42, 21, 0, 0, 36, 20, 0, 0, 6, 0, 0, 0, 80, 15, 0, 0, 25, 5, 0, 0, 0, 
    63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 38, 24, 8, 0, 16, 10, 0, 0, 0, 5, 0, 0, 71, 25, 0, 0, 4, 0, 0, 0, 0, 
    66, 0, 0, 1, 0, 0, 0, 0, 0, 0, 30, 43, 16, 1, 0, 0, 0, 10, 0, 0, 34, 1, 0, 68, 35, 0, 0, 0, 0, 0, 0, 0, 
    64, 0, 3, 20, 0, 0, 0, 0, 0, 0, 57, 35, 0, 0, 0, 0, 6, 42, 0, 0, 50, 20, 0, 53, 31, 0, 0, 0, 0, 0, 0, 0, 
    57, 0, 25, 35, 0, 0, 0, 0, 0, 16, 68, 16, 0, 0, 0, 0, 38, 44, 0, 0, 49, 13, 0, 24, 19, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 45, 38, 0, 0, 0, 0, 0, 42, 55, 0, 0, 0, 0, 17, 55, 9, 0, 0, 17, 0, 0, 6, 15, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 58, 44, 0, 0, 0, 0, 0, 53, 23, 0, 0, 0, 0, 45, 38, 0, 0, 0, 0, 0, 0, 17, 16, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 64, 51, 0, 0, 0, 0, 28, 38, 0, 0, 0, 0, 10, 30, 0, 0, 0, 0, 0, 0, 0, 36, 6, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 66, 52, 0, 0, 0, 0, 11, 3, 0, 0, 0, 0, 24, 11, 0, 0, 0, 0, 0, 0, 0, 40, 4, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 53, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 23, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 36, 27, 0, 6, 0, 0, 0, 0, 0, 2, 0, 1, 12, 0, 0, 0, 0, 0, 0, 9, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 0, 20, 18, 0, 13, 0, 0, 0, 0, 0, 5, 27, 9, 0, 2, 0, 0, 0, 3, 0, 11, 18, 6, 0, 0, 0, 0, 0, 0, 5, 0, 
    52, 0, 12, 13, 0, 0, 0, 0, 0, 0, 0, 0, 42, 20, 5, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 41, 0, 
    61, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 20, 14, 8, 0, 0, 0, 0, 0, 0, 0, 9, 14, 0, 0, 0, 0, 0, 0, 47, 0, 
    72, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 43, 0, 
    81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 1, 0, 0, 33, 0, 
    84, 0, 0, 0, 0, 0, 12, 1, 0, 0, 6, 10, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 11, 0, 
    79, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 5, 25, 18, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 0, 0, 
    68, 0, 0, 12, 0, 0, 7, 3, 0, 0, 0, 0, 36, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 0, 0, 0, 
    61, 0, 23, 3, 0, 0, 0, 12, 0, 0, 0, 0, 22, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 3, 0, 0, 0, 
    78, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 
    86, 4, 20, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 5, 0, 0, 9, 0, 0, 0, 0, 0, 0, 31, 2, 0, 0, 0, 
    91, 0, 12, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 8, 0, 0, 0, 0, 0, 0, 0, 0, 50, 21, 0, 0, 0, 
    82, 0, 0, 52, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 33, 0, 0, 0, 0, 0, 0, 0, 0, 71, 12, 0, 0, 0, 
    77, 0, 0, 47, 72, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 26, 0, 0, 0, 0, 0, 0, 0, 14, 45, 0, 0, 0, 0, 
    75, 0, 0, 7, 68, 73, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 9, 0, 0, 0, 0, 0, 29, 10, 18, 26, 0, 0, 
    66, 0, 0, 0, 26, 76, 64, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 0, 0, 0, 11, 0, 26, 33, 0, 0, 
    49, 0, 13, 0, 0, 31, 71, 64, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 8, 12, 0, 0, 0, 0, 12, 8, 0, 0, 
    35, 0, 41, 17, 0, 12, 61, 78, 43, 24, 20, 4, 0, 0, 1, 2, 0, 0, 16, 9, 10, 29, 36, 43, 6, 0, 0, 16, 10, 5, 0, 0, 
    
    -- channel=67
    38, 0, 5, 33, 40, 32, 26, 22, 18, 28, 50, 61, 40, 20, 18, 20, 11, 3, 0, 0, 0, 0, 2, 4, 0, 0, 3, 36, 17, 10, 8, 12, 
    94, 80, 74, 82, 82, 83, 92, 107, 103, 102, 101, 101, 107, 97, 98, 115, 126, 138, 157, 157, 140, 118, 118, 119, 117, 99, 117, 142, 125, 100, 91, 88, 
    93, 95, 80, 80, 91, 102, 104, 106, 100, 100, 100, 113, 131, 126, 119, 134, 135, 126, 134, 144, 136, 117, 111, 121, 126, 101, 85, 92, 79, 70, 88, 94, 
    98, 92, 83, 87, 107, 111, 107, 103, 96, 100, 106, 126, 138, 133, 111, 110, 124, 109, 92, 106, 126, 118, 110, 113, 123, 85, 47, 62, 73, 82, 91, 67, 
    113, 98, 100, 89, 124, 114, 106, 111, 101, 101, 109, 119, 120, 106, 94, 93, 119, 137, 126, 132, 154, 128, 103, 116, 112, 78, 58, 84, 114, 103, 74, 48, 
    128, 135, 158, 145, 124, 107, 100, 115, 114, 102, 96, 85, 82, 83, 90, 113, 142, 138, 113, 138, 160, 134, 103, 112, 113, 93, 83, 103, 112, 93, 99, 93, 
    127, 140, 156, 148, 118, 96, 87, 98, 115, 107, 85, 79, 99, 112, 131, 158, 165, 151, 111, 84, 116, 123, 112, 113, 133, 101, 87, 95, 92, 98, 132, 141, 
    113, 123, 109, 92, 73, 90, 104, 82, 86, 95, 94, 115, 139, 156, 173, 160, 134, 114, 125, 78, 62, 106, 118, 133, 148, 138, 99, 98, 98, 104, 119, 111, 
    99, 100, 101, 77, 61, 54, 95, 104, 64, 54, 92, 129, 148, 167, 156, 115, 74, 78, 96, 97, 81, 93, 131, 156, 151, 144, 120, 107, 107, 110, 105, 87, 
    99, 98, 114, 115, 95, 70, 60, 113, 121, 80, 96, 119, 120, 116, 102, 82, 92, 110, 102, 103, 120, 131, 174, 189, 165, 127, 116, 106, 107, 105, 102, 87, 
    100, 103, 121, 130, 121, 94, 53, 74, 128, 143, 141, 135, 105, 58, 18, 34, 90, 128, 134, 132, 143, 161, 161, 159, 163, 133, 119, 105, 101, 93, 84, 87, 
    110, 101, 128, 140, 141, 115, 76, 38, 60, 117, 128, 117, 94, 68, 61, 47, 66, 99, 120, 132, 129, 140, 116, 106, 129, 132, 133, 122, 101, 90, 76, 69, 
    109, 95, 117, 139, 148, 148, 102, 55, 43, 78, 86, 85, 77, 79, 115, 141, 133, 119, 106, 88, 80, 77, 87, 110, 146, 138, 122, 133, 123, 91, 54, 37, 
    90, 75, 81, 107, 126, 150, 131, 101, 97, 99, 102, 88, 81, 68, 62, 89, 111, 112, 106, 86, 71, 59, 57, 72, 120, 140, 109, 116, 120, 88, 62, 43, 
    108, 97, 104, 104, 114, 127, 144, 117, 101, 73, 101, 133, 106, 83, 75, 51, 40, 54, 74, 97, 98, 99, 77, 44, 61, 92, 124, 114, 121, 123, 120, 86, 
    123, 115, 122, 122, 108, 102, 125, 121, 96, 51, 17, 99, 133, 100, 86, 82, 71, 51, 38, 45, 54, 65, 102, 93, 42, 38, 90, 122, 118, 135, 135, 92, 
    113, 100, 92, 111, 103, 109, 111, 138, 126, 128, 44, 0, 70, 82, 62, 71, 88, 96, 81, 50, 45, 39, 56, 102, 101, 74, 57, 113, 113, 86, 103, 81, 
    104, 92, 81, 90, 119, 142, 150, 147, 140, 136, 116, 0, 4, 78, 82, 74, 59, 65, 89, 103, 101, 104, 78, 67, 103, 117, 134, 114, 127, 81, 80, 92, 
    99, 89, 94, 114, 120, 136, 158, 137, 133, 111, 140, 119, 29, 59, 87, 69, 77, 62, 43, 49, 68, 84, 96, 85, 80, 97, 139, 150, 157, 129, 60, 45, 
    100, 94, 128, 144, 142, 132, 135, 133, 135, 130, 106, 180, 130, 36, 43, 46, 55, 80, 75, 58, 68, 84, 86, 84, 83, 84, 71, 97, 112, 115, 106, 60, 
    108, 117, 150, 130, 122, 116, 114, 133, 132, 163, 116, 107, 175, 110, 43, 62, 57, 51, 86, 89, 65, 70, 85, 82, 85, 83, 65, 68, 62, 67, 114, 113, 
    124, 122, 130, 124, 97, 99, 113, 113, 99, 102, 138, 70, 81, 118, 85, 61, 67, 63, 63, 96, 100, 81, 88, 93, 80, 84, 89, 90, 82, 91, 122, 118, 
    130, 107, 75, 76, 99, 100, 112, 129, 102, 79, 108, 131, 62, 74, 102, 82, 70, 75, 69, 72, 83, 78, 72, 69, 77, 86, 92, 81, 106, 145, 159, 119, 
    104, 63, 28, 17, 42, 82, 94, 120, 136, 130, 105, 112, 122, 83, 88, 98, 84, 79, 76, 70, 68, 51, 63, 84, 97, 110, 114, 111, 120, 159, 155, 104, 
    103, 86, 93, 93, 86, 79, 89, 97, 123, 140, 125, 74, 80, 113, 88, 101, 105, 92, 73, 62, 62, 63, 51, 84, 106, 107, 127, 160, 161, 155, 153, 122, 
    146, 171, 222, 221, 170, 126, 100, 111, 125, 116, 124, 133, 101, 104, 120, 132, 156, 142, 105, 66, 56, 85, 78, 70, 83, 94, 108, 158, 171, 160, 177, 138, 
    139, 155, 211, 257, 243, 188, 151, 115, 119, 126, 121, 157, 185, 164, 152, 143, 146, 157, 123, 81, 75, 70, 92, 78, 70, 100, 134, 125, 155, 173, 164, 134, 
    112, 119, 147, 215, 274, 247, 194, 149, 108, 114, 134, 136, 150, 167, 147, 101, 64, 76, 108, 93, 85, 79, 67, 92, 116, 129, 126, 123, 159, 131, 101, 90, 
    109, 106, 114, 132, 206, 261, 219, 179, 144, 108, 110, 134, 139, 146, 148, 126, 96, 78, 92, 102, 88, 90, 92, 97, 117, 126, 111, 137, 147, 128, 74, 42, 
    123, 121, 119, 85, 114, 202, 255, 219, 189, 148, 105, 99, 121, 137, 147, 149, 147, 156, 142, 116, 123, 131, 137, 121, 87, 64, 78, 95, 105, 142, 139, 104, 
    146, 161, 151, 124, 89, 138, 225, 270, 234, 213, 184, 130, 100, 111, 119, 100, 75, 89, 143, 165, 169, 174, 150, 106, 57, 28, 29, 40, 57, 109, 148, 97, 
    181, 162, 163, 172, 137, 125, 166, 237, 284, 280, 284, 273, 244, 221, 209, 202, 178, 140, 138, 171, 174, 167, 152, 151, 162, 154, 158, 166, 190, 210, 210, 148, 
    
    -- channel=68
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 2, 19, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 4, 0, 0, 65, 23, 0, 0, 0, 0, 24, 
    0, 16, 24, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 3, 0, 0, 82, 40, 0, 0, 0, 11, 26, 
    0, 27, 25, 2, 0, 0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 9, 0, 0, 0, 92, 58, 0, 0, 19, 35, 28, 
    0, 22, 19, 1, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 5, 95, 76, 0, 6, 38, 46, 46, 
    0, 10, 1, 0, 0, 0, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 10, 108, 101, 24, 22, 43, 56, 51, 
    0, 1, 0, 0, 0, 2, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 12, 110, 117, 46, 41, 63, 79, 38, 
    0, 2, 0, 0, 7, 26, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 7, 99, 116, 60, 61, 90, 93, 2, 
    0, 3, 0, 0, 44, 61, 36, 5, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 77, 105, 69, 76, 104, 79, 0, 
    0, 12, 0, 0, 61, 97, 65, 6, 0, 0, 0, 14, 27, 36, 0, 0, 0, 0, 0, 0, 0, 7, 13, 0, 0, 65, 89, 74, 88, 103, 56, 0, 
    0, 26, 0, 0, 56, 97, 102, 40, 0, 0, 0, 34, 48, 59, 11, 0, 0, 12, 8, 0, 2, 16, 19, 0, 0, 69, 78, 78, 97, 99, 38, 0, 
    0, 28, 0, 0, 41, 71, 107, 82, 0, 0, 19, 36, 53, 56, 16, 19, 45, 38, 24, 30, 31, 38, 24, 0, 0, 65, 66, 64, 87, 97, 37, 0, 
    0, 36, 0, 0, 28, 49, 85, 100, 46, 23, 40, 43, 51, 53, 28, 47, 64, 56, 53, 56, 64, 63, 39, 16, 15, 64, 58, 47, 78, 99, 37, 0, 
    0, 37, 0, 0, 24, 31, 53, 98, 92, 70, 55, 49, 55, 59, 42, 55, 66, 65, 66, 62, 73, 78, 67, 67, 52, 68, 49, 37, 71, 95, 28, 0, 
    0, 32, 0, 0, 29, 25, 35, 95, 117, 100, 81, 54, 34, 53, 64, 72, 78, 81, 72, 66, 70, 76, 76, 101, 104, 86, 52, 39, 75, 81, 0, 0, 
    0, 28, 0, 0, 35, 39, 38, 85, 106, 110, 115, 71, 21, 56, 78, 87, 95, 93, 90, 88, 90, 86, 77, 101, 127, 128, 75, 46, 80, 72, 0, 0, 
    0, 24, 0, 2, 30, 49, 38, 69, 74, 95, 148, 116, 45, 66, 89, 99, 105, 103, 100, 94, 97, 94, 78, 92, 118, 145, 91, 61, 78, 62, 0, 0, 
    0, 25, 19, 26, 38, 49, 32, 49, 55, 62, 116, 142, 102, 79, 89, 115, 111, 108, 110, 115, 116, 110, 100, 91, 100, 121, 96, 46, 43, 40, 0, 10, 
    0, 34, 41, 49, 38, 33, 13, 20, 40, 53, 65, 110, 141, 111, 99, 122, 125, 127, 121, 122, 126, 99, 92, 104, 106, 99, 72, 32, 10, 12, 0, 51, 
    0, 49, 55, 42, 27, 25, 0, 0, 24, 42, 38, 58, 108, 113, 113, 131, 135, 137, 134, 140, 146, 115, 96, 107, 106, 97, 67, 25, 7, 0, 2, 87, 
    0, 67, 50, 14, 18, 23, 0, 0, 20, 21, 41, 39, 49, 94, 124, 150, 159, 142, 138, 144, 142, 111, 97, 104, 102, 86, 65, 29, 18, 2, 19, 102, 
    0, 75, 25, 0, 13, 23, 0, 0, 35, 10, 33, 57, 29, 61, 130, 152, 161, 160, 147, 135, 131, 109, 103, 107, 100, 76, 60, 34, 18, 31, 40, 90, 
    0, 71, 19, 8, 51, 33, 0, 0, 28, 42, 23, 51, 48, 62, 120, 149, 152, 153, 159, 136, 113, 109, 110, 99, 93, 69, 52, 22, 17, 43, 39, 82, 
    0, 65, 46, 70, 88, 56, 18, 0, 14, 60, 45, 27, 63, 88, 118, 134, 149, 144, 153, 146, 114, 109, 129, 108, 90, 66, 36, 9, 17, 35, 20, 81, 
    0, 43, 43, 91, 121, 91, 50, 9, 15, 42, 44, 35, 65, 109, 119, 121, 128, 120, 133, 142, 118, 126, 145, 116, 88, 68, 37, 0, 0, 16, 11, 79, 
    0, 31, 27, 45, 86, 105, 79, 44, 31, 27, 15, 31, 64, 84, 102, 100, 83, 68, 98, 135, 124, 128, 145, 124, 91, 79, 45, 0, 0, 7, 12, 54, 
    0, 25, 0, 0, 2, 57, 84, 72, 55, 38, 11, 6, 42, 55, 69, 79, 55, 33, 59, 121, 137, 126, 136, 122, 88, 78, 41, 0, 0, 10, 0, 35, 
    0, 30, 0, 0, 0, 0, 41, 82, 84, 59, 34, 5, 2, 16, 34, 53, 50, 26, 48, 107, 127, 125, 123, 113, 86, 64, 0, 0, 0, 0, 12, 57, 
    0, 31, 15, 0, 0, 0, 0, 41, 93, 99, 71, 36, 9, 4, 8, 17, 42, 34, 43, 96, 112, 113, 127, 99, 64, 43, 0, 0, 0, 0, 27, 90, 
    0, 26, 0, 0, 0, 0, 0, 0, 47, 96, 102, 78, 53, 36, 22, 18, 41, 44, 35, 57, 82, 75, 81, 71, 57, 39, 0, 0, 0, 0, 48, 126, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 41, 80, 93, 91, 82, 60, 56, 75, 61, 26, 26, 42, 35, 47, 52, 66, 72, 37, 33, 15, 12, 69, 128, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 20, 0, 0, 18, 18, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 6, 56, 
    
    -- channel=69
    36, 46, 34, 24, 35, 39, 41, 54, 49, 24, 20, 33, 46, 47, 41, 54, 75, 81, 91, 95, 91, 75, 61, 82, 95, 68, 57, 53, 57, 61, 51, 15, 
    97, 94, 71, 60, 82, 95, 107, 111, 95, 44, 41, 77, 102, 105, 91, 112, 145, 154, 150, 166, 161, 123, 107, 163, 184, 114, 93, 102, 98, 97, 93, 28, 
    115, 109, 88, 88, 114, 113, 119, 116, 89, 41, 48, 84, 110, 102, 88, 117, 141, 142, 128, 138, 148, 117, 110, 169, 192, 115, 87, 89, 100, 114, 98, 28, 
    120, 134, 100, 109, 130, 123, 121, 118, 85, 40, 48, 73, 100, 87, 82, 112, 130, 134, 133, 142, 152, 122, 115, 176, 200, 128, 104, 114, 144, 144, 111, 30, 
    116, 145, 115, 148, 131, 127, 118, 115, 80, 42, 44, 65, 83, 83, 84, 122, 146, 138, 130, 131, 145, 134, 127, 175, 214, 160, 147, 163, 171, 154, 121, 33, 
    116, 140, 116, 138, 135, 121, 106, 104, 64, 41, 48, 80, 99, 120, 129, 128, 131, 146, 131, 96, 127, 126, 138, 195, 230, 189, 174, 175, 181, 160, 137, 56, 
    106, 111, 116, 115, 116, 117, 102, 93, 45, 47, 81, 121, 153, 172, 146, 117, 120, 128, 107, 85, 110, 130, 161, 219, 238, 213, 189, 181, 196, 166, 124, 33, 
    100, 78, 114, 128, 136, 116, 93, 92, 46, 59, 116, 165, 196, 178, 123, 90, 95, 121, 84, 89, 139, 149, 185, 233, 257, 211, 206, 193, 203, 139, 73, 7, 
    96, 85, 131, 169, 167, 142, 97, 78, 67, 101, 148, 184, 187, 143, 94, 76, 103, 140, 143, 122, 160, 183, 201, 240, 274, 218, 205, 199, 193, 103, 45, 0, 
    98, 102, 155, 199, 197, 150, 125, 82, 82, 152, 177, 187, 173, 112, 70, 94, 148, 171, 178, 182, 201, 206, 197, 238, 258, 223, 206, 200, 182, 87, 31, 0, 
    100, 98, 158, 201, 220, 178, 130, 99, 117, 162, 181, 177, 140, 99, 109, 142, 177, 186, 186, 203, 216, 202, 190, 222, 226, 220, 212, 201, 173, 72, 27, 0, 
    90, 99, 146, 190, 220, 215, 157, 126, 140, 160, 178, 164, 121, 110, 145, 192, 199, 199, 202, 191, 192, 164, 155, 213, 245, 230, 210, 204, 180, 72, 34, 0, 
    89, 85, 128, 170, 204, 218, 198, 162, 173, 181, 180, 162, 138, 145, 161, 165, 173, 184, 186, 171, 152, 149, 155, 208, 233, 220, 216, 204, 173, 84, 51, 0, 
    94, 94, 138, 159, 186, 209, 223, 210, 188, 171, 162, 169, 143, 137, 158, 159, 151, 144, 143, 156, 145, 153, 162, 189, 196, 188, 210, 215, 179, 100, 80, 26, 
    109, 122, 144, 165, 173, 206, 214, 221, 188, 164, 121, 129, 160, 160, 156, 163, 155, 143, 146, 147, 143, 150, 166, 181, 179, 177, 183, 222, 173, 103, 120, 50, 
    115, 132, 148, 166, 167, 197, 207, 208, 190, 169, 146, 118, 137, 166, 169, 161, 162, 172, 167, 153, 147, 155, 154, 179, 190, 174, 177, 197, 163, 95, 113, 32, 
    114, 133, 156, 168, 174, 191, 220, 208, 227, 180, 140, 145, 123, 148, 176, 182, 177, 163, 164, 182, 171, 185, 199, 185, 173, 169, 199, 174, 141, 84, 100, 43, 
    123, 146, 165, 189, 179, 184, 196, 196, 207, 206, 141, 164, 160, 161, 175, 173, 182, 186, 185, 183, 178, 166, 174, 197, 188, 160, 141, 181, 137, 112, 147, 42, 
    137, 171, 170, 185, 179, 172, 158, 190, 178, 201, 179, 169, 193, 170, 164, 177, 168, 181, 195, 177, 170, 188, 181, 180, 164, 152, 125, 133, 122, 122, 175, 49, 
    150, 181, 171, 182, 149, 142, 149, 170, 174, 179, 214, 156, 167, 199, 173, 189, 197, 185, 193, 196, 172, 172, 180, 174, 158, 125, 118, 100, 128, 149, 179, 80, 
    158, 169, 153, 163, 131, 130, 151, 152, 181, 149, 170, 186, 147, 190, 216, 190, 194, 204, 192, 184, 178, 173, 177, 176, 162, 121, 120, 122, 147, 180, 210, 88, 
    152, 148, 139, 149, 157, 138, 150, 156, 162, 178, 128, 174, 191, 186, 214, 220, 197, 192, 204, 174, 165, 179, 175, 159, 158, 142, 136, 143, 171, 199, 227, 90, 
    138, 132, 163, 169, 156, 152, 154, 164, 161, 189, 179, 150, 209, 217, 211, 216, 214, 192, 182, 177, 171, 158, 168, 169, 164, 159, 147, 171, 200, 217, 219, 84, 
    143, 157, 186, 212, 219, 190, 182, 186, 183, 166, 193, 182, 178, 217, 222, 208, 206, 199, 178, 164, 175, 180, 169, 165, 168, 164, 155, 187, 217, 215, 218, 91, 
    153, 214, 267, 280, 266, 240, 214, 220, 209, 172, 156, 203, 211, 188, 211, 194, 193, 199, 189, 176, 185, 172, 180, 163, 159, 152, 148, 176, 204, 218, 211, 90, 
    169, 222, 250, 277, 284, 273, 266, 244, 217, 205, 185, 184, 230, 219, 193, 177, 173, 190, 189, 181, 199, 182, 179, 161, 145, 127, 128, 163, 193, 211, 200, 92, 
    143, 163, 180, 227, 275, 292, 278, 277, 244, 215, 232, 221, 204, 216, 185, 150, 135, 153, 182, 182, 192, 200, 155, 153, 160, 118, 93, 164, 175, 194, 186, 62, 
    129, 113, 125, 160, 216, 278, 286, 271, 275, 255, 231, 232, 222, 211, 184, 145, 137, 164, 173, 190, 184, 187, 184, 159, 129, 103, 99, 139, 168, 204, 168, 48, 
    137, 112, 88, 100, 142, 209, 291, 296, 280, 276, 259, 238, 239, 234, 222, 193, 174, 200, 199, 177, 188, 181, 166, 163, 127, 76, 100, 132, 186, 200, 193, 99, 
    137, 113, 93, 86, 107, 159, 232, 303, 300, 283, 284, 278, 257, 247, 253, 237, 197, 167, 179, 176, 169, 182, 173, 156, 121, 98, 121, 127, 181, 233, 220, 83, 
    125, 106, 124, 100, 93, 115, 173, 246, 309, 301, 290, 296, 289, 263, 255, 239, 216, 183, 152, 148, 160, 155, 143, 147, 141, 151, 161, 158, 214, 266, 230, 82, 
    68, 74, 78, 78, 84, 75, 106, 151, 195, 241, 246, 242, 244, 246, 252, 239, 208, 188, 175, 123, 107, 98, 127, 173, 185, 190, 184, 200, 208, 231, 199, 99, 
    
    -- channel=70
    32, 56, 55, 40, 28, 40, 39, 41, 51, 66, 31, 20, 42, 50, 45, 28, 35, 46, 50, 44, 54, 63, 43, 13, 58, 93, 27, 38, 54, 37, 40, 85, 
    13, 46, 58, 29, 23, 39, 28, 29, 46, 56, 23, 11, 28, 46, 36, 9, 26, 34, 28, 20, 33, 56, 28, 0, 34, 96, 27, 18, 34, 31, 38, 74, 
    20, 32, 59, 23, 27, 39, 30, 30, 52, 51, 21, 15, 22, 43, 35, 4, 27, 46, 29, 16, 30, 58, 25, 0, 31, 101, 34, 19, 31, 39, 46, 66, 
    27, 24, 59, 19, 35, 36, 31, 30, 57, 46, 25, 19, 22, 29, 35, 11, 16, 41, 39, 24, 28, 57, 22, 0, 25, 92, 42, 18, 27, 47, 47, 86, 
    17, 22, 44, 31, 34, 32, 31, 23, 61, 44, 29, 20, 26, 25, 33, 27, 21, 30, 41, 30, 11, 53, 26, 0, 17, 80, 42, 19, 21, 47, 46, 104, 
    9, 32, 14, 34, 32, 32, 38, 19, 57, 41, 25, 22, 33, 33, 39, 39, 22, 20, 54, 34, 0, 44, 35, 0, 12, 71, 38, 30, 18, 49, 41, 84, 
    12, 48, 4, 27, 34, 31, 43, 31, 51, 26, 14, 28, 34, 41, 56, 43, 13, 0, 58, 49, 0, 34, 33, 0, 2, 67, 37, 34, 16, 60, 41, 60, 
    23, 45, 9, 28, 46, 34, 31, 49, 56, 9, 10, 32, 35, 57, 62, 34, 16, 15, 35, 50, 15, 23, 31, 8, 0, 51, 35, 28, 18, 73, 48, 55, 
    35, 38, 0, 21, 46, 63, 27, 36, 55, 13, 17, 35, 48, 67, 49, 21, 24, 43, 29, 25, 25, 26, 40, 14, 15, 36, 29, 25, 28, 79, 44, 54, 
    40, 38, 0, 7, 29, 70, 56, 21, 19, 18, 26, 38, 62, 66, 36, 15, 21, 38, 37, 26, 25, 46, 44, 0, 28, 36, 24, 27, 36, 85, 39, 50, 
    47, 33, 0, 1, 18, 45, 81, 42, 0, 17, 30, 34, 56, 49, 39, 31, 28, 31, 37, 40, 28, 49, 42, 0, 28, 37, 20, 30, 41, 93, 42, 42, 
    48, 31, 0, 0, 7, 25, 66, 62, 23, 33, 37, 32, 43, 23, 17, 34, 42, 40, 39, 37, 35, 37, 42, 3, 27, 48, 16, 18, 49, 93, 43, 52, 
    43, 40, 0, 3, 4, 8, 38, 53, 49, 39, 41, 29, 40, 32, 8, 16, 27, 30, 36, 30, 38, 32, 40, 4, 17, 52, 20, 7, 52, 82, 40, 79, 
    41, 43, 11, 12, 18, 0, 22, 34, 46, 30, 29, 27, 37, 40, 36, 27, 25, 27, 23, 24, 31, 25, 38, 23, 24, 31, 29, 14, 50, 71, 30, 89, 
    34, 34, 14, 16, 28, 0, 10, 26, 35, 53, 31, 6, 30, 32, 33, 37, 43, 40, 26, 23, 28, 6, 18, 37, 44, 30, 15, 23, 52, 58, 7, 90, 
    25, 35, 11, 12, 27, 17, 6, 25, 9, 60, 84, 0, 11, 32, 25, 27, 31, 37, 43, 34, 44, 23, 2, 8, 41, 60, 11, 22, 65, 46, 0, 103, 
    19, 33, 25, 10, 28, 17, 17, 20, 4, 6, 89, 44, 5, 19, 30, 30, 23, 23, 29, 33, 37, 41, 27, 0, 16, 43, 44, 15, 63, 58, 0, 103, 
    18, 19, 35, 21, 33, 4, 22, 12, 25, 0, 19, 78, 29, 2, 25, 22, 32, 31, 18, 26, 27, 20, 38, 23, 16, 17, 37, 17, 40, 64, 2, 99, 
    17, 13, 35, 22, 38, 18, 12, 16, 22, 29, 0, 29, 58, 10, 19, 20, 21, 28, 30, 33, 34, 18, 26, 33, 29, 44, 15, 26, 20, 28, 23, 118, 
    15, 22, 31, 16, 39, 35, 1, 29, 7, 36, 16, 0, 30, 37, 14, 29, 24, 13, 22, 37, 31, 23, 26, 34, 28, 56, 32, 37, 21, 6, 15, 122, 
    21, 36, 13, 28, 43, 37, 7, 31, 24, 0, 59, 2, 0, 24, 22, 20, 26, 27, 10, 29, 34, 24, 22, 36, 29, 44, 42, 26, 23, 25, 9, 115, 
    23, 45, 6, 27, 46, 42, 13, 17, 49, 11, 24, 53, 0, 0, 24, 26, 16, 33, 24, 20, 22, 26, 21, 34, 36, 39, 39, 11, 14, 27, 21, 117, 
    19, 36, 23, 34, 44, 53, 22, 3, 34, 52, 9, 20, 23, 6, 6, 32, 18, 19, 35, 28, 19, 31, 25, 33, 36, 37, 41, 17, 10, 20, 32, 117, 
    15, 22, 23, 46, 56, 61, 47, 14, 19, 40, 34, 2, 7, 26, 6, 27, 22, 15, 32, 30, 13, 38, 24, 29, 32, 41, 34, 11, 21, 22, 36, 118, 
    6, 6, 0, 23, 56, 69, 59, 37, 36, 24, 19, 26, 8, 19, 20, 22, 17, 11, 30, 32, 4, 33, 37, 27, 31, 54, 35, 0, 26, 25, 35, 109, 
    0, 4, 0, 0, 28, 55, 64, 49, 47, 46, 11, 12, 22, 16, 30, 26, 8, 0, 18, 30, 20, 13, 40, 36, 31, 50, 49, 0, 22, 34, 33, 101, 
    4, 39, 0, 0, 0, 23, 45, 60, 54, 54, 40, 12, 11, 20, 33, 43, 19, 0, 10, 25, 23, 20, 31, 32, 42, 47, 35, 2, 28, 34, 35, 102, 
    12, 60, 35, 0, 0, 2, 17, 45, 62, 55, 49, 40, 29, 30, 34, 56, 51, 5, 7, 25, 13, 30, 41, 30, 43, 48, 15, 30, 15, 29, 65, 103, 
    14, 59, 54, 38, 0, 0, 3, 13, 40, 62, 56, 47, 45, 45, 33, 43, 44, 27, 11, 20, 15, 20, 38, 35, 47, 43, 22, 36, 0, 16, 72, 125, 
    17, 60, 36, 68, 25, 0, 0, 0, 13, 39, 58, 56, 48, 50, 40, 47, 44, 21, 4, 21, 12, 14, 24, 29, 60, 52, 33, 31, 7, 1, 55, 126, 
    28, 48, 10, 59, 59, 20, 0, 0, 6, 10, 24, 44, 52, 51, 39, 52, 77, 55, 11, 29, 12, 13, 18, 21, 54, 49, 38, 30, 28, 13, 59, 127, 
    21, 38, 8, 28, 49, 38, 8, 0, 0, 0, 0, 0, 9, 20, 9, 3, 30, 51, 29, 24, 18, 9, 5, 0, 12, 17, 16, 6, 6, 6, 27, 93, 
    
    -- channel=71
    110, 38, 3, 20, 50, 62, 44, 44, 40, 18, 12, 76, 77, 35, 28, 41, 57, 42, 21, 21, 29, 8, 6, 56, 77, 0, 0, 60, 34, 22, 48, 17, 
    145, 44, 0, 6, 59, 62, 31, 47, 36, 0, 11, 88, 80, 31, 15, 42, 76, 34, 15, 33, 44, 6, 0, 75, 98, 0, 0, 75, 52, 30, 40, 0, 
    157, 33, 3, 3, 66, 42, 21, 48, 26, 0, 21, 86, 67, 35, 14, 50, 89, 26, 5, 39, 52, 9, 0, 86, 103, 0, 0, 77, 59, 29, 13, 0, 
    171, 24, 19, 0, 60, 23, 28, 46, 16, 0, 30, 76, 59, 48, 35, 50, 76, 28, 7, 35, 48, 11, 0, 94, 102, 0, 0, 62, 57, 24, 1, 0, 
    169, 15, 30, 0, 43, 21, 36, 39, 17, 0, 39, 71, 68, 56, 48, 47, 56, 37, 20, 19, 41, 41, 2, 89, 105, 0, 0, 41, 50, 29, 0, 0, 
    160, 19, 20, 35, 39, 32, 32, 22, 25, 0, 55, 78, 69, 48, 39, 18, 27, 56, 37, 0, 42, 86, 8, 74, 116, 0, 0, 26, 39, 24, 0, 0, 
    149, 23, 15, 79, 38, 34, 26, 6, 18, 2, 84, 85, 49, 28, 5, 0, 26, 81, 64, 0, 40, 106, 12, 58, 114, 5, 0, 21, 25, 15, 0, 0, 
    143, 17, 29, 106, 33, 4, 15, 18, 4, 15, 105, 76, 23, 6, 0, 0, 60, 87, 52, 4, 48, 84, 12, 47, 81, 18, 0, 20, 19, 0, 0, 0, 
    147, 5, 52, 112, 33, 0, 0, 29, 17, 27, 99, 45, 0, 0, 0, 27, 91, 69, 18, 27, 52, 42, 5, 28, 62, 21, 0, 21, 14, 0, 0, 20, 
    156, 0, 63, 122, 38, 0, 0, 0, 36, 61, 72, 21, 0, 0, 0, 61, 88, 39, 7, 34, 46, 17, 0, 19, 83, 8, 0, 26, 9, 0, 0, 40, 
    157, 0, 63, 128, 49, 11, 0, 0, 41, 91, 50, 21, 5, 0, 12, 58, 42, 10, 12, 23, 18, 13, 0, 32, 92, 0, 0, 35, 1, 0, 0, 43, 
    153, 0, 64, 124, 57, 35, 0, 0, 19, 67, 20, 15, 3, 0, 36, 50, 5, 0, 6, 5, 0, 0, 0, 38, 79, 0, 0, 46, 7, 0, 0, 40, 
    160, 0, 58, 110, 54, 54, 28, 0, 1, 13, 0, 0, 3, 0, 28, 34, 6, 1, 2, 0, 2, 0, 1, 15, 46, 0, 0, 47, 19, 0, 0, 35, 
    164, 0, 48, 85, 44, 49, 60, 8, 0, 0, 0, 0, 2, 0, 10, 7, 3, 1, 2, 8, 7, 2, 18, 0, 9, 0, 1, 34, 18, 0, 0, 31, 
    171, 0, 45, 70, 41, 35, 74, 23, 4, 0, 0, 0, 32, 5, 3, 2, 0, 0, 0, 7, 4, 7, 40, 14, 0, 0, 6, 32, 0, 0, 1, 44, 
    172, 0, 43, 70, 47, 33, 56, 24, 8, 24, 0, 0, 63, 33, 2, 0, 0, 0, 0, 0, 0, 0, 19, 34, 15, 0, 0, 28, 0, 0, 29, 62, 
    168, 18, 38, 54, 46, 26, 40, 28, 17, 43, 0, 0, 29, 36, 10, 1, 0, 0, 0, 0, 0, 0, 0, 15, 25, 0, 0, 4, 0, 0, 27, 68, 
    172, 30, 47, 27, 29, 7, 49, 27, 34, 29, 46, 0, 0, 9, 22, 0, 3, 0, 0, 5, 0, 0, 0, 0, 18, 0, 0, 0, 21, 0, 29, 48, 
    184, 32, 40, 1, 18, 0, 54, 41, 44, 18, 30, 66, 0, 0, 33, 3, 2, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 15, 27, 32, 52, 13, 
    197, 20, 24, 3, 27, 1, 44, 59, 25, 41, 9, 49, 51, 0, 15, 12, 0, 0, 7, 0, 0, 0, 10, 0, 0, 0, 0, 28, 28, 50, 72, 0, 
    203, 0, 8, 37, 29, 0, 37, 74, 10, 38, 47, 3, 70, 64, 15, 2, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 25, 41, 59, 47, 0, 
    201, 0, 1, 72, 24, 0, 29, 70, 31, 13, 53, 13, 37, 80, 33, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 17, 60, 49, 13, 0, 
    193, 0, 42, 65, 0, 0, 3, 56, 59, 12, 8, 40, 42, 52, 27, 1, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 17, 57, 31, 15, 0, 
    200, 25, 55, 31, 0, 0, 0, 32, 54, 17, 7, 39, 57, 38, 6, 8, 0, 0, 0, 0, 3, 20, 0, 0, 0, 0, 0, 25, 49, 20, 31, 0, 
    198, 34, 61, 35, 0, 0, 0, 0, 22, 0, 27, 56, 42, 26, 0, 0, 0, 12, 18, 0, 0, 23, 0, 0, 0, 0, 0, 22, 70, 25, 26, 0, 
    194, 30, 48, 68, 36, 0, 0, 0, 0, 0, 15, 53, 35, 15, 0, 0, 0, 44, 52, 2, 0, 9, 0, 0, 0, 0, 0, 15, 99, 22, 18, 0, 
    180, 20, 4, 73, 93, 34, 0, 0, 0, 0, 0, 28, 32, 23, 10, 0, 0, 58, 83, 13, 0, 0, 0, 0, 0, 0, 0, 43, 97, 16, 14, 0, 
    171, 12, 0, 41, 103, 100, 38, 11, 0, 0, 0, 0, 14, 19, 15, 8, 1, 31, 72, 20, 0, 8, 0, 0, 0, 0, 0, 71, 69, 48, 24, 0, 
    174, 6, 0, 18, 56, 120, 88, 46, 5, 0, 0, 0, 0, 0, 0, 12, 0, 15, 44, 21, 4, 12, 0, 0, 0, 0, 22, 74, 38, 92, 31, 0, 
    171, 0, 0, 33, 12, 77, 102, 81, 43, 6, 0, 0, 0, 0, 0, 11, 0, 0, 24, 28, 1, 12, 0, 2, 7, 0, 32, 47, 29, 92, 14, 0, 
    153, 0, 7, 71, 0, 26, 73, 102, 78, 32, 12, 0, 0, 0, 0, 7, 0, 0, 0, 30, 11, 43, 42, 42, 29, 0, 8, 19, 35, 41, 3, 0, 
    113, 0, 27, 71, 8, 18, 46, 72, 66, 33, 29, 27, 7, 0, 0, 10, 0, 0, 0, 28, 14, 42, 48, 48, 40, 2, 14, 26, 36, 20, 12, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    
    -- channel=73
    6, 8, 14, 7, 7, 19, 34, 49, 47, 29, 18, 6, 10, 15, 14, 18, 15, 15, 12, 15, 20, 18, 26, 21, 17, 0, 0, 0, 0, 9, 16, 11, 
    17, 31, 27, 15, 11, 30, 53, 70, 66, 47, 19, 2, 17, 21, 23, 22, 11, 15, 14, 17, 32, 31, 35, 19, 21, 7, 0, 0, 12, 20, 31, 36, 
    26, 52, 33, 16, 15, 41, 60, 72, 63, 39, 7, 0, 19, 22, 17, 11, 12, 18, 19, 22, 35, 34, 31, 16, 18, 11, 0, 11, 29, 34, 42, 33, 
    31, 60, 35, 21, 27, 51, 63, 74, 59, 31, 0, 0, 14, 23, 16, 11, 24, 32, 30, 28, 35, 32, 26, 16, 25, 25, 10, 29, 47, 50, 52, 23, 
    33, 46, 34, 18, 38, 55, 64, 72, 50, 24, 0, 0, 12, 25, 26, 24, 40, 50, 42, 30, 29, 23, 24, 23, 33, 39, 29, 45, 61, 60, 54, 23, 
    32, 30, 32, 9, 38, 53, 61, 63, 39, 18, 0, 1, 15, 26, 33, 34, 42, 52, 41, 29, 21, 18, 25, 30, 42, 51, 50, 57, 70, 59, 45, 32, 
    31, 30, 27, 12, 34, 47, 50, 42, 28, 13, 0, 5, 19, 22, 23, 21, 21, 35, 40, 27, 18, 17, 28, 26, 49, 61, 59, 64, 75, 59, 44, 26, 
    31, 42, 31, 34, 46, 46, 42, 21, 16, 6, 0, 14, 21, 14, 12, 4, 1, 13, 43, 21, 11, 15, 23, 19, 48, 64, 61, 69, 77, 66, 44, 9, 
    32, 49, 42, 61, 72, 52, 41, 16, 5, 0, 4, 24, 18, 12, 7, 0, 0, 14, 34, 18, 9, 12, 11, 15, 34, 58, 64, 76, 80, 70, 38, 0, 
    37, 48, 49, 73, 95, 76, 42, 20, 7, 0, 15, 27, 18, 15, 4, 0, 10, 31, 23, 13, 17, 11, 9, 7, 21, 47, 69, 85, 89, 68, 26, 0, 
    36, 42, 44, 71, 97, 101, 62, 30, 16, 13, 23, 16, 8, 6, 5, 18, 31, 32, 17, 15, 15, 12, 14, 3, 21, 43, 73, 96, 93, 55, 10, 0, 
    27, 28, 34, 62, 92, 104, 90, 54, 23, 24, 14, 0, 0, 0, 0, 19, 25, 15, 1, 0, 0, 0, 3, 0, 17, 39, 74, 96, 80, 44, 4, 0, 
    27, 25, 32, 56, 80, 98, 101, 68, 21, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 34, 66, 88, 71, 47, 13, 0, 
    30, 33, 34, 55, 62, 86, 90, 68, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 48, 75, 75, 54, 20, 9, 
    33, 41, 39, 55, 59, 69, 83, 68, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 36, 65, 74, 45, 17, 12, 
    36, 40, 43, 59, 70, 67, 84, 70, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 54, 65, 40, 12, 9, 
    35, 43, 45, 66, 71, 78, 77, 75, 33, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 41, 61, 34, 8, 17, 
    34, 54, 52, 66, 63, 76, 64, 73, 35, 21, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 51, 30, 20, 33, 
    39, 64, 61, 62, 51, 52, 55, 54, 51, 21, 29, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 37, 44, 38, 44, 
    51, 69, 65, 55, 44, 41, 49, 40, 51, 41, 14, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 41, 54, 64, 64, 
    55, 67, 62, 35, 39, 46, 43, 47, 41, 57, 29, 16, 15, 0, 2, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 46, 60, 62, 89, 75, 
    51, 56, 39, 19, 30, 37, 42, 64, 50, 50, 63, 26, 15, 13, 4, 7, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 5, 49, 70, 84, 92, 70, 
    46, 50, 23, 18, 23, 18, 36, 64, 72, 55, 62, 46, 13, 5, 0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 28, 69, 97, 87, 68, 
    45, 51, 36, 23, 14, 9, 18, 48, 70, 72, 53, 47, 24, 0, 0, 0, 0, 4, 9, 0, 0, 0, 0, 0, 0, 0, 0, 15, 62, 92, 86, 70, 
    41, 43, 41, 30, 14, 4, 7, 23, 43, 56, 58, 52, 37, 9, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 12, 53, 81, 79, 68, 
    38, 34, 32, 23, 16, 4, 0, 5, 19, 23, 41, 58, 37, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 49, 69, 64, 53, 
    35, 21, 9, 2, 8, 6, 1, 0, 7, 11, 13, 34, 30, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 64, 44, 29, 
    30, 21, 0, 0, 0, 0, 4, 6, 3, 3, 1, 7, 7, 3, 6, 13, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 55, 54, 23, 26, 
    29, 27, 0, 0, 0, 0, 0, 6, 10, 4, 2, 8, 3, 3, 12, 17, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 36, 21, 12, 19, 
    26, 24, 4, 0, 0, 0, 0, 0, 6, 14, 15, 18, 16, 12, 14, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 36, 10, 13, 17, 13, 
    12, 14, 0, 0, 0, 0, 0, 0, 0, 10, 20, 26, 28, 26, 19, 11, 0, 0, 0, 0, 0, 0, 0, 15, 32, 39, 42, 49, 23, 32, 32, 26, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 25, 24, 27, 22, 20, 24, 24, 
    
    -- channel=74
    61, 38, 3, 0, 24, 40, 41, 47, 31, 0, 0, 27, 51, 38, 26, 50, 78, 85, 77, 83, 80, 46, 39, 101, 123, 28, 6, 37, 27, 35, 46, 0, 
    123, 85, 28, 28, 73, 82, 78, 86, 55, 0, 0, 62, 90, 62, 43, 85, 122, 108, 95, 118, 125, 72, 64, 168, 197, 39, 9, 76, 74, 80, 76, 0, 
    136, 104, 45, 62, 103, 89, 85, 94, 45, 0, 2, 62, 78, 49, 31, 91, 132, 104, 89, 117, 130, 71, 66, 184, 210, 49, 22, 99, 113, 101, 61, 0, 
    151, 131, 76, 88, 111, 88, 91, 99, 34, 0, 0, 38, 49, 46, 46, 94, 126, 101, 91, 115, 128, 68, 76, 198, 230, 91, 59, 132, 149, 118, 82, 0, 
    145, 117, 96, 94, 102, 86, 89, 93, 23, 0, 0, 35, 60, 72, 79, 109, 128, 111, 88, 80, 108, 84, 90, 207, 253, 137, 105, 155, 172, 144, 105, 0, 
    135, 86, 76, 87, 99, 95, 80, 74, 12, 0, 21, 73, 99, 114, 108, 80, 84, 116, 80, 39, 99, 110, 106, 220, 280, 178, 138, 165, 189, 145, 94, 0, 
    116, 52, 72, 101, 100, 103, 74, 51, 0, 0, 75, 124, 137, 129, 76, 27, 44, 110, 85, 24, 107, 136, 128, 222, 292, 199, 158, 177, 200, 133, 47, 0, 
    102, 42, 97, 158, 131, 98, 78, 55, 3, 37, 129, 158, 150, 102, 24, 3, 69, 121, 89, 60, 138, 164, 156, 230, 279, 206, 173, 191, 201, 91, 0, 0, 
    104, 51, 133, 198, 174, 105, 67, 60, 38, 96, 172, 166, 126, 51, 0, 37, 118, 140, 113, 119, 171, 178, 161, 214, 259, 210, 188, 199, 183, 46, 0, 0, 
    110, 59, 156, 227, 206, 134, 69, 48, 65, 134, 173, 161, 122, 41, 26, 104, 161, 147, 141, 174, 197, 166, 125, 189, 245, 206, 197, 200, 169, 21, 0, 0, 
    112, 49, 154, 230, 228, 181, 91, 56, 109, 162, 162, 155, 111, 78, 120, 179, 186, 164, 168, 177, 177, 151, 119, 202, 248, 200, 201, 204, 160, 6, 0, 0, 
    99, 33, 136, 207, 225, 216, 149, 105, 151, 179, 158, 153, 113, 94, 151, 188, 176, 169, 166, 160, 152, 133, 121, 213, 248, 185, 185, 207, 158, 5, 0, 0, 
    109, 42, 130, 188, 202, 230, 200, 162, 169, 167, 145, 146, 128, 131, 165, 166, 150, 151, 155, 157, 149, 141, 147, 202, 222, 178, 185, 216, 161, 28, 9, 0, 
    120, 66, 131, 173, 174, 220, 228, 203, 166, 135, 137, 148, 138, 142, 160, 162, 151, 140, 142, 151, 146, 160, 174, 192, 190, 169, 179, 214, 162, 45, 49, 0, 
    135, 79, 129, 164, 160, 202, 236, 218, 204, 160, 105, 121, 150, 154, 162, 171, 166, 155, 150, 155, 142, 165, 199, 206, 191, 163, 185, 204, 131, 29, 75, 0, 
    141, 93, 135, 174, 175, 200, 230, 205, 211, 203, 103, 106, 164, 180, 181, 175, 173, 177, 178, 186, 179, 174, 194, 223, 213, 170, 180, 189, 101, 24, 99, 1, 
    146, 119, 147, 182, 175, 190, 201, 201, 208, 224, 148, 124, 174, 190, 194, 198, 189, 178, 180, 179, 173, 181, 197, 219, 206, 179, 159, 170, 99, 14, 100, 6, 
    162, 151, 172, 186, 161, 163, 171, 180, 190, 207, 206, 169, 167, 189, 190, 194, 204, 206, 210, 210, 191, 182, 182, 203, 205, 147, 114, 125, 106, 60, 140, 9, 
    185, 181, 167, 160, 132, 125, 152, 169, 187, 173, 205, 219, 178, 192, 214, 209, 210, 212, 217, 201, 181, 191, 194, 184, 173, 127, 98, 95, 99, 113, 174, 16, 
    205, 170, 148, 140, 113, 98, 140, 150, 158, 164, 159, 190, 196, 203, 226, 234, 223, 220, 236, 215, 180, 191, 201, 177, 159, 115, 91, 100, 120, 155, 205, 18, 
    208, 130, 126, 138, 119, 95, 136, 156, 132, 158, 154, 159, 207, 239, 248, 240, 232, 223, 224, 205, 179, 180, 191, 172, 157, 115, 96, 122, 155, 196, 219, 10, 
    191, 96, 112, 153, 129, 92, 131, 161, 150, 159, 161, 153, 214, 257, 262, 249, 237, 229, 213, 189, 185, 189, 191, 176, 157, 135, 119, 147, 191, 204, 195, 5, 
    177, 123, 190, 209, 159, 116, 125, 167, 172, 161, 150, 165, 217, 255, 259, 241, 236, 224, 200, 189, 192, 186, 190, 180, 157, 141, 134, 168, 208, 199, 181, 3, 
    209, 198, 259, 260, 206, 159, 147, 180, 181, 150, 158, 184, 225, 239, 248, 236, 223, 227, 205, 179, 212, 210, 189, 174, 155, 130, 122, 171, 191, 190, 189, 6, 
    209, 217, 284, 285, 253, 205, 176, 190, 182, 142, 166, 218, 237, 232, 222, 201, 188, 215, 215, 194, 222, 219, 181, 163, 155, 121, 95, 149, 178, 187, 170, 0, 
    204, 180, 225, 271, 273, 251, 218, 199, 183, 160, 171, 200, 212, 208, 181, 134, 134, 195, 222, 210, 217, 217, 185, 163, 146, 105, 54, 126, 180, 161, 146, 0, 
    177, 113, 121, 195, 258, 259, 253, 238, 204, 179, 185, 195, 193, 191, 166, 115, 109, 191, 234, 215, 221, 213, 179, 161, 139, 65, 37, 130, 171, 142, 120, 0, 
    159, 73, 39, 90, 191, 251, 267, 265, 245, 207, 182, 188, 192, 188, 174, 144, 137, 189, 228, 211, 204, 213, 185, 146, 95, 36, 58, 115, 163, 181, 148, 0, 
    167, 71, 22, 31, 99, 200, 261, 285, 277, 250, 219, 205, 201, 190, 182, 161, 146, 178, 205, 197, 206, 204, 158, 126, 76, 34, 75, 108, 150, 221, 184, 0, 
    161, 52, 35, 28, 46, 120, 208, 269, 284, 275, 260, 245, 229, 207, 212, 204, 154, 137, 164, 155, 150, 152, 136, 138, 113, 92, 132, 139, 186, 274, 191, 0, 
    118, 24, 57, 65, 26, 54, 125, 215, 261, 269, 270, 272, 262, 237, 239, 245, 200, 143, 137, 123, 127, 145, 162, 196, 181, 163, 170, 184, 231, 268, 203, 0, 
    33, 0, 3, 18, 0, 0, 20, 76, 106, 114, 121, 118, 102, 84, 89, 94, 57, 21, 32, 26, 14, 32, 53, 83, 80, 60, 64, 81, 92, 93, 62, 0, 
    
    -- channel=75
    33, 46, 51, 49, 30, 29, 36, 37, 47, 70, 47, 28, 31, 36, 44, 31, 23, 33, 40, 36, 42, 51, 41, 11, 26, 65, 39, 51, 60, 38, 37, 83, 
    12, 42, 54, 35, 17, 30, 34, 32, 50, 72, 42, 22, 30, 45, 49, 25, 25, 35, 42, 29, 30, 53, 36, 0, 11, 78, 42, 30, 33, 21, 37, 90, 
    14, 37, 55, 22, 17, 37, 33, 31, 57, 69, 38, 30, 36, 57, 54, 16, 19, 29, 24, 14, 23, 55, 30, 0, 9, 76, 29, 7, 11, 23, 51, 87, 
    22, 16, 43, 14, 26, 39, 33, 32, 64, 66, 45, 44, 42, 50, 40, 8, 22, 43, 34, 22, 26, 55, 26, 0, 0, 58, 20, 6, 14, 34, 37, 70, 
    31, 28, 55, 27, 35, 39, 37, 37, 72, 62, 45, 33, 24, 21, 24, 13, 17, 33, 42, 44, 35, 49, 18, 0, 0, 45, 24, 8, 12, 28, 24, 88, 
    27, 44, 54, 46, 32, 31, 40, 36, 77, 59, 33, 10, 9, 11, 22, 41, 45, 32, 46, 51, 15, 36, 21, 0, 0, 36, 21, 10, 0, 32, 50, 112, 
    28, 57, 22, 26, 26, 33, 46, 38, 74, 47, 11, 3, 12, 22, 53, 71, 47, 22, 57, 47, 0, 25, 18, 0, 0, 37, 20, 14, 0, 49, 64, 97, 
    30, 54, 0, 1, 12, 28, 45, 44, 56, 14, 0, 11, 17, 43, 76, 58, 10, 0, 47, 44, 0, 7, 2, 0, 0, 39, 22, 15, 7, 74, 74, 81, 
    35, 44, 0, 2, 18, 30, 32, 52, 51, 0, 0, 11, 30, 70, 69, 24, 0, 12, 17, 14, 0, 9, 17, 0, 0, 24, 16, 11, 19, 91, 72, 76, 
    41, 41, 0, 0, 15, 44, 32, 38, 44, 13, 15, 23, 39, 53, 25, 0, 3, 25, 11, 0, 0, 26, 44, 3, 0, 16, 11, 14, 29, 90, 62, 74, 
    43, 44, 0, 0, 7, 30, 48, 27, 0, 4, 23, 27, 45, 36, 0, 0, 0, 5, 11, 13, 13, 39, 30, 0, 0, 18, 12, 18, 31, 89, 61, 73, 
    57, 50, 0, 8, 10, 15, 44, 20, 0, 0, 12, 10, 33, 34, 26, 24, 20, 16, 20, 22, 19, 28, 22, 0, 0, 21, 15, 21, 34, 90, 55, 60, 
    43, 37, 0, 6, 6, 7, 26, 24, 14, 17, 17, 10, 26, 13, 0, 24, 40, 34, 24, 14, 23, 16, 16, 0, 7, 27, 6, 2, 37, 77, 33, 62, 
    38, 37, 1, 7, 13, 0, 14, 21, 33, 30, 31, 17, 21, 17, 6, 4, 11, 19, 22, 21, 29, 18, 15, 0, 8, 27, 14, 1, 38, 67, 33, 87, 
    41, 39, 16, 16, 22, 0, 7, 15, 7, 3, 22, 29, 28, 20, 21, 12, 5, 8, 6, 9, 20, 13, 10, 7, 10, 9, 12, 10, 49, 78, 34, 92, 
    34, 30, 9, 9, 13, 0, 0, 18, 7, 23, 33, 1, 9, 7, 1, 13, 24, 17, 3, 0, 0, 0, 0, 13, 17, 17, 2, 19, 61, 62, 0, 85, 
    25, 23, 3, 0, 19, 15, 12, 20, 1, 16, 57, 0, 0, 5, 5, 3, 3, 11, 23, 24, 28, 18, 0, 0, 24, 44, 17, 21, 61, 51, 0, 103, 
    15, 12, 11, 0, 28, 18, 29, 17, 12, 0, 32, 30, 0, 1, 17, 14, 5, 0, 0, 0, 5, 13, 19, 0, 10, 32, 58, 42, 58, 50, 0, 86, 
    8, 2, 27, 26, 44, 23, 28, 11, 11, 6, 0, 41, 23, 0, 0, 0, 6, 11, 0, 8, 19, 5, 11, 14, 19, 33, 35, 37, 40, 39, 0, 89, 
    6, 16, 42, 25, 41, 34, 15, 24, 23, 34, 0, 15, 43, 3, 0, 0, 0, 0, 3, 12, 15, 4, 4, 16, 21, 45, 21, 30, 13, 0, 1, 113, 
    12, 41, 34, 15, 31, 32, 5, 25, 17, 15, 29, 0, 0, 9, 0, 2, 4, 0, 3, 26, 21, 12, 14, 24, 19, 39, 37, 31, 3, 0, 0, 112, 
    28, 52, 14, 19, 33, 31, 13, 18, 19, 0, 30, 17, 0, 0, 1, 0, 0, 11, 0, 15, 21, 12, 4, 16, 16, 24, 29, 9, 1, 19, 14, 109, 
    26, 28, 0, 0, 7, 22, 11, 7, 27, 20, 12, 32, 0, 0, 0, 8, 1, 13, 20, 11, 1, 12, 8, 14, 21, 27, 25, 0, 4, 19, 19, 107, 
    1, 0, 0, 0, 0, 12, 4, 0, 15, 41, 12, 0, 0, 1, 0, 7, 6, 4, 18, 17, 0, 5, 4, 18, 25, 32, 31, 18, 22, 14, 15, 103, 
    11, 9, 0, 13, 12, 8, 7, 0, 9, 22, 16, 0, 0, 3, 2, 20, 25, 16, 18, 9, 0, 15, 17, 20, 23, 31, 30, 18, 31, 13, 28, 113, 
    10, 19, 8, 13, 19, 17, 6, 2, 14, 10, 1, 20, 18, 10, 28, 45, 39, 18, 15, 10, 0, 13, 24, 14, 19, 47, 52, 7, 21, 26, 40, 102, 
    12, 37, 18, 12, 18, 20, 16, 3, 0, 11, 0, 0, 13, 11, 23, 32, 16, 0, 0, 10, 8, 0, 21, 26, 30, 60, 61, 0, 19, 34, 30, 92, 
    13, 58, 40, 20, 8, 10, 3, 11, 4, 2, 8, 1, 0, 3, 10, 19, 5, 0, 0, 14, 10, 12, 15, 21, 55, 69, 28, 20, 27, 1, 3, 77, 
    13, 57, 48, 30, 0, 6, 0, 0, 7, 3, 0, 0, 1, 4, 5, 31, 38, 8, 0, 13, 3, 14, 37, 36, 50, 50, 21, 42, 0, 0, 34, 91, 
    20, 66, 49, 52, 19, 2, 6, 2, 5, 15, 8, 0, 0, 4, 0, 0, 16, 25, 20, 32, 39, 46, 47, 29, 28, 13, 0, 5, 0, 0, 39, 117, 
    41, 78, 30, 48, 44, 23, 6, 4, 2, 9, 19, 11, 1, 2, 0, 0, 0, 0, 0, 34, 26, 15, 2, 0, 10, 7, 1, 0, 0, 0, 23, 103, 
    76, 89, 55, 83, 98, 81, 49, 39, 69, 83, 92, 111, 129, 129, 113, 120, 144, 133, 92, 92, 78, 78, 86, 91, 116, 115, 108, 98, 107, 101, 121, 160, 
    
    -- channel=76
    13, 0, 8, 19, 25, 11, 9, 10, 9, 14, 33, 32, 15, 9, 10, 16, 12, 1, 0, 0, 0, 0, 7, 18, 0, 0, 20, 15, 7, 12, 8, 0, 
    6, 0, 0, 8, 8, 0, 0, 0, 0, 3, 23, 25, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 24, 22, 6, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 24, 22, 10, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 25, 23, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 24, 17, 2, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 3, 0, 0, 0, 0, 0, 0, 16, 21, 2, 0, 0, 0, 0, 6, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 7, 0, 0, 0, 0, 0, 0, 17, 11, 0, 0, 0, 0, 5, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 15, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 24, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 21, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 21, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 6, 22, 18, 6, 18, 31, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=77
    0, 48, 28, 0, 0, 2, 40, 48, 36, 0, 0, 0, 4, 38, 34, 49, 70, 107, 121, 126, 120, 98, 75, 105, 138, 116, 71, 7, 28, 40, 38, 0, 
    65, 166, 125, 76, 69, 105, 146, 146, 123, 52, 0, 9, 89, 122, 112, 128, 160, 205, 213, 220, 229, 201, 174, 222, 289, 235, 152, 77, 118, 143, 142, 58, 
    87, 216, 156, 130, 121, 160, 174, 164, 127, 50, 0, 16, 95, 112, 97, 122, 167, 212, 205, 205, 223, 197, 175, 234, 315, 261, 172, 102, 165, 193, 167, 50, 
    110, 264, 196, 193, 163, 190, 185, 181, 128, 46, 0, 0, 57, 84, 84, 119, 173, 208, 198, 199, 222, 187, 179, 248, 351, 314, 234, 182, 242, 252, 217, 54, 
    112, 253, 218, 208, 184, 193, 181, 186, 113, 39, 0, 0, 50, 95, 118, 158, 200, 221, 202, 181, 198, 167, 189, 278, 387, 380, 324, 266, 305, 301, 263, 95, 
    99, 208, 192, 170, 180, 193, 181, 173, 84, 30, 0, 34, 103, 163, 180, 177, 176, 195, 174, 155, 157, 150, 215, 316, 425, 451, 399, 321, 348, 319, 286, 109, 
    72, 150, 152, 133, 185, 202, 181, 149, 57, 28, 30, 115, 201, 224, 190, 139, 100, 140, 159, 141, 144, 168, 254, 333, 457, 483, 443, 364, 388, 333, 263, 58, 
    52, 129, 142, 177, 247, 235, 195, 140, 68, 61, 97, 208, 267, 229, 158, 75, 59, 127, 181, 167, 186, 242, 300, 362, 465, 485, 458, 398, 414, 312, 191, 0, 
    52, 144, 180, 252, 341, 285, 214, 142, 96, 126, 192, 283, 278, 198, 99, 42, 89, 187, 231, 223, 262, 307, 323, 373, 436, 470, 461, 420, 409, 270, 128, 0, 
    65, 172, 216, 313, 413, 358, 251, 152, 122, 169, 254, 319, 288, 199, 111, 102, 193, 263, 275, 286, 334, 336, 316, 346, 387, 454, 456, 425, 401, 235, 88, 0, 
    76, 185, 213, 316, 440, 422, 309, 200, 165, 208, 293, 325, 285, 240, 208, 253, 321, 331, 324, 331, 352, 333, 301, 333, 386, 452, 449, 431, 398, 211, 58, 0, 
    68, 165, 180, 283, 420, 444, 388, 295, 248, 271, 318, 321, 285, 267, 281, 334, 372, 364, 348, 347, 339, 317, 281, 342, 406, 437, 431, 423, 383, 212, 68, 0, 
    76, 168, 176, 263, 378, 437, 433, 393, 346, 337, 325, 320, 298, 300, 324, 355, 365, 354, 346, 347, 337, 330, 313, 374, 414, 421, 418, 415, 378, 241, 112, 0, 
    84, 197, 193, 261, 335, 407, 436, 457, 408, 353, 318, 318, 308, 314, 323, 345, 347, 332, 331, 335, 336, 355, 359, 397, 403, 405, 390, 409, 378, 258, 160, 10, 
    103, 223, 213, 265, 317, 374, 421, 467, 455, 382, 320, 297, 288, 324, 348, 362, 362, 356, 345, 342, 334, 365, 391, 430, 436, 405, 399, 406, 357, 238, 172, 23, 
    111, 233, 231, 283, 332, 376, 421, 440, 457, 422, 341, 306, 280, 348, 388, 394, 400, 396, 386, 394, 385, 388, 407, 459, 472, 436, 418, 394, 326, 212, 157, 27, 
    110, 250, 253, 310, 337, 385, 395, 421, 435, 458, 398, 352, 324, 368, 408, 431, 433, 418, 413, 410, 405, 406, 414, 458, 469, 463, 401, 386, 304, 178, 148, 38, 
    123, 292, 306, 351, 346, 367, 346, 376, 379, 420, 438, 412, 398, 398, 405, 439, 440, 450, 463, 463, 453, 438, 414, 435, 451, 418, 353, 314, 263, 196, 216, 84, 
    149, 343, 338, 362, 308, 296, 291, 322, 354, 363, 419, 443, 442, 438, 434, 462, 470, 474, 475, 464, 447, 432, 421, 428, 413, 355, 306, 239, 221, 223, 263, 143, 
    174, 359, 342, 327, 261, 244, 252, 265, 321, 326, 337, 389, 408, 437, 470, 497, 505, 504, 509, 501, 471, 438, 430, 426, 401, 328, 272, 215, 231, 253, 329, 203, 
    185, 344, 309, 265, 253, 237, 239, 263, 292, 309, 294, 333, 376, 446, 515, 539, 536, 513, 516, 491, 460, 431, 425, 410, 393, 323, 276, 255, 274, 318, 397, 225, 
    174, 303, 254, 245, 270, 242, 244, 271, 294, 307, 311, 316, 371, 448, 537, 560, 557, 534, 514, 470, 447, 426, 428, 412, 390, 343, 307, 306, 331, 383, 405, 204, 
    158, 304, 307, 340, 361, 292, 263, 288, 316, 333, 325, 332, 380, 459, 538, 548, 554, 532, 499, 461, 436, 419, 431, 411, 391, 347, 316, 329, 377, 411, 388, 193, 
    179, 376, 428, 484, 472, 386, 321, 325, 346, 353, 337, 343, 411, 464, 525, 527, 535, 524, 498, 460, 454, 443, 458, 420, 387, 332, 299, 329, 362, 393, 373, 197, 
    181, 410, 498, 567, 568, 489, 412, 377, 363, 346, 338, 372, 442, 481, 492, 480, 472, 476, 481, 473, 477, 473, 468, 417, 376, 316, 279, 295, 313, 369, 350, 189, 
    181, 372, 431, 504, 557, 562, 504, 448, 396, 351, 344, 378, 426, 445, 429, 387, 360, 387, 440, 478, 485, 493, 466, 418, 367, 306, 229, 236, 262, 334, 322, 145, 
    146, 266, 272, 324, 438, 519, 544, 514, 462, 402, 375, 379, 399, 402, 380, 325, 278, 325, 401, 473, 501, 484, 451, 414, 356, 272, 188, 182, 240, 315, 265, 107, 
    121, 210, 157, 143, 266, 396, 510, 549, 536, 478, 415, 375, 367, 367, 356, 320, 296, 329, 395, 455, 476, 472, 450, 404, 313, 215, 152, 148, 263, 310, 288, 151, 
    127, 211, 133, 52, 120, 249, 411, 535, 581, 557, 498, 440, 403, 379, 368, 342, 332, 345, 386, 426, 455, 457, 428, 365, 259, 170, 132, 159, 254, 311, 363, 203, 
    119, 196, 135, 32, 66, 130, 281, 433, 543, 585, 573, 534, 491, 447, 428, 403, 367, 333, 336, 338, 368, 363, 348, 324, 266, 228, 221, 236, 299, 395, 420, 230, 
    76, 153, 117, 67, 81, 74, 149, 295, 432, 535, 573, 579, 566, 527, 499, 478, 441, 368, 316, 278, 295, 290, 314, 356, 361, 365, 334, 340, 389, 461, 450, 236, 
    0, 11, 0, 0, 5, 0, 0, 73, 171, 246, 286, 311, 313, 285, 265, 261, 233, 168, 116, 85, 76, 71, 110, 172, 210, 216, 197, 207, 229, 250, 224, 99, 
    
    -- channel=78
    0, 0, 2, 12, 28, 18, 12, 10, 1, 0, 17, 27, 19, 16, 9, 17, 17, 5, 4, 7, 1, 0, 7, 27, 0, 0, 21, 0, 0, 15, 6, 0, 
    55, 66, 59, 67, 67, 61, 82, 82, 69, 49, 52, 61, 69, 70, 67, 83, 95, 111, 118, 128, 122, 98, 94, 121, 114, 89, 105, 98, 102, 91, 67, 30, 
    59, 78, 66, 81, 79, 83, 94, 85, 65, 50, 51, 61, 78, 74, 76, 102, 113, 126, 134, 130, 116, 94, 99, 124, 125, 100, 117, 96, 86, 75, 66, 38, 
    57, 106, 83, 94, 86, 97, 91, 80, 62, 50, 44, 57, 79, 81, 85, 99, 94, 90, 93, 99, 106, 94, 100, 126, 136, 110, 103, 73, 80, 89, 101, 53, 
    56, 85, 65, 95, 94, 100, 80, 75, 56, 53, 51, 75, 90, 96, 79, 86, 107, 109, 94, 88, 107, 102, 108, 125, 136, 109, 104, 105, 119, 118, 102, 15, 
    68, 86, 92, 93, 107, 97, 74, 77, 51, 52, 61, 82, 89, 96, 91, 84, 89, 106, 94, 91, 124, 100, 104, 142, 143, 123, 134, 129, 138, 104, 70, 23, 
    64, 87, 127, 110, 97, 81, 70, 74, 48, 59, 75, 86, 109, 120, 97, 90, 105, 103, 68, 89, 110, 93, 122, 155, 144, 132, 140, 125, 127, 91, 95, 59, 
    64, 85, 112, 103, 107, 92, 74, 68, 64, 83, 87, 111, 154, 138, 113, 120, 119, 106, 75, 76, 100, 120, 151, 165, 172, 138, 138, 123, 121, 83, 80, 35, 
    54, 83, 93, 93, 100, 99, 88, 55, 55, 89, 107, 148, 154, 120, 117, 104, 82, 87, 130, 112, 98, 132, 141, 169, 184, 161, 145, 130, 117, 68, 57, 11, 
    49, 82, 106, 114, 122, 94, 98, 82, 63, 83, 110, 136, 131, 127, 117, 90, 91, 122, 138, 132, 140, 146, 148, 192, 173, 159, 145, 126, 113, 72, 56, 5, 
    50, 81, 107, 120, 136, 119, 86, 98, 124, 119, 132, 132, 101, 94, 95, 103, 143, 161, 145, 143, 156, 149, 180, 210, 166, 156, 147, 125, 113, 63, 46, 4, 
    33, 79, 100, 111, 134, 133, 102, 108, 127, 130, 152, 136, 92, 69, 52, 76, 116, 135, 150, 153, 152, 146, 134, 144, 157, 163, 146, 125, 111, 61, 58, 21, 
    59, 93, 105, 117, 139, 139, 128, 98, 92, 123, 134, 113, 98, 114, 130, 117, 111, 122, 132, 127, 113, 125, 115, 145, 162, 153, 163, 150, 113, 82, 75, 7, 
    48, 73, 92, 109, 122, 143, 138, 127, 115, 115, 102, 112, 107, 101, 116, 133, 136, 121, 103, 91, 83, 93, 102, 140, 147, 139, 146, 143, 119, 85, 55, 0, 
    47, 85, 89, 102, 113, 145, 138, 145, 149, 137, 112, 101, 100, 102, 96, 107, 110, 107, 116, 116, 103, 101, 96, 105, 124, 142, 132, 142, 115, 69, 79, 32, 
    69, 107, 114, 118, 123, 132, 142, 132, 116, 79, 96, 131, 114, 122, 132, 107, 87, 101, 116, 125, 123, 131, 106, 94, 106, 106, 132, 130, 110, 103, 125, 34, 
    69, 104, 114, 121, 106, 105, 127, 131, 143, 110, 75, 118, 106, 98, 107, 121, 137, 117, 88, 85, 77, 92, 128, 137, 90, 78, 115, 123, 107, 94, 81, 3, 
    69, 106, 106, 127, 113, 128, 122, 139, 136, 143, 90, 62, 88, 102, 96, 105, 113, 127, 147, 145, 139, 123, 104, 116, 124, 114, 66, 104, 94, 78, 120, 51, 
    72, 117, 97, 104, 112, 126, 120, 135, 129, 129, 125, 72, 98, 127, 122, 126, 102, 103, 116, 106, 101, 126, 122, 113, 112, 99, 118, 117, 103, 93, 115, 33, 
    71, 105, 98, 131, 118, 107, 123, 105, 112, 106, 138, 119, 80, 102, 105, 102, 122, 124, 109, 111, 121, 122, 121, 115, 105, 86, 110, 90, 118, 135, 101, 31, 
    69, 101, 124, 130, 109, 108, 119, 108, 139, 133, 105, 158, 130, 101, 120, 109, 112, 121, 116, 103, 104, 101, 104, 107, 110, 89, 68, 78, 105, 111, 136, 71, 
    64, 110, 126, 97, 109, 109, 105, 113, 120, 145, 100, 105, 146, 126, 115, 128, 121, 103, 126, 119, 105, 114, 126, 116, 116, 104, 99, 115, 96, 97, 147, 77, 
    76, 124, 144, 150, 145, 129, 127, 121, 98, 104, 132, 95, 111, 130, 133, 120, 121, 112, 101, 114, 124, 106, 107, 109, 107, 108, 114, 119, 117, 150, 163, 77, 
    96, 134, 110, 120, 153, 154, 157, 155, 128, 107, 134, 149, 113, 117, 144, 127, 126, 126, 110, 103, 110, 110, 115, 105, 114, 121, 109, 106, 136, 164, 160, 79, 
    61, 92, 108, 145, 167, 178, 166, 164, 157, 146, 115, 123, 145, 125, 127, 112, 108, 109, 104, 109, 118, 91, 101, 108, 126, 123, 114, 135, 143, 161, 144, 66, 
    84, 141, 164, 182, 180, 183, 194, 187, 172, 165, 142, 100, 111, 126, 106, 103, 109, 116, 106, 105, 110, 108, 108, 119, 110, 83, 96, 148, 143, 145, 145, 90, 
    90, 130, 153, 171, 178, 190, 191, 207, 203, 172, 174, 183, 165, 154, 143, 143, 141, 136, 118, 105, 110, 135, 106, 91, 89, 80, 89, 137, 126, 150, 165, 74, 
    76, 89, 116, 147, 178, 195, 209, 192, 196, 203, 190, 185, 190, 175, 160, 131, 117, 130, 110, 108, 117, 106, 115, 111, 81, 86, 115, 90, 123, 184, 157, 71, 
    72, 93, 98, 115, 156, 167, 199, 208, 195, 202, 214, 203, 197, 193, 176, 129, 96, 105, 120, 114, 121, 111, 94, 104, 109, 104, 88, 85, 169, 137, 102, 72, 
    69, 83, 86, 68, 111, 150, 170, 200, 202, 186, 193, 210, 210, 203, 210, 205, 178, 134, 116, 97, 80, 84, 102, 122, 117, 112, 112, 146, 170, 159, 155, 72, 
    62, 92, 121, 81, 88, 113, 160, 190, 213, 210, 193, 186, 197, 200, 206, 195, 182, 180, 157, 117, 134, 152, 153, 140, 104, 99, 107, 107, 121, 181, 185, 95, 
    32, 71, 57, 27, 29, 41, 83, 113, 104, 114, 105, 72, 50, 51, 55, 34, 5, 9, 45, 53, 52, 23, 1, 0, 0, 9, 11, 19, 32, 55, 46, 8, 
    
    -- channel=79
    26, 8, 8, 20, 25, 14, 0, 0, 0, 0, 23, 30, 12, 5, 8, 10, 4, 0, 0, 0, 0, 0, 0, 11, 0, 0, 17, 17, 10, 17, 12, 0, 
    36, 0, 0, 1, 4, 0, 0, 0, 0, 0, 1, 20, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 3, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 13, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 29, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 30, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 17, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    29, 0, 0, 0, 0, 0, 0, 0, 6, 6, 4, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    28, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 17, 6, 11, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 21, 20, 1, 7, 14, 5, 4, 7, 8, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 14, 18, 14, 8, 9, 7, 6, 17, 15, 12, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 24, 9, 13, 3, 0, 6, 4, 7, 0, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 12, 3, 3, 8, 0, 0, 2, 2, 0, 8, 8, 0, 0, 0, 0, 0, 0, 0, 12, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 4, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 2, 0, 0, 0, 0, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    27, 0, 0, 10, 31, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    30, 0, 0, 0, 12, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 17, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 15, 8, 29, 3, 20, 38, 40, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 11, 18, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=80
    157, 134, 119, 105, 115, 118, 121, 118, 116, 124, 114, 118, 123, 125, 117, 107, 117, 119, 114, 110, 117, 117, 121, 111, 114, 116, 114, 106, 127, 115, 116, 148, 
    111, 138, 117, 65, 75, 96, 98, 95, 90, 114, 102, 100, 107, 120, 112, 86, 105, 122, 115, 93, 98, 106, 114, 110, 107, 107, 93, 73, 109, 114, 103, 179, 
    104, 97, 83, 84, 100, 93, 83, 94, 95, 111, 104, 111, 111, 111, 120, 99, 110, 130, 117, 92, 94, 101, 104, 115, 110, 97, 85, 81, 100, 109, 104, 187, 
    72, 69, 72, 104, 116, 91, 86, 96, 87, 103, 104, 106, 116, 109, 104, 109, 115, 149, 140, 94, 88, 95, 92, 93, 91, 95, 96, 104, 104, 99, 101, 191, 
    55, 71, 67, 107, 115, 85, 87, 95, 86, 94, 98, 96, 110, 115, 95, 107, 128, 141, 158, 110, 86, 100, 104, 87, 82, 92, 97, 112, 115, 90, 88, 200, 
    56, 86, 64, 100, 103, 82, 83, 90, 91, 89, 92, 99, 109, 120, 107, 84, 110, 117, 146, 135, 85, 90, 115, 95, 85, 87, 92, 101, 108, 94, 86, 203, 
    63, 91, 66, 80, 94, 87, 85, 86, 86, 83, 99, 96, 98, 113, 121, 84, 90, 98, 113, 128, 93, 76, 122, 104, 94, 102, 93, 92, 96, 95, 89, 205, 
    86, 88, 62, 71, 91, 87, 85, 80, 82, 78, 98, 96, 91, 98, 116, 98, 86, 83, 90, 107, 123, 93, 129, 115, 94, 116, 107, 90, 91, 90, 88, 206, 
    85, 78, 59, 81, 89, 86, 82, 70, 86, 90, 97, 94, 96, 94, 106, 103, 90, 77, 89, 95, 128, 93, 119, 121, 97, 109, 104, 88, 87, 92, 87, 206, 
    55, 71, 79, 79, 80, 84, 91, 79, 82, 93, 94, 84, 89, 97, 93, 100, 99, 84, 76, 81, 105, 75, 106, 134, 98, 94, 87, 92, 90, 97, 89, 206, 
    55, 73, 81, 63, 70, 89, 95, 86, 75, 77, 89, 91, 84, 75, 48, 77, 109, 104, 75, 76, 90, 72, 93, 139, 101, 96, 95, 96, 90, 95, 91, 204, 
    69, 53, 81, 84, 74, 81, 80, 74, 86, 83, 85, 67, 62, 60, 23, 37, 99, 124, 80, 78, 84, 82, 116, 134, 96, 91, 105, 99, 89, 90, 87, 205, 
    64, 3, 75, 88, 61, 57, 70, 74, 97, 84, 57, 16, 44, 85, 85, 68, 75, 127, 77, 64, 91, 93, 134, 123, 86, 87, 103, 103, 90, 91, 88, 202, 
    64, 0, 46, 56, 52, 64, 73, 87, 99, 64, 36, 19, 59, 91, 112, 134, 57, 78, 70, 49, 90, 105, 127, 120, 102, 93, 100, 104, 89, 93, 93, 198, 
    74, 32, 37, 39, 57, 70, 57, 83, 93, 39, 33, 66, 90, 73, 61, 96, 45, 45, 57, 61, 93, 117, 125, 113, 102, 89, 96, 111, 92, 95, 96, 191, 
    90, 97, 39, 15, 51, 74, 63, 53, 65, 33, 40, 73, 100, 55, 27, 43, 35, 42, 42, 71, 100, 116, 114, 105, 98, 85, 78, 107, 114, 91, 93, 189, 
    98, 121, 43, 8, 48, 77, 92, 38, 30, 34, 32, 41, 94, 66, 23, 36, 47, 47, 35, 55, 75, 117, 119, 117, 107, 73, 54, 78, 138, 109, 80, 186, 
    84, 106, 51, 22, 46, 64, 106, 41, 0, 62, 59, 44, 80, 71, 36, 51, 49, 65, 47, 46, 78, 141, 149, 138, 114, 57, 43, 58, 129, 141, 79, 175, 
    75, 92, 39, 28, 46, 51, 114, 77, 0, 99, 103, 24, 55, 100, 80, 112, 54, 76, 89, 86, 123, 149, 148, 135, 99, 59, 30, 54, 107, 157, 91, 166, 
    79, 116, 49, 10, 31, 49, 109, 138, 0, 39, 92, 17, 71, 132, 57, 109, 99, 92, 121, 114, 138, 124, 107, 120, 85, 63, 27, 36, 90, 172, 109, 155, 
    82, 114, 54, 3, 17, 40, 92, 195, 47, 0, 46, 49, 91, 112, 7, 48, 135, 142, 138, 101, 110, 96, 87, 132, 104, 65, 21, 10, 62, 183, 134, 150, 
    71, 94, 61, 20, 26, 53, 101, 204, 152, 59, 42, 62, 93, 116, 51, 45, 105, 144, 156, 101, 92, 97, 87, 131, 122, 71, 11, 0, 43, 169, 156, 156, 
    62, 101, 84, 34, 31, 78, 132, 174, 141, 119, 108, 98, 92, 109, 86, 82, 102, 112, 140, 124, 109, 112, 84, 92, 107, 86, 47, 0, 32, 154, 174, 162, 
    66, 96, 94, 58, 34, 79, 135, 130, 101, 106, 132, 116, 103, 85, 87, 124, 146, 123, 119, 121, 115, 125, 106, 84, 91, 92, 88, 14, 15, 128, 188, 174, 
    86, 83, 69, 83, 61, 48, 78, 99, 135, 109, 108, 84, 95, 96, 114, 151, 154, 128, 120, 112, 113, 121, 119, 111, 87, 75, 100, 60, 19, 69, 169, 206, 
    86, 76, 59, 89, 104, 47, 20, 69, 157, 84, 80, 95, 88, 108, 119, 125, 135, 126, 129, 124, 127, 125, 114, 124, 89, 71, 121, 105, 62, 42, 85, 226, 
    66, 79, 74, 74, 99, 87, 60, 23, 107, 97, 78, 122, 84, 83, 105, 114, 120, 123, 127, 122, 126, 130, 112, 115, 102, 97, 127, 101, 71, 89, 47, 206, 
    63, 88, 73, 54, 79, 97, 120, 49, 57, 129, 103, 103, 62, 65, 100, 123, 109, 107, 108, 103, 112, 122, 101, 102, 114, 115, 106, 78, 49, 124, 107, 193, 
    57, 107, 89, 52, 77, 100, 114, 90, 75, 103, 98, 95, 67, 69, 88, 118, 103, 85, 93, 99, 110, 105, 84, 94, 107, 104, 99, 95, 84, 108, 103, 206, 
    61, 114, 89, 64, 79, 105, 95, 76, 105, 91, 62, 87, 87, 80, 79, 98, 99, 91, 107, 99, 95, 93, 81, 89, 100, 93, 97, 114, 116, 82, 57, 216, 
    69, 83, 66, 76, 78, 80, 85, 74, 85, 77, 71, 91, 95, 95, 88, 85, 102, 106, 113, 91, 81, 91, 83, 80, 96, 89, 94, 114, 106, 72, 64, 221, 
    16, 45, 50, 79, 83, 62, 61, 61, 73, 57, 64, 77, 80, 91, 96, 73, 76, 77, 79, 74, 61, 67, 62, 54, 71, 75, 70, 79, 77, 60, 62, 211, 
    
    -- channel=81
    28, 71, 47, 71, 87, 81, 72, 73, 82, 74, 69, 64, 61, 51, 49, 49, 41, 33, 17, 12, 7, 9, 7, 4, 1, 0, 3, 23, 24, 19, 10, 0, 
    45, 161, 144, 143, 133, 133, 128, 132, 137, 133, 135, 121, 116, 107, 94, 93, 87, 81, 57, 35, 31, 42, 48, 49, 47, 51, 59, 63, 58, 59, 45, 0, 
    55, 189, 175, 171, 158, 142, 132, 142, 150, 144, 146, 134, 128, 120, 112, 105, 98, 72, 46, 25, 19, 36, 47, 53, 59, 64, 67, 66, 62, 58, 52, 9, 
    61, 193, 182, 180, 164, 148, 142, 154, 161, 155, 156, 153, 144, 129, 121, 115, 107, 95, 61, 37, 21, 31, 43, 51, 57, 63, 74, 71, 63, 62, 62, 10, 
    64, 189, 186, 173, 175, 163, 152, 164, 165, 162, 169, 161, 154, 143, 129, 125, 124, 119, 94, 65, 51, 54, 64, 66, 62, 70, 74, 74, 73, 70, 71, 18, 
    66, 189, 176, 172, 185, 170, 164, 172, 170, 177, 176, 174, 166, 158, 141, 136, 135, 136, 124, 110, 97, 89, 79, 73, 56, 56, 64, 65, 71, 74, 76, 22, 
    55, 182, 163, 177, 182, 173, 169, 175, 181, 186, 184, 180, 171, 162, 147, 143, 140, 151, 149, 143, 119, 103, 84, 80, 61, 51, 51, 52, 64, 75, 80, 22, 
    46, 175, 172, 171, 179, 175, 173, 180, 179, 187, 182, 173, 163, 162, 147, 138, 131, 139, 140, 148, 137, 133, 115, 106, 72, 53, 55, 63, 71, 76, 82, 22, 
    46, 177, 154, 169, 183, 182, 177, 177, 177, 185, 184, 181, 169, 161, 151, 145, 140, 134, 131, 138, 140, 150, 128, 115, 83, 56, 65, 66, 71, 75, 80, 19, 
    31, 143, 140, 178, 183, 183, 183, 182, 190, 195, 188, 173, 167, 169, 171, 170, 165, 142, 124, 125, 131, 146, 134, 112, 79, 49, 59, 61, 67, 72, 80, 23, 
    0, 96, 131, 166, 165, 171, 188, 195, 188, 186, 178, 187, 202, 208, 197, 179, 176, 155, 128, 119, 132, 135, 110, 84, 55, 44, 54, 60, 66, 70, 78, 18, 
    0, 80, 128, 185, 194, 211, 218, 201, 188, 183, 186, 213, 229, 217, 178, 156, 142, 114, 120, 117, 127, 126, 90, 63, 47, 31, 42, 48, 55, 63, 73, 16, 
    0, 72, 127, 193, 200, 213, 215, 205, 188, 181, 191, 225, 230, 215, 179, 143, 153, 139, 149, 147, 139, 125, 78, 44, 18, 18, 37, 45, 53, 58, 62, 7, 
    0, 73, 122, 174, 203, 225, 225, 204, 195, 202, 212, 226, 217, 205, 187, 176, 181, 177, 193, 180, 170, 132, 78, 45, 18, 26, 39, 48, 57, 51, 55, 1, 
    6, 70, 98, 157, 202, 230, 220, 206, 203, 221, 231, 243, 233, 224, 209, 215, 227, 210, 223, 215, 188, 151, 99, 53, 25, 29, 47, 66, 75, 60, 46, 0, 
    12, 83, 105, 136, 188, 219, 201, 193, 204, 234, 251, 265, 238, 218, 208, 220, 242, 234, 239, 227, 217, 172, 107, 43, 13, 22, 58, 95, 93, 74, 46, 0, 
    20, 101, 110, 144, 196, 223, 203, 195, 199, 227, 244, 225, 211, 221, 206, 201, 208, 210, 214, 204, 185, 128, 69, 12, 0, 17, 57, 108, 116, 86, 48, 0, 
    27, 112, 122, 142, 195, 233, 202, 176, 180, 190, 225, 215, 219, 215, 173, 137, 166, 150, 148, 128, 95, 62, 25, 0, 0, 16, 66, 118, 140, 107, 56, 0, 
    28, 106, 114, 141, 201, 238, 216, 167, 157, 146, 212, 223, 197, 184, 170, 158, 182, 142, 98, 68, 40, 28, 13, 0, 4, 18, 69, 129, 161, 134, 70, 0, 
    28, 115, 129, 156, 204, 241, 223, 144, 99, 77, 139, 167, 167, 162, 157, 147, 158, 116, 68, 31, 13, 22, 14, 0, 2, 13, 66, 136, 191, 157, 94, 0, 
    35, 132, 133, 140, 183, 225, 205, 116, 47, 1, 58, 84, 88, 92, 97, 97, 125, 89, 37, 14, 0, 0, 3, 2, 14, 22, 74, 135, 194, 179, 116, 0, 
    42, 138, 130, 135, 169, 197, 176, 105, 49, 2, 18, 36, 40, 44, 53, 61, 81, 59, 11, 0, 0, 0, 0, 0, 11, 26, 58, 116, 171, 180, 128, 6, 
    38, 138, 125, 133, 155, 174, 165, 124, 89, 49, 22, 21, 39, 57, 61, 46, 19, 0, 0, 0, 0, 0, 0, 0, 0, 9, 34, 89, 140, 160, 134, 25, 
    25, 125, 123, 130, 147, 161, 172, 174, 131, 83, 55, 59, 55, 60, 55, 30, 13, 0, 0, 0, 0, 0, 0, 0, 0, 6, 29, 60, 87, 128, 129, 49, 
    24, 131, 133, 132, 129, 145, 168, 176, 154, 146, 113, 105, 88, 72, 67, 61, 35, 5, 0, 0, 0, 0, 0, 0, 0, 0, 8, 24, 34, 83, 106, 47, 
    29, 129, 123, 136, 144, 145, 147, 166, 154, 162, 115, 87, 92, 99, 105, 90, 61, 36, 13, 3, 0, 0, 0, 0, 0, 3, 4, 22, 40, 66, 105, 28, 
    30, 122, 126, 129, 138, 146, 122, 135, 145, 142, 128, 104, 105, 108, 117, 104, 84, 62, 53, 52, 41, 27, 25, 29, 39, 34, 38, 51, 59, 62, 72, 13, 
    30, 118, 115, 117, 129, 140, 118, 107, 107, 124, 105, 99, 121, 116, 127, 116, 99, 91, 86, 78, 63, 62, 69, 71, 77, 74, 70, 68, 67, 62, 72, 13, 
    22, 96, 112, 121, 133, 133, 124, 124, 110, 121, 132, 114, 118, 116, 126, 118, 110, 99, 88, 79, 77, 87, 96, 100, 107, 105, 96, 88, 76, 75, 105, 33, 
    21, 119, 138, 134, 135, 135, 128, 127, 125, 132, 133, 132, 134, 117, 113, 106, 100, 98, 89, 90, 91, 97, 108, 117, 121, 121, 111, 102, 90, 90, 97, 37, 
    33, 131, 147, 135, 124, 110, 104, 117, 124, 134, 120, 122, 122, 110, 104, 96, 91, 97, 98, 99, 99, 109, 121, 127, 130, 126, 117, 111, 111, 109, 110, 44, 
    0, 7, 9, 4, 1, 0, 2, 4, 1, 4, 10, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    33, 0, 19, 31, 12, 8, 18, 22, 14, 6, 15, 17, 13, 12, 13, 24, 12, 0, 4, 20, 23, 18, 14, 18, 16, 22, 30, 33, 6, 4, 15, 0, 
    58, 0, 18, 24, 13, 17, 36, 32, 27, 19, 23, 27, 24, 21, 25, 40, 20, 0, 0, 29, 37, 29, 24, 22, 24, 28, 31, 37, 12, 7, 18, 0, 
    66, 9, 18, 3, 0, 22, 42, 22, 26, 21, 19, 25, 23, 25, 29, 34, 18, 0, 1, 33, 42, 33, 30, 23, 27, 29, 29, 25, 13, 20, 27, 0, 
    81, 14, 13, 0, 0, 28, 38, 19, 27, 23, 22, 21, 15, 23, 35, 35, 25, 3, 0, 24, 42, 39, 31, 29, 39, 33, 24, 16, 15, 28, 29, 0, 
    92, 0, 11, 5, 0, 26, 34, 21, 28, 26, 20, 22, 18, 17, 30, 39, 31, 15, 0, 6, 35, 37, 19, 28, 41, 32, 28, 19, 17, 32, 32, 0, 
    87, 0, 23, 13, 0, 23, 28, 24, 28, 26, 17, 17, 25, 15, 19, 42, 36, 30, 7, 0, 19, 27, 5, 17, 39, 34, 31, 33, 27, 29, 31, 0, 
    68, 0, 36, 10, 0, 17, 25, 29, 25, 23, 11, 18, 28, 16, 13, 38, 42, 38, 21, 0, 10, 26, 11, 13, 31, 26, 32, 45, 37, 29, 31, 0, 
    62, 0, 25, 10, 8, 16, 22, 29, 25, 17, 9, 26, 32, 20, 16, 31, 38, 40, 36, 23, 8, 29, 12, 0, 23, 25, 35, 43, 35, 31, 30, 0, 
    69, 1, 23, 17, 11, 15, 17, 27, 26, 19, 18, 27, 26, 21, 26, 30, 22, 27, 37, 41, 15, 34, 15, 0, 12, 31, 34, 35, 33, 28, 29, 0, 
    70, 14, 37, 17, 12, 15, 13, 28, 25, 13, 16, 29, 28, 18, 32, 23, 0, 3, 35, 49, 30, 41, 11, 0, 8, 39, 32, 29, 33, 28, 31, 0, 
    62, 58, 46, 6, 24, 28, 15, 20, 19, 14, 29, 41, 24, 0, 16, 18, 0, 0, 30, 48, 30, 32, 1, 0, 25, 38, 28, 29, 34, 30, 32, 0, 
    71, 107, 49, 4, 34, 19, 7, 16, 6, 16, 45, 49, 2, 0, 0, 0, 0, 0, 28, 42, 22, 12, 0, 0, 28, 35, 27, 31, 39, 35, 32, 0, 
    84, 123, 41, 14, 35, 10, 4, 3, 0, 25, 58, 41, 0, 0, 0, 0, 3, 6, 16, 27, 1, 0, 0, 0, 32, 37, 29, 31, 39, 32, 32, 0, 
    87, 86, 42, 52, 32, 0, 0, 0, 0, 32, 42, 6, 0, 0, 0, 0, 15, 6, 0, 10, 0, 0, 0, 0, 23, 30, 32, 29, 33, 28, 29, 0, 
    71, 38, 61, 76, 28, 0, 0, 0, 3, 33, 22, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 30, 45, 27, 13, 15, 31, 0, 
    64, 9, 61, 86, 31, 0, 0, 14, 28, 29, 0, 0, 0, 7, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 13, 44, 60, 27, 0, 0, 28, 0, 
    65, 12, 64, 79, 28, 0, 0, 13, 54, 13, 0, 2, 0, 0, 24, 14, 3, 0, 0, 0, 0, 0, 0, 0, 21, 60, 75, 39, 0, 0, 18, 0, 
    77, 15, 54, 77, 31, 0, 0, 0, 77, 8, 0, 29, 2, 0, 9, 24, 16, 12, 0, 4, 0, 0, 0, 13, 30, 71, 79, 51, 0, 0, 0, 0, 
    78, 14, 59, 83, 37, 0, 0, 0, 78, 29, 0, 28, 0, 0, 27, 24, 0, 0, 0, 11, 2, 0, 18, 17, 32, 66, 82, 62, 0, 0, 0, 0, 
    78, 12, 58, 83, 39, 0, 0, 0, 47, 67, 24, 37, 0, 0, 49, 31, 0, 0, 0, 18, 16, 15, 31, 12, 28, 63, 94, 78, 0, 0, 0, 0, 
    81, 7, 41, 81, 49, 0, 0, 0, 9, 89, 46, 36, 10, 0, 69, 55, 0, 0, 0, 22, 27, 25, 38, 14, 24, 59, 92, 92, 13, 0, 0, 0, 
    85, 6, 29, 70, 48, 0, 0, 0, 0, 55, 39, 31, 23, 18, 67, 62, 0, 0, 3, 31, 37, 25, 37, 28, 29, 51, 83, 95, 38, 0, 0, 0, 
    81, 4, 30, 58, 46, 0, 0, 0, 0, 0, 17, 35, 31, 25, 40, 22, 8, 23, 18, 28, 34, 23, 37, 44, 38, 51, 66, 87, 60, 0, 0, 0, 
    71, 19, 43, 40, 33, 15, 0, 0, 0, 0, 17, 23, 24, 28, 26, 4, 0, 17, 24, 23, 26, 19, 31, 43, 46, 59, 40, 63, 81, 5, 0, 0, 
    71, 33, 41, 23, 24, 30, 21, 0, 0, 1, 22, 12, 20, 33, 18, 0, 0, 5, 12, 18, 19, 15, 22, 28, 47, 60, 23, 43, 88, 51, 0, 0, 
    76, 38, 45, 29, 17, 27, 27, 20, 0, 0, 12, 16, 38, 39, 13, 1, 0, 4, 6, 13, 12, 9, 23, 22, 32, 39, 15, 39, 77, 51, 5, 0, 
    86, 32, 29, 46, 26, 7, 13, 44, 16, 0, 0, 7, 40, 41, 14, 2, 5, 16, 14, 10, 3, 5, 27, 24, 16, 20, 13, 34, 55, 15, 22, 0, 
    88, 16, 23, 59, 32, 0, 0, 48, 35, 0, 18, 26, 37, 39, 16, 2, 16, 25, 14, 10, 12, 13, 31, 25, 9, 12, 20, 31, 38, 2, 28, 0, 
    84, 17, 28, 53, 24, 9, 11, 32, 30, 3, 21, 21, 29, 35, 24, 11, 21, 25, 14, 20, 28, 28, 38, 29, 15, 17, 22, 17, 25, 30, 35, 0, 
    88, 23, 30, 33, 17, 15, 24, 34, 14, 18, 34, 13, 16, 27, 25, 24, 27, 25, 18, 28, 38, 37, 40, 35, 22, 21, 22, 9, 15, 44, 50, 0, 
    91, 41, 32, 13, 9, 28, 40, 41, 19, 19, 30, 18, 26, 24, 17, 31, 35, 31, 24, 32, 42, 35, 35, 37, 21, 19, 23, 16, 20, 38, 35, 0, 
    75, 58, 50, 33, 33, 50, 53, 51, 42, 50, 46, 40, 45, 40, 34, 49, 51, 50, 46, 47, 53, 50, 51, 54, 42, 40, 45, 41, 41, 49, 46, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    115, 62, 36, 35, 63, 82, 73, 67, 73, 76, 77, 83, 86, 83, 72, 75, 80, 77, 81, 79, 76, 69, 62, 61, 66, 67, 63, 61, 62, 53, 51, 50, 
    115, 58, 56, 60, 84, 92, 85, 87, 88, 80, 76, 76, 74, 78, 74, 62, 72, 70, 80, 92, 88, 77, 63, 49, 31, 27, 34, 53, 72, 70, 57, 54, 
    118, 82, 89, 93, 88, 82, 80, 79, 85, 83, 74, 73, 71, 66, 70, 67, 63, 72, 60, 77, 91, 85, 77, 76, 64, 51, 48, 55, 62, 67, 58, 45, 
    118, 96, 118, 113, 93, 85, 82, 79, 82, 81, 83, 81, 83, 82, 85, 88, 72, 51, 33, 27, 55, 59, 54, 65, 74, 77, 70, 64, 55, 51, 59, 55, 
    110, 95, 106, 105, 87, 82, 90, 94, 88, 85, 86, 95, 87, 79, 79, 92, 98, 70, 38, 8, 12, 34, 29, 35, 50, 61, 76, 74, 61, 51, 52, 54, 
    120, 103, 95, 101, 89, 87, 88, 89, 90, 85, 86, 88, 83, 73, 66, 77, 97, 92, 68, 42, 25, 55, 65, 61, 68, 72, 81, 84, 75, 67, 62, 57, 
    140, 90, 104, 100, 104, 96, 90, 92, 87, 89, 97, 91, 82, 86, 85, 80, 86, 93, 87, 78, 67, 69, 79, 70, 73, 78, 66, 68, 71, 67, 69, 61, 
    121, 89, 89, 97, 98, 91, 94, 103, 104, 95, 93, 95, 86, 85, 91, 83, 86, 100, 107, 89, 71, 56, 55, 50, 68, 68, 55, 48, 55, 62, 65, 60, 
    120, 110, 90, 90, 84, 83, 92, 93, 101, 98, 91, 86, 80, 75, 63, 48, 49, 74, 99, 100, 86, 79, 84, 76, 78, 77, 74, 76, 73, 70, 64, 61, 
    162, 131, 103, 92, 102, 98, 87, 83, 81, 105, 113, 97, 64, 58, 64, 54, 40, 56, 78, 87, 86, 91, 105, 116, 93, 92, 84, 88, 87, 77, 68, 57, 
    155, 134, 95, 81, 89, 93, 91, 88, 95, 118, 121, 85, 42, 42, 71, 117, 124, 84, 75, 72, 64, 81, 100, 103, 99, 92, 84, 78, 76, 74, 72, 65, 
    95, 101, 90, 59, 41, 52, 71, 84, 100, 106, 95, 82, 78, 78, 81, 92, 140, 121, 76, 75, 65, 72, 79, 72, 77, 92, 98, 88, 77, 75, 73, 68, 
    47, 72, 126, 106, 86, 83, 91, 81, 79, 80, 77, 84, 108, 110, 68, 13, 0, 26, 26, 31, 62, 66, 69, 70, 68, 80, 84, 77, 74, 75, 78, 72, 
    48, 59, 110, 121, 94, 85, 91, 95, 66, 55, 64, 73, 80, 92, 71, 24, 0, 10, 19, 30, 38, 46, 52, 50, 58, 68, 68, 53, 52, 74, 75, 70, 
    80, 51, 81, 96, 86, 79, 84, 103, 92, 67, 66, 69, 52, 49, 65, 57, 63, 70, 74, 63, 43, 38, 48, 60, 76, 80, 71, 49, 26, 55, 80, 67, 
    86, 36, 35, 71, 93, 82, 79, 100, 110, 84, 103, 111, 91, 72, 88, 105, 98, 93, 98, 98, 87, 79, 85, 100, 97, 99, 86, 64, 40, 36, 76, 80, 
    87, 40, 40, 50, 62, 65, 64, 83, 119, 107, 115, 128, 102, 85, 115, 130, 148, 126, 122, 148, 161, 157, 129, 100, 89, 85, 93, 74, 55, 37, 65, 83, 
    88, 55, 74, 86, 71, 58, 65, 82, 142, 140, 67, 70, 70, 81, 97, 88, 93, 135, 139, 157, 162, 137, 95, 59, 53, 62, 76, 74, 38, 32, 57, 81, 
    94, 53, 61, 91, 84, 64, 58, 66, 123, 192, 118, 76, 98, 92, 63, 25, 0, 37, 92, 99, 82, 54, 40, 34, 47, 72, 82, 77, 44, 16, 40, 75, 
    85, 32, 38, 65, 79, 80, 88, 86, 97, 180, 226, 184, 152, 118, 110, 114, 88, 52, 54, 72, 71, 55, 57, 55, 55, 73, 97, 91, 60, 28, 24, 58, 
    85, 41, 58, 84, 95, 93, 107, 101, 55, 68, 140, 190, 180, 142, 117, 134, 158, 137, 94, 78, 99, 108, 108, 90, 51, 50, 84, 114, 95, 61, 38, 57, 
    96, 58, 52, 70, 94, 95, 90, 59, 14, 3, 8, 39, 66, 77, 62, 86, 122, 146, 139, 106, 94, 97, 109, 119, 101, 78, 85, 117, 131, 84, 45, 53, 
    112, 70, 49, 40, 77, 99, 57, 13, 12, 30, 19, 0, 0, 1, 34, 60, 84, 100, 105, 102, 89, 85, 88, 106, 123, 105, 90, 108, 140, 111, 41, 24, 
    106, 62, 58, 50, 60, 94, 83, 38, 23, 34, 30, 22, 38, 35, 42, 46, 32, 26, 38, 53, 67, 74, 79, 79, 81, 88, 85, 103, 134, 145, 82, 11, 
    87, 43, 50, 61, 55, 64, 111, 134, 76, 35, 49, 43, 52, 44, 26, 22, 17, 13, 20, 27, 33, 42, 53, 53, 53, 79, 91, 84, 92, 104, 131, 82, 
    96, 58, 70, 65, 43, 38, 66, 121, 138, 86, 106, 109, 64, 42, 28, 27, 35, 27, 16, 10, 9, 6, 8, 9, 18, 41, 54, 42, 30, 38, 72, 108, 
    90, 60, 74, 82, 73, 64, 64, 65, 93, 103, 58, 53, 52, 58, 54, 46, 38, 37, 25, 19, 19, 17, 11, 7, 9, 12, 17, 26, 52, 71, 44, 41, 
    101, 55, 48, 56, 72, 68, 63, 54, 53, 68, 60, 31, 31, 53, 60, 51, 37, 40, 47, 47, 42, 36, 34, 35, 32, 32, 32, 44, 70, 74, 54, 24, 
    101, 60, 29, 27, 41, 47, 35, 33, 35, 23, 29, 42, 53, 63, 73, 75, 61, 61, 62, 57, 55, 49, 50, 52, 45, 44, 48, 53, 49, 44, 41, 46, 
    79, 33, 31, 42, 58, 70, 58, 51, 57, 65, 58, 58, 61, 67, 83, 96, 90, 70, 54, 47, 52, 58, 58, 59, 55, 50, 56, 50, 42, 41, 54, 61, 
    156, 143, 150, 154, 154, 157, 164, 157, 156, 158, 173, 167, 157, 145, 136, 138, 148, 141, 131, 125, 129, 138, 138, 143, 144, 140, 136, 135, 124, 120, 130, 125, 
    
    -- channel=84
    0, 17, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 72, 26, 13, 22, 41, 38, 40, 42, 39, 37, 25, 27, 24, 17, 7, 12, 28, 13, 0, 0, 7, 11, 9, 5, 3, 5, 8, 25, 35, 14, 5, 
    0, 72, 40, 49, 52, 42, 31, 47, 48, 42, 45, 35, 33, 29, 26, 18, 19, 17, 4, 0, 0, 0, 8, 15, 17, 14, 17, 21, 27, 27, 16, 17, 
    0, 70, 55, 66, 63, 40, 29, 49, 46, 45, 51, 43, 42, 34, 25, 26, 24, 23, 11, 0, 0, 0, 4, 14, 17, 24, 34, 34, 29, 19, 16, 22, 
    0, 74, 67, 58, 67, 44, 32, 50, 46, 48, 55, 47, 46, 43, 29, 27, 28, 30, 30, 13, 0, 0, 16, 23, 17, 28, 35, 36, 34, 21, 20, 31, 
    0, 88, 62, 48, 70, 49, 43, 53, 49, 56, 59, 54, 49, 51, 41, 23, 22, 34, 42, 44, 18, 9, 28, 30, 16, 22, 27, 26, 28, 28, 28, 35, 
    0, 94, 46, 47, 68, 56, 52, 52, 54, 63, 66, 57, 50, 59, 53, 32, 21, 37, 47, 58, 40, 23, 29, 34, 20, 22, 19, 11, 19, 31, 33, 37, 
    0, 84, 44, 53, 63, 58, 55, 53, 55, 67, 68, 56, 52, 64, 56, 41, 29, 37, 45, 56, 58, 43, 31, 41, 21, 18, 17, 10, 21, 30, 34, 38, 
    0, 75, 44, 56, 62, 61, 55, 50, 54, 66, 65, 59, 64, 70, 61, 52, 50, 47, 43, 46, 58, 51, 32, 50, 30, 9, 15, 15, 23, 30, 34, 35, 
    0, 58, 39, 59, 67, 63, 60, 53, 55, 63, 59, 53, 67, 80, 73, 73, 82, 65, 39, 36, 53, 52, 43, 62, 35, 0, 9, 18, 22, 28, 34, 36, 
    0, 17, 18, 61, 60, 55, 62, 62, 58, 55, 43, 51, 81, 107, 94, 87, 107, 87, 45, 34, 57, 55, 45, 54, 18, 0, 9, 13, 15, 22, 31, 34, 
    0, 0, 7, 82, 67, 68, 80, 72, 73, 60, 36, 49, 98, 132, 99, 80, 89, 68, 45, 37, 61, 65, 54, 41, 3, 0, 1, 2, 5, 15, 28, 34, 
    0, 0, 9, 84, 66, 84, 94, 87, 86, 61, 31, 58, 113, 140, 109, 85, 78, 58, 60, 53, 73, 78, 57, 29, 0, 0, 0, 0, 1, 13, 24, 27, 
    0, 0, 16, 59, 75, 112, 110, 98, 96, 68, 53, 88, 119, 112, 90, 105, 87, 64, 90, 77, 96, 90, 56, 29, 0, 0, 0, 0, 3, 11, 20, 19, 
    0, 4, 14, 32, 78, 122, 109, 98, 94, 77, 84, 125, 128, 98, 76, 112, 123, 102, 117, 114, 119, 103, 69, 31, 0, 0, 0, 1, 21, 20, 13, 12, 
    0, 44, 23, 13, 72, 121, 108, 84, 79, 91, 115, 144, 133, 101, 77, 107, 138, 131, 130, 131, 138, 119, 83, 27, 0, 0, 0, 17, 48, 39, 10, 4, 
    0, 61, 35, 27, 79, 123, 119, 85, 57, 90, 132, 122, 117, 124, 93, 97, 116, 117, 117, 114, 116, 107, 71, 10, 0, 0, 0, 21, 72, 66, 14, 0, 
    0, 65, 52, 38, 82, 128, 129, 87, 37, 79, 142, 100, 105, 137, 95, 61, 79, 76, 84, 72, 68, 71, 34, 0, 0, 0, 0, 19, 83, 95, 30, 0, 
    0, 68, 50, 34, 86, 137, 149, 108, 32, 51, 133, 89, 95, 139, 95, 67, 87, 68, 62, 40, 29, 27, 0, 0, 0, 0, 0, 16, 87, 122, 57, 0, 
    0, 82, 55, 31, 83, 144, 158, 127, 30, 0, 69, 74, 101, 132, 74, 63, 110, 80, 53, 14, 0, 0, 0, 0, 0, 0, 0, 11, 98, 146, 89, 0, 
    0, 90, 65, 32, 71, 135, 149, 130, 43, 0, 0, 34, 60, 79, 40, 41, 108, 91, 41, 0, 0, 0, 0, 0, 0, 0, 0, 5, 93, 162, 116, 0, 
    0, 96, 79, 45, 66, 119, 132, 112, 45, 0, 0, 0, 8, 28, 16, 13, 58, 55, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 150, 128, 11, 
    0, 103, 83, 53, 61, 100, 119, 91, 39, 5, 0, 0, 0, 8, 10, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 116, 127, 31, 
    0, 91, 75, 68, 68, 79, 99, 93, 61, 40, 24, 20, 16, 14, 16, 20, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 113, 56, 
    0, 77, 66, 82, 76, 59, 68, 86, 93, 73, 40, 53, 52, 44, 43, 44, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 77, 70, 
    0, 69, 63, 84, 91, 67, 53, 72, 88, 81, 45, 55, 55, 55, 66, 54, 33, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 55, 
    0, 70, 76, 74, 81, 90, 66, 44, 57, 83, 66, 55, 50, 51, 77, 70, 49, 30, 19, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 18, 31, 23, 
    0, 79, 81, 59, 71, 98, 83, 42, 29, 80, 62, 40, 53, 55, 85, 86, 62, 42, 42, 41, 30, 22, 10, 11, 26, 21, 11, 4, 3, 35, 41, 13, 
    0, 75, 81, 56, 76, 96, 81, 62, 51, 72, 68, 57, 64, 57, 78, 83, 70, 49, 52, 54, 42, 37, 32, 39, 53, 48, 37, 34, 28, 30, 41, 39, 
    0, 73, 80, 70, 88, 93, 80, 67, 72, 76, 63, 78, 82, 59, 64, 66, 61, 53, 54, 53, 43, 43, 46, 53, 65, 66, 57, 55, 45, 28, 30, 57, 
    0, 63, 78, 84, 91, 76, 68, 70, 73, 75, 62, 75, 74, 61, 59, 47, 44, 49, 52, 51, 44, 50, 57, 59, 72, 75, 67, 65, 57, 44, 49, 66, 
    0, 0, 11, 24, 25, 4, 0, 6, 10, 4, 0, 9, 7, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 3, 1, 0, 0, 0, 21, 
    
    -- channel=85
    48, 58, 61, 47, 48, 60, 62, 64, 61, 63, 65, 59, 58, 58, 49, 49, 49, 45, 37, 26, 24, 27, 25, 25, 20, 28, 32, 33, 27, 30, 21, 0, 
    122, 103, 98, 119, 128, 113, 111, 114, 122, 113, 109, 107, 99, 87, 91, 98, 89, 67, 52, 56, 55, 53, 50, 50, 47, 44, 47, 67, 58, 51, 47, 0, 
    126, 138, 140, 151, 130, 118, 122, 119, 126, 117, 115, 111, 105, 92, 86, 93, 80, 72, 50, 48, 52, 54, 55, 52, 54, 58, 67, 72, 58, 56, 59, 0, 
    140, 159, 164, 156, 131, 128, 127, 126, 130, 124, 128, 118, 110, 106, 99, 101, 98, 65, 47, 35, 42, 55, 56, 55, 67, 75, 75, 69, 62, 55, 58, 3, 
    155, 157, 160, 156, 132, 131, 135, 137, 142, 137, 133, 135, 127, 114, 110, 105, 107, 85, 55, 46, 43, 55, 52, 52, 61, 64, 71, 66, 62, 65, 66, 3, 
    158, 143, 161, 150, 139, 143, 140, 143, 148, 144, 145, 138, 133, 117, 112, 115, 112, 114, 89, 72, 68, 67, 65, 60, 62, 66, 64, 68, 68, 72, 77, 4, 
    152, 141, 163, 150, 153, 147, 146, 151, 149, 150, 147, 144, 134, 124, 115, 124, 125, 125, 113, 98, 103, 99, 87, 74, 61, 59, 60, 67, 71, 73, 78, 5, 
    136, 149, 141, 158, 156, 148, 147, 152, 160, 156, 144, 150, 142, 127, 115, 122, 125, 127, 132, 124, 110, 110, 86, 69, 60, 52, 57, 58, 63, 72, 75, 5, 
    123, 136, 151, 158, 148, 149, 149, 154, 159, 160, 149, 140, 132, 129, 116, 117, 112, 114, 118, 126, 105, 117, 108, 85, 65, 57, 57, 68, 74, 74, 75, 5, 
    120, 139, 158, 144, 150, 157, 152, 159, 153, 152, 151, 151, 139, 128, 124, 123, 110, 104, 105, 117, 113, 130, 118, 89, 72, 71, 70, 74, 79, 76, 78, 1, 
    95, 140, 142, 142, 157, 165, 159, 154, 159, 164, 170, 168, 152, 127, 134, 147, 136, 109, 108, 112, 105, 118, 109, 73, 76, 66, 70, 67, 70, 71, 76, 5, 
    59, 120, 141, 147, 151, 146, 155, 164, 157, 159, 168, 177, 171, 161, 163, 138, 133, 131, 115, 115, 112, 102, 84, 50, 47, 58, 64, 65, 70, 73, 73, 2, 
    44, 111, 139, 155, 169, 175, 180, 167, 140, 153, 179, 202, 194, 173, 154, 130, 101, 96, 109, 112, 111, 90, 55, 38, 46, 57, 57, 60, 66, 66, 70, 2, 
    55, 110, 136, 182, 189, 184, 174, 168, 147, 156, 183, 204, 182, 164, 141, 108, 123, 110, 128, 142, 107, 91, 54, 32, 35, 44, 56, 59, 60, 63, 61, 0, 
    67, 99, 132, 167, 183, 179, 172, 160, 163, 182, 198, 196, 168, 151, 161, 141, 162, 170, 172, 163, 136, 95, 50, 36, 32, 48, 69, 70, 60, 50, 57, 0, 
    79, 76, 99, 154, 181, 173, 169, 166, 179, 207, 206, 185, 169, 172, 188, 191, 193, 193, 193, 181, 151, 101, 62, 48, 39, 61, 84, 85, 75, 49, 49, 0, 
    79, 69, 105, 151, 171, 171, 150, 157, 190, 212, 193, 206, 189, 175, 180, 186, 197, 193, 186, 176, 158, 116, 76, 42, 34, 56, 99, 112, 82, 60, 45, 0, 
    91, 76, 102, 162, 180, 169, 141, 151, 190, 208, 185, 187, 162, 145, 160, 172, 158, 165, 161, 154, 136, 80, 46, 19, 13, 56, 100, 134, 93, 55, 44, 0, 
    95, 86, 114, 160, 185, 187, 143, 123, 164, 177, 171, 165, 168, 144, 139, 125, 116, 94, 101, 91, 62, 24, 6, 0, 12, 57, 109, 143, 124, 53, 36, 0, 
    98, 82, 107, 149, 183, 188, 148, 95, 129, 129, 172, 199, 162, 108, 119, 117, 134, 87, 43, 39, 24, 12, 12, 13, 27, 56, 121, 158, 147, 76, 36, 0, 
    101, 77, 102, 162, 194, 188, 151, 64, 79, 99, 105, 149, 135, 103, 130, 133, 114, 87, 42, 23, 23, 38, 45, 30, 30, 48, 105, 168, 175, 94, 45, 0, 
    110, 96, 106, 147, 175, 177, 138, 43, 24, 47, 53, 63, 64, 60, 93, 102, 72, 51, 33, 35, 29, 30, 36, 27, 34, 51, 105, 160, 187, 115, 57, 0, 
    115, 96, 102, 125, 152, 156, 116, 58, 24, 14, 34, 37, 35, 27, 46, 48, 48, 36, 12, 18, 18, 14, 24, 26, 34, 58, 96, 138, 165, 129, 61, 0, 
    106, 96, 99, 116, 132, 140, 127, 93, 71, 56, 42, 31, 46, 55, 57, 46, 16, 1, 0, 0, 0, 0, 10, 22, 25, 47, 56, 101, 140, 127, 78, 3, 
    97, 96, 94, 105, 126, 129, 137, 153, 126, 91, 66, 60, 58, 77, 62, 27, 4, 0, 0, 0, 0, 0, 0, 6, 22, 41, 42, 69, 108, 109, 86, 26, 
    90, 102, 117, 106, 104, 127, 138, 144, 132, 116, 99, 103, 84, 71, 57, 45, 30, 23, 13, 10, 0, 0, 0, 1, 21, 39, 31, 41, 69, 92, 64, 14, 
    100, 102, 101, 111, 108, 112, 126, 134, 118, 139, 105, 76, 84, 86, 83, 74, 52, 47, 36, 27, 19, 16, 24, 25, 35, 42, 24, 33, 59, 75, 91, 0, 
    102, 90, 91, 113, 114, 103, 88, 122, 111, 84, 106, 81, 88, 100, 92, 77, 70, 61, 56, 54, 55, 48, 55, 59, 57, 55, 53, 67, 83, 60, 83, 2, 
    96, 90, 89, 102, 98, 100, 80, 87, 105, 81, 76, 83, 104, 106, 96, 79, 78, 80, 75, 70, 67, 68, 82, 86, 80, 75, 79, 80, 82, 65, 62, 4, 
    100, 77, 87, 101, 100, 88, 88, 97, 91, 100, 108, 96, 98, 101, 99, 88, 91, 90, 78, 67, 68, 83, 95, 96, 93, 89, 87, 77, 67, 72, 95, 13, 
    97, 100, 112, 110, 101, 95, 105, 113, 104, 106, 122, 111, 105, 98, 90, 84, 83, 84, 73, 74, 83, 89, 97, 104, 97, 96, 90, 83, 78, 87, 98, 8, 
    75, 119, 131, 117, 104, 96, 89, 100, 107, 117, 108, 102, 97, 91, 87, 86, 77, 83, 86, 91, 96, 98, 106, 112, 108, 105, 100, 92, 96, 105, 104, 27, 
    
    -- channel=86
    79, 62, 46, 37, 50, 54, 48, 48, 48, 56, 47, 50, 52, 56, 49, 40, 53, 54, 47, 37, 42, 43, 45, 41, 41, 40, 38, 35, 55, 46, 42, 73, 
    51, 53, 56, 41, 42, 39, 38, 48, 42, 52, 47, 47, 46, 51, 51, 37, 46, 49, 42, 28, 31, 36, 40, 44, 36, 34, 31, 26, 39, 43, 36, 80, 
    36, 45, 47, 49, 53, 37, 38, 42, 40, 53, 48, 50, 54, 48, 49, 49, 47, 60, 46, 26, 27, 32, 36, 41, 40, 41, 35, 35, 34, 36, 37, 84, 
    23, 41, 35, 53, 56, 40, 42, 43, 41, 48, 48, 49, 55, 53, 45, 52, 53, 63, 63, 31, 23, 30, 33, 28, 29, 36, 37, 42, 39, 30, 36, 90, 
    22, 43, 24, 50, 54, 41, 42, 44, 43, 44, 47, 48, 51, 57, 45, 38, 59, 63, 77, 54, 27, 37, 45, 30, 26, 28, 33, 39, 44, 35, 31, 93, 
    32, 46, 22, 48, 50, 42, 42, 41, 43, 44, 50, 46, 52, 60, 53, 31, 47, 56, 68, 69, 39, 37, 53, 38, 33, 33, 31, 33, 39, 38, 32, 96, 
    43, 32, 31, 40, 45, 44, 42, 40, 44, 42, 53, 47, 48, 53, 60, 41, 39, 45, 51, 59, 52, 28, 51, 43, 32, 41, 30, 28, 34, 33, 32, 96, 
    35, 33, 32, 32, 43, 42, 40, 38, 46, 43, 46, 47, 47, 44, 52, 44, 40, 37, 43, 45, 60, 34, 56, 53, 35, 40, 36, 32, 32, 33, 32, 95, 
    24, 41, 27, 36, 42, 41, 43, 33, 42, 46, 45, 43, 46, 44, 43, 47, 44, 32, 33, 39, 55, 37, 59, 64, 38, 36, 38, 37, 32, 37, 30, 96, 
    24, 23, 31, 38, 37, 43, 46, 40, 40, 43, 46, 43, 41, 44, 35, 52, 55, 41, 26, 32, 44, 33, 49, 68, 33, 35, 33, 32, 31, 36, 33, 96, 
    9, 3, 40, 34, 25, 41, 45, 45, 45, 38, 38, 38, 46, 43, 19, 39, 62, 53, 29, 32, 38, 36, 46, 52, 30, 34, 34, 32, 29, 32, 33, 95, 
    0, 0, 44, 36, 28, 38, 41, 41, 47, 34, 30, 32, 51, 48, 27, 18, 31, 53, 29, 30, 41, 39, 53, 44, 27, 26, 36, 36, 29, 33, 31, 92, 
    0, 0, 34, 32, 39, 41, 42, 47, 48, 30, 31, 29, 40, 40, 46, 40, 3, 42, 34, 22, 48, 44, 55, 48, 27, 23, 33, 36, 30, 33, 31, 89, 
    22, 0, 5, 18, 34, 36, 35, 49, 45, 25, 31, 36, 34, 31, 41, 65, 26, 38, 38, 33, 48, 48, 53, 42, 32, 26, 31, 39, 32, 33, 30, 85, 
    39, 19, 0, 8, 31, 41, 31, 33, 41, 26, 31, 45, 48, 28, 26, 42, 34, 32, 34, 46, 48, 57, 54, 40, 36, 23, 26, 48, 42, 32, 31, 84, 
    41, 40, 2, 0, 28, 41, 40, 15, 24, 27, 33, 36, 57, 36, 19, 28, 27, 25, 25, 36, 49, 66, 50, 42, 31, 15, 18, 43, 64, 35, 26, 83, 
    35, 49, 16, 0, 22, 37, 54, 13, 3, 37, 29, 12, 45, 43, 20, 21, 23, 29, 20, 25, 40, 61, 48, 40, 27, 6, 11, 27, 69, 54, 21, 77, 
    30, 45, 14, 6, 24, 33, 62, 25, 0, 53, 29, 6, 39, 50, 18, 27, 11, 30, 23, 16, 30, 44, 45, 42, 28, 8, 2, 22, 56, 73, 25, 68, 
    30, 45, 4, 0, 23, 33, 61, 55, 0, 34, 47, 14, 40, 55, 15, 59, 32, 28, 34, 22, 39, 39, 42, 48, 25, 15, 0, 16, 52, 86, 32, 61, 
    31, 48, 15, 0, 14, 30, 57, 92, 0, 0, 34, 19, 38, 49, 9, 51, 73, 52, 47, 31, 44, 39, 37, 51, 26, 9, 0, 8, 46, 97, 47, 58, 
    30, 49, 26, 1, 13, 25, 47, 96, 25, 0, 0, 8, 29, 42, 0, 4, 51, 63, 57, 27, 29, 30, 26, 50, 36, 10, 0, 0, 31, 94, 64, 60, 
    28, 48, 25, 4, 13, 29, 51, 76, 54, 32, 9, 6, 12, 32, 12, 11, 25, 38, 56, 35, 26, 27, 14, 34, 43, 23, 0, 0, 20, 81, 75, 64, 
    28, 42, 33, 16, 9, 33, 57, 63, 60, 55, 48, 38, 29, 27, 31, 38, 34, 28, 38, 40, 34, 35, 17, 14, 30, 24, 19, 0, 3, 66, 84, 67, 
    29, 28, 34, 36, 14, 21, 50, 65, 66, 39, 49, 45, 47, 35, 40, 50, 52, 40, 36, 34, 34, 35, 28, 21, 15, 19, 35, 1, 0, 40, 88, 84, 
    30, 29, 26, 40, 34, 10, 21, 49, 73, 37, 48, 36, 32, 37, 43, 54, 63, 50, 45, 37, 36, 35, 32, 36, 17, 19, 40, 14, 0, 5, 57, 112, 
    27, 34, 27, 29, 46, 30, 7, 4, 68, 49, 39, 49, 28, 41, 53, 53, 56, 48, 47, 43, 47, 45, 34, 39, 29, 23, 40, 28, 18, 22, 13, 103, 
    20, 35, 28, 22, 43, 47, 39, 0, 32, 60, 26, 41, 25, 33, 49, 55, 45, 45, 49, 49, 51, 50, 40, 44, 45, 37, 40, 33, 23, 56, 16, 80, 
    21, 43, 25, 13, 36, 41, 49, 26, 20, 47, 37, 44, 23, 24, 38, 55, 41, 39, 47, 44, 44, 44, 38, 44, 47, 46, 43, 36, 24, 39, 38, 95, 
    18, 46, 29, 23, 32, 40, 40, 35, 41, 31, 32, 45, 32, 27, 32, 47, 43, 37, 41, 34, 37, 38, 33, 38, 44, 42, 42, 45, 36, 26, 31, 110, 
    17, 38, 33, 36, 32, 40, 40, 32, 43, 39, 32, 40, 37, 33, 29, 34, 43, 39, 40, 32, 31, 37, 32, 33, 45, 38, 40, 47, 43, 31, 25, 107, 
    22, 33, 33, 37, 31, 26, 31, 31, 36, 27, 31, 36, 39, 42, 36, 25, 36, 38, 42, 36, 29, 37, 34, 31, 43, 39, 37, 46, 46, 32, 29, 104, 
    0, 1, 6, 16, 17, 4, 1, 5, 14, 5, 4, 8, 12, 22, 25, 11, 8, 11, 15, 13, 7, 9, 8, 5, 10, 14, 9, 12, 15, 10, 7, 69, 
    
    -- channel=87
    122, 0, 0, 20, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 9, 19, 8, 4, 3, 12, 14, 22, 24, 15, 0, 9, 0, 
    174, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 30, 17, 10, 6, 9, 14, 19, 21, 13, 0, 5, 0, 
    183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 37, 26, 15, 10, 5, 11, 7, 4, 0, 1, 13, 0, 
    184, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 35, 17, 10, 17, 15, 0, 0, 0, 2, 17, 0, 
    189, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 37, 9, 0, 16, 13, 0, 0, 0, 0, 14, 0, 
    192, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 6, 4, 0, 3, 2, 0, 5, 0, 
    192, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 14, 3, 4, 0, 
    193, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 14, 13, 5, 5, 0, 
    180, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 8, 5, 4, 1, 0, 
    165, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 11, 6, 7, 10, 1, 0, 
    143, 18, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 7, 0, 0, 0, 0, 0, 37, 11, 5, 12, 13, 6, 0, 
    108, 79, 81, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 1, 39, 17, 8, 14, 17, 7, 0, 
    90, 108, 78, 0, 0, 0, 0, 0, 0, 0, 10, 12, 0, 0, 0, 0, 0, 24, 0, 15, 1, 0, 0, 0, 13, 39, 28, 15, 14, 16, 6, 0, 
    104, 74, 53, 11, 17, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 17, 34, 34, 18, 8, 13, 5, 0, 
    123, 19, 28, 55, 28, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 16, 30, 45, 27, 0, 0, 10, 0, 
    143, 0, 6, 69, 33, 0, 0, 0, 10, 9, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 13, 37, 62, 38, 0, 0, 10, 0, 
    147, 0, 0, 54, 31, 0, 0, 0, 36, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 52, 82, 45, 0, 0, 0, 9, 
    151, 0, 0, 46, 25, 0, 0, 0, 37, 50, 0, 0, 16, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 12, 28, 62, 87, 55, 0, 0, 0, 15, 
    153, 0, 0, 56, 35, 0, 0, 0, 2, 99, 0, 0, 10, 0, 0, 23, 0, 0, 0, 0, 6, 0, 15, 22, 21, 60, 74, 68, 6, 0, 0, 15, 
    160, 0, 0, 52, 42, 0, 0, 0, 0, 107, 32, 0, 0, 0, 0, 43, 0, 0, 0, 0, 28, 13, 29, 18, 1, 54, 75, 79, 21, 0, 0, 2, 
    166, 0, 0, 33, 41, 0, 0, 0, 0, 78, 78, 31, 16, 0, 0, 48, 0, 0, 0, 0, 35, 26, 38, 27, 0, 40, 71, 86, 36, 0, 0, 0, 
    172, 0, 0, 19, 38, 0, 0, 0, 0, 46, 46, 39, 41, 25, 23, 40, 0, 0, 0, 0, 38, 33, 37, 46, 16, 28, 52, 80, 57, 0, 0, 0, 
    174, 0, 0, 7, 24, 1, 0, 0, 0, 2, 1, 24, 33, 30, 18, 5, 0, 0, 24, 23, 40, 36, 34, 55, 46, 37, 45, 55, 73, 0, 0, 0, 
    165, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 2, 5, 0, 3, 0, 0, 7, 36, 36, 40, 38, 39, 56, 62, 59, 43, 21, 68, 38, 0, 0, 
    161, 0, 5, 0, 0, 0, 18, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 21, 26, 37, 37, 42, 54, 53, 67, 37, 3, 56, 58, 5, 0, 
    154, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 6, 14, 27, 24, 34, 48, 37, 51, 33, 15, 62, 44, 10, 0, 
    158, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 22, 0, 0, 0, 0, 2, 0, 5, 5, 17, 32, 17, 17, 16, 18, 43, 24, 0, 0, 
    160, 0, 0, 11, 15, 0, 0, 0, 18, 0, 0, 7, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 0, 0, 3, 10, 10, 0, 0, 
    157, 0, 0, 15, 7, 0, 0, 0, 4, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 15, 0, 
    155, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    110, 12, 4, 0, 0, 5, 18, 13, 5, 0, 12, 2, 0, 0, 0, 2, 17, 8, 8, 2, 7, 11, 2, 7, 5, 0, 0, 3, 0, 3, 10, 0, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 3, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    90, 28, 36, 62, 65, 50, 52, 56, 57, 44, 41, 42, 40, 30, 25, 38, 33, 13, 0, 6, 11, 9, 3, 0, 0, 2, 16, 34, 22, 6, 7, 0, 
    168, 77, 94, 119, 108, 91, 96, 100, 104, 88, 83, 81, 69, 58, 54, 74, 68, 29, 11, 27, 42, 43, 39, 37, 39, 43, 53, 70, 51, 28, 34, 0, 
    188, 122, 144, 127, 95, 96, 111, 108, 110, 99, 91, 89, 78, 68, 67, 68, 60, 20, 0, 11, 36, 42, 44, 44, 50, 60, 66, 61, 44, 42, 50, 0, 
    204, 143, 150, 122, 93, 104, 121, 114, 116, 113, 105, 100, 86, 72, 75, 81, 68, 34, 0, 2, 34, 46, 42, 43, 61, 69, 65, 54, 41, 47, 58, 0, 
    220, 137, 144, 133, 102, 113, 125, 119, 125, 120, 115, 113, 98, 79, 75, 87, 84, 62, 24, 15, 49, 67, 51, 50, 62, 66, 63, 56, 49, 59, 70, 0, 
    217, 122, 141, 145, 121, 124, 126, 127, 131, 131, 124, 119, 110, 92, 77, 91, 97, 89, 70, 51, 66, 80, 52, 41, 54, 54, 52, 56, 57, 64, 73, 0, 
    198, 113, 143, 152, 129, 127, 131, 136, 139, 139, 129, 120, 114, 103, 84, 96, 108, 107, 99, 82, 70, 80, 58, 39, 46, 37, 38, 55, 63, 66, 73, 0, 
    192, 115, 148, 148, 132, 130, 130, 142, 142, 135, 123, 121, 114, 102, 85, 88, 95, 106, 111, 108, 85, 91, 73, 39, 39, 41, 45, 60, 67, 68, 74, 0, 
    178, 120, 148, 145, 140, 135, 130, 136, 140, 141, 131, 124, 115, 108, 105, 101, 93, 93, 104, 113, 90, 101, 95, 40, 35, 47, 54, 63, 68, 66, 71, 0, 
    153, 123, 145, 147, 145, 141, 137, 141, 144, 140, 130, 127, 124, 125, 141, 137, 105, 84, 95, 111, 101, 112, 98, 29, 28, 53, 56, 56, 64, 69, 72, 0, 
    107, 118, 145, 128, 137, 150, 142, 143, 136, 136, 143, 166, 167, 147, 161, 168, 123, 83, 96, 114, 104, 102, 66, 11, 25, 58, 52, 50, 60, 65, 71, 0, 
    60, 143, 177, 148, 166, 169, 156, 152, 131, 129, 160, 202, 197, 164, 143, 121, 104, 79, 95, 122, 109, 89, 45, 0, 20, 46, 41, 43, 57, 65, 67, 0, 
    49, 157, 173, 157, 183, 185, 170, 151, 120, 136, 186, 221, 200, 158, 145, 111, 116, 115, 116, 141, 115, 72, 19, 0, 18, 39, 40, 42, 51, 56, 58, 0, 
    82, 136, 156, 183, 205, 181, 173, 160, 137, 169, 211, 206, 167, 151, 154, 129, 156, 169, 165, 166, 122, 69, 23, 5, 16, 35, 49, 45, 48, 48, 47, 0, 
    99, 92, 131, 197, 211, 179, 167, 165, 164, 205, 230, 206, 164, 164, 192, 178, 193, 207, 196, 184, 138, 78, 32, 13, 16, 40, 75, 71, 45, 38, 42, 0, 
    124, 58, 107, 196, 205, 172, 150, 164, 198, 234, 228, 201, 166, 166, 209, 216, 214, 209, 212, 202, 156, 84, 26, 3, 8, 48, 100, 107, 54, 24, 38, 0, 
    130, 67, 120, 197, 210, 184, 137, 152, 224, 221, 186, 196, 185, 164, 178, 190, 192, 188, 187, 171, 133, 55, 0, 0, 0, 52, 122, 135, 72, 14, 27, 0, 
    146, 74, 118, 199, 212, 190, 130, 117, 219, 212, 165, 203, 193, 126, 133, 131, 142, 137, 115, 105, 69, 5, 0, 0, 0, 60, 137, 160, 101, 11, 11, 0, 
    149, 69, 115, 200, 225, 211, 145, 68, 169, 206, 154, 199, 187, 115, 143, 147, 118, 93, 53, 40, 15, 0, 0, 0, 3, 61, 140, 187, 140, 20, 0, 0, 
    160, 79, 118, 204, 232, 215, 151, 23, 61, 149, 152, 182, 150, 78, 130, 159, 107, 51, 2, 6, 5, 1, 16, 0, 0, 54, 146, 209, 182, 44, 0, 0, 
    169, 82, 109, 190, 224, 204, 135, 0, 0, 76, 93, 102, 88, 51, 109, 138, 79, 23, 0, 0, 2, 10, 31, 9, 5, 49, 137, 217, 211, 70, 0, 0, 
    182, 95, 104, 164, 201, 179, 104, 0, 0, 39, 45, 42, 43, 38, 81, 96, 41, 0, 0, 0, 0, 0, 10, 14, 12, 46, 111, 197, 215, 94, 0, 0, 
    178, 96, 101, 142, 176, 157, 97, 38, 22, 22, 20, 36, 48, 53, 55, 33, 0, 0, 0, 0, 0, 0, 0, 1, 10, 41, 79, 148, 198, 117, 0, 0, 
    157, 92, 117, 128, 139, 157, 137, 100, 61, 38, 30, 42, 52, 54, 50, 11, 0, 0, 0, 0, 0, 0, 0, 0, 12, 45, 46, 84, 152, 135, 37, 0, 
    153, 101, 124, 117, 109, 132, 156, 156, 97, 81, 88, 68, 63, 71, 55, 14, 0, 0, 0, 0, 0, 0, 0, 0, 4, 39, 18, 30, 91, 116, 76, 0, 
    148, 108, 128, 124, 114, 123, 135, 158, 107, 79, 92, 74, 83, 93, 70, 41, 16, 6, 0, 0, 0, 0, 0, 0, 11, 32, 11, 25, 89, 90, 73, 0, 
    160, 101, 101, 126, 124, 111, 101, 128, 137, 96, 81, 68, 91, 114, 93, 56, 37, 39, 37, 28, 18, 9, 25, 36, 36, 37, 23, 44, 86, 68, 64, 0, 
    165, 89, 85, 128, 129, 91, 69, 103, 108, 74, 83, 88, 105, 123, 102, 69, 59, 67, 60, 51, 45, 43, 61, 68, 56, 49, 52, 61, 72, 51, 64, 0, 
    153, 85, 93, 129, 124, 96, 81, 102, 109, 85, 96, 100, 104, 112, 104, 80, 71, 77, 65, 60, 64, 71, 87, 92, 77, 73, 74, 64, 64, 64, 88, 0, 
    156, 101, 114, 128, 112, 97, 98, 110, 104, 105, 128, 112, 95, 93, 87, 82, 78, 78, 65, 64, 79, 86, 96, 104, 94, 88, 84, 65, 52, 78, 113, 0, 
    161, 124, 131, 109, 80, 88, 103, 115, 98, 100, 114, 103, 93, 83, 68, 71, 77, 78, 71, 77, 94, 97, 102, 113, 103, 91, 92, 82, 77, 96, 110, 0, 
    56, 32, 33, 17, 5, 10, 18, 20, 16, 18, 24, 13, 7, 0, 0, 0, 2, 1, 2, 2, 10, 13, 14, 22, 16, 9, 8, 4, 3, 12, 16, 0, 
    
    -- channel=91
    50, 54, 26, 14, 34, 46, 42, 38, 41, 49, 43, 48, 50, 49, 46, 43, 54, 58, 54, 51, 54, 54, 55, 54, 61, 58, 48, 41, 57, 50, 47, 74, 
    16, 26, 17, 8, 18, 25, 23, 26, 21, 28, 23, 26, 30, 38, 35, 22, 34, 47, 50, 40, 40, 38, 38, 35, 29, 25, 26, 26, 45, 47, 42, 85, 
    9, 12, 14, 17, 26, 18, 17, 24, 16, 26, 23, 23, 23, 26, 28, 25, 36, 51, 53, 44, 42, 41, 41, 42, 33, 28, 26, 30, 42, 42, 34, 83, 
    0, 17, 18, 30, 32, 14, 15, 18, 12, 22, 19, 20, 27, 27, 26, 29, 27, 42, 47, 37, 35, 35, 39, 42, 39, 37, 35, 39, 38, 34, 35, 89, 
    0, 22, 15, 26, 26, 12, 17, 20, 14, 18, 21, 20, 24, 29, 25, 27, 28, 32, 45, 31, 16, 17, 26, 23, 25, 33, 36, 40, 37, 27, 28, 91, 
    0, 33, 8, 19, 20, 11, 16, 17, 14, 15, 18, 17, 19, 25, 22, 14, 27, 30, 40, 33, 11, 18, 38, 33, 32, 34, 38, 40, 39, 33, 28, 93, 
    14, 32, 8, 18, 20, 18, 16, 9, 11, 14, 20, 13, 21, 28, 28, 13, 15, 20, 31, 39, 32, 27, 45, 39, 38, 44, 40, 35, 35, 34, 31, 95, 
    21, 14, 13, 16, 19, 18, 16, 12, 15, 18, 25, 16, 22, 28, 37, 28, 25, 25, 27, 26, 32, 11, 28, 36, 36, 41, 28, 23, 28, 30, 30, 94, 
    10, 22, 15, 12, 13, 13, 16, 14, 19, 16, 12, 11, 23, 23, 22, 20, 24, 24, 26, 22, 36, 17, 31, 44, 38, 36, 33, 31, 30, 33, 30, 95, 
    22, 29, 13, 13, 14, 14, 15, 5, 8, 12, 17, 17, 23, 20, 6, 11, 22, 22, 18, 21, 33, 20, 39, 64, 44, 37, 38, 40, 35, 35, 28, 93, 
    40, 17, 18, 26, 21, 18, 13, 12, 18, 16, 14, 1, 2, 10, 6, 22, 33, 30, 13, 14, 25, 26, 50, 73, 43, 35, 35, 35, 33, 34, 32, 95, 
    25, 0, 9, 2, 0, 0, 8, 13, 26, 15, 3, 0, 13, 21, 14, 43, 61, 53, 23, 18, 24, 32, 53, 56, 42, 40, 44, 39, 32, 32, 32, 96, 
    5, 0, 18, 11, 3, 8, 8, 14, 31, 9, 0, 0, 26, 29, 18, 18, 4, 19, 7, 6, 28, 39, 61, 58, 43, 36, 39, 37, 33, 36, 36, 94, 
    0, 0, 16, 5, 8, 14, 13, 19, 17, 0, 0, 5, 30, 23, 16, 26, 0, 0, 0, 0, 28, 39, 53, 51, 41, 33, 30, 32, 33, 38, 38, 93, 
    19, 21, 3, 0, 4, 13, 11, 20, 12, 0, 0, 5, 9, 0, 0, 19, 2, 4, 4, 12, 24, 34, 48, 46, 47, 35, 20, 24, 30, 38, 37, 89, 
    20, 30, 2, 0, 9, 21, 22, 11, 6, 0, 0, 13, 23, 5, 0, 8, 9, 9, 8, 15, 21, 45, 56, 59, 57, 32, 13, 22, 38, 39, 39, 89, 
    17, 33, 0, 0, 0, 11, 25, 4, 0, 6, 28, 20, 26, 14, 7, 24, 22, 19, 17, 29, 49, 79, 75, 70, 57, 26, 10, 16, 50, 47, 36, 90, 
    6, 33, 15, 0, 0, 10, 40, 19, 0, 28, 18, 0, 9, 35, 27, 35, 33, 43, 44, 53, 72, 91, 73, 59, 43, 14, 0, 3, 41, 61, 38, 85, 
    8, 39, 14, 0, 1, 6, 34, 39, 0, 37, 15, 0, 22, 42, 0, 3, 0, 32, 51, 50, 63, 60, 47, 48, 37, 19, 0, 0, 26, 69, 45, 81, 
    5, 30, 0, 0, 0, 12, 36, 73, 15, 42, 49, 15, 42, 57, 10, 34, 30, 35, 57, 47, 49, 39, 38, 56, 44, 29, 0, 0, 20, 71, 46, 73, 
    1, 33, 16, 0, 0, 21, 47, 100, 42, 13, 53, 58, 67, 64, 21, 43, 74, 70, 67, 52, 59, 54, 45, 57, 38, 20, 0, 0, 16, 76, 59, 73, 
    0, 34, 22, 0, 8, 27, 50, 84, 45, 7, 14, 32, 47, 51, 16, 21, 61, 79, 81, 55, 52, 56, 49, 59, 47, 28, 3, 0, 16, 73, 69, 75, 
    6, 37, 21, 3, 8, 30, 44, 42, 34, 42, 32, 15, 9, 14, 15, 43, 64, 65, 75, 66, 57, 58, 48, 52, 59, 43, 22, 0, 15, 59, 71, 75, 
    16, 32, 19, 13, 13, 23, 23, 18, 35, 42, 42, 35, 30, 23, 36, 52, 56, 48, 49, 54, 57, 63, 51, 42, 41, 30, 39, 18, 15, 48, 67, 72, 
    7, 12, 15, 30, 24, 16, 26, 29, 35, 9, 18, 27, 38, 33, 36, 47, 54, 46, 46, 48, 53, 58, 54, 49, 31, 28, 57, 38, 19, 40, 69, 93, 
    8, 19, 14, 22, 25, 7, 15, 27, 51, 32, 43, 44, 23, 20, 30, 40, 50, 45, 43, 38, 39, 43, 36, 37, 26, 29, 51, 26, 1, 10, 43, 117, 
    2, 25, 28, 21, 30, 29, 23, 3, 36, 38, 26, 38, 19, 22, 34, 39, 44, 40, 36, 34, 40, 40, 25, 25, 25, 22, 30, 20, 13, 39, 19, 92, 
    0, 33, 28, 11, 28, 42, 48, 12, 24, 59, 24, 17, 8, 16, 31, 39, 30, 29, 36, 40, 39, 34, 23, 27, 33, 29, 27, 23, 28, 59, 26, 75, 
    10, 41, 17, 0, 22, 30, 28, 16, 17, 22, 18, 27, 16, 17, 26, 38, 32, 31, 41, 38, 33, 27, 21, 26, 30, 30, 28, 32, 28, 26, 20, 93, 
    0, 24, 10, 11, 21, 28, 23, 17, 31, 18, 7, 23, 23, 26, 32, 39, 38, 33, 34, 27, 27, 25, 21, 22, 29, 26, 29, 37, 33, 21, 17, 102, 
    0, 14, 15, 32, 40, 40, 35, 24, 34, 33, 31, 35, 30, 32, 34, 33, 36, 30, 30, 24, 19, 21, 19, 17, 28, 27, 29, 30, 24, 15, 17, 100, 
    62, 99, 103, 109, 99, 84, 88, 97, 103, 89, 91, 98, 101, 106, 100, 85, 88, 93, 99, 97, 92, 97, 97, 97, 104, 103, 99, 104, 104, 98, 97, 140, 
    
    -- channel=92
    0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 9, 6, 5, 9, 9, 11, 11, 6, 0, 1, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    44, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 
    27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 20, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 17, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 9, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 7, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 8, 13, 3, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 3, 10, 17, 17, 23, 22, 8, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 19, 19, 20, 20, 26, 31, 26, 10, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 20, 20, 22, 26, 30, 35, 18, 0, 4, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 12, 19, 18, 21, 14, 1, 3, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 0, 1, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=93
    22, 117, 74, 79, 107, 120, 117, 113, 119, 111, 104, 92, 95, 80, 68, 72, 70, 63, 31, 15, 14, 21, 15, 6, 0, 4, 15, 44, 50, 46, 21, 0, 
    134, 259, 205, 230, 238, 237, 230, 234, 247, 229, 221, 204, 194, 175, 161, 172, 170, 146, 97, 76, 81, 99, 100, 96, 95, 94, 109, 138, 140, 123, 99, 1, 
    158, 312, 296, 300, 266, 246, 242, 258, 264, 244, 243, 223, 208, 193, 181, 175, 171, 128, 77, 52, 59, 87, 103, 110, 117, 126, 144, 149, 139, 128, 119, 20, 
    174, 343, 339, 315, 274, 251, 253, 272, 274, 268, 266, 250, 231, 208, 195, 196, 187, 148, 83, 50, 50, 79, 100, 116, 134, 153, 166, 155, 136, 126, 128, 30, 
    188, 346, 346, 310, 287, 269, 268, 283, 289, 286, 284, 275, 258, 228, 210, 209, 203, 187, 134, 95, 89, 106, 122, 133, 137, 156, 165, 158, 144, 141, 153, 44, 
    188, 345, 330, 303, 311, 291, 286, 298, 300, 308, 302, 294, 275, 253, 226, 219, 218, 228, 206, 176, 159, 160, 151, 142, 130, 136, 144, 145, 147, 157, 167, 50, 
    177, 345, 302, 317, 322, 303, 303, 309, 315, 328, 316, 302, 286, 275, 244, 235, 236, 254, 253, 238, 208, 203, 169, 152, 131, 117, 119, 124, 143, 163, 173, 54, 
    175, 323, 302, 325, 319, 310, 307, 318, 325, 331, 316, 302, 289, 284, 252, 235, 229, 248, 260, 269, 244, 239, 191, 167, 132, 112, 113, 124, 148, 163, 175, 54, 
    155, 308, 307, 319, 322, 319, 309, 318, 321, 331, 321, 309, 297, 287, 268, 252, 243, 241, 244, 258, 247, 256, 222, 187, 142, 110, 120, 137, 155, 161, 174, 49, 
    125, 292, 288, 320, 334, 327, 323, 323, 328, 330, 319, 312, 308, 305, 309, 303, 287, 248, 226, 237, 251, 271, 249, 193, 142, 103, 128, 141, 151, 160, 173, 51, 
    75, 224, 251, 314, 322, 322, 332, 333, 327, 328, 323, 347, 366, 365, 368, 360, 335, 272, 232, 232, 253, 260, 221, 162, 109, 96, 122, 127, 138, 150, 167, 49, 
    9, 162, 260, 353, 350, 357, 369, 358, 335, 323, 323, 381, 427, 430, 379, 335, 307, 240, 230, 239, 257, 250, 189, 116, 73, 75, 94, 103, 121, 140, 160, 45, 
    0, 143, 268, 360, 368, 403, 404, 374, 336, 322, 341, 428, 472, 447, 377, 313, 298, 249, 266, 284, 277, 247, 153, 81, 51, 60, 78, 92, 110, 127, 144, 33, 
    5, 164, 276, 357, 410, 441, 426, 390, 360, 359, 394, 453, 447, 405, 362, 331, 339, 322, 358, 351, 323, 259, 153, 90, 50, 58, 78, 90, 111, 117, 126, 18, 
    38, 177, 242, 329, 415, 446, 421, 398, 383, 412, 456, 481, 434, 399, 400, 416, 440, 437, 445, 424, 379, 281, 178, 102, 56, 68, 100, 124, 134, 119, 108, 7, 
    79, 181, 214, 304, 401, 434, 398, 388, 403, 464, 497, 498, 435, 408, 427, 468, 504, 493, 491, 474, 424, 315, 203, 95, 51, 70, 124, 186, 176, 137, 99, 0, 
    91, 200, 236, 322, 411, 443, 388, 376, 411, 458, 487, 474, 435, 426, 418, 436, 459, 454, 455, 433, 389, 285, 162, 51, 12, 51, 139, 234, 227, 160, 98, 0, 
    108, 220, 259, 335, 418, 453, 385, 342, 387, 420, 465, 438, 424, 405, 370, 323, 355, 342, 339, 310, 256, 168, 70, 0, 0, 43, 158, 265, 280, 187, 105, 0, 
    113, 226, 261, 333, 436, 487, 420, 306, 336, 356, 411, 414, 412, 386, 351, 299, 322, 274, 222, 173, 109, 59, 11, 0, 2, 51, 170, 292, 333, 231, 119, 0, 
    125, 243, 261, 338, 447, 503, 440, 268, 221, 227, 318, 382, 375, 318, 298, 302, 322, 237, 137, 78, 34, 29, 24, 11, 21, 56, 177, 314, 396, 294, 152, 0, 
    136, 255, 264, 332, 429, 486, 424, 227, 115, 85, 171, 239, 243, 212, 239, 278, 288, 205, 88, 33, 8, 28, 48, 37, 41, 62, 173, 323, 432, 346, 185, 0, 
    152, 283, 280, 317, 395, 437, 367, 197, 71, 27, 73, 102, 111, 114, 155, 186, 190, 126, 34, 2, 0, 0, 17, 21, 34, 66, 152, 298, 411, 368, 211, 0, 
    153, 293, 270, 294, 358, 380, 327, 209, 110, 71, 60, 57, 76, 99, 111, 106, 71, 13, 0, 0, 0, 0, 0, 0, 6, 56, 114, 236, 349, 349, 222, 23, 
    131, 273, 265, 289, 326, 348, 333, 281, 209, 161, 106, 106, 113, 126, 129, 96, 26, 0, 0, 0, 0, 0, 0, 0, 0, 34, 74, 158, 246, 297, 236, 59, 
    122, 261, 273, 295, 295, 306, 333, 351, 295, 246, 190, 195, 182, 175, 161, 115, 46, 0, 0, 0, 0, 0, 0, 0, 0, 9, 40, 82, 126, 211, 225, 80, 
    112, 258, 280, 302, 296, 297, 311, 350, 297, 267, 223, 205, 207, 203, 199, 164, 108, 65, 26, 6, 0, 0, 0, 0, 0, 23, 34, 52, 102, 158, 205, 66, 
    126, 257, 265, 284, 290, 299, 273, 290, 295, 286, 253, 197, 209, 230, 246, 208, 161, 125, 102, 85, 63, 40, 38, 45, 67, 72, 61, 76, 123, 150, 180, 37, 
    130, 252, 252, 267, 288, 293, 241, 236, 240, 244, 223, 195, 235, 258, 271, 236, 200, 175, 164, 157, 136, 119, 126, 139, 146, 130, 121, 130, 155, 158, 163, 28, 
    119, 237, 248, 259, 289, 284, 245, 242, 246, 245, 234, 229, 254, 257, 267, 244, 219, 202, 193, 185, 168, 171, 191, 207, 208, 197, 186, 173, 172, 163, 183, 65, 
    119, 247, 269, 282, 294, 273, 257, 262, 260, 265, 274, 277, 269, 246, 241, 230, 215, 212, 195, 184, 185, 199, 221, 239, 241, 239, 221, 198, 168, 171, 213, 98, 
    119, 266, 299, 294, 270, 247, 248, 269, 266, 271, 267, 269, 257, 231, 213, 200, 192, 199, 191, 195, 207, 221, 242, 258, 261, 256, 242, 223, 209, 217, 240, 103, 
    22, 106, 125, 116, 95, 78, 81, 94, 96, 97, 95, 92, 81, 65, 48, 37, 35, 45, 49, 55, 61, 68, 79, 90, 94, 90, 78, 71, 66, 70, 78, 0, 
    
    -- channel=94
    0, 0, 36, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 119, 89, 86, 99, 102, 96, 90, 104, 108, 107, 105, 102, 88, 88, 95, 85, 72, 55, 52, 47, 48, 53, 56, 68, 66, 52, 49, 44, 40, 35, 1, 
    72, 117, 102, 118, 118, 118, 109, 108, 117, 109, 110, 112, 110, 106, 98, 91, 79, 69, 62, 55, 46, 42, 41, 39, 41, 39, 48, 55, 52, 50, 54, 10, 
    77, 115, 122, 123, 120, 121, 113, 120, 119, 114, 120, 114, 103, 103, 96, 92, 101, 87, 76, 64, 53, 51, 49, 44, 40, 43, 50, 53, 60, 58, 44, 2, 
    85, 126, 139, 134, 128, 119, 114, 118, 121, 125, 118, 117, 120, 112, 108, 108, 99, 93, 71, 67, 67, 63, 62, 68, 64, 57, 57, 58, 57, 58, 57, 9, 
    76, 117, 142, 127, 124, 126, 125, 127, 129, 129, 129, 131, 131, 120, 119, 123, 104, 99, 82, 69, 68, 53, 45, 48, 47, 52, 54, 56, 52, 52, 59, 8, 
    60, 124, 130, 117, 125, 122, 127, 136, 129, 131, 129, 133, 123, 113, 108, 122, 125, 119, 100, 74, 66, 73, 66, 65, 57, 49, 57, 61, 58, 58, 58, 8, 
    72, 139, 111, 126, 130, 128, 127, 126, 129, 132, 126, 127, 125, 116, 102, 107, 109, 106, 107, 108, 99, 121, 99, 81, 69, 59, 68, 65, 61, 63, 62, 12, 
    80, 99, 115, 132, 130, 133, 128, 132, 132, 139, 144, 133, 124, 121, 119, 117, 111, 110, 107, 107, 93, 101, 85, 78, 71, 59, 46, 48, 58, 57, 61, 10, 
    49, 100, 123, 116, 121, 127, 133, 147, 147, 137, 127, 123, 122, 112, 114, 105, 101, 103, 105, 99, 95, 104, 89, 70, 72, 55, 50, 54, 59, 59, 66, 11, 
    48, 121, 99, 101, 118, 127, 135, 129, 129, 132, 145, 152, 142, 108, 92, 84, 88, 92, 103, 101, 97, 95, 83, 71, 77, 58, 66, 69, 66, 61, 58, 8, 
    77, 112, 101, 145, 160, 143, 135, 133, 131, 147, 157, 141, 105, 93, 99, 79, 69, 77, 89, 86, 86, 84, 83, 81, 57, 47, 52, 56, 62, 61, 60, 9, 
    63, 82, 81, 109, 104, 114, 136, 133, 125, 143, 148, 132, 114, 114, 113, 134, 145, 110, 105, 95, 77, 73, 56, 41, 43, 55, 57, 58, 61, 53, 55, 10, 
    39, 71, 97, 123, 122, 132, 130, 125, 134, 141, 131, 132, 134, 127, 104, 84, 107, 87, 97, 105, 81, 77, 57, 44, 43, 49, 60, 60, 59, 55, 55, 9, 
    9, 59, 117, 125, 130, 134, 130, 120, 122, 126, 131, 147, 153, 142, 119, 86, 72, 81, 97, 87, 96, 81, 52, 41, 28, 42, 61, 62, 62, 53, 53, 9, 
    30, 73, 91, 102, 112, 117, 117, 129, 123, 132, 135, 128, 108, 116, 120, 114, 111, 117, 113, 112, 103, 63, 46, 29, 27, 51, 62, 58, 56, 56, 47, 5, 
    37, 58, 86, 111, 122, 131, 118, 130, 138, 125, 112, 128, 121, 123, 120, 110, 119, 118, 116, 102, 72, 50, 49, 35, 41, 53, 63, 71, 50, 55, 51, 2, 
    45, 55, 63, 94, 117, 117, 92, 108, 131, 114, 154, 170, 129, 98, 109, 118, 113, 96, 95, 90, 82, 70, 59, 45, 42, 57, 76, 90, 71, 46, 50, 8, 
    38, 58, 85, 99, 110, 123, 107, 95, 127, 107, 133, 116, 94, 107, 152, 138, 140, 104, 94, 101, 89, 77, 50, 24, 27, 43, 76, 89, 87, 45, 46, 7, 
    46, 81, 105, 111, 115, 114, 93, 60, 107, 77, 66, 97, 99, 87, 77, 42, 65, 79, 63, 63, 49, 35, 14, 4, 21, 39, 78, 99, 88, 53, 53, 12, 
    47, 62, 63, 94, 112, 110, 88, 45, 85, 102, 74, 77, 80, 70, 72, 65, 43, 47, 45, 33, 9, 6, 17, 22, 40, 58, 76, 95, 97, 53, 43, 9, 
    44, 65, 78, 99, 106, 112, 99, 67, 64, 73, 101, 102, 85, 66, 87, 97, 77, 52, 28, 35, 36, 33, 34, 22, 24, 39, 68, 95, 103, 69, 51, 14, 
    43, 72, 83, 90, 104, 108, 102, 88, 40, 6, 35, 64, 76, 69, 55, 41, 59, 62, 34, 26, 28, 28, 36, 31, 17, 35, 62, 97, 101, 86, 58, 19, 
    41, 80, 70, 75, 95, 104, 107, 80, 43, 51, 33, 15, 17, 29, 28, 49, 60, 53, 43, 29, 17, 10, 24, 39, 48, 55, 46, 73, 95, 82, 62, 28, 
    60, 93, 67, 62, 88, 99, 77, 73, 90, 111, 69, 50, 39, 48, 59, 49, 28, 22, 15, 17, 14, 12, 12, 19, 40, 33, 27, 60, 83, 74, 49, 6, 
    42, 67, 78, 88, 88, 104, 105, 103, 79, 65, 39, 52, 74, 64, 52, 41, 29, 24, 19, 25, 24, 22, 28, 28, 33, 35, 46, 68, 85, 96, 68, 0, 
    46, 73, 71, 76, 65, 69, 99, 128, 96, 101, 113, 81, 71, 51, 51, 52, 46, 40, 36, 29, 18, 20, 31, 30, 36, 56, 56, 42, 38, 37, 89, 27, 
    50, 67, 78, 85, 71, 69, 65, 92, 92, 65, 91, 80, 75, 71, 69, 60, 68, 56, 37, 30, 36, 38, 38, 34, 40, 44, 44, 43, 43, 40, 68, 19, 
    31, 61, 83, 82, 77, 88, 84, 76, 86, 99, 70, 48, 67, 77, 74, 62, 60, 54, 46, 52, 54, 52, 58, 60, 61, 57, 58, 60, 76, 87, 57, 0, 
    63, 79, 70, 61, 76, 71, 65, 65, 60, 72, 74, 72, 75, 75, 72, 65, 62, 68, 71, 67, 58, 61, 72, 74, 70, 71, 67, 66, 66, 58, 56, 2, 
    45, 71, 65, 62, 62, 55, 57, 69, 68, 63, 64, 69, 76, 80, 82, 81, 71, 75, 66, 62, 70, 73, 81, 83, 74, 73, 72, 74, 70, 71, 73, 15, 
    0, 0, 5, 15, 26, 32, 17, 8, 13, 34, 30, 23, 13, 9, 17, 26, 17, 7, 0, 1, 3, 2, 6, 7, 4, 6, 7, 0, 0, 0, 1, 0, 
    
    -- channel=95
    35, 54, 69, 65, 58, 66, 74, 77, 73, 72, 78, 78, 75, 76, 74, 71, 59, 52, 56, 60, 61, 62, 61, 63, 60, 62, 64, 62, 51, 57, 57, 42, 
    93, 51, 44, 65, 87, 85, 85, 80, 85, 86, 82, 92, 93, 87, 85, 84, 73, 57, 54, 66, 70, 65, 64, 59, 68, 66, 64, 66, 64, 49, 56, 42, 
    98, 39, 50, 64, 72, 81, 82, 81, 81, 83, 83, 92, 92, 98, 93, 91, 86, 71, 67, 68, 71, 67, 67, 65, 67, 66, 71, 69, 66, 56, 61, 40, 
    100, 37, 58, 53, 64, 77, 81, 83, 80, 85, 84, 89, 89, 97, 101, 96, 98, 78, 66, 66, 71, 69, 70, 72, 71, 73, 70, 66, 67, 67, 62, 41, 
    94, 40, 51, 53, 59, 69, 83, 80, 79, 87, 78, 86, 92, 90, 98, 105, 92, 88, 61, 61, 74, 73, 71, 76, 80, 77, 71, 69, 63, 67, 70, 41, 
    88, 33, 48, 53, 54, 70, 81, 77, 79, 77, 78, 85, 90, 88, 91, 104, 96, 85, 69, 54, 74, 78, 75, 77, 83, 84, 77, 75, 69, 66, 72, 41, 
    82, 35, 42, 53, 57, 67, 77, 78, 73, 74, 76, 87, 92, 90, 86, 94, 102, 84, 76, 62, 70, 88, 78, 72, 81, 77, 81, 80, 74, 69, 67, 42, 
    86, 34, 35, 62, 56, 66, 74, 72, 74, 74, 84, 88, 95, 90, 84, 87, 95, 87, 86, 84, 75, 84, 75, 62, 74, 75, 77, 78, 75, 71, 68, 43, 
    97, 15, 57, 57, 56, 66, 69, 75, 73, 73, 88, 85, 82, 79, 81, 77, 77, 82, 88, 89, 82, 72, 69, 55, 64, 76, 68, 73, 75, 68, 70, 43, 
    86, 40, 61, 50, 60, 64, 68, 73, 75, 74, 78, 75, 68, 55, 60, 53, 53, 66, 88, 88, 83, 67, 63, 40, 56, 69, 71, 71, 69, 68, 69, 42, 
    92, 66, 54, 58, 65, 64, 68, 63, 72, 74, 75, 55, 34, 22, 29, 32, 29, 45, 75, 83, 75, 60, 61, 42, 52, 65, 70, 69, 68, 71, 66, 45, 
    104, 62, 62, 55, 57, 54, 50, 58, 58, 65, 62, 36, 6, 1, 21, 32, 24, 38, 57, 66, 59, 51, 50, 49, 44, 68, 66, 68, 73, 72, 71, 44, 
    90, 73, 71, 45, 44, 49, 47, 46, 49, 55, 50, 24, 4, 0, 3, 31, 41, 27, 34, 46, 37, 40, 44, 38, 55, 69, 65, 67, 73, 71, 72, 48, 
    66, 81, 78, 44, 39, 34, 28, 31, 40, 39, 34, 20, 20, 17, 24, 10, 23, 29, 13, 28, 21, 26, 37, 36, 50, 58, 66, 68, 69, 72, 70, 47, 
    64, 75, 87, 50, 41, 22, 28, 31, 27, 24, 27, 16, 23, 34, 38, 16, 0, 15, 4, 0, 17, 13, 25, 36, 42, 57, 66, 61, 62, 65, 68, 47, 
    82, 74, 70, 67, 45, 23, 26, 40, 24, 15, 18, 12, 18, 42, 46, 23, 0, 5, 0, 2, 1, 0, 22, 32, 46, 58, 64, 54, 44, 56, 61, 45, 
    101, 65, 69, 71, 43, 24, 20, 31, 34, 12, 7, 25, 30, 30, 42, 30, 17, 12, 14, 17, 5, 11, 23, 36, 53, 59, 65, 59, 27, 34, 59, 43, 
    107, 74, 64, 64, 43, 17, 13, 24, 44, 11, 16, 32, 32, 21, 40, 55, 38, 33, 32, 32, 31, 31, 29, 50, 53, 66, 71, 53, 27, 8, 44, 48, 
    107, 76, 74, 62, 29, 7, 4, 6, 47, 31, 8, 24, 40, 30, 51, 45, 49, 50, 43, 46, 42, 45, 47, 54, 61, 67, 78, 49, 21, 0, 26, 47, 
    108, 75, 68, 62, 30, 0, 0, 0, 48, 69, 7, 30, 42, 35, 53, 63, 42, 69, 58, 56, 54, 51, 58, 62, 66, 75, 74, 56, 6, 0, 6, 44, 
    108, 70, 60, 69, 35, 0, 0, 0, 23, 93, 48, 32, 45, 46, 64, 94, 44, 47, 59, 57, 58, 53, 64, 63, 59, 80, 73, 54, 12, 0, 0, 38, 
    105, 65, 67, 67, 37, 10, 7, 19, 21, 64, 77, 55, 56, 55, 74, 92, 65, 45, 43, 52, 61, 53, 61, 62, 56, 72, 79, 64, 22, 0, 0, 30, 
    106, 67, 68, 65, 50, 21, 13, 30, 34, 55, 68, 71, 74, 75, 73, 73, 70, 59, 48, 43, 54, 51, 58, 70, 58, 69, 73, 75, 41, 7, 0, 24, 
    108, 77, 69, 65, 56, 34, 24, 21, 39, 77, 71, 70, 79, 89, 78, 75, 55, 47, 56, 49, 50, 47, 49, 61, 67, 68, 65, 70, 73, 33, 4, 16, 
    113, 79, 81, 66, 57, 57, 35, 24, 40, 56, 60, 70, 76, 78, 82, 63, 46, 52, 56, 57, 54, 52, 47, 52, 69, 66, 67, 67, 81, 62, 23, 1, 
    110, 73, 87, 77, 50, 52, 59, 48, 32, 32, 62, 68, 85, 76, 68, 61, 56, 54, 55, 53, 52, 48, 53, 56, 59, 70, 71, 65, 71, 72, 49, 5, 
    108, 78, 77, 75, 62, 46, 59, 72, 43, 25, 63, 58, 70, 77, 71, 68, 67, 60, 58, 53, 53, 57, 63, 64, 58, 71, 71, 61, 73, 51, 68, 42, 
    107, 70, 74, 76, 68, 59, 56, 62, 80, 37, 58, 74, 71, 84, 77, 67, 73, 67, 61, 61, 69, 70, 70, 72, 67, 67, 70, 72, 74, 66, 51, 50, 
    104, 74, 71, 76, 76, 66, 70, 61, 67, 73, 54, 71, 78, 88, 81, 73, 69, 74, 72, 77, 78, 78, 80, 80, 72, 69, 73, 72, 73, 82, 54, 34, 
    112, 77, 66, 75, 84, 71, 73, 76, 68, 62, 72, 81, 74, 83, 82, 77, 72, 78, 81, 81, 83, 84, 84, 82, 73, 74, 73, 71, 73, 70, 75, 43, 
    104, 82, 70, 76, 72, 75, 78, 76, 73, 62, 73, 80, 76, 78, 76, 80, 77, 81, 79, 77, 88, 83, 81, 81, 74, 72, 75, 74, 68, 73, 77, 43, 
    92, 65, 61, 59, 54, 65, 64, 59, 56, 60, 61, 63, 60, 58, 57, 65, 71, 65, 63, 63, 66, 65, 64, 63, 62, 55, 62, 56, 56, 59, 62, 40, 
    
    -- channel=96
    166, 150, 156, 152, 153, 162, 162, 160, 164, 165, 161, 157, 155, 158, 162, 156, 153, 141, 112, 142, 136, 138, 136, 149, 129, 117, 120, 122, 136, 138, 138, 154, 
    144, 145, 158, 151, 146, 159, 166, 159, 165, 171, 169, 160, 153, 156, 168, 165, 156, 136, 98, 136, 165, 147, 140, 145, 119, 103, 102, 118, 141, 145, 139, 178, 
    141, 158, 173, 164, 153, 159, 169, 159, 161, 166, 164, 158, 150, 152, 161, 160, 153, 146, 148, 142, 143, 152, 141, 119, 114, 129, 115, 105, 135, 148, 142, 181, 
    144, 159, 169, 157, 156, 156, 165, 157, 155, 157, 156, 152, 145, 149, 154, 154, 149, 145, 146, 148, 139, 143, 141, 115, 123, 141, 119, 104, 131, 148, 141, 181, 
    139, 138, 143, 140, 156, 159, 158, 153, 149, 149, 150, 147, 142, 146, 149, 149, 146, 145, 142, 148, 132, 117, 122, 121, 128, 134, 113, 115, 130, 146, 137, 180, 
    118, 127, 137, 147, 155, 153, 151, 149, 147, 146, 148, 145, 142, 145, 145, 147, 143, 144, 143, 139, 94, 75, 96, 124, 138, 124, 105, 117, 125, 142, 140, 183, 
    115, 142, 152, 152, 148, 142, 148, 147, 147, 143, 143, 143, 143, 146, 141, 146, 141, 142, 145, 125, 65, 72, 97, 102, 139, 121, 103, 118, 130, 150, 147, 187, 
    129, 147, 147, 142, 144, 140, 147, 143, 145, 141, 140, 141, 139, 145, 137, 144, 138, 135, 138, 112, 83, 114, 122, 84, 115, 130, 125, 136, 141, 152, 145, 185, 
    132, 141, 143, 138, 143, 139, 146, 141, 141, 140, 140, 142, 127, 132, 122, 131, 126, 124, 128, 113, 117, 145, 136, 86, 105, 135, 141, 144, 141, 146, 143, 184, 
    130, 138, 144, 139, 144, 137, 143, 140, 139, 135, 128, 128, 104, 116, 115, 127, 135, 133, 130, 123, 113, 124, 110, 75, 111, 134, 133, 142, 140, 141, 141, 184, 
    131, 139, 145, 139, 145, 138, 140, 140, 137, 128, 109, 118, 106, 127, 118, 103, 92, 64, 48, 94, 83, 101, 102, 52, 95, 126, 136, 135, 135, 138, 139, 183, 
    134, 139, 145, 139, 144, 139, 140, 140, 134, 128, 114, 108, 60, 43, 28, 0, 0, 0, 0, 40, 46, 98, 160, 76, 65, 80, 132, 141, 128, 136, 138, 180, 
    136, 138, 143, 137, 142, 140, 139, 141, 130, 116, 79, 30, 0, 0, 0, 0, 16, 29, 28, 16, 0, 36, 197, 172, 81, 35, 71, 150, 129, 132, 139, 178, 
    137, 137, 143, 136, 140, 143, 135, 138, 108, 68, 31, 20, 27, 71, 91, 86, 86, 120, 104, 0, 0, 0, 120, 223, 133, 57, 31, 112, 134, 127, 137, 176, 
    135, 135, 143, 137, 136, 148, 138, 112, 69, 54, 84, 86, 75, 108, 134, 124, 82, 131, 106, 0, 0, 0, 16, 176, 178, 100, 60, 85, 124, 133, 132, 166, 
    134, 133, 143, 140, 130, 123, 127, 74, 71, 93, 101, 68, 67, 106, 134, 148, 88, 74, 12, 0, 0, 0, 0, 86, 167, 157, 103, 92, 90, 117, 132, 149, 
    134, 133, 140, 137, 114, 59, 75, 80, 79, 99, 60, 51, 73, 85, 77, 66, 1, 0, 0, 0, 0, 0, 13, 105, 126, 168, 148, 81, 21, 56, 158, 157, 
    132, 134, 135, 130, 120, 52, 48, 75, 64, 99, 93, 71, 97, 1, 0, 0, 0, 0, 0, 0, 0, 19, 132, 170, 104, 119, 133, 23, 0, 2, 182, 180, 
    131, 136, 130, 109, 125, 75, 52, 42, 85, 117, 115, 76, 107, 0, 0, 0, 0, 0, 0, 0, 0, 68, 190, 141, 65, 44, 26, 0, 0, 0, 165, 194, 
    133, 131, 82, 40, 92, 99, 67, 52, 119, 120, 104, 52, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 114, 97, 12, 0, 0, 0, 10, 9, 137, 197, 
    137, 83, 0, 0, 87, 147, 81, 59, 125, 127, 110, 62, 38, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 45, 4, 0, 0, 8, 18, 54, 147, 194, 
    130, 15, 0, 0, 94, 161, 88, 86, 132, 131, 110, 93, 48, 0, 0, 0, 0, 15, 89, 125, 88, 0, 0, 0, 12, 6, 5, 20, 58, 125, 161, 175, 
    110, 22, 21, 8, 41, 145, 95, 113, 137, 120, 68, 51, 24, 0, 0, 0, 0, 109, 147, 129, 94, 84, 0, 0, 8, 39, 30, 62, 121, 164, 132, 152, 
    99, 76, 124, 53, 0, 104, 113, 120, 131, 105, 23, 7, 0, 0, 0, 0, 17, 170, 126, 99, 92, 114, 59, 0, 0, 46, 49, 119, 152, 134, 102, 151, 
    106, 92, 100, 61, 0, 78, 135, 124, 105, 77, 24, 29, 0, 0, 0, 0, 61, 179, 98, 95, 106, 99, 102, 0, 0, 25, 90, 148, 135, 106, 97, 158, 
    114, 88, 67, 63, 0, 67, 148, 121, 82, 47, 31, 45, 0, 0, 0, 0, 75, 168, 74, 65, 106, 111, 118, 40, 0, 17, 126, 155, 123, 106, 105, 158, 
    116, 89, 65, 65, 0, 47, 129, 87, 26, 0, 0, 0, 0, 0, 0, 0, 57, 165, 76, 31, 66, 109, 114, 91, 0, 32, 143, 155, 123, 109, 105, 150, 
    116, 99, 60, 58, 2, 35, 90, 59, 9, 0, 0, 0, 0, 0, 0, 0, 61, 164, 87, 44, 42, 115, 134, 122, 56, 74, 142, 144, 119, 108, 98, 145, 
    113, 111, 75, 63, 50, 82, 117, 99, 77, 71, 70, 70, 67, 68, 74, 73, 88, 136, 62, 65, 89, 99, 131, 123, 113, 115, 127, 121, 116, 111, 97, 143, 
    100, 106, 111, 103, 103, 117, 125, 117, 102, 102, 107, 106, 105, 104, 108, 111, 113, 121, 59, 35, 80, 94, 131, 143, 126, 120, 121, 118, 114, 107, 98, 141, 
    93, 99, 109, 108, 100, 75, 69, 96, 95, 89, 90, 91, 97, 101, 105, 110, 112, 116, 100, 60, 63, 115, 142, 135, 122, 118, 118, 115, 110, 98, 98, 143, 
    74, 76, 59, 38, 35, 31, 45, 91, 85, 64, 59, 60, 69, 75, 76, 83, 90, 98, 98, 82, 81, 111, 118, 111, 109, 110, 110, 105, 98, 90, 96, 144, 
    
    -- channel=97
    9, 48, 50, 50, 53, 57, 60, 60, 57, 52, 41, 33, 31, 30, 25, 18, 11, 6, 10, 14, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 99, 96, 99, 100, 103, 105, 102, 96, 90, 79, 70, 67, 66, 63, 55, 44, 35, 26, 37, 51, 24, 24, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 98, 96, 99, 95, 92, 79, 72, 63, 57, 50, 45, 43, 43, 41, 36, 29, 21, 14, 16, 19, 16, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 93, 92, 96, 81, 67, 52, 43, 35, 31, 27, 24, 24, 23, 23, 20, 17, 13, 10, 9, 13, 23, 26, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 79, 73, 59, 44, 37, 26, 19, 14, 13, 12, 13, 13, 11, 12, 12, 15, 12, 13, 14, 25, 42, 59, 36, 7, 0, 0, 1, 12, 9, 2, 0, 
    0, 43, 33, 26, 20, 18, 8, 4, 3, 6, 8, 9, 9, 8, 13, 15, 19, 15, 17, 20, 29, 42, 51, 38, 11, 9, 16, 22, 22, 10, 0, 0, 
    0, 13, 10, 6, 4, 5, 2, 3, 4, 5, 6, 9, 11, 11, 18, 22, 26, 24, 31, 35, 29, 24, 26, 13, 9, 23, 23, 13, 15, 2, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 4, 4, 7, 9, 12, 19, 24, 39, 43, 52, 51, 52, 45, 24, 12, 0, 0, 2, 21, 8, 8, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 3, 6, 10, 17, 27, 45, 56, 65, 54, 54, 51, 50, 44, 28, 20, 13, 12, 11, 12, 5, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 5, 11, 22, 34, 52, 59, 75, 75, 97, 128, 159, 156, 134, 85, 51, 33, 11, 22, 20, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 1, 5, 9, 20, 36, 82, 135, 186, 209, 230, 250, 252, 226, 209, 182, 141, 78, 2, 16, 25, 29, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 2, 2, 7, 15, 39, 89, 154, 186, 194, 181, 170, 164, 157, 160, 209, 232, 215, 117, 6, 5, 25, 26, 22, 0, 0, 0, 
    0, 0, 0, 3, 2, 4, 3, 3, 15, 35, 79, 106, 110, 109, 115, 91, 73, 68, 66, 97, 188, 283, 297, 184, 45, 0, 0, 20, 16, 0, 0, 0, 
    0, 3, 2, 6, 2, 0, 1, 6, 25, 50, 63, 60, 75, 84, 68, 31, 15, 0, 14, 72, 180, 298, 339, 251, 119, 9, 0, 0, 1, 0, 0, 0, 
    0, 6, 3, 6, 3, 8, 20, 38, 37, 45, 41, 65, 67, 57, 37, 0, 0, 15, 84, 174, 255, 317, 344, 284, 174, 34, 0, 0, 0, 13, 21, 0, 
    0, 7, 3, 6, 7, 30, 51, 62, 59, 55, 77, 52, 45, 57, 79, 107, 169, 216, 278, 302, 316, 350, 329, 248, 140, 27, 0, 0, 19, 84, 88, 8, 
    0, 6, 2, 5, 3, 23, 40, 53, 64, 71, 41, 22, 20, 65, 130, 236, 308, 310, 326, 335, 358, 345, 269, 149, 74, 23, 0, 29, 99, 161, 139, 47, 
    0, 2, 0, 16, 21, 50, 46, 61, 61, 38, 13, 7, 13, 93, 177, 283, 343, 344, 350, 362, 375, 338, 256, 167, 76, 44, 93, 132, 165, 196, 169, 79, 
    0, 0, 22, 72, 109, 103, 39, 22, 20, 17, 0, 0, 7, 98, 175, 291, 348, 342, 348, 357, 357, 339, 300, 233, 158, 148, 178, 190, 194, 214, 173, 78, 
    0, 8, 73, 169, 200, 139, 58, 18, 3, 0, 0, 0, 0, 84, 165, 288, 328, 322, 306, 271, 227, 228, 255, 264, 247, 233, 235, 238, 230, 198, 132, 37, 
    0, 22, 100, 191, 201, 158, 81, 12, 0, 0, 0, 0, 0, 101, 181, 288, 317, 290, 234, 140, 81, 110, 169, 227, 275, 274, 256, 229, 194, 135, 54, 0, 
    0, 14, 51, 114, 139, 129, 95, 13, 0, 0, 0, 0, 52, 140, 203, 290, 308, 246, 163, 61, 29, 24, 71, 148, 217, 245, 221, 186, 132, 46, 5, 0, 
    0, 0, 2, 66, 112, 116, 107, 18, 0, 0, 0, 28, 86, 152, 216, 312, 303, 217, 130, 25, 0, 0, 0, 62, 141, 206, 203, 143, 66, 6, 0, 0, 
    0, 0, 0, 46, 75, 96, 108, 22, 0, 0, 12, 49, 114, 187, 257, 314, 281, 195, 113, 7, 6, 7, 0, 8, 78, 165, 174, 104, 32, 0, 0, 0, 
    0, 0, 0, 33, 69, 91, 103, 29, 0, 3, 48, 86, 150, 201, 253, 297, 263, 192, 107, 16, 28, 18, 0, 0, 37, 113, 132, 70, 0, 0, 0, 0, 
    0, 0, 0, 29, 76, 93, 108, 67, 43, 84, 144, 186, 229, 251, 286, 313, 275, 199, 107, 34, 57, 62, 29, 0, 9, 51, 76, 31, 0, 0, 0, 0, 
    0, 0, 0, 21, 75, 86, 100, 66, 47, 76, 112, 140, 160, 170, 196, 204, 178, 125, 74, 29, 60, 42, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 26, 28, 25, 2, 0, 0, 22, 43, 57, 62, 67, 69, 60, 36, 24, 5, 45, 52, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 34, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 21, 31, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 20, 44, 66, 80, 72, 47, 25, 10, 18, 25, 27, 26, 21, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    36, 41, 38, 45, 55, 50, 48, 55, 54, 49, 50, 53, 56, 53, 46, 47, 51, 57, 65, 24, 18, 34, 36, 33, 54, 36, 18, 26, 22, 28, 36, 16, 
    59, 84, 81, 90, 102, 96, 94, 103, 100, 94, 93, 94, 98, 95, 83, 82, 86, 94, 104, 56, 37, 63, 58, 60, 69, 37, 29, 36, 32, 44, 57, 28, 
    67, 102, 95, 96, 96, 90, 94, 101, 101, 96, 93, 92, 95, 91, 83, 81, 83, 82, 77, 68, 62, 67, 72, 73, 52, 15, 19, 34, 35, 47, 61, 31, 
    71, 109, 98, 90, 82, 84, 92, 97, 97, 93, 89, 86, 88, 85, 81, 78, 77, 75, 73, 69, 76, 83, 63, 45, 28, 8, 22, 38, 40, 53, 61, 32, 
    70, 98, 83, 81, 77, 81, 88, 89, 89, 87, 83, 80, 80, 78, 78, 74, 73, 71, 70, 69, 96, 90, 30, 13, 10, 12, 41, 40, 42, 49, 53, 30, 
    63, 83, 73, 74, 75, 79, 82, 82, 82, 81, 79, 75, 74, 74, 76, 70, 68, 70, 66, 74, 113, 73, 0, 0, 8, 19, 45, 38, 45, 44, 48, 28, 
    58, 70, 65, 73, 76, 77, 75, 76, 76, 77, 77, 72, 73, 74, 77, 71, 69, 71, 64, 76, 105, 37, 0, 6, 9, 21, 40, 42, 50, 48, 52, 28, 
    51, 69, 69, 75, 74, 74, 70, 73, 72, 76, 77, 74, 80, 76, 74, 68, 64, 65, 61, 74, 74, 4, 0, 31, 27, 24, 46, 52, 54, 57, 63, 31, 
    50, 69, 71, 76, 74, 75, 72, 73, 72, 77, 83, 80, 80, 66, 63, 63, 61, 65, 68, 67, 45, 0, 0, 30, 35, 38, 57, 62, 60, 63, 65, 31, 
    49, 68, 70, 76, 75, 76, 74, 75, 74, 81, 89, 78, 81, 65, 58, 71, 71, 71, 63, 18, 0, 0, 0, 12, 39, 39, 52, 58, 62, 62, 63, 31, 
    47, 70, 72, 77, 75, 75, 74, 75, 75, 81, 92, 90, 103, 73, 41, 46, 41, 34, 24, 0, 0, 0, 0, 0, 30, 46, 40, 30, 51, 60, 61, 31, 
    48, 74, 73, 77, 75, 73, 73, 74, 77, 92, 107, 93, 81, 38, 3, 12, 14, 11, 1, 0, 24, 0, 0, 0, 5, 49, 36, 14, 30, 54, 57, 32, 
    50, 77, 74, 76, 74, 71, 72, 73, 92, 106, 84, 62, 63, 21, 0, 0, 1, 0, 0, 47, 109, 0, 0, 0, 0, 47, 54, 4, 15, 45, 54, 32, 
    51, 79, 73, 74, 75, 69, 74, 84, 105, 83, 48, 46, 40, 0, 0, 0, 13, 4, 15, 123, 142, 0, 0, 0, 0, 0, 58, 10, 8, 36, 48, 29, 
    51, 78, 72, 72, 79, 82, 77, 79, 85, 51, 24, 22, 21, 0, 0, 0, 42, 40, 58, 116, 67, 0, 0, 0, 0, 0, 19, 24, 28, 33, 16, 4, 
    51, 77, 73, 74, 86, 95, 68, 56, 52, 14, 0, 31, 25, 0, 7, 14, 28, 25, 25, 31, 0, 0, 0, 0, 0, 0, 0, 46, 78, 23, 0, 0, 
    51, 75, 74, 79, 85, 93, 58, 39, 24, 0, 0, 31, 13, 38, 85, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 72, 88, 1, 0, 0, 
    51, 74, 80, 99, 78, 51, 38, 22, 0, 0, 0, 33, 14, 88, 134, 18, 0, 0, 0, 0, 0, 0, 0, 0, 10, 40, 24, 55, 49, 0, 0, 0, 
    50, 80, 115, 129, 20, 0, 4, 34, 0, 0, 0, 47, 24, 118, 136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 34, 15, 11, 0, 0, 0, 0, 
    49, 108, 175, 113, 0, 0, 0, 23, 0, 0, 16, 55, 45, 128, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 148, 193, 57, 0, 0, 0, 4, 0, 0, 30, 61, 63, 129, 78, 0, 0, 0, 0, 0, 0, 36, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 161, 140, 23, 0, 0, 0, 0, 0, 0, 51, 65, 48, 108, 53, 0, 0, 0, 0, 0, 2, 37, 90, 67, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 139, 73, 29, 34, 0, 0, 0, 0, 23, 72, 60, 28, 90, 36, 0, 0, 0, 0, 0, 4, 12, 79, 114, 29, 0, 0, 0, 0, 0, 16, 0, 
    68, 110, 45, 32, 78, 0, 0, 0, 0, 39, 75, 45, 32, 73, 1, 0, 0, 0, 0, 13, 3, 0, 18, 108, 80, 0, 0, 0, 0, 6, 35, 0, 
    62, 100, 63, 29, 76, 0, 0, 0, 20, 53, 58, 15, 34, 58, 0, 0, 0, 0, 0, 18, 0, 0, 0, 70, 110, 17, 0, 0, 0, 27, 38, 0, 
    54, 91, 75, 31, 64, 0, 0, 0, 37, 55, 32, 0, 11, 16, 0, 0, 0, 0, 0, 36, 0, 0, 0, 27, 104, 34, 0, 0, 0, 34, 41, 4, 
    48, 74, 74, 38, 49, 0, 0, 0, 31, 37, 16, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 1, 73, 32, 0, 0, 13, 33, 43, 8, 
    49, 60, 64, 37, 36, 0, 0, 0, 27, 29, 18, 0, 0, 0, 0, 0, 0, 0, 4, 49, 2, 0, 0, 0, 36, 29, 0, 0, 21, 31, 40, 4, 
    53, 47, 51, 35, 22, 0, 0, 2, 12, 16, 15, 11, 11, 7, 1, 1, 0, 0, 35, 47, 14, 0, 0, 0, 18, 23, 15, 21, 27, 31, 38, 0, 
    56, 42, 37, 32, 19, 7, 0, 0, 0, 13, 16, 11, 8, 5, 6, 7, 9, 7, 43, 54, 16, 0, 0, 0, 17, 23, 23, 25, 29, 33, 31, 0, 
    58, 42, 43, 32, 8, 0, 0, 0, 0, 8, 5, 0, 0, 0, 0, 0, 0, 0, 14, 40, 30, 0, 0, 2, 20, 22, 19, 22, 28, 31, 22, 0, 
    44, 40, 42, 32, 9, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 2, 7, 17, 15, 0, 2, 18, 21, 20, 19, 22, 25, 27, 21, 0, 
    
    -- channel=99
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    97, 46, 63, 79, 96, 108, 113, 116, 119, 114, 107, 103, 105, 107, 105, 96, 93, 92, 101, 118, 126, 92, 82, 80, 53, 71, 99, 106, 79, 59, 54, 61, 
    146, 92, 100, 96, 97, 111, 109, 104, 103, 98, 91, 88, 89, 93, 93, 86, 84, 79, 70, 70, 80, 76, 66, 72, 76, 85, 85, 84, 73, 57, 51, 56, 
    156, 102, 94, 82, 81, 89, 91, 84, 82, 81, 77, 75, 74, 78, 78, 75, 72, 70, 62, 64, 66, 56, 47, 63, 71, 67, 50, 45, 56, 47, 47, 53, 
    138, 83, 88, 83, 84, 82, 76, 70, 72, 74, 69, 65, 63, 67, 69, 66, 63, 62, 59, 63, 55, 21, 27, 39, 56, 58, 37, 40, 45, 42, 43, 51, 
    138, 93, 98, 99, 91, 81, 69, 63, 66, 66, 59, 52, 50, 53, 57, 58, 54, 54, 51, 55, 43, 37, 57, 66, 53, 45, 40, 44, 45, 48, 44, 55, 
    134, 99, 89, 74, 65, 60, 59, 55, 56, 54, 48, 41, 37, 37, 42, 46, 49, 50, 48, 54, 58, 81, 118, 121, 87, 43, 49, 57, 68, 66, 57, 62, 
    101, 64, 53, 48, 47, 43, 45, 42, 45, 44, 40, 39, 36, 30, 32, 36, 40, 44, 44, 50, 62, 84, 105, 102, 86, 61, 56, 67, 71, 67, 57, 60, 
    81, 42, 38, 38, 41, 39, 40, 37, 40, 40, 36, 33, 35, 32, 33, 34, 37, 50, 50, 54, 59, 53, 54, 50, 60, 57, 58, 59, 60, 59, 54, 56, 
    77, 38, 37, 37, 40, 38, 41, 39, 40, 41, 37, 37, 47, 49, 53, 50, 40, 23, 1, 0, 9, 7, 16, 40, 54, 55, 60, 64, 60, 59, 54, 55, 
    77, 36, 36, 36, 39, 38, 43, 43, 44, 44, 51, 59, 51, 28, 1, 0, 0, 0, 0, 0, 0, 0, 0, 63, 107, 86, 47, 54, 61, 58, 55, 57, 
    80, 36, 34, 34, 38, 38, 42, 44, 46, 45, 34, 22, 4, 0, 0, 0, 22, 56, 96, 107, 37, 0, 0, 0, 113, 132, 85, 27, 50, 58, 56, 58, 
    82, 36, 36, 34, 36, 38, 43, 46, 45, 24, 11, 21, 45, 86, 155, 211, 238, 242, 255, 243, 161, 61, 0, 0, 25, 108, 121, 78, 45, 59, 58, 60, 
    82, 36, 36, 35, 35, 39, 44, 50, 29, 29, 59, 102, 134, 150, 161, 178, 181, 148, 121, 89, 58, 52, 16, 0, 0, 54, 106, 124, 87, 72, 69, 64, 
    82, 36, 36, 35, 39, 37, 23, 33, 34, 72, 91, 100, 82, 67, 63, 57, 61, 52, 0, 0, 0, 15, 29, 0, 0, 0, 67, 101, 99, 57, 50, 68, 
    83, 38, 37, 37, 40, 33, 7, 5, 46, 54, 83, 57, 51, 52, 29, 0, 0, 0, 0, 0, 0, 15, 40, 83, 63, 6, 23, 61, 39, 0, 0, 38, 
    81, 36, 37, 39, 45, 58, 72, 56, 38, 56, 68, 102, 107, 86, 0, 0, 0, 0, 0, 0, 4, 28, 91, 143, 136, 83, 12, 6, 0, 0, 0, 12, 
    79, 34, 38, 37, 26, 63, 114, 114, 84, 93, 105, 123, 114, 92, 37, 0, 0, 37, 61, 60, 46, 46, 65, 87, 66, 15, 0, 0, 0, 0, 0, 15, 
    81, 38, 30, 0, 0, 0, 57, 80, 89, 101, 106, 81, 55, 34, 56, 75, 91, 93, 79, 68, 61, 32, 0, 0, 0, 0, 0, 0, 0, 44, 58, 48, 
    80, 41, 0, 0, 0, 0, 42, 71, 76, 84, 87, 85, 78, 54, 48, 60, 64, 49, 54, 105, 150, 130, 26, 0, 0, 0, 0, 21, 42, 65, 101, 94, 
    80, 31, 0, 6, 2, 6, 27, 54, 80, 80, 82, 82, 88, 91, 68, 50, 48, 46, 109, 188, 240, 262, 220, 82, 0, 2, 36, 51, 66, 115, 134, 115, 
    79, 35, 75, 151, 136, 50, 29, 58, 82, 86, 70, 31, 11, 28, 56, 50, 46, 74, 138, 153, 148, 158, 211, 201, 94, 59, 70, 89, 132, 150, 137, 101, 
    78, 56, 103, 163, 175, 76, 33, 65, 72, 69, 45, 14, 0, 0, 18, 35, 41, 81, 100, 86, 55, 59, 98, 174, 155, 88, 76, 105, 135, 129, 91, 64, 
    83, 62, 50, 49, 66, 51, 32, 59, 74, 52, 34, 48, 56, 40, 32, 26, 42, 62, 67, 60, 52, 67, 77, 110, 135, 70, 48, 84, 96, 80, 57, 56, 
    88, 61, 44, 35, 44, 55, 42, 54, 59, 37, 17, 27, 39, 46, 51, 60, 62, 56, 57, 44, 22, 30, 51, 87, 120, 93, 67, 80, 84, 76, 73, 72, 
    83, 59, 55, 55, 61, 63, 40, 34, 29, 5, 0, 0, 0, 20, 48, 57, 47, 37, 47, 52, 22, 5, 32, 60, 112, 130, 111, 98, 90, 88, 87, 81, 
    73, 50, 50, 43, 54, 63, 48, 19, 14, 14, 15, 11, 15, 42, 74, 81, 76, 52, 45, 54, 54, 26, 29, 58, 101, 152, 141, 105, 86, 82, 81, 74, 
    69, 41, 47, 61, 68, 104, 111, 108, 119, 152, 191, 217, 226, 229, 231, 231, 218, 169, 99, 70, 79, 101, 71, 86, 100, 134, 138, 107, 80, 75, 76, 73, 
    65, 37, 43, 75, 115, 139, 137, 126, 133, 148, 161, 171, 180, 186, 188, 187, 184, 166, 130, 106, 59, 41, 62, 60, 83, 87, 88, 81, 76, 73, 70, 71, 
    68, 41, 39, 42, 56, 59, 39, 21, 29, 43, 42, 40, 41, 47, 52, 55, 61, 68, 83, 105, 109, 79, 75, 83, 76, 71, 70, 71, 72, 71, 67, 67, 
    73, 53, 39, 11, 0, 0, 0, 0, 13, 24, 26, 22, 20, 20, 20, 21, 24, 33, 43, 61, 87, 103, 98, 83, 67, 61, 63, 64, 64, 63, 68, 69, 
    107, 95, 91, 81, 75, 76, 88, 94, 82, 79, 76, 80, 83, 79, 74, 69, 67, 68, 67, 66, 68, 67, 66, 72, 76, 75, 73, 74, 78, 83, 88, 89, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 10, 10, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 12, 15, 15, 11, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 33, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 10, 14, 10, 6, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 42, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 5, 2, 0, 0, 0, 0, 0, 0, 0, 1, 6, 3, 0, 0, 0, 0, 0, 0, 0, 10, 47, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 8, 14, 7, 9, 2, 6, 0, 0, 22, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 2, 0, 1, 2, 4, 6, 19, 30, 22, 17, 7, 10, 3, 8, 30, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 4, 3, 3, 2, 4, 7, 17, 33, 32, 42, 51, 72, 84, 89, 67, 36, 1, 0, 8, 10, 0, 0, 0, 0, 0, 
    0, 0, 2, 3, 0, 5, 0, 4, 3, 1, 0, 5, 17, 52, 94, 104, 113, 125, 140, 166, 160, 131, 128, 56, 0, 0, 15, 18, 0, 0, 0, 0, 
    0, 0, 3, 7, 2, 5, 0, 2, 0, 0, 5, 27, 53, 88, 124, 120, 114, 118, 129, 153, 151, 167, 231, 130, 0, 0, 3, 32, 20, 0, 0, 0, 
    0, 0, 4, 10, 7, 6, 1, 0, 0, 0, 22, 46, 56, 84, 117, 101, 81, 81, 80, 69, 68, 176, 306, 224, 48, 0, 0, 28, 37, 0, 0, 0, 
    0, 4, 6, 11, 8, 7, 4, 0, 0, 8, 41, 49, 53, 84, 93, 48, 7, 0, 9, 0, 15, 179, 314, 288, 153, 0, 0, 0, 23, 0, 0, 0, 
    0, 8, 7, 11, 4, 6, 16, 11, 4, 29, 48, 48, 34, 54, 55, 4, 0, 0, 7, 8, 85, 219, 289, 305, 234, 55, 0, 0, 0, 0, 8, 0, 
    0, 11, 10, 11, 0, 1, 28, 35, 40, 48, 51, 15, 14, 49, 51, 45, 54, 68, 106, 129, 194, 265, 277, 282, 213, 74, 0, 0, 0, 25, 77, 20, 
    0, 13, 9, 6, 0, 0, 17, 44, 51, 61, 27, 0, 0, 28, 29, 98, 163, 170, 197, 234, 272, 281, 280, 228, 118, 51, 29, 0, 0, 81, 161, 85, 
    0, 13, 7, 2, 1, 24, 20, 34, 43, 53, 20, 0, 0, 0, 10, 148, 248, 257, 272, 285, 290, 300, 302, 212, 66, 31, 73, 53, 60, 134, 210, 137, 
    0, 6, 2, 9, 65, 98, 33, 4, 26, 42, 0, 0, 0, 0, 16, 192, 282, 271, 268, 271, 273, 297, 314, 229, 107, 84, 117, 127, 136, 166, 208, 145, 
    0, 0, 0, 51, 164, 172, 67, 6, 22, 23, 0, 0, 0, 0, 42, 209, 266, 250, 247, 237, 198, 194, 241, 246, 190, 164, 176, 188, 186, 170, 175, 102, 
    0, 0, 0, 100, 214, 207, 96, 8, 15, 0, 0, 0, 0, 0, 63, 215, 250, 236, 243, 188, 94, 66, 111, 187, 231, 227, 215, 194, 174, 156, 114, 29, 
    0, 0, 0, 100, 159, 171, 115, 22, 10, 0, 0, 0, 0, 14, 82, 219, 239, 239, 233, 114, 22, 0, 0, 68, 184, 232, 204, 173, 156, 107, 38, 0, 
    0, 0, 10, 66, 62, 122, 129, 38, 0, 0, 0, 0, 30, 51, 111, 233, 243, 254, 196, 33, 0, 0, 0, 0, 94, 196, 190, 160, 121, 42, 0, 0, 
    0, 0, 16, 31, 0, 82, 139, 50, 0, 0, 0, 0, 61, 81, 154, 241, 248, 256, 148, 0, 0, 2, 0, 0, 9, 135, 174, 154, 79, 0, 0, 0, 
    0, 0, 0, 19, 7, 71, 143, 58, 0, 0, 0, 42, 78, 87, 170, 237, 247, 247, 119, 0, 21, 19, 0, 0, 0, 70, 160, 135, 30, 0, 0, 0, 
    0, 0, 0, 16, 23, 69, 141, 75, 0, 4, 61, 118, 132, 138, 204, 239, 250, 243, 112, 0, 41, 64, 40, 0, 0, 12, 120, 92, 0, 0, 0, 0, 
    0, 0, 0, 8, 29, 61, 122, 69, 4, 18, 65, 112, 126, 131, 166, 178, 194, 197, 96, 0, 40, 68, 45, 0, 0, 0, 46, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 30, 61, 23, 0, 0, 23, 53, 67, 73, 82, 87, 97, 106, 42, 0, 34, 67, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 2, 0, 0, 20, 40, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 1, 1, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 10, 26, 37, 40, 39, 44, 29, 0, 0, 4, 7, 5, 1, 0, 0, 0, 0, 0, 0, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=101
    21, 33, 38, 44, 53, 60, 62, 64, 64, 59, 53, 47, 47, 48, 44, 38, 33, 31, 34, 42, 56, 27, 23, 14, 9, 5, 6, 21, 7, 0, 0, 0, 
    74, 74, 78, 76, 81, 85, 84, 83, 80, 74, 64, 58, 58, 59, 52, 44, 40, 46, 60, 41, 37, 30, 27, 22, 17, 19, 22, 12, 8, 0, 0, 0, 
    88, 82, 78, 74, 70, 62, 58, 54, 49, 43, 37, 33, 35, 37, 33, 28, 24, 24, 15, 16, 24, 15, 18, 27, 14, 0, 2, 8, 3, 0, 0, 0, 
    83, 65, 61, 57, 51, 47, 34, 28, 24, 21, 17, 16, 18, 19, 20, 17, 14, 15, 9, 8, 22, 24, 14, 13, 10, 0, 0, 13, 5, 0, 0, 0, 
    71, 54, 48, 50, 39, 31, 16, 10, 11, 11, 8, 6, 7, 7, 11, 11, 9, 11, 11, 6, 23, 42, 26, 25, 10, 0, 6, 16, 14, 0, 0, 0, 
    57, 49, 42, 28, 13, 7, 3, 0, 1, 2, 1, 0, 0, 2, 7, 10, 9, 10, 12, 16, 42, 58, 52, 40, 27, 13, 17, 18, 23, 11, 3, 0, 
    41, 19, 7, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 7, 15, 18, 20, 21, 29, 60, 59, 47, 38, 26, 30, 31, 35, 28, 11, 3, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 5, 11, 11, 16, 22, 26, 25, 25, 43, 54, 30, 19, 25, 20, 23, 29, 22, 12, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 15, 25, 25, 27, 29, 41, 45, 45, 52, 37, 12, 3, 17, 21, 14, 8, 7, 7, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 25, 48, 61, 60, 58, 66, 69, 63, 49, 18, 10, 8, 33, 45, 23, 5, 0, 6, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 1, 6, 21, 43, 79, 83, 79, 74, 85, 107, 128, 125, 128, 88, 29, 21, 37, 43, 34, 0, 0, 1, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 2, 15, 40, 53, 80, 105, 137, 166, 194, 222, 224, 196, 213, 187, 93, 42, 16, 35, 39, 31, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 12, 33, 45, 81, 151, 184, 174, 172, 171, 160, 133, 144, 218, 214, 133, 52, 0, 32, 43, 29, 16, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 4, 27, 48, 81, 122, 133, 103, 75, 49, 38, 34, 32, 102, 208, 235, 179, 83, 12, 1, 43, 20, 18, 5, 0, 0, 
    12, 0, 0, 0, 0, 1, 6, 7, 40, 66, 81, 63, 64, 44, 18, 10, 23, 22, 53, 133, 212, 265, 230, 117, 45, 20, 12, 18, 15, 17, 0, 0, 
    13, 0, 0, 0, 7, 18, 30, 47, 56, 65, 29, 64, 75, 61, 55, 45, 56, 63, 112, 208, 270, 272, 239, 135, 71, 35, 0, 13, 45, 41, 10, 0, 
    12, 0, 0, 0, 15, 44, 61, 87, 74, 46, 67, 80, 74, 76, 124, 130, 164, 220, 274, 299, 290, 261, 199, 127, 60, 0, 9, 29, 80, 97, 53, 0, 
    10, 0, 0, 14, 30, 43, 58, 63, 73, 52, 57, 57, 55, 95, 187, 255, 298, 304, 303, 291, 282, 248, 142, 31, 20, 15, 12, 68, 136, 166, 78, 0, 
    8, 0, 17, 55, 31, 25, 42, 69, 61, 26, 13, 37, 40, 142, 242, 276, 280, 272, 267, 264, 275, 228, 128, 57, 49, 65, 89, 150, 188, 184, 79, 7, 
    5, 1, 67, 112, 82, 67, 38, 48, 24, 6, 6, 30, 46, 165, 247, 249, 245, 247, 240, 236, 258, 252, 201, 170, 153, 163, 184, 182, 176, 166, 76, 13, 
    2, 24, 125, 180, 165, 82, 40, 41, 6, 2, 0, 29, 54, 148, 222, 237, 242, 237, 193, 181, 181, 187, 200, 230, 230, 208, 195, 191, 170, 123, 65, 1, 
    2, 56, 141, 183, 168, 92, 52, 35, 0, 0, 0, 31, 56, 153, 211, 234, 242, 197, 117, 74, 46, 92, 151, 193, 228, 208, 195, 168, 119, 75, 19, 0, 
    9, 57, 90, 113, 104, 76, 53, 14, 0, 0, 21, 53, 92, 200, 236, 231, 231, 134, 50, 12, 13, 40, 108, 156, 186, 182, 153, 112, 60, 10, 0, 0, 
    14, 26, 20, 54, 109, 88, 56, 12, 0, 9, 55, 89, 130, 206, 225, 244, 217, 94, 42, 29, 29, 4, 31, 117, 145, 159, 131, 62, 14, 0, 8, 0, 
    8, 10, 19, 55, 127, 101, 49, 11, 15, 36, 80, 95, 134, 205, 237, 251, 194, 77, 43, 35, 31, 19, 11, 67, 126, 150, 111, 36, 4, 6, 18, 0, 
    1, 4, 30, 56, 117, 104, 55, 21, 37, 70, 102, 113, 161, 207, 227, 226, 168, 69, 50, 58, 57, 31, 0, 35, 104, 127, 76, 17, 0, 3, 11, 0, 
    0, 0, 28, 56, 103, 100, 55, 50, 73, 118, 155, 173, 211, 233, 230, 232, 183, 96, 72, 73, 60, 55, 28, 24, 74, 76, 40, 6, 0, 0, 2, 0, 
    5, 5, 22, 43, 97, 94, 69, 68, 92, 126, 145, 150, 157, 166, 168, 166, 126, 56, 64, 85, 81, 38, 20, 0, 30, 28, 0, 0, 0, 0, 1, 0, 
    12, 5, 25, 33, 53, 52, 35, 23, 22, 33, 40, 41, 44, 46, 44, 43, 32, 1, 26, 44, 71, 40, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    20, 15, 15, 22, 22, 10, 0, 0, 0, 0, 4, 4, 4, 2, 0, 0, 0, 0, 20, 37, 31, 42, 21, 0, 0, 0, 0, 0, 0, 0, 12, 0, 
    27, 23, 24, 26, 31, 39, 45, 35, 28, 25, 23, 26, 27, 24, 17, 9, 2, 0, 7, 30, 35, 7, 0, 0, 0, 0, 0, 0, 0, 9, 15, 0, 
    16, 34, 41, 62, 82, 102, 99, 67, 48, 43, 52, 56, 54, 53, 49, 43, 37, 29, 23, 23, 23, 11, 4, 0, 0, 0, 0, 1, 4, 14, 19, 0, 
    
    -- channel=102
    73, 57, 59, 53, 52, 57, 58, 54, 58, 58, 55, 51, 48, 50, 55, 51, 46, 41, 30, 52, 57, 51, 44, 53, 34, 29, 29, 38, 50, 45, 40, 59, 
    62, 63, 70, 66, 63, 72, 76, 72, 75, 76, 73, 68, 63, 65, 71, 69, 63, 59, 53, 37, 52, 62, 44, 41, 44, 40, 28, 35, 50, 52, 49, 73, 
    56, 65, 74, 71, 69, 68, 74, 68, 67, 68, 68, 63, 59, 61, 64, 64, 61, 59, 61, 53, 47, 57, 52, 41, 46, 51, 35, 26, 45, 51, 49, 74, 
    50, 63, 75, 71, 71, 65, 69, 64, 59, 61, 61, 58, 55, 58, 58, 59, 57, 56, 54, 56, 45, 43, 58, 50, 48, 51, 32, 28, 39, 51, 51, 74, 
    47, 61, 67, 63, 62, 62, 63, 58, 55, 56, 58, 56, 53, 53, 54, 57, 55, 56, 53, 54, 36, 36, 55, 56, 52, 40, 27, 37, 39, 56, 52, 76, 
    41, 56, 55, 54, 52, 53, 57, 54, 55, 54, 55, 55, 53, 53, 52, 57, 54, 55, 54, 47, 25, 36, 39, 40, 58, 43, 37, 41, 48, 59, 50, 78, 
    37, 52, 51, 52, 54, 50, 56, 52, 55, 53, 53, 53, 52, 55, 51, 54, 51, 51, 54, 42, 30, 41, 30, 18, 50, 53, 41, 39, 47, 54, 48, 77, 
    41, 52, 51, 49, 52, 49, 54, 50, 52, 52, 51, 49, 42, 51, 51, 55, 53, 54, 55, 46, 47, 48, 34, 14, 35, 45, 40, 43, 46, 53, 52, 77, 
    44, 50, 52, 47, 51, 48, 52, 50, 50, 49, 47, 49, 40, 52, 54, 57, 52, 48, 47, 47, 50, 48, 40, 19, 31, 40, 45, 51, 47, 52, 53, 77, 
    45, 48, 51, 47, 51, 47, 50, 49, 47, 45, 40, 47, 36, 47, 41, 39, 40, 39, 46, 66, 46, 48, 45, 13, 29, 47, 50, 54, 48, 50, 51, 76, 
    46, 47, 51, 47, 51, 48, 50, 49, 47, 44, 35, 35, 23, 38, 37, 32, 37, 34, 40, 70, 49, 70, 77, 8, 12, 33, 62, 56, 48, 48, 49, 74, 
    47, 46, 51, 47, 51, 49, 48, 50, 44, 36, 29, 26, 17, 24, 30, 24, 22, 11, 3, 4, 0, 64, 113, 50, 6, 0, 37, 66, 47, 46, 47, 73, 
    48, 46, 51, 48, 51, 50, 46, 50, 35, 28, 27, 18, 9, 13, 7, 0, 0, 4, 0, 0, 0, 8, 95, 109, 35, 0, 0, 52, 49, 45, 47, 71, 
    48, 47, 52, 48, 48, 52, 43, 40, 25, 31, 26, 13, 7, 25, 24, 12, 0, 29, 9, 0, 0, 0, 42, 122, 80, 15, 0, 18, 41, 41, 46, 71, 
    48, 47, 53, 48, 42, 45, 48, 28, 29, 24, 30, 16, 20, 36, 41, 38, 9, 28, 19, 0, 0, 0, 5, 85, 93, 51, 21, 7, 16, 42, 56, 67, 
    47, 46, 50, 47, 36, 24, 47, 36, 29, 38, 25, 16, 27, 31, 27, 47, 30, 23, 17, 3, 0, 0, 19, 46, 50, 77, 39, 5, 0, 46, 80, 65, 
    47, 46, 46, 43, 36, 10, 20, 33, 30, 51, 17, 9, 25, 0, 0, 37, 27, 18, 7, 0, 0, 17, 43, 34, 17, 44, 40, 2, 0, 27, 96, 74, 
    46, 46, 41, 32, 52, 24, 8, 11, 32, 34, 25, 10, 30, 0, 0, 0, 0, 0, 0, 0, 0, 37, 67, 42, 13, 11, 31, 13, 0, 0, 91, 85, 
    46, 41, 18, 26, 75, 46, 17, 4, 35, 29, 27, 6, 28, 0, 0, 0, 0, 0, 0, 0, 0, 23, 84, 60, 18, 15, 19, 17, 3, 0, 73, 82, 
    47, 21, 0, 35, 76, 64, 20, 6, 44, 32, 23, 1, 1, 0, 0, 0, 0, 0, 5, 0, 0, 0, 32, 55, 28, 16, 8, 9, 10, 22, 51, 67, 
    43, 0, 0, 15, 53, 77, 26, 20, 41, 31, 26, 11, 0, 0, 0, 0, 0, 13, 23, 0, 0, 0, 0, 6, 23, 12, 3, 6, 24, 33, 35, 60, 
    35, 0, 0, 0, 11, 72, 30, 35, 36, 30, 15, 20, 15, 0, 0, 0, 0, 47, 27, 18, 18, 0, 0, 0, 6, 9, 1, 18, 30, 30, 30, 58, 
    29, 15, 17, 0, 0, 56, 40, 37, 36, 29, 0, 13, 7, 0, 0, 0, 13, 71, 28, 34, 26, 31, 0, 0, 0, 9, 13, 38, 31, 33, 31, 58, 
    29, 24, 33, 13, 0, 41, 54, 34, 29, 24, 0, 3, 0, 0, 0, 0, 32, 77, 28, 32, 28, 32, 23, 0, 0, 12, 36, 48, 35, 33, 29, 60, 
    31, 24, 23, 20, 0, 30, 59, 33, 19, 14, 8, 10, 0, 0, 0, 0, 39, 77, 22, 23, 41, 37, 37, 0, 0, 4, 49, 48, 32, 28, 26, 57, 
    31, 27, 17, 13, 0, 18, 57, 28, 12, 5, 9, 20, 0, 0, 0, 0, 41, 79, 16, 5, 38, 48, 42, 12, 0, 0, 47, 42, 29, 25, 24, 53, 
    34, 31, 13, 15, 0, 12, 43, 25, 6, 0, 0, 1, 0, 0, 0, 0, 25, 72, 17, 1, 14, 49, 39, 34, 0, 0, 35, 38, 30, 25, 24, 53, 
    35, 35, 14, 12, 0, 9, 22, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 6, 15, 11, 25, 46, 34, 15, 12, 27, 33, 30, 27, 22, 52, 
    34, 38, 30, 15, 8, 10, 21, 20, 10, 5, 4, 2, 2, 1, 4, 4, 6, 20, 0, 0, 27, 32, 48, 36, 32, 29, 32, 31, 30, 27, 24, 50, 
    29, 33, 36, 30, 26, 23, 33, 44, 31, 25, 28, 29, 31, 30, 30, 31, 30, 32, 16, 0, 10, 33, 37, 39, 35, 33, 33, 32, 30, 26, 29, 51, 
    25, 26, 26, 28, 34, 28, 31, 44, 31, 25, 26, 26, 32, 33, 33, 35, 35, 38, 32, 16, 12, 28, 33, 34, 34, 34, 34, 31, 31, 28, 29, 51, 
    10, 16, 14, 12, 15, 17, 19, 30, 26, 20, 19, 19, 21, 25, 26, 29, 31, 33, 33, 27, 25, 34, 36, 33, 32, 32, 33, 31, 27, 26, 26, 43, 
    
    -- channel=103
    73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 12, 0, 0, 0, 
    91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 41, 25, 0, 0, 0, 
    88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 21, 53, 30, 0, 0, 0, 
    88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 25, 44, 19, 0, 0, 0, 
    94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 8, 29, 36, 1, 0, 0, 0, 
    93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 16, 9, 23, 17, 0, 0, 0, 0, 
    84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 35, 59, 4, 0, 0, 0, 0, 0, 0, 
    73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 65, 0, 0, 0, 0, 0, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 45, 42, 0, 0, 0, 0, 0, 0, 0, 
    73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 40, 0, 0, 0, 0, 0, 0, 0, 
    73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 25, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 44, 36, 13, 0, 0, 0, 0, 0, 
    72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 19, 26, 0, 0, 7, 6, 14, 18, 45, 70, 0, 0, 11, 59, 70, 0, 0, 0, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 12, 34, 36, 4, 19, 47, 41, 33, 78, 159, 133, 0, 0, 0, 46, 95, 43, 0, 0, 0, 0, 
    74, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 27, 48, 37, 0, 15, 54, 61, 37, 118, 207, 125, 0, 0, 0, 0, 80, 73, 11, 10, 5, 0, 
    78, 0, 0, 0, 0, 0, 0, 0, 8, 19, 18, 27, 46, 20, 0, 18, 54, 91, 72, 124, 154, 71, 13, 0, 0, 0, 37, 59, 61, 52, 6, 0, 
    79, 0, 0, 0, 0, 0, 10, 0, 21, 11, 8, 38, 52, 26, 41, 72, 60, 76, 60, 79, 64, 30, 0, 0, 0, 0, 0, 46, 105, 88, 0, 0, 
    80, 0, 0, 0, 0, 4, 41, 30, 27, 15, 0, 51, 54, 55, 125, 102, 22, 28, 32, 29, 14, 0, 0, 0, 0, 34, 0, 54, 120, 87, 0, 0, 
    79, 0, 0, 0, 4, 0, 44, 57, 47, 16, 7, 65, 71, 77, 194, 122, 10, 19, 24, 24, 18, 0, 0, 0, 3, 65, 38, 52, 89, 60, 0, 0, 
    77, 0, 1, 41, 11, 0, 15, 69, 59, 0, 28, 70, 85, 94, 212, 108, 9, 27, 35, 30, 25, 11, 0, 0, 1, 56, 48, 46, 46, 29, 0, 0, 
    73, 0, 57, 89, 0, 0, 0, 66, 50, 0, 42, 70, 99, 125, 202, 81, 17, 33, 18, 0, 14, 59, 39, 0, 0, 37, 36, 30, 19, 3, 0, 0, 
    73, 2, 99, 99, 0, 0, 0, 51, 34, 0, 55, 78, 104, 145, 200, 65, 25, 24, 0, 0, 35, 90, 131, 101, 30, 7, 9, 20, 1, 0, 0, 0, 
    76, 17, 90, 60, 45, 0, 0, 36, 13, 19, 76, 100, 97, 124, 178, 56, 25, 0, 0, 0, 56, 71, 118, 178, 92, 8, 10, 10, 0, 0, 0, 23, 
    76, 29, 59, 30, 114, 68, 0, 12, 8, 42, 86, 115, 87, 113, 151, 44, 17, 0, 0, 17, 50, 47, 72, 160, 157, 40, 9, 0, 0, 0, 38, 36, 
    73, 25, 31, 29, 116, 101, 0, 0, 24, 66, 94, 116, 89, 128, 124, 28, 8, 0, 0, 64, 42, 33, 42, 103, 176, 86, 6, 0, 0, 31, 52, 28, 
    71, 22, 40, 50, 93, 108, 0, 0, 46, 89, 101, 92, 74, 134, 97, 30, 9, 0, 0, 76, 40, 22, 26, 59, 157, 126, 2, 0, 0, 50, 49, 25, 
    72, 30, 55, 62, 83, 109, 0, 0, 72, 108, 104, 73, 56, 101, 65, 31, 6, 0, 0, 89, 69, 10, 0, 29, 115, 139, 8, 0, 15, 55, 49, 32, 
    75, 32, 56, 69, 76, 94, 3, 0, 71, 92, 86, 61, 46, 61, 44, 34, 20, 0, 0, 85, 68, 18, 0, 23, 69, 113, 26, 0, 39, 55, 55, 42, 
    79, 27, 36, 59, 59, 70, 18, 28, 77, 87, 89, 78, 68, 70, 63, 58, 49, 6, 14, 109, 58, 35, 6, 11, 46, 81, 43, 34, 53, 57, 61, 49, 
    87, 23, 23, 34, 46, 59, 44, 50, 63, 71, 75, 72, 72, 72, 68, 64, 61, 46, 49, 113, 69, 28, 9, 0, 40, 58, 50, 50, 55, 59, 63, 47, 
    93, 24, 21, 28, 46, 53, 54, 40, 28, 52, 63, 57, 55, 51, 50, 49, 47, 46, 55, 86, 76, 42, 17, 15, 45, 51, 51, 52, 55, 60, 62, 40, 
    101, 32, 39, 48, 53, 47, 48, 31, 21, 57, 66, 58, 55, 46, 45, 43, 39, 38, 43, 65, 80, 51, 20, 35, 51, 51, 50, 51, 56, 59, 57, 32, 
    84, 41, 52, 61, 63, 56, 53, 41, 34, 62, 66, 60, 58, 51, 49, 48, 45, 43, 43, 52, 61, 50, 35, 45, 51, 52, 51, 50, 54, 56, 52, 40, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 13, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 3, 2, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 16, 10, 6, 4, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 7, 5, 11, 13, 10, 8, 3, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 6, 9, 9, 10, 10, 8, 6, 1, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 6, 5, 6, 4, 1, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 7, 8, 7, 7, 6, 3, 0, 0, 16, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 70, 91, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 39, 64, 104, 142, 152, 102, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 65, 62, 54, 52, 64, 100, 147, 191, 158, 62, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 55, 64, 42, 21, 9, 29, 75, 139, 211, 206, 123, 51, 16, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 39, 46, 21, 7, 16, 50, 103, 179, 230, 229, 177, 95, 32, 11, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 42, 66, 64, 66, 91, 120, 163, 219, 235, 211, 170, 99, 15, 0, 5, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 32, 27, 11, 22, 64, 98, 124, 140, 154, 176, 206, 222, 206, 162, 100, 28, 0, 0, 15, 61, 72, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 51, 59, 64, 40, 35, 45, 84, 126, 177, 197, 203, 212, 217, 214, 187, 127, 41, 0, 0, 16, 57, 104, 120, 32, 0, 
    0, 0, 0, 0, 0, 14, 55, 73, 68, 55, 30, 41, 63, 97, 155, 211, 223, 225, 223, 218, 212, 200, 137, 65, 39, 62, 97, 120, 139, 131, 61, 4, 
    0, 0, 0, 0, 53, 91, 88, 76, 60, 35, 16, 30, 72, 116, 178, 223, 233, 230, 214, 196, 180, 185, 174, 146, 140, 159, 175, 172, 155, 119, 62, 6, 
    0, 0, 0, 51, 148, 133, 105, 70, 50, 19, 8, 30, 79, 136, 194, 227, 233, 216, 187, 149, 116, 128, 174, 192, 205, 212, 202, 180, 142, 95, 33, 0, 
    0, 0, 0, 105, 165, 143, 114, 66, 40, 11, 23, 58, 104, 153, 204, 229, 224, 190, 154, 93, 62, 67, 118, 176, 204, 210, 194, 159, 114, 59, 0, 0, 
    0, 0, 0, 86, 149, 147, 115, 64, 29, 16, 48, 91, 136, 171, 212, 233, 212, 172, 114, 50, 43, 41, 56, 126, 175, 195, 177, 133, 81, 16, 0, 0, 
    0, 0, 0, 58, 132, 149, 117, 65, 32, 36, 72, 119, 162, 185, 219, 233, 205, 159, 85, 47, 48, 44, 37, 76, 143, 172, 160, 116, 44, 0, 0, 0, 
    0, 0, 0, 60, 126, 150, 121, 68, 46, 67, 104, 142, 167, 186, 222, 228, 203, 149, 82, 64, 58, 52, 40, 45, 107, 148, 144, 92, 13, 0, 0, 0, 
    0, 0, 0, 68, 125, 157, 135, 96, 87, 121, 157, 180, 184, 204, 225, 226, 205, 149, 92, 82, 85, 74, 53, 33, 72, 114, 115, 64, 0, 0, 0, 0, 
    0, 0, 0, 55, 115, 153, 140, 113, 115, 145, 170, 180, 178, 188, 196, 195, 182, 137, 91, 84, 98, 81, 57, 28, 38, 70, 71, 32, 0, 0, 0, 0, 
    0, 0, 0, 24, 77, 110, 105, 89, 93, 112, 123, 129, 128, 132, 134, 133, 125, 97, 70, 69, 88, 85, 52, 28, 14, 29, 28, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 40, 67, 64, 58, 62, 67, 68, 69, 69, 73, 71, 66, 57, 45, 33, 55, 68, 67, 42, 17, 1, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 74, 74, 68, 65, 63, 63, 63, 58, 53, 44, 38, 26, 16, 11, 38, 56, 49, 36, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 101, 127, 130, 122, 111, 106, 110, 109, 99, 87, 75, 66, 53, 41, 36, 45, 63, 60, 38, 11, 5, 5, 6, 6, 7, 10, 8, 4, 
    0, 0, 0, 48, 87, 105, 108, 101, 87, 83, 88, 88, 80, 70, 61, 56, 47, 38, 34, 36, 42, 37, 19, 6, 3, 4, 6, 5, 5, 5, 4, 1, 
    
    -- channel=106
    47, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    104, 23, 12, 5, 15, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    101, 8, 3, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    91, 7, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    85, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 42, 25, 0, 0, 0, 0, 19, 6, 0, 0, 0, 
    62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 55, 24, 9, 1, 0, 17, 17, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 44, 25, 0, 16, 21, 3, 10, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 8, 12, 7, 21, 22, 0, 0, 16, 25, 2, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 25, 22, 15, 8, 15, 19, 23, 11, 0, 0, 23, 27, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 33, 42, 45, 59, 84, 119, 141, 103, 61, 33, 9, 33, 38, 3, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 42, 101, 146, 162, 182, 199, 221, 231, 193, 186, 158, 43, 9, 21, 32, 15, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 11, 60, 106, 159, 182, 176, 180, 187, 191, 187, 180, 261, 268, 97, 0, 0, 29, 51, 3, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 8, 51, 78, 111, 162, 160, 120, 111, 118, 102, 86, 165, 327, 356, 178, 2, 0, 15, 60, 18, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 33, 63, 78, 103, 125, 94, 40, 15, 33, 20, 33, 193, 371, 392, 273, 85, 0, 0, 37, 18, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 26, 45, 65, 59, 74, 88, 43, 0, 0, 33, 73, 137, 284, 391, 387, 329, 156, 9, 0, 2, 7, 25, 30, 0, 0, 
    28, 0, 0, 0, 0, 30, 51, 60, 82, 52, 42, 74, 85, 69, 100, 141, 195, 239, 290, 371, 396, 378, 297, 129, 25, 0, 0, 15, 104, 117, 19, 0, 
    29, 0, 0, 0, 0, 34, 69, 85, 78, 42, 33, 59, 48, 109, 235, 287, 308, 343, 379, 390, 381, 323, 190, 51, 13, 6, 0, 80, 190, 204, 50, 0, 
    28, 0, 0, 25, 29, 44, 70, 82, 70, 26, 9, 49, 46, 162, 342, 387, 371, 376, 383, 382, 384, 315, 130, 13, 57, 92, 100, 168, 245, 248, 76, 0, 
    25, 0, 44, 125, 83, 25, 40, 79, 47, 0, 0, 35, 57, 213, 390, 388, 354, 360, 367, 367, 374, 324, 180, 112, 152, 185, 202, 235, 254, 238, 80, 0, 
    18, 18, 157, 236, 149, 35, 32, 65, 9, 0, 0, 17, 64, 234, 373, 354, 334, 341, 301, 251, 253, 286, 266, 230, 245, 267, 268, 255, 233, 182, 44, 0, 
    18, 63, 216, 276, 174, 47, 32, 40, 0, 0, 0, 24, 80, 250, 360, 336, 333, 293, 181, 114, 123, 186, 273, 304, 298, 274, 255, 236, 173, 84, 0, 0, 
    26, 71, 159, 188, 168, 74, 37, 20, 0, 0, 9, 70, 123, 272, 356, 331, 322, 208, 67, 22, 46, 85, 189, 292, 284, 245, 226, 171, 83, 0, 0, 0, 
    31, 57, 80, 103, 180, 111, 32, 0, 0, 0, 48, 108, 156, 296, 361, 340, 299, 120, 0, 0, 9, 14, 88, 228, 266, 227, 185, 100, 3, 0, 0, 0, 
    23, 23, 20, 64, 187, 140, 32, 0, 0, 15, 91, 143, 200, 315, 355, 336, 263, 60, 0, 39, 27, 0, 13, 137, 235, 220, 148, 30, 0, 0, 0, 0, 
    8, 2, 26, 69, 178, 151, 23, 0, 10, 69, 135, 158, 218, 322, 339, 324, 235, 42, 17, 61, 37, 14, 0, 63, 194, 206, 97, 0, 0, 0, 0, 0, 
    0, 0, 43, 73, 163, 163, 50, 27, 90, 166, 220, 230, 278, 342, 337, 326, 232, 49, 30, 101, 95, 39, 0, 15, 135, 159, 40, 0, 0, 0, 0, 0, 
    0, 0, 47, 76, 146, 145, 57, 46, 100, 156, 191, 197, 224, 250, 243, 242, 180, 38, 36, 94, 91, 33, 0, 0, 50, 67, 0, 0, 0, 0, 0, 0, 
    10, 0, 23, 49, 86, 79, 19, 17, 56, 89, 109, 111, 115, 122, 121, 118, 79, 0, 33, 101, 87, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 4, 14, 17, 30, 28, 7, 5, 12, 23, 30, 32, 34, 35, 29, 24, 11, 0, 10, 71, 74, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 11, 10, 19, 30, 37, 35, 11, 0, 1, 8, 9, 7, 2, 0, 0, 0, 0, 1, 35, 31, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 32, 46, 70, 84, 92, 86, 46, 28, 41, 49, 50, 47, 41, 34, 24, 11, 0, 1, 32, 47, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 31, 36, 29, 0, 0, 0, 5, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    33, 39, 50, 55, 56, 61, 64, 64, 68, 71, 72, 72, 70, 70, 73, 73, 71, 66, 67, 98, 71, 71, 70, 63, 58, 66, 77, 71, 66, 63, 63, 73, 
    0, 24, 32, 34, 31, 35, 40, 39, 42, 45, 46, 45, 41, 42, 48, 49, 47, 39, 42, 52, 47, 51, 49, 42, 57, 65, 60, 54, 49, 49, 51, 74, 
    0, 36, 39, 34, 33, 38, 44, 43, 45, 46, 48, 46, 43, 43, 47, 48, 48, 44, 52, 49, 42, 49, 46, 36, 61, 72, 53, 36, 40, 49, 51, 75, 
    0, 33, 36, 36, 45, 42, 46, 46, 45, 47, 50, 48, 45, 45, 47, 48, 48, 45, 49, 51, 38, 32, 40, 48, 65, 68, 50, 31, 35, 47, 50, 76, 
    0, 37, 48, 52, 57, 48, 49, 49, 47, 47, 48, 46, 45, 46, 45, 46, 45, 42, 43, 44, 21, 19, 46, 56, 57, 56, 40, 29, 27, 45, 50, 76, 
    16, 53, 52, 51, 51, 47, 49, 49, 47, 44, 45, 45, 42, 42, 41, 43, 42, 42, 45, 36, 15, 44, 69, 65, 54, 39, 31, 34, 39, 53, 52, 76, 
    21, 51, 49, 46, 45, 42, 45, 46, 46, 42, 43, 44, 42, 42, 38, 41, 39, 38, 39, 23, 23, 71, 77, 53, 53, 41, 36, 44, 49, 55, 52, 77, 
    24, 47, 46, 44, 46, 43, 45, 44, 44, 41, 41, 41, 36, 38, 31, 31, 28, 31, 36, 25, 44, 82, 67, 36, 43, 44, 40, 45, 47, 52, 51, 77, 
    27, 45, 46, 44, 47, 45, 46, 45, 44, 40, 35, 29, 20, 31, 33, 41, 42, 40, 41, 36, 56, 67, 47, 25, 31, 44, 49, 51, 47, 50, 51, 77, 
    28, 44, 46, 44, 47, 44, 46, 46, 44, 39, 34, 39, 33, 40, 31, 25, 8, 0, 0, 0, 18, 42, 47, 30, 30, 41, 48, 52, 48, 49, 52, 78, 
    27, 43, 46, 43, 46, 44, 45, 45, 43, 38, 34, 31, 0, 0, 0, 0, 0, 0, 0, 22, 0, 2, 36, 28, 46, 47, 42, 44, 47, 50, 52, 78, 
    26, 43, 46, 43, 45, 44, 44, 46, 41, 30, 9, 0, 0, 8, 29, 39, 51, 54, 67, 75, 17, 21, 59, 29, 37, 39, 49, 49, 45, 49, 52, 77, 
    24, 43, 46, 44, 45, 45, 45, 46, 28, 11, 16, 30, 32, 51, 67, 69, 61, 57, 57, 15, 0, 1, 66, 61, 41, 26, 35, 69, 56, 52, 52, 77, 
    23, 41, 45, 44, 45, 49, 47, 38, 17, 28, 46, 37, 26, 49, 56, 49, 40, 54, 33, 0, 0, 0, 32, 74, 52, 30, 24, 61, 62, 52, 53, 77, 
    25, 43, 46, 43, 41, 39, 32, 17, 29, 47, 46, 26, 26, 57, 67, 53, 19, 18, 0, 0, 0, 0, 0, 78, 80, 42, 33, 41, 37, 26, 37, 70, 
    25, 43, 46, 42, 34, 26, 31, 19, 31, 37, 42, 30, 39, 47, 11, 0, 0, 0, 0, 0, 0, 0, 13, 98, 101, 78, 54, 30, 0, 3, 40, 62, 
    25, 42, 45, 42, 40, 35, 52, 45, 39, 63, 47, 42, 62, 30, 0, 0, 0, 0, 0, 0, 0, 6, 74, 96, 64, 75, 45, 0, 0, 0, 64, 65, 
    26, 44, 40, 23, 27, 24, 29, 36, 55, 75, 54, 33, 41, 0, 0, 0, 0, 0, 0, 0, 0, 16, 60, 50, 11, 7, 3, 0, 0, 2, 84, 79, 
    26, 42, 11, 0, 27, 47, 42, 31, 61, 70, 62, 35, 39, 0, 0, 0, 0, 0, 0, 0, 0, 14, 39, 2, 0, 0, 0, 0, 0, 4, 91, 95, 
    28, 19, 0, 0, 44, 60, 39, 31, 72, 68, 57, 41, 46, 0, 0, 0, 0, 0, 11, 41, 47, 43, 51, 15, 0, 0, 0, 1, 9, 33, 98, 100, 
    27, 0, 0, 17, 64, 76, 42, 41, 81, 67, 52, 30, 17, 0, 0, 0, 0, 11, 69, 72, 46, 25, 29, 28, 6, 4, 13, 20, 43, 82, 95, 86, 
    20, 0, 27, 58, 68, 85, 46, 55, 72, 60, 34, 10, 0, 0, 0, 0, 0, 57, 87, 57, 35, 13, 0, 12, 33, 31, 24, 44, 82, 91, 70, 73, 
    16, 15, 48, 19, 10, 68, 53, 69, 67, 49, 16, 19, 16, 0, 0, 0, 0, 88, 74, 59, 58, 53, 3, 0, 21, 25, 27, 67, 82, 68, 46, 67, 
    19, 36, 61, 24, 0, 54, 64, 64, 53, 34, 4, 15, 0, 0, 0, 0, 30, 99, 54, 41, 38, 51, 44, 0, 4, 24, 46, 84, 73, 53, 43, 73, 
    27, 42, 55, 41, 0, 48, 77, 64, 39, 20, 1, 7, 0, 0, 0, 0, 42, 92, 43, 38, 46, 49, 54, 9, 0, 33, 77, 92, 68, 53, 50, 79, 
    31, 39, 41, 37, 0, 38, 65, 34, 1, 0, 0, 0, 0, 0, 0, 0, 33, 83, 36, 22, 32, 40, 53, 31, 0, 43, 94, 89, 63, 53, 49, 76, 
    33, 42, 35, 32, 3, 37, 71, 45, 27, 26, 37, 51, 38, 35, 45, 47, 80, 108, 41, 24, 52, 79, 73, 60, 22, 61, 99, 81, 60, 53, 49, 74, 
    34, 42, 39, 52, 40, 67, 88, 72, 59, 53, 56, 65, 67, 68, 70, 70, 90, 115, 51, 28, 32, 57, 63, 65, 44, 56, 74, 69, 59, 53, 46, 72, 
    32, 42, 39, 49, 53, 60, 57, 44, 41, 39, 38, 38, 40, 41, 45, 46, 53, 68, 40, 47, 46, 48, 76, 69, 59, 60, 62, 59, 56, 52, 44, 71, 
    34, 46, 49, 42, 33, 25, 27, 40, 44, 43, 43, 41, 42, 43, 46, 47, 49, 52, 34, 34, 65, 81, 84, 70, 59, 59, 59, 56, 53, 48, 46, 72, 
    31, 36, 33, 26, 21, 16, 29, 51, 43, 32, 32, 33, 35, 34, 35, 38, 41, 44, 39, 25, 28, 53, 61, 58, 54, 53, 54, 52, 49, 44, 48, 73, 
    63, 75, 79, 86, 95, 93, 92, 96, 82, 77, 78, 79, 82, 83, 84, 84, 84, 81, 76, 71, 74, 84, 76, 68, 67, 70, 69, 67, 67, 68, 70, 83, 
    
    -- channel=108
    37, 4, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 0, 0, 0, 11, 0, 12, 5, 0, 3, 12, 27, 26, 18, 17, 0, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 22, 7, 7, 0, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 19, 40, 25, 6, 5, 0, 
    52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 39, 22, 4, 4, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 23, 25, 11, 0, 2, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 16, 13, 2, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 12, 10, 5, 0, 0, 0, 0, 
    46, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 25, 5, 1, 0, 0, 0, 0, 0, 
    44, 6, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 37, 31, 7, 0, 0, 2, 2, 1, 0, 
    42, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 23, 6, 5, 2, 2, 3, 2, 0, 
    41, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 9, 7, 5, 3, 4, 3, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 19, 6, 4, 6, 6, 4, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 27, 19, 0, 10, 14, 7, 0, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 25, 5, 10, 23, 15, 0, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 21, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 16, 12, 15, 13, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 15, 10, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 15, 24, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 6, 18, 24, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    36, 0, 0, 0, 0, 0, 0, 0, 12, 21, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 9, 0, 0, 0, 0, 0, 0, 0, 16, 9, 
    36, 0, 0, 0, 0, 0, 0, 0, 13, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 0, 0, 0, 0, 0, 17, 24, 5, 
    36, 0, 0, 0, 0, 0, 0, 0, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 0, 0, 0, 0, 9, 27, 23, 2, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 21, 31, 24, 5, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 0, 0, 2, 27, 33, 28, 12, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 18, 9, 18, 30, 32, 29, 16, 
    29, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 18, 28, 31, 29, 32, 32, 30, 27, 16, 
    26, 0, 0, 0, 0, 0, 0, 2, 13, 18, 17, 15, 15, 15, 15, 16, 20, 22, 23, 18, 0, 0, 5, 17, 30, 32, 33, 33, 32, 29, 24, 16, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 1, 2, 3, 3, 5, 10, 14, 16, 15, 4, 0, 6, 20, 28, 28, 28, 29, 28, 24, 20, 14, 
    28, 9, 0, 0, 0, 0, 0, 0, 1, 7, 7, 6, 7, 8, 8, 10, 13, 17, 20, 20, 18, 17, 24, 32, 31, 29, 30, 31, 30, 27, 25, 21, 
    
    -- channel=109
    0, 35, 35, 36, 36, 38, 37, 34, 28, 23, 12, 4, 3, 3, 0, 0, 0, 0, 7, 28, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 102, 93, 89, 88, 88, 83, 76, 69, 62, 49, 40, 41, 41, 33, 21, 9, 17, 50, 65, 45, 10, 8, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    21, 91, 81, 81, 74, 70, 52, 44, 38, 32, 23, 17, 18, 18, 14, 4, 0, 0, 0, 1, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    11, 79, 76, 80, 66, 50, 24, 17, 13, 9, 5, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 16, 17, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 72, 70, 64, 43, 23, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 70, 96, 68, 5, 0, 0, 0, 14, 0, 0, 0, 
    0, 51, 45, 30, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 58, 114, 140, 90, 21, 7, 10, 27, 31, 7, 0, 0, 
    0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 10, 9, 18, 20, 23, 39, 81, 114, 106, 58, 29, 31, 31, 30, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 30, 50, 50, 57, 56, 57, 69, 80, 73, 25, 2, 13, 35, 24, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 20, 37, 64, 76, 91, 81, 80, 78, 81, 89, 87, 60, 10, 1, 12, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 34, 52, 92, 107, 133, 142, 171, 213, 256, 246, 220, 140, 72, 55, 32, 27, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 46, 91, 171, 238, 304, 336, 367, 417, 458, 452, 435, 351, 235, 127, 28, 47, 34, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 34, 96, 172, 270, 349, 398, 412, 428, 457, 475, 479, 528, 531, 423, 208, 28, 27, 61, 50, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 76, 146, 226, 316, 369, 378, 345, 321, 301, 289, 342, 501, 660, 604, 315, 67, 0, 44, 57, 31, 0, 0, 0, 
    0, 0, 0, 5, 4, 0, 0, 11, 56, 115, 190, 239, 275, 273, 218, 125, 87, 56, 82, 214, 469, 724, 733, 473, 186, 14, 0, 31, 20, 0, 0, 0, 
    0, 4, 2, 7, 9, 21, 30, 62, 92, 156, 167, 177, 183, 163, 97, 11, 12, 52, 161, 344, 597, 782, 789, 590, 327, 73, 0, 0, 22, 22, 1, 0, 
    0, 8, 5, 11, 19, 61, 97, 138, 171, 154, 141, 134, 155, 175, 185, 194, 274, 352, 472, 628, 767, 827, 761, 578, 335, 90, 0, 0, 70, 147, 120, 0, 
    0, 9, 7, 13, 20, 73, 130, 182, 185, 155, 126, 101, 107, 190, 298, 444, 582, 652, 747, 818, 849, 797, 660, 428, 205, 83, 48, 80, 208, 342, 266, 73, 
    0, 6, 12, 53, 68, 123, 145, 172, 174, 144, 81, 66, 75, 220, 425, 680, 816, 835, 856, 861, 865, 795, 586, 311, 151, 138, 184, 258, 386, 491, 363, 134, 
    0, 7, 67, 159, 196, 191, 123, 129, 124, 81, 5, 19, 61, 263, 509, 753, 831, 817, 815, 822, 837, 784, 607, 408, 295, 309, 380, 451, 509, 532, 381, 147, 
    0, 39, 176, 340, 411, 298, 152, 108, 67, 22, 0, 0, 61, 288, 520, 726, 774, 759, 725, 684, 642, 642, 627, 578, 532, 537, 567, 571, 548, 483, 324, 90, 
    0, 76, 260, 494, 527, 346, 186, 85, 32, 0, 0, 0, 68, 305, 524, 710, 751, 698, 605, 466, 348, 386, 515, 614, 672, 656, 616, 567, 483, 366, 190, 0, 
    0, 86, 249, 438, 441, 322, 219, 80, 8, 0, 0, 23, 139, 360, 551, 709, 728, 611, 449, 212, 110, 144, 289, 474, 605, 632, 573, 477, 363, 195, 39, 0, 
    0, 74, 173, 269, 318, 295, 233, 73, 0, 0, 0, 97, 241, 436, 595, 733, 708, 523, 292, 56, 19, 23, 100, 295, 465, 551, 498, 371, 213, 38, 0, 0, 
    0, 34, 80, 141, 253, 283, 244, 77, 0, 0, 70, 188, 340, 494, 643, 747, 674, 447, 220, 56, 58, 28, 24, 149, 322, 454, 433, 276, 87, 0, 0, 0, 
    0, 0, 59, 130, 256, 288, 239, 80, 0, 43, 160, 258, 380, 518, 662, 732, 636, 407, 204, 81, 88, 64, 13, 65, 219, 365, 361, 189, 11, 0, 0, 0, 
    0, 0, 64, 139, 255, 298, 256, 142, 102, 198, 330, 417, 509, 608, 695, 726, 625, 403, 216, 134, 169, 143, 63, 26, 137, 249, 248, 99, 0, 0, 0, 0, 
    0, 0, 62, 132, 246, 280, 250, 167, 152, 246, 353, 423, 482, 528, 565, 579, 514, 337, 200, 134, 187, 153, 75, 0, 37, 93, 90, 0, 0, 0, 0, 0, 
    0, 0, 41, 97, 169, 189, 158, 104, 105, 171, 235, 277, 302, 318, 328, 330, 288, 174, 123, 121, 188, 168, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 38, 59, 83, 80, 56, 25, 20, 32, 48, 63, 73, 81, 81, 76, 58, 10, 14, 65, 134, 119, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 41, 50, 56, 57, 47, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 59, 65, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 61, 85, 120, 146, 165, 163, 128, 88, 56, 64, 77, 75, 67, 54, 37, 16, 0, 0, 9, 48, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 50, 92, 117, 114, 78, 35, 14, 24, 34, 32, 24, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 10, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 103, 114, 126, 135, 139, 146, 151, 146, 140, 131, 123, 120, 118, 113, 106, 99, 89, 94, 109, 84, 74, 75, 48, 27, 18, 41, 36, 25, 28, 33, 2, 
    64, 133, 136, 142, 137, 130, 127, 123, 116, 108, 101, 95, 94, 93, 92, 86, 81, 72, 63, 64, 66, 58, 56, 49, 32, 28, 35, 35, 26, 28, 32, 0, 
    79, 138, 127, 117, 105, 106, 98, 91, 85, 78, 73, 70, 69, 69, 71, 68, 66, 59, 54, 49, 62, 70, 52, 38, 35, 18, 13, 21, 24, 30, 30, 0, 
    63, 105, 85, 80, 81, 80, 71, 65, 63, 61, 59, 56, 54, 54, 58, 58, 58, 54, 57, 53, 63, 57, 29, 38, 34, 16, 23, 25, 37, 33, 29, 0, 
    38, 76, 77, 77, 72, 60, 51, 50, 51, 52, 49, 45, 44, 47, 53, 54, 53, 50, 52, 53, 49, 21, 19, 25, 20, 32, 31, 26, 33, 29, 33, 0, 
    45, 71, 61, 53, 47, 47, 43, 44, 44, 45, 43, 38, 38, 39, 48, 52, 57, 58, 62, 60, 48, 38, 46, 40, 21, 30, 31, 41, 45, 42, 40, 0, 
    30, 43, 37, 35, 33, 37, 35, 37, 39, 40, 40, 40, 46, 47, 55, 61, 66, 61, 58, 54, 44, 44, 44, 44, 31, 28, 44, 53, 51, 41, 38, 2, 
    14, 27, 26, 29, 30, 32, 30, 33, 36, 38, 45, 52, 59, 51, 46, 42, 50, 54, 59, 53, 44, 45, 31, 34, 30, 33, 39, 42, 43, 38, 34, 1, 
    10, 26, 25, 29, 29, 32, 30, 31, 35, 37, 40, 36, 48, 58, 67, 78, 103, 123, 126, 95, 68, 34, 2, 17, 32, 40, 41, 36, 41, 37, 30, 0, 
    9, 26, 25, 29, 30, 32, 31, 33, 37, 36, 41, 60, 106, 122, 125, 114, 93, 63, 32, 14, 62, 56, 26, 32, 20, 36, 45, 36, 35, 34, 28, 0, 
    10, 28, 25, 29, 29, 32, 33, 35, 37, 45, 71, 84, 65, 22, 0, 0, 0, 9, 19, 30, 49, 26, 16, 49, 47, 46, 20, 27, 31, 30, 26, 0, 
    11, 31, 27, 28, 28, 31, 34, 34, 48, 55, 32, 5, 15, 42, 61, 81, 105, 112, 119, 140, 130, 73, 36, 20, 30, 41, 34, 4, 20, 21, 22, 0, 
    11, 33, 29, 29, 27, 26, 33, 38, 45, 18, 19, 64, 93, 87, 91, 88, 76, 53, 70, 105, 98, 99, 73, 17, 18, 23, 36, 18, 18, 21, 20, 0, 
    10, 32, 29, 30, 31, 40, 49, 42, 22, 34, 72, 74, 48, 26, 17, 14, 35, 42, 75, 75, 65, 105, 94, 13, 0, 17, 17, 34, 39, 43, 32, 0, 
    11, 32, 27, 31, 36, 42, 27, 27, 41, 67, 37, 25, 20, 39, 70, 85, 105, 97, 60, 45, 93, 112, 72, 16, 4, 0, 0, 26, 53, 33, 15, 0, 
    11, 30, 27, 29, 27, 27, 11, 23, 40, 1, 25, 30, 23, 49, 59, 16, 1, 6, 34, 82, 111, 80, 46, 77, 60, 0, 13, 47, 39, 19, 4, 1, 
    7, 25, 28, 45, 48, 62, 68, 48, 17, 18, 42, 56, 60, 88, 50, 37, 77, 98, 121, 127, 120, 107, 116, 93, 52, 44, 26, 22, 24, 48, 13, 0, 
    6, 27, 56, 72, 26, 21, 22, 27, 22, 32, 15, 27, 19, 67, 85, 113, 133, 138, 132, 111, 107, 98, 69, 48, 35, 16, 0, 12, 57, 75, 21, 0, 
    4, 41, 80, 42, 9, 27, 24, 19, 5, 12, 7, 6, 0, 49, 81, 103, 109, 102, 68, 50, 60, 59, 25, 18, 23, 30, 55, 66, 67, 54, 30, 11, 
    5, 44, 33, 10, 41, 23, 14, 4, 0, 9, 7, 25, 45, 77, 74, 90, 99, 69, 43, 87, 117, 108, 78, 50, 55, 62, 60, 60, 44, 30, 50, 20, 
    6, 27, 13, 59, 60, 16, 18, 4, 12, 10, 18, 33, 40, 77, 75, 93, 95, 49, 73, 91, 68, 84, 111, 76, 55, 58, 71, 55, 34, 57, 53, 1, 
    4, 22, 64, 125, 84, 25, 17, 0, 8, 7, 16, 0, 0, 54, 84, 100, 87, 50, 68, 6, 0, 5, 58, 92, 75, 82, 67, 39, 57, 49, 23, 0, 
    3, 19, 32, 33, 49, 18, 12, 14, 13, 13, 21, 18, 56, 80, 69, 85, 67, 44, 42, 13, 29, 15, 8, 62, 65, 53, 35, 29, 33, 10, 6, 0, 
    3, 17, 10, 2, 42, 22, 7, 8, 11, 15, 26, 41, 67, 61, 75, 96, 75, 42, 31, 9, 2, 4, 6, 34, 56, 35, 20, 19, 9, 1, 11, 0, 
    5, 15, 18, 19, 43, 33, 25, 34, 39, 47, 52, 58, 77, 92, 112, 112, 76, 33, 31, 23, 20, 17, 2, 14, 49, 38, 23, 17, 7, 10, 20, 2, 
    3, 6, 15, 20, 37, 25, 0, 0, 0, 0, 0, 0, 0, 16, 26, 28, 18, 4, 28, 15, 0, 0, 0, 0, 31, 25, 19, 14, 4, 6, 12, 0, 
    4, 10, 7, 0, 9, 4, 2, 0, 4, 29, 50, 58, 61, 65, 68, 69, 53, 14, 21, 23, 45, 34, 22, 3, 22, 39, 31, 7, 0, 4, 10, 0, 
    8, 10, 15, 24, 29, 45, 55, 50, 52, 61, 69, 75, 79, 80, 78, 73, 69, 45, 26, 3, 19, 20, 0, 2, 6, 10, 6, 2, 3, 6, 12, 0, 
    4, 7, 7, 25, 43, 47, 26, 2, 0, 2, 3, 5, 7, 8, 8, 7, 9, 9, 20, 30, 0, 0, 0, 8, 3, 1, 0, 4, 7, 11, 11, 0, 
    13, 22, 23, 21, 11, 1, 0, 0, 2, 7, 4, 4, 6, 9, 11, 7, 6, 5, 11, 31, 44, 37, 22, 6, 4, 6, 4, 5, 8, 12, 12, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    112, 174, 178, 183, 185, 186, 189, 190, 187, 185, 184, 180, 177, 173, 170, 169, 165, 161, 144, 116, 117, 128, 125, 116, 113, 83, 63, 74, 87, 105, 115, 88, 
    191, 248, 251, 250, 253, 256, 256, 258, 255, 248, 240, 234, 231, 228, 221, 213, 209, 199, 170, 176, 137, 153, 158, 142, 105, 73, 66, 75, 111, 134, 147, 103, 
    216, 260, 251, 242, 243, 247, 249, 248, 247, 237, 228, 221, 218, 216, 211, 202, 197, 192, 175, 166, 170, 161, 154, 133, 85, 50, 49, 89, 126, 146, 154, 107, 
    219, 242, 232, 222, 223, 233, 235, 232, 229, 219, 210, 204, 203, 202, 198, 190, 184, 180, 175, 165, 167, 154, 124, 95, 77, 52, 66, 108, 139, 153, 153, 108, 
    196, 213, 204, 204, 211, 212, 217, 213, 209, 201, 194, 189, 190, 190, 187, 181, 177, 174, 175, 169, 154, 123, 70, 54, 58, 62, 89, 114, 143, 147, 147, 106, 
    173, 184, 189, 188, 193, 193, 197, 194, 191, 189, 185, 182, 185, 185, 182, 177, 176, 173, 173, 169, 140, 82, 37, 22, 42, 75, 98, 126, 143, 148, 149, 104, 
    163, 175, 178, 180, 182, 187, 184, 183, 182, 184, 184, 183, 186, 186, 183, 177, 173, 169, 166, 156, 111, 57, 13, 30, 58, 89, 119, 148, 148, 152, 150, 105, 
    153, 171, 177, 181, 180, 182, 179, 180, 182, 183, 186, 183, 181, 176, 172, 170, 165, 160, 158, 139, 92, 41, 10, 50, 96, 118, 153, 159, 157, 156, 155, 109, 
    145, 173, 178, 183, 182, 183, 180, 181, 183, 184, 185, 177, 167, 159, 154, 161, 158, 154, 148, 118, 71, 29, 11, 61, 110, 143, 157, 160, 161, 159, 155, 108, 
    144, 176, 181, 185, 184, 185, 183, 181, 183, 182, 180, 161, 143, 139, 130, 131, 119, 107, 84, 48, 17, 0, 0, 52, 98, 117, 132, 144, 154, 155, 151, 106, 
    147, 180, 184, 185, 183, 183, 182, 181, 180, 179, 168, 144, 113, 84, 59, 52, 35, 20, 2, 0, 0, 0, 0, 26, 70, 78, 95, 119, 141, 152, 149, 104, 
    152, 185, 185, 184, 182, 180, 180, 177, 175, 164, 143, 109, 59, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 61, 58, 88, 118, 143, 145, 103, 
    155, 186, 184, 182, 182, 178, 178, 171, 164, 143, 96, 54, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 48, 69, 50, 85, 122, 137, 101, 
    156, 185, 182, 181, 182, 175, 174, 162, 145, 99, 61, 43, 15, 0, 0, 0, 14, 13, 13, 9, 0, 0, 0, 0, 0, 22, 63, 56, 53, 95, 119, 93, 
    154, 182, 182, 181, 179, 162, 151, 133, 96, 61, 41, 24, 11, 1, 0, 9, 37, 30, 6, 0, 0, 0, 0, 0, 0, 2, 34, 58, 43, 63, 88, 74, 
    154, 181, 183, 176, 166, 139, 100, 76, 48, 32, 4, 19, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 49, 43, 24, 41, 55, 
    155, 180, 182, 167, 140, 104, 63, 22, 18, 0, 11, 19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 37, 39, 13, 0, 0, 20, 
    155, 179, 177, 150, 101, 52, 33, 1, 0, 0, 0, 16, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 57, 7, 0, 0, 0, 0, 0, 
    158, 176, 161, 111, 31, 0, 3, 6, 0, 2, 4, 27, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    157, 168, 136, 35, 0, 0, 0, 2, 4, 2, 30, 32, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    154, 156, 90, 0, 0, 0, 0, 2, 10, 16, 35, 30, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    152, 132, 62, 1, 0, 0, 0, 0, 19, 19, 36, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 16, 25, 
    144, 112, 65, 4, 0, 0, 0, 0, 16, 26, 34, 1, 0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 19, 22, 0, 0, 0, 0, 0, 4, 34, 50, 
    134, 113, 61, 0, 0, 0, 0, 0, 12, 23, 12, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 10, 1, 33, 0, 0, 0, 0, 0, 27, 60, 55, 
    125, 109, 52, 0, 0, 0, 0, 0, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 4, 15, 19, 27, 0, 0, 0, 1, 51, 69, 56, 
    115, 97, 54, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 13, 32, 0, 0, 0, 20, 58, 67, 53, 
    103, 90, 59, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 12, 32, 24, 0, 0, 35, 58, 60, 49, 
    94, 88, 66, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 0, 8, 26, 45, 23, 18, 43, 53, 54, 44, 
    92, 84, 62, 44, 7, 7, 0, 0, 6, 6, 4, 2, 0, 0, 0, 0, 7, 9, 8, 22, 0, 4, 0, 26, 34, 47, 40, 41, 46, 44, 45, 40, 
    86, 77, 53, 32, 11, 1, 0, 0, 5, 10, 11, 8, 9, 12, 17, 20, 24, 30, 27, 49, 11, 0, 20, 20, 38, 44, 43, 44, 43, 41, 38, 37, 
    80, 61, 40, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 16, 22, 21, 7, 6, 18, 35, 38, 36, 37, 37, 35, 33, 32, 
    70, 55, 40, 20, 2, 0, 0, 0, 0, 6, 11, 8, 9, 11, 15, 18, 20, 25, 28, 29, 30, 28, 29, 40, 43, 41, 41, 42, 42, 40, 41, 37, 
    
    -- channel=112
    117, 93, 95, 92, 93, 89, 91, 91, 90, 91, 103, 100, 97, 94, 95, 99, 100, 101, 101, 103, 102, 102, 105, 106, 108, 109, 110, 109, 115, 114, 117, 130, 
    52, 65, 72, 67, 65, 58, 55, 60, 68, 66, 79, 89, 82, 73, 72, 82, 84, 84, 80, 86, 88, 89, 95, 97, 102, 104, 104, 102, 111, 113, 114, 147, 
    52, 66, 73, 73, 64, 62, 63, 60, 84, 81, 70, 83, 94, 89, 80, 81, 82, 84, 82, 91, 96, 95, 102, 104, 108, 108, 106, 101, 107, 106, 101, 154, 
    53, 67, 71, 77, 60, 67, 94, 62, 77, 89, 75, 68, 88, 106, 97, 91, 92, 86, 88, 98, 104, 100, 105, 103, 101, 98, 94, 89, 92, 93, 90, 166, 
    52, 67, 69, 79, 62, 73, 115, 66, 64, 97, 101, 86, 85, 104, 110, 107, 112, 93, 90, 91, 97, 92, 88, 87, 85, 80, 80, 80, 83, 87, 90, 174, 
    55, 68, 67, 79, 74, 75, 95, 83, 87, 108, 112, 107, 100, 104, 115, 111, 110, 88, 79, 72, 71, 76, 73, 79, 80, 74, 76, 80, 85, 92, 98, 177, 
    60, 73, 69, 77, 89, 95, 87, 89, 110, 108, 110, 110, 115, 116, 117, 112, 98, 70, 63, 73, 69, 73, 71, 77, 83, 78, 79, 88, 95, 101, 105, 175, 
    63, 78, 75, 80, 105, 130, 108, 75, 107, 117, 118, 120, 121, 117, 105, 107, 113, 87, 66, 74, 76, 73, 81, 85, 87, 85, 85, 90, 96, 102, 106, 178, 
    68, 80, 77, 81, 89, 118, 119, 81, 108, 113, 111, 119, 111, 108, 106, 100, 117, 116, 92, 76, 77, 80, 98, 102, 81, 81, 88, 93, 98, 100, 102, 187, 
    70, 66, 56, 48, 35, 91, 131, 105, 111, 96, 78, 98, 94, 100, 115, 107, 110, 115, 115, 102, 91, 88, 92, 102, 84, 81, 92, 94, 95, 93, 92, 195, 
    45, 30, 21, 16, 11, 111, 145, 104, 117, 104, 62, 78, 78, 85, 120, 114, 109, 115, 118, 118, 110, 99, 89, 97, 87, 81, 88, 87, 86, 87, 90, 202, 
    10, 15, 13, 14, 15, 130, 160, 81, 109, 126, 73, 64, 84, 76, 112, 118, 104, 115, 116, 116, 119, 115, 96, 98, 89, 72, 82, 86, 85, 85, 87, 200, 
    0, 17, 20, 20, 21, 105, 175, 80, 69, 108, 83, 61, 99, 94, 93, 115, 96, 106, 112, 110, 112, 123, 106, 93, 98, 72, 72, 82, 80, 82, 86, 195, 
    0, 20, 27, 29, 29, 67, 159, 127, 56, 65, 68, 63, 92, 113, 100, 110, 90, 97, 109, 107, 106, 122, 115, 83, 98, 87, 64, 77, 81, 87, 94, 189, 
    3, 29, 33, 34, 33, 42, 98, 147, 104, 72, 60, 70, 95, 114, 111, 107, 89, 90, 102, 105, 106, 121, 121, 88, 88, 104, 72, 77, 91, 98, 102, 185, 
    14, 36, 35, 31, 27, 30, 41, 77, 128, 140, 102, 58, 91, 106, 97, 92, 79, 81, 92, 105, 110, 119, 121, 104, 82, 112, 94, 86, 99, 98, 94, 184, 
    17, 32, 28, 22, 24, 51, 63, 17, 93, 141, 112, 47, 61, 115, 96, 83, 73, 76, 90, 105, 115, 117, 117, 117, 85, 106, 110, 88, 90, 84, 87, 187, 
    11, 25, 25, 24, 29, 56, 102, 0, 9, 89, 71, 86, 34, 108, 111, 85, 80, 76, 87, 102, 110, 113, 111, 120, 95, 95, 105, 77, 86, 101, 116, 188, 
    11, 23, 16, 0, 0, 0, 69, 34, 0, 59, 56, 122, 26, 69, 126, 98, 83, 79, 83, 96, 102, 107, 112, 119, 105, 88, 105, 90, 106, 129, 134, 178, 
    0, 0, 0, 0, 0, 0, 0, 91, 0, 21, 27, 129, 67, 46, 122, 108, 86, 81, 83, 89, 95, 101, 112, 118, 111, 94, 119, 120, 119, 126, 118, 171, 
    0, 0, 0, 0, 0, 0, 0, 86, 77, 33, 16, 106, 110, 53, 99, 112, 92, 85, 86, 86, 89, 95, 111, 120, 117, 105, 124, 134, 113, 113, 114, 172, 
    0, 0, 0, 0, 77, 44, 22, 81, 86, 57, 53, 97, 110, 81, 88, 97, 94, 88, 87, 84, 89, 102, 117, 126, 121, 106, 104, 129, 120, 107, 116, 175, 
    0, 0, 0, 0, 122, 113, 65, 85, 71, 74, 97, 107, 103, 107, 105, 71, 79, 91, 92, 91, 99, 109, 113, 118, 117, 106, 86, 109, 134, 114, 111, 177, 
    0, 0, 0, 31, 93, 83, 48, 89, 116, 108, 111, 109, 93, 102, 128, 89, 73, 99, 101, 96, 96, 91, 96, 113, 121, 109, 87, 85, 130, 132, 110, 175, 
    0, 44, 58, 52, 46, 50, 56, 82, 127, 136, 116, 101, 73, 73, 120, 129, 88, 91, 96, 82, 80, 80, 84, 110, 134, 114, 91, 78, 105, 138, 122, 172, 
    14, 55, 50, 51, 59, 66, 70, 63, 73, 106, 115, 88, 60, 74, 107, 125, 96, 86, 90, 68, 68, 81, 80, 91, 126, 130, 102, 89, 80, 116, 138, 178, 
    34, 57, 65, 69, 73, 64, 59, 58, 64, 78, 101, 110, 89, 88, 98, 114, 105, 88, 86, 52, 49, 83, 96, 94, 103, 129, 118, 104, 83, 90, 134, 193, 
    53, 75, 72, 62, 60, 65, 74, 85, 100, 99, 93, 116, 116, 88, 83, 103, 115, 99, 92, 62, 50, 87, 109, 108, 103, 115, 120, 115, 103, 86, 108, 201, 
    63, 68, 64, 66, 76, 93, 107, 115, 120, 102, 81, 97, 118, 96, 92, 104, 119, 108, 106, 98, 76, 85, 102, 107, 108, 120, 124, 116, 112, 100, 92, 195, 
    57, 73, 84, 95, 107, 118, 124, 119, 115, 90, 78, 95, 108, 99, 110, 121, 124, 116, 112, 117, 104, 92, 96, 103, 117, 132, 127, 114, 113, 114, 98, 184, 
    66, 102, 115, 118, 117, 114, 118, 116, 116, 91, 82, 97, 100, 114, 118, 121, 125, 119, 113, 118, 118, 108, 110, 112, 118, 129, 126, 116, 113, 119, 114, 176, 
    78, 111, 114, 104, 102, 102, 106, 108, 111, 88, 73, 90, 83, 109, 115, 109, 114, 109, 103, 110, 115, 104, 108, 108, 103, 111, 117, 113, 106, 109, 112, 168, 
    
    -- channel=113
    4, 61, 58, 57, 54, 56, 60, 63, 65, 69, 69, 68, 62, 50, 44, 39, 36, 33, 30, 25, 21, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 103, 99, 96, 93, 95, 98, 102, 98, 108, 119, 121, 115, 104, 88, 78, 75, 68, 62, 55, 49, 39, 31, 23, 13, 7, 2, 1, 1, 3, 1, 0, 
    10, 104, 99, 96, 95, 93, 86, 87, 86, 111, 122, 124, 123, 116, 103, 86, 72, 61, 55, 51, 46, 38, 29, 28, 27, 28, 29, 31, 31, 31, 28, 0, 
    9, 100, 98, 94, 95, 87, 76, 82, 84, 103, 104, 104, 112, 112, 106, 93, 77, 66, 56, 58, 59, 60, 58, 61, 60, 60, 58, 59, 57, 55, 48, 5, 
    5, 95, 94, 91, 91, 80, 74, 77, 74, 88, 95, 95, 102, 110, 109, 99, 87, 83, 83, 93, 96, 93, 91, 88, 87, 84, 81, 79, 72, 62, 51, 4, 
    2, 88, 88, 86, 81, 66, 54, 50, 55, 85, 89, 89, 93, 98, 106, 111, 109, 104, 103, 112, 117, 112, 110, 108, 104, 94, 83, 76, 66, 56, 46, 2, 
    0, 82, 83, 81, 73, 48, 31, 36, 52, 74, 80, 82, 85, 91, 103, 112, 110, 111, 108, 114, 124, 128, 128, 116, 98, 87, 80, 76, 69, 60, 50, 4, 
    0, 83, 85, 88, 90, 78, 62, 50, 47, 79, 91, 98, 105, 109, 112, 116, 112, 111, 113, 117, 122, 128, 125, 115, 103, 87, 82, 78, 71, 64, 58, 11, 
    8, 103, 119, 136, 154, 144, 107, 61, 47, 80, 98, 111, 127, 131, 130, 126, 120, 121, 114, 113, 120, 127, 133, 127, 113, 97, 90, 87, 85, 84, 82, 26, 
    36, 159, 177, 193, 208, 181, 135, 74, 50, 77, 91, 106, 139, 148, 146, 139, 124, 127, 126, 120, 120, 127, 132, 130, 121, 110, 108, 108, 105, 100, 95, 34, 
    64, 201, 213, 224, 236, 202, 154, 88, 51, 75, 91, 109, 141, 155, 145, 144, 134, 130, 132, 131, 126, 126, 129, 126, 127, 119, 118, 119, 115, 111, 106, 41, 
    76, 226, 234, 239, 241, 211, 158, 95, 58, 86, 110, 129, 149, 159, 154, 146, 139, 135, 139, 134, 130, 125, 125, 125, 126, 128, 121, 123, 122, 115, 104, 38, 
    74, 229, 229, 227, 226, 212, 168, 105, 64, 77, 111, 136, 156, 161, 154, 144, 141, 136, 140, 135, 130, 124, 121, 125, 126, 127, 120, 117, 115, 103, 87, 26, 
    65, 214, 214, 214, 215, 213, 192, 144, 95, 82, 90, 100, 124, 143, 139, 136, 143, 143, 150, 146, 136, 126, 121, 122, 124, 123, 115, 102, 99, 86, 70, 17, 
    59, 205, 207, 211, 217, 223, 216, 191, 142, 102, 82, 85, 112, 144, 145, 139, 149, 158, 169, 159, 146, 132, 123, 119, 120, 118, 111, 89, 81, 74, 71, 23, 
    61, 208, 216, 225, 232, 228, 211, 199, 172, 148, 120, 122, 131, 144, 144, 137, 149, 162, 170, 165, 150, 136, 128, 118, 119, 114, 110, 92, 88, 90, 80, 22, 
    70, 223, 230, 236, 244, 246, 232, 238, 225, 237, 214, 151, 155, 150, 159, 148, 146, 163, 171, 168, 157, 143, 135, 124, 121, 113, 115, 107, 95, 83, 59, 0, 
    79, 238, 254, 278, 305, 331, 317, 297, 274, 257, 259, 202, 193, 162, 168, 154, 147, 158, 168, 168, 162, 152, 143, 131, 123, 117, 115, 106, 76, 54, 32, 0, 
    105, 299, 329, 355, 372, 383, 369, 334, 300, 271, 276, 222, 211, 160, 166, 167, 150, 156, 165, 169, 166, 161, 154, 142, 129, 118, 105, 87, 51, 32, 23, 0, 
    146, 370, 384, 388, 376, 366, 341, 315, 280, 239, 256, 217, 196, 156, 166, 170, 155, 158, 166, 170, 170, 167, 160, 146, 129, 115, 97, 75, 43, 20, 13, 0, 
    167, 399, 409, 409, 365, 314, 250, 232, 228, 200, 207, 184, 177, 150, 152, 161, 153, 159, 168, 170, 168, 163, 152, 137, 123, 110, 95, 75, 48, 24, 14, 0, 
    169, 420, 420, 400, 333, 267, 204, 197, 206, 168, 148, 143, 149, 138, 127, 128, 126, 148, 157, 157, 152, 146, 143, 141, 130, 112, 96, 79, 62, 42, 22, 0, 
    157, 392, 358, 315, 265, 234, 193, 176, 160, 129, 107, 111, 121, 120, 109, 104, 91, 103, 125, 132, 137, 147, 152, 144, 125, 99, 84, 83, 77, 58, 33, 0, 
    106, 285, 255, 241, 229, 209, 169, 152, 134, 115, 105, 94, 103, 113, 108, 86, 78, 97, 120, 134, 142, 151, 156, 149, 130, 102, 75, 76, 81, 73, 50, 0, 
    55, 217, 207, 190, 167, 148, 141, 146, 148, 133, 114, 112, 112, 115, 110, 96, 81, 87, 113, 135, 150, 167, 173, 161, 136, 108, 82, 68, 79, 80, 64, 3, 
    31, 160, 143, 134, 130, 135, 139, 138, 131, 123, 105, 88, 85, 86, 102, 108, 101, 99, 116, 143, 161, 177, 177, 161, 145, 117, 86, 68, 69, 78, 72, 15, 
    16, 114, 116, 125, 131, 131, 125, 115, 100, 88, 85, 82, 80, 84, 95, 102, 105, 103, 112, 131, 143, 158, 165, 154, 141, 124, 97, 64, 57, 67, 72, 21, 
    11, 112, 114, 115, 113, 107, 95, 78, 63, 61, 71, 80, 79, 75, 82, 96, 89, 83, 85, 93, 103, 122, 140, 142, 135, 116, 88, 57, 47, 52, 61, 16, 
    15, 107, 98, 88, 78, 71, 62, 52, 42, 44, 54, 72, 86, 83, 75, 70, 60, 56, 55, 59, 67, 84, 103, 109, 102, 86, 66, 45, 35, 36, 41, 1, 
    4, 76, 61, 50, 47, 47, 44, 37, 27, 32, 45, 67, 84, 81, 70, 57, 42, 36, 37, 43, 46, 50, 58, 65, 62, 55, 44, 30, 23, 24, 25, 0, 
    0, 37, 30, 30, 27, 27, 23, 21, 20, 28, 39, 58, 79, 71, 65, 48, 28, 26, 28, 30, 32, 33, 32, 36, 36, 33, 27, 18, 14, 13, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=114
    50, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 2, 2, 1, 3, 6, 9, 13, 10, 10, 13, 0, 
    72, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 13, 7, 6, 9, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 6, 8, 10, 5, 4, 7, 0, 
    70, 0, 0, 0, 0, 0, 0, 4, 13, 0, 0, 7, 0, 0, 0, 0, 0, 0, 5, 0, 0, 2, 3, 3, 2, 4, 7, 7, 3, 1, 2, 0, 
    69, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 8, 8, 0, 0, 0, 0, 10, 9, 0, 0, 0, 1, 1, 0, 4, 4, 0, 0, 0, 0, 0, 
    67, 0, 0, 0, 0, 0, 0, 13, 8, 0, 0, 5, 8, 6, 7, 7, 3, 15, 13, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    65, 0, 0, 0, 0, 0, 0, 19, 7, 0, 3, 7, 7, 13, 17, 16, 12, 17, 18, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    65, 0, 0, 0, 0, 0, 0, 13, 17, 4, 11, 8, 4, 11, 13, 10, 11, 18, 20, 8, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 6, 0, 
    71, 2, 3, 0, 0, 0, 0, 0, 20, 11, 19, 9, 4, 4, 0, 2, 7, 8, 13, 13, 8, 3, 0, 0, 0, 4, 0, 0, 0, 4, 6, 0, 
    85, 0, 0, 0, 0, 0, 0, 0, 18, 11, 32, 20, 5, 0, 0, 0, 8, 8, 3, 9, 12, 11, 6, 0, 1, 7, 0, 0, 4, 7, 9, 0, 
    99, 0, 0, 0, 0, 0, 0, 0, 20, 4, 33, 28, 3, 0, 0, 0, 2, 7, 1, 4, 11, 13, 14, 4, 3, 11, 8, 7, 8, 8, 7, 0, 
    109, 0, 0, 0, 0, 0, 0, 0, 27, 1, 22, 26, 0, 0, 0, 0, 2, 5, 0, 2, 8, 7, 13, 14, 8, 14, 17, 11, 7, 5, 3, 0, 
    111, 0, 0, 0, 0, 0, 0, 0, 24, 22, 21, 22, 0, 0, 0, 0, 4, 2, 0, 0, 4, 0, 7, 20, 10, 11, 21, 15, 6, 1, 0, 0, 
    106, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 27, 2, 0, 0, 0, 10, 3, 0, 0, 0, 0, 0, 24, 12, 3, 18, 17, 2, 0, 0, 0, 
    101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 19, 0, 0, 5, 16, 4, 0, 0, 0, 0, 0, 18, 19, 0, 4, 12, 3, 0, 1, 0, 
    100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 12, 0, 0, 11, 19, 6, 0, 0, 0, 0, 0, 6, 21, 0, 0, 11, 7, 0, 0, 0, 
    104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 19, 5, 0, 0, 0, 0, 0, 0, 15, 6, 0, 8, 7, 0, 0, 0, 
    110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 0, 0, 0, 0, 0, 0, 5, 11, 0, 1, 2, 0, 7, 0, 
    128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 7, 5, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 5, 9, 18, 0, 
    148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 7, 22, 29, 0, 
    160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 23, 29, 0, 
    166, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 19, 3, 0, 0, 0, 0, 0, 0, 0, 0, 12, 3, 0, 12, 25, 0, 
    154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 1, 24, 15, 0, 2, 1, 0, 0, 0, 0, 0, 27, 20, 0, 0, 19, 0, 
    124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 30, 11, 0, 0, 23, 16, 4, 7, 8, 1, 0, 0, 0, 0, 30, 35, 6, 0, 9, 0, 
    105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 26, 11, 0, 0, 9, 17, 9, 17, 16, 0, 0, 0, 0, 0, 18, 39, 26, 1, 0, 0, 
    84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 20, 1, 0, 0, 10, 10, 22, 17, 0, 0, 0, 0, 0, 8, 29, 39, 19, 0, 0, 
    75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 18, 0, 0, 10, 11, 23, 21, 0, 0, 0, 0, 0, 0, 22, 41, 35, 5, 0, 
    72, 0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 5, 0, 20, 23, 0, 0, 16, 16, 22, 25, 0, 0, 0, 0, 0, 0, 22, 37, 41, 25, 0, 
    69, 0, 0, 0, 0, 0, 0, 4, 12, 34, 50, 22, 0, 13, 11, 3, 10, 20, 21, 20, 26, 18, 4, 0, 0, 0, 0, 26, 37, 38, 37, 0, 
    62, 0, 0, 3, 10, 12, 11, 16, 24, 46, 55, 27, 7, 8, 0, 8, 19, 29, 32, 22, 23, 30, 23, 14, 10, 4, 10, 30, 39, 36, 38, 0, 
    52, 3, 7, 16, 24, 26, 26, 28, 27, 45, 55, 31, 18, 7, 0, 14, 26, 35, 38, 29, 25, 33, 30, 25, 26, 22, 22, 33, 40, 37, 34, 0, 
    44, 24, 29, 39, 43, 45, 44, 42, 39, 51, 58, 44, 41, 25, 24, 37, 43, 49, 51, 44, 39, 45, 41, 41, 46, 43, 41, 45, 49, 46, 41, 8, 
    
    -- channel=115
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 17, 22, 27, 29, 30, 33, 38, 44, 
    94, 85, 85, 85, 89, 84, 81, 91, 99, 117, 132, 119, 100, 99, 98, 93, 85, 83, 84, 87, 89, 88, 88, 87, 87, 84, 80, 76, 73, 68, 64, 57, 
    95, 88, 88, 87, 90, 86, 92, 114, 117, 121, 138, 139, 116, 104, 109, 110, 99, 91, 88, 92, 93, 92, 87, 83, 79, 71, 62, 55, 50, 45, 43, 43, 
    95, 86, 85, 83, 86, 90, 94, 110, 127, 130, 146, 164, 163, 142, 129, 123, 112, 101, 91, 87, 81, 75, 67, 59, 53, 46, 38, 35, 37, 41, 47, 51, 
    99, 92, 90, 87, 89, 97, 94, 95, 132, 157, 171, 182, 193, 196, 181, 159, 127, 92, 73, 63, 58, 48, 46, 44, 47, 51, 51, 52, 58, 63, 69, 68, 
    100, 95, 96, 93, 90, 103, 114, 119, 134, 166, 174, 173, 180, 194, 196, 183, 155, 107, 68, 52, 59, 64, 65, 68, 70, 73, 74, 76, 82, 87, 90, 80, 
    100, 94, 96, 94, 92, 99, 121, 150, 161, 169, 182, 182, 186, 187, 185, 175, 159, 149, 132, 107, 94, 97, 97, 99, 90, 84, 84, 88, 89, 87, 84, 74, 
    99, 93, 89, 84, 74, 55, 69, 126, 168, 183, 181, 173, 173, 173, 174, 181, 175, 168, 173, 164, 137, 124, 119, 111, 101, 78, 69, 74, 76, 75, 71, 61, 
    88, 74, 64, 51, 27, 5, 26, 89, 153, 170, 159, 136, 127, 132, 147, 172, 187, 180, 172, 174, 175, 167, 151, 121, 92, 74, 65, 67, 69, 70, 67, 57, 
    59, 32, 20, 12, 10, 18, 56, 105, 144, 164, 169, 150, 134, 131, 138, 163, 183, 186, 185, 183, 187, 190, 177, 147, 107, 81, 69, 64, 61, 61, 62, 58, 
    50, 16, 21, 32, 49, 64, 84, 123, 139, 149, 168, 175, 163, 169, 163, 168, 183, 183, 185, 192, 191, 195, 199, 180, 142, 102, 76, 65, 66, 70, 75, 67, 
    79, 52, 62, 74, 84, 80, 63, 101, 132, 120, 122, 148, 160, 174, 191, 181, 178, 172, 172, 183, 188, 187, 194, 189, 154, 126, 100, 79, 75, 76, 80, 72, 
    99, 79, 82, 87, 94, 83, 50, 59, 126, 127, 112, 127, 145, 152, 177, 186, 173, 162, 159, 170, 180, 184, 188, 187, 157, 127, 114, 93, 82, 84, 90, 83, 
    109, 93, 93, 91, 91, 79, 47, 21, 72, 142, 168, 172, 173, 173, 172, 181, 171, 160, 154, 162, 175, 183, 189, 188, 174, 139, 126, 112, 99, 100, 100, 86, 
    110, 96, 91, 84, 76, 69, 52, 15, 0, 57, 145, 189, 184, 185, 184, 176, 165, 152, 150, 153, 169, 184, 189, 190, 186, 159, 137, 130, 112, 97, 87, 70, 
    102, 82, 74, 68, 64, 70, 83, 82, 32, 5, 29, 86, 116, 120, 149, 166, 167, 159, 154, 158, 168, 183, 187, 186, 185, 168, 138, 124, 101, 80, 68, 62, 
    94, 72, 65, 62, 62, 65, 77, 113, 97, 27, 6, 8, 75, 89, 115, 162, 179, 182, 175, 172, 175, 179, 184, 184, 182, 172, 139, 109, 85, 72, 86, 89, 
    92, 65, 60, 50, 32, 11, 0, 16, 82, 50, 27, 40, 80, 107, 104, 146, 178, 179, 178, 174, 172, 173, 179, 184, 182, 175, 149, 125, 112, 106, 111, 103, 
    72, 31, 13, 0, 0, 0, 0, 0, 69, 134, 86, 59, 78, 134, 130, 151, 176, 178, 176, 175, 171, 170, 176, 184, 184, 178, 161, 140, 129, 112, 97, 80, 
    32, 0, 0, 0, 18, 77, 96, 79, 92, 156, 155, 120, 100, 145, 165, 158, 172, 176, 176, 176, 173, 170, 176, 184, 187, 178, 156, 122, 101, 83, 73, 70, 
    53, 2, 22, 43, 81, 163, 225, 222, 184, 174, 192, 184, 162, 158, 180, 173, 166, 169, 172, 171, 168, 174, 186, 192, 191, 174, 138, 91, 68, 69, 69, 69, 
    93, 53, 58, 68, 93, 135, 200, 222, 218, 203, 209, 219, 209, 187, 187, 189, 175, 173, 178, 177, 175, 179, 185, 187, 178, 159, 127, 83, 55, 66, 73, 67, 
    106, 85, 109, 133, 127, 89, 85, 104, 139, 193, 219, 230, 215, 178, 148, 172, 203, 200, 201, 194, 181, 171, 165, 161, 153, 140, 119, 96, 67, 61, 77, 71, 
    164, 160, 178, 184, 158, 109, 83, 96, 100, 130, 186, 203, 185, 141, 101, 105, 165, 201, 200, 189, 166, 148, 149, 150, 146, 140, 122, 108, 88, 61, 68, 75, 
    192, 196, 173, 141, 121, 114, 114, 113, 95, 73, 87, 127, 137, 133, 115, 98, 109, 143, 158, 156, 142, 134, 147, 154, 134, 115, 119, 114, 107, 77, 58, 69, 
    134, 134, 121, 116, 112, 109, 100, 89, 84, 78, 64, 68, 109, 142, 147, 133, 130, 153, 166, 160, 141, 127, 145, 166, 159, 122, 100, 107, 109, 102, 74, 61, 
    117, 112, 114, 108, 97, 88, 89, 101, 117, 127, 120, 105, 117, 153, 158, 141, 140, 159, 173, 174, 171, 161, 165, 180, 182, 156, 120, 103, 105, 112, 97, 62, 
    110, 102, 92, 87, 95, 109, 122, 130, 132, 127, 113, 98, 88, 105, 126, 142, 143, 149, 161, 172, 192, 199, 189, 179, 174, 160, 137, 113, 103, 106, 108, 80, 
    92, 83, 90, 106, 124, 136, 135, 128, 115, 101, 91, 88, 89, 90, 105, 120, 129, 134, 139, 144, 160, 181, 179, 164, 154, 145, 129, 112, 99, 97, 105, 95, 
    109, 104, 117, 126, 129, 122, 107, 96, 91, 91, 94, 96, 97, 99, 109, 107, 103, 103, 106, 109, 117, 134, 144, 147, 141, 127, 111, 101, 97, 93, 98, 96, 
    131, 127, 123, 114, 101, 92, 86, 83, 87, 91, 98, 98, 102, 101, 99, 101, 93, 90, 93, 95, 97, 104, 109, 112, 112, 103, 93, 93, 96, 93, 91, 85, 
    138, 138, 127, 117, 118, 119, 123, 125, 122, 121, 133, 142, 140, 145, 130, 126, 127, 125, 127, 130, 126, 122, 123, 120, 121, 122, 120, 120, 121, 122, 118, 106, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 4, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 35, 34, 32, 26, 27, 37, 44, 30, 11, 0, 0, 6, 12, 12, 14, 16, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 35, 34, 33, 25, 22, 33, 27, 2, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 32, 32, 24, 19, 32, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 7, 4, 10, 
    0, 28, 27, 29, 24, 16, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 10, 9, 9, 11, 12, 16, 24, 24, 19, 13, 16, 
    0, 21, 20, 23, 24, 14, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 25, 25, 23, 26, 31, 26, 26, 30, 26, 18, 9, 10, 
    0, 14, 12, 16, 24, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 26, 25, 30, 32, 30, 31, 32, 24, 13, 3, 1, 
    0, 11, 11, 15, 30, 33, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 24, 29, 34, 27, 16, 7, 0, 1, 
    0, 20, 26, 39, 54, 65, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 22, 34, 27, 17, 11, 7, 13, 
    0, 51, 62, 75, 85, 102, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 34, 32, 25, 20, 16, 26, 
    0, 87, 99, 110, 118, 141, 124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 26, 36, 34, 33, 31, 40, 
    0, 119, 129, 134, 133, 154, 135, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 39, 45, 44, 39, 46, 
    0, 131, 136, 135, 131, 146, 142, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 32, 46, 46, 40, 42, 
    0, 125, 128, 129, 124, 131, 143, 97, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 38, 40, 31, 29, 
    0, 114, 117, 119, 118, 124, 135, 128, 69, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 25, 20, 20, 
    0, 104, 111, 117, 121, 125, 122, 108, 92, 84, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 14, 18, 
    0, 105, 114, 121, 130, 142, 139, 103, 86, 127, 101, 26, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 6, 
    0, 117, 131, 146, 166, 191, 200, 146, 91, 123, 134, 96, 69, 27, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 157, 177, 197, 217, 234, 251, 219, 135, 120, 135, 123, 101, 19, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 213, 230, 244, 257, 255, 234, 234, 164, 85, 91, 111, 96, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 262, 277, 287, 290, 239, 146, 143, 117, 41, 33, 55, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 294, 296, 295, 293, 211, 81, 62, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 280, 265, 250, 243, 176, 69, 43, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 8, 0, 0, 
    0, 221, 200, 185, 173, 137, 80, 64, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 0, 0, 
    0, 153, 135, 116, 100, 89, 77, 69, 64, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 
    0, 83, 69, 65, 63, 64, 61, 54, 47, 44, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 2, 
    0, 45, 44, 46, 45, 42, 39, 37, 31, 24, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 
    0, 35, 33, 31, 26, 24, 22, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 27, 23, 20, 12, 5, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    37, 60, 58, 57, 56, 58, 59, 62, 65, 74, 81, 77, 64, 58, 52, 50, 48, 43, 41, 41, 36, 33, 30, 26, 22, 17, 13, 12, 9, 7, 4, 0, 
    98, 112, 108, 107, 107, 113, 109, 109, 123, 134, 139, 141, 129, 112, 102, 93, 87, 82, 83, 80, 74, 67, 58, 52, 47, 40, 36, 34, 29, 24, 20, 0, 
    99, 111, 107, 103, 105, 110, 102, 107, 123, 130, 142, 146, 145, 133, 117, 102, 90, 82, 80, 76, 70, 63, 57, 52, 46, 42, 38, 37, 34, 34, 35, 0, 
    97, 111, 107, 101, 106, 106, 91, 101, 112, 130, 150, 158, 155, 152, 145, 127, 102, 81, 76, 74, 72, 64, 58, 56, 56, 57, 58, 60, 59, 58, 57, 6, 
    95, 108, 108, 102, 106, 100, 81, 103, 117, 132, 141, 151, 156, 151, 152, 146, 123, 100, 83, 79, 79, 82, 81, 85, 85, 87, 85, 81, 77, 73, 68, 10, 
    92, 105, 105, 100, 97, 85, 74, 105, 128, 124, 130, 139, 148, 153, 156, 153, 134, 126, 117, 114, 112, 115, 116, 109, 101, 98, 94, 90, 83, 75, 66, 7, 
    88, 102, 103, 97, 84, 70, 68, 83, 111, 131, 135, 139, 141, 147, 151, 159, 161, 154, 149, 145, 142, 135, 128, 115, 107, 98, 90, 82, 74, 66, 58, 4, 
    86, 97, 101, 100, 84, 59, 42, 67, 107, 131, 138, 135, 132, 138, 148, 155, 163, 170, 163, 149, 150, 152, 148, 128, 100, 88, 81, 77, 73, 69, 67, 9, 
    89, 102, 106, 107, 103, 77, 54, 83, 107, 130, 141, 143, 146, 149, 151, 158, 157, 161, 170, 166, 162, 167, 157, 137, 112, 92, 87, 86, 83, 78, 75, 12, 
    106, 117, 129, 142, 160, 133, 83, 91, 107, 127, 148, 161, 170, 172, 162, 161, 166, 166, 166, 171, 171, 172, 172, 155, 137, 112, 98, 92, 90, 92, 92, 20, 
    135, 163, 179, 193, 207, 155, 86, 79, 106, 125, 144, 161, 178, 178, 175, 170, 166, 168, 167, 168, 174, 176, 179, 170, 148, 127, 113, 108, 106, 104, 100, 21, 
    167, 197, 203, 205, 211, 149, 87, 75, 98, 121, 144, 160, 177, 182, 167, 171, 170, 165, 161, 165, 169, 170, 175, 173, 160, 135, 123, 118, 110, 104, 97, 20, 
    178, 200, 201, 201, 202, 154, 89, 78, 83, 120, 155, 179, 179, 185, 174, 170, 175, 167, 161, 163, 166, 163, 170, 174, 166, 149, 127, 119, 111, 103, 93, 17, 
    174, 195, 191, 189, 189, 168, 107, 88, 83, 91, 130, 177, 186, 180, 185, 176, 180, 173, 165, 161, 165, 161, 163, 177, 168, 156, 133, 118, 107, 93, 82, 12, 
    167, 184, 180, 181, 184, 179, 141, 107, 108, 85, 93, 131, 157, 153, 162, 172, 185, 183, 173, 169, 166, 163, 163, 174, 170, 155, 135, 112, 98, 85, 73, 7, 
    163, 182, 182, 183, 187, 188, 176, 155, 142, 108, 92, 96, 122, 144, 152, 172, 190, 196, 192, 180, 173, 167, 165, 168, 171, 152, 137, 113, 91, 75, 72, 12, 
    168, 186, 191, 198, 206, 200, 180, 179, 173, 135, 104, 137, 136, 154, 152, 167, 195, 198, 196, 184, 173, 170, 168, 165, 170, 155, 138, 118, 98, 87, 80, 18, 
    175, 202, 209, 215, 217, 204, 176, 195, 195, 213, 189, 155, 152, 152, 160, 172, 188, 198, 193, 187, 179, 174, 175, 167, 171, 161, 143, 126, 103, 84, 67, 4, 
    194, 215, 222, 233, 246, 261, 240, 249, 249, 222, 237, 170, 167, 161, 169, 173, 186, 196, 195, 190, 186, 182, 180, 172, 170, 165, 139, 116, 81, 50, 33, 0, 
    224, 247, 270, 295, 301, 304, 297, 257, 269, 240, 244, 181, 186, 177, 166, 178, 187, 193, 195, 192, 190, 187, 183, 177, 170, 163, 127, 89, 50, 30, 29, 0, 
    265, 311, 321, 319, 284, 266, 277, 238, 238, 234, 233, 193, 179, 187, 169, 175, 189, 194, 195, 193, 191, 186, 182, 178, 166, 153, 117, 78, 49, 31, 32, 0, 
    294, 321, 320, 302, 238, 216, 205, 179, 172, 196, 208, 188, 174, 173, 155, 159, 183, 193, 196, 192, 185, 182, 177, 166, 152, 137, 113, 86, 63, 40, 34, 0, 
    291, 311, 306, 286, 208, 173, 159, 155, 158, 161, 170, 165, 166, 158, 130, 118, 145, 181, 188, 188, 177, 166, 162, 157, 146, 131, 120, 95, 73, 55, 39, 0, 
    258, 294, 275, 232, 166, 145, 160, 150, 142, 126, 117, 137, 155, 145, 109, 110, 120, 140, 161, 165, 163, 165, 171, 167, 140, 113, 109, 102, 84, 68, 48, 0, 
    210, 210, 178, 162, 155, 153, 153, 136, 106, 101, 106, 111, 137, 149, 123, 101, 113, 134, 156, 173, 180, 177, 174, 166, 146, 117, 92, 98, 89, 77, 62, 0, 
    144, 147, 149, 152, 147, 132, 122, 126, 123, 105, 105, 117, 132, 152, 146, 121, 124, 143, 164, 184, 194, 189, 188, 180, 154, 129, 103, 87, 94, 86, 73, 11, 
    116, 137, 132, 125, 122, 126, 128, 128, 126, 118, 106, 103, 104, 109, 128, 130, 131, 145, 158, 181, 198, 197, 191, 185, 171, 135, 103, 85, 91, 91, 76, 19, 
    106, 112, 110, 118, 127, 130, 123, 111, 96, 88, 90, 82, 84, 99, 114, 110, 114, 127, 138, 158, 172, 174, 174, 170, 161, 135, 101, 78, 75, 84, 77, 18, 
    97, 108, 111, 113, 115, 109, 93, 74, 59, 63, 86, 93, 86, 95, 98, 98, 90, 93, 101, 112, 124, 131, 137, 141, 138, 120, 90, 67, 61, 68, 74, 12, 
    91, 106, 99, 90, 80, 69, 58, 51, 49, 61, 81, 91, 93, 97, 85, 75, 61, 64, 71, 71, 80, 95, 104, 105, 100, 85, 68, 57, 52, 51, 59, 5, 
    72, 79, 63, 50, 48, 47, 49, 52, 48, 59, 77, 84, 89, 89, 72, 57, 50, 51, 56, 60, 62, 67, 70, 67, 61, 54, 50, 48, 45, 42, 44, 0, 
    33, 39, 34, 38, 40, 45, 42, 41, 41, 53, 62, 68, 81, 69, 66, 55, 43, 44, 49, 48, 47, 49, 46, 47, 46, 42, 40, 39, 39, 35, 33, 2, 
    
    -- channel=118
    41, 43, 46, 42, 42, 39, 42, 44, 43, 41, 50, 52, 48, 45, 44, 46, 45, 44, 41, 44, 43, 42, 43, 42, 42, 42, 40, 38, 42, 40, 40, 53, 
    14, 24, 27, 25, 21, 20, 22, 18, 23, 24, 27, 40, 40, 33, 26, 29, 31, 31, 28, 31, 31, 30, 32, 31, 33, 32, 32, 30, 35, 35, 35, 60, 
    14, 23, 26, 27, 19, 24, 31, 8, 25, 34, 27, 32, 45, 45, 36, 34, 33, 30, 28, 32, 33, 32, 33, 33, 35, 34, 34, 33, 36, 37, 35, 70, 
    14, 24, 25, 29, 19, 27, 40, 9, 24, 38, 35, 30, 36, 48, 48, 43, 42, 31, 30, 32, 37, 35, 35, 36, 37, 35, 36, 34, 35, 35, 34, 74, 
    13, 23, 23, 29, 23, 26, 39, 24, 23, 37, 42, 39, 35, 43, 49, 48, 51, 39, 35, 32, 37, 38, 35, 37, 36, 32, 33, 32, 32, 33, 33, 72, 
    15, 23, 22, 27, 31, 30, 25, 26, 32, 39, 47, 48, 49, 47, 50, 53, 50, 40, 36, 37, 32, 33, 31, 36, 34, 29, 28, 29, 30, 32, 33, 71, 
    16, 26, 23, 26, 37, 38, 23, 16, 36, 43, 49, 51, 52, 51, 52, 57, 54, 36, 26, 34, 31, 31, 35, 35, 35, 31, 28, 30, 33, 36, 37, 74, 
    17, 27, 25, 29, 35, 51, 47, 18, 36, 45, 51, 56, 52, 53, 53, 49, 58, 49, 34, 30, 32, 34, 41, 40, 33, 35, 33, 33, 35, 37, 39, 82, 
    19, 27, 27, 29, 30, 62, 66, 29, 40, 44, 47, 57, 54, 57, 60, 49, 54, 59, 53, 40, 34, 35, 42, 50, 38, 36, 35, 35, 36, 37, 39, 91, 
    22, 26, 26, 25, 22, 66, 63, 35, 45, 43, 29, 43, 46, 54, 64, 54, 54, 59, 59, 54, 46, 42, 41, 50, 44, 37, 38, 37, 38, 38, 38, 95, 
    18, 21, 19, 18, 15, 68, 65, 28, 47, 51, 22, 30, 41, 40, 60, 57, 54, 60, 60, 58, 58, 52, 43, 47, 43, 36, 39, 38, 37, 36, 37, 96, 
    5, 15, 14, 13, 12, 60, 81, 22, 35, 55, 35, 29, 50, 39, 48, 59, 51, 59, 60, 57, 60, 63, 48, 47, 48, 33, 34, 37, 36, 36, 36, 93, 
    0, 12, 15, 13, 13, 41, 86, 41, 14, 37, 40, 32, 50, 57, 46, 56, 48, 55, 57, 55, 57, 64, 56, 43, 54, 38, 29, 35, 34, 34, 34, 84, 
    0, 12, 14, 15, 15, 25, 65, 72, 27, 22, 21, 25, 40, 57, 50, 53, 45, 49, 55, 54, 55, 62, 60, 42, 47, 49, 29, 33, 35, 34, 34, 79, 
    0, 14, 15, 15, 15, 21, 37, 63, 67, 51, 18, 12, 39, 48, 48, 47, 44, 48, 53, 57, 56, 60, 61, 49, 40, 56, 37, 33, 36, 36, 36, 83, 
    1, 17, 17, 16, 17, 25, 24, 16, 63, 75, 54, 19, 40, 54, 46, 43, 41, 47, 51, 56, 57, 58, 60, 58, 40, 55, 48, 35, 40, 38, 37, 84, 
    5, 18, 17, 16, 17, 30, 43, 0, 31, 70, 59, 46, 23, 60, 53, 39, 40, 41, 48, 54, 57, 59, 59, 62, 45, 49, 54, 40, 45, 41, 37, 74, 
    4, 16, 15, 13, 16, 28, 68, 21, 0, 61, 41, 70, 8, 48, 62, 43, 43, 42, 45, 51, 55, 58, 59, 62, 51, 45, 56, 42, 42, 42, 38, 69, 
    3, 15, 14, 12, 13, 11, 48, 68, 0, 26, 30, 84, 19, 22, 63, 50, 44, 44, 44, 48, 52, 56, 60, 62, 56, 46, 59, 46, 40, 41, 40, 73, 
    4, 11, 8, 8, 14, 0, 1, 67, 25, 7, 19, 67, 42, 14, 56, 57, 47, 46, 45, 47, 50, 54, 60, 62, 60, 51, 61, 55, 41, 42, 40, 72, 
    0, 3, 0, 7, 39, 0, 0, 27, 34, 20, 20, 41, 48, 29, 46, 54, 49, 47, 46, 47, 50, 52, 56, 61, 60, 54, 56, 61, 45, 40, 42, 72, 
    0, 0, 0, 12, 60, 22, 3, 23, 27, 29, 26, 35, 44, 45, 43, 34, 42, 46, 46, 45, 47, 50, 53, 62, 62, 55, 43, 54, 56, 41, 41, 74, 
    0, 0, 0, 4, 44, 48, 31, 48, 44, 31, 34, 40, 42, 53, 59, 27, 25, 40, 43, 43, 45, 48, 55, 63, 64, 54, 37, 40, 61, 49, 39, 76, 
    0, 0, 3, 4, 21, 33, 26, 39, 58, 49, 41, 43, 36, 47, 65, 48, 25, 36, 42, 41, 44, 46, 49, 61, 66, 50, 38, 29, 50, 60, 44, 75, 
    0, 7, 14, 16, 17, 18, 21, 25, 45, 62, 58, 45, 34, 37, 48, 58, 40, 38, 45, 39, 43, 47, 44, 53, 69, 60, 42, 31, 32, 57, 57, 76, 
    0, 17, 18, 18, 20, 19, 24, 25, 30, 43, 55, 49, 32, 29, 39, 53, 43, 36, 42, 32, 39, 50, 46, 45, 57, 68, 53, 40, 26, 40, 61, 84, 
    9, 20, 21, 21, 24, 27, 28, 28, 29, 27, 30, 45, 37, 26, 34, 52, 50, 39, 41, 28, 26, 43, 49, 47, 48, 60, 59, 46, 34, 29, 49, 94, 
    13, 25, 27, 26, 27, 31, 33, 33, 35, 29, 24, 40, 49, 35, 39, 47, 51, 44, 43, 32, 20, 31, 46, 51, 52, 56, 54, 46, 42, 32, 34, 93, 
    21, 30, 29, 28, 29, 34, 37, 37, 38, 29, 26, 37, 46, 41, 46, 44, 48, 43, 41, 42, 31, 30, 40, 48, 52, 55, 50, 43, 42, 39, 30, 83, 
    21, 31, 32, 32, 34, 38, 42, 40, 40, 28, 27, 36, 40, 46, 45, 46, 49, 43, 41, 46, 43, 37, 38, 40, 44, 50, 47, 40, 40, 43, 37, 73, 
    18, 32, 36, 35, 38, 39, 40, 40, 42, 30, 27, 37, 34, 50, 46, 44, 46, 43, 42, 46, 46, 39, 42, 39, 39, 46, 46, 41, 38, 42, 42, 71, 
    10, 22, 24, 22, 22, 23, 23, 26, 28, 19, 13, 20, 18, 27, 31, 26, 26, 26, 24, 26, 29, 25, 27, 27, 24, 26, 29, 29, 26, 26, 28, 55, 
    
    -- channel=119
    128, 27, 25, 24, 30, 31, 34, 25, 19, 20, 22, 12, 15, 21, 26, 24, 22, 26, 29, 32, 28, 30, 32, 31, 33, 35, 37, 40, 40, 35, 40, 33, 
    161, 33, 31, 28, 36, 41, 38, 30, 32, 27, 27, 22, 14, 15, 25, 31, 28, 28, 30, 33, 27, 31, 33, 31, 35, 36, 40, 44, 44, 36, 41, 23, 
    161, 32, 33, 28, 34, 43, 26, 23, 51, 26, 15, 26, 19, 5, 9, 23, 24, 27, 32, 32, 24, 30, 34, 33, 37, 37, 39, 39, 37, 31, 34, 11, 
    159, 33, 33, 29, 30, 42, 18, 14, 61, 20, 4, 20, 22, 9, 2, 12, 15, 20, 36, 35, 29, 28, 32, 30, 29, 29, 32, 30, 28, 24, 24, 0, 
    156, 34, 36, 32, 26, 36, 19, 15, 49, 18, 6, 15, 19, 13, 1, 6, 14, 19, 37, 30, 27, 21, 23, 23, 18, 21, 26, 20, 18, 17, 17, 0, 
    152, 34, 37, 36, 24, 19, 18, 35, 39, 14, 10, 10, 9, 8, 6, 4, 7, 18, 36, 23, 16, 18, 19, 18, 8, 12, 21, 18, 17, 17, 18, 0, 
    147, 34, 36, 36, 24, 10, 15, 42, 42, 14, 13, 9, 6, 3, 6, 4, 0, 5, 30, 30, 18, 20, 14, 9, 8, 16, 22, 21, 19, 18, 17, 0, 
    144, 35, 36, 40, 33, 15, 0, 17, 45, 18, 19, 13, 3, 4, 2, 0, 0, 0, 13, 26, 23, 21, 14, 2, 9, 22, 20, 17, 17, 16, 16, 0, 
    150, 41, 43, 42, 34, 10, 0, 0, 37, 17, 26, 20, 2, 2, 0, 0, 0, 0, 0, 8, 19, 20, 13, 1, 4, 22, 15, 12, 13, 11, 11, 0, 
    174, 39, 38, 32, 27, 0, 0, 0, 33, 9, 31, 41, 12, 5, 0, 0, 0, 0, 0, 0, 2, 7, 9, 7, 4, 18, 12, 4, 3, 2, 3, 0, 
    204, 29, 27, 23, 21, 0, 0, 0, 44, 8, 25, 56, 20, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 6, 17, 13, 0, 0, 0, 0, 0, 
    230, 24, 20, 16, 15, 0, 0, 0, 54, 20, 16, 46, 21, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 11, 17, 2, 0, 0, 0, 0, 
    237, 19, 17, 13, 16, 2, 0, 0, 32, 41, 24, 29, 16, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 7, 17, 0, 14, 9, 0, 0, 0, 0, 
    232, 21, 21, 17, 20, 14, 0, 0, 0, 25, 22, 32, 23, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 1, 21, 0, 7, 20, 4, 3, 9, 0, 
    225, 25, 25, 24, 25, 18, 0, 0, 0, 0, 0, 48, 47, 0, 0, 2, 7, 12, 0, 0, 0, 0, 0, 0, 16, 8, 0, 22, 17, 15, 18, 0, 
    220, 28, 26, 24, 21, 8, 0, 0, 5, 0, 0, 23, 43, 0, 0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 6, 16, 0, 18, 24, 15, 11, 0, 
    222, 24, 21, 20, 21, 11, 0, 0, 56, 0, 0, 0, 11, 2, 0, 0, 9, 13, 3, 0, 0, 0, 0, 0, 0, 19, 0, 10, 20, 0, 0, 0, 
    231, 25, 27, 29, 28, 14, 0, 0, 32, 9, 0, 0, 0, 25, 0, 0, 5, 11, 8, 0, 0, 0, 0, 0, 0, 15, 7, 0, 11, 0, 0, 0, 
    258, 31, 27, 20, 14, 2, 0, 0, 0, 22, 0, 0, 0, 35, 0, 0, 0, 11, 9, 1, 0, 0, 0, 0, 0, 7, 7, 0, 5, 0, 0, 0, 
    298, 17, 11, 7, 0, 0, 1, 0, 0, 10, 7, 0, 0, 18, 7, 0, 0, 10, 6, 3, 0, 0, 0, 0, 0, 0, 7, 0, 0, 8, 8, 0, 
    339, 8, 6, 0, 0, 0, 14, 7, 0, 8, 19, 0, 0, 4, 12, 0, 0, 5, 1, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 8, 10, 0, 
    361, 2, 0, 0, 0, 0, 15, 18, 0, 10, 10, 0, 0, 3, 0, 0, 15, 4, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 8, 0, 
    353, 0, 0, 0, 0, 0, 2, 2, 0, 0, 4, 8, 16, 22, 0, 0, 27, 20, 5, 8, 9, 1, 0, 0, 0, 0, 8, 21, 0, 0, 0, 0, 
    310, 0, 0, 3, 0, 0, 2, 4, 0, 0, 0, 12, 31, 37, 2, 0, 20, 34, 16, 17, 18, 10, 2, 0, 0, 0, 6, 22, 9, 0, 0, 0, 
    255, 10, 13, 12, 17, 20, 22, 18, 5, 0, 0, 0, 24, 32, 3, 0, 3, 30, 20, 22, 31, 12, 0, 0, 0, 0, 0, 14, 18, 0, 0, 0, 
    197, 17, 23, 26, 29, 27, 26, 20, 14, 0, 0, 0, 6, 22, 14, 2, 0, 19, 24, 26, 39, 10, 0, 0, 0, 0, 0, 2, 13, 17, 0, 0, 
    170, 27, 31, 29, 28, 22, 18, 11, 8, 8, 14, 11, 0, 9, 24, 15, 0, 8, 21, 23, 41, 17, 0, 0, 0, 0, 0, 0, 7, 18, 6, 0, 
    160, 27, 28, 24, 20, 11, 4, 3, 6, 10, 26, 22, 0, 4, 25, 7, 0, 0, 13, 14, 32, 28, 5, 0, 0, 0, 0, 0, 5, 9, 13, 0, 
    154, 20, 17, 12, 10, 8, 3, 2, 5, 13, 33, 25, 0, 0, 12, 0, 0, 0, 7, 10, 16, 25, 17, 4, 0, 0, 0, 0, 6, 4, 9, 0, 
    144, 10, 9, 9, 12, 10, 4, 2, 7, 16, 36, 23, 0, 0, 0, 0, 0, 0, 8, 8, 3, 13, 15, 6, 0, 0, 0, 0, 9, 5, 5, 0, 
    123, 13, 12, 11, 14, 9, 6, 4, 7, 14, 36, 21, 1, 3, 0, 0, 0, 0, 6, 6, 0, 5, 11, 2, 3, 0, 0, 0, 8, 10, 7, 0, 
    82, 22, 23, 20, 24, 20, 18, 18, 19, 19, 33, 27, 13, 18, 0, 7, 12, 11, 16, 15, 11, 15, 20, 13, 16, 17, 11, 12, 18, 22, 20, 19, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    
    -- channel=121
    23, 40, 38, 35, 31, 33, 37, 36, 27, 9, 0, 0, 1, 15, 24, 28, 25, 22, 19, 17, 19, 20, 21, 19, 16, 12, 9, 6, 4, 2, 0, 0, 
    38, 57, 56, 49, 45, 46, 49, 45, 25, 0, 0, 0, 0, 6, 18, 25, 28, 29, 27, 22, 22, 21, 22, 19, 16, 12, 9, 7, 7, 5, 3, 0, 
    38, 57, 56, 48, 44, 41, 36, 29, 5, 0, 0, 0, 0, 0, 0, 0, 6, 17, 18, 12, 7, 3, 4, 2, 1, 1, 1, 2, 3, 1, 0, 0, 
    38, 56, 56, 48, 41, 36, 26, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 54, 54, 47, 37, 31, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 48, 48, 44, 31, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 40, 40, 38, 27, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 34, 35, 35, 32, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 36, 40, 45, 47, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 48, 55, 60, 61, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 62, 68, 72, 74, 54, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 72, 75, 78, 81, 70, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 76, 76, 77, 79, 77, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 79, 76, 74, 74, 73, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 75, 73, 69, 67, 62, 51, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 67, 65, 64, 60, 51, 37, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 60, 58, 58, 59, 54, 32, 24, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 62, 64, 71, 81, 85, 61, 32, 32, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 85, 91, 102, 113, 119, 108, 57, 45, 24, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 118, 125, 130, 130, 127, 115, 73, 32, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    102, 148, 153, 150, 122, 94, 64, 44, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    119, 165, 164, 150, 111, 57, 19, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    118, 159, 150, 133, 102, 45, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    102, 131, 121, 109, 90, 54, 32, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    78, 96, 87, 76, 65, 52, 36, 25, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 56, 52, 49, 43, 35, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 29, 29, 26, 18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    77, 65, 60, 58, 60, 67, 71, 68, 65, 69, 71, 61, 53, 50, 48, 44, 39, 35, 35, 31, 24, 19, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    134, 108, 101, 96, 104, 114, 109, 106, 107, 107, 112, 109, 98, 88, 85, 79, 71, 65, 63, 58, 49, 42, 32, 24, 17, 12, 12, 16, 12, 7, 8, 0, 
    134, 108, 102, 94, 103, 108, 82, 92, 107, 101, 103, 111, 105, 89, 81, 74, 64, 58, 59, 52, 41, 37, 34, 31, 31, 32, 34, 38, 35, 30, 31, 0, 
    131, 105, 102, 92, 100, 101, 64, 77, 100, 84, 80, 90, 93, 83, 76, 73, 58, 55, 59, 61, 57, 56, 56, 56, 55, 58, 61, 63, 59, 53, 48, 0, 
    126, 100, 102, 91, 91, 87, 57, 68, 88, 68, 62, 72, 78, 71, 63, 67, 66, 73, 84, 86, 85, 82, 85, 83, 80, 83, 83, 77, 67, 56, 46, 0, 
    119, 93, 96, 90, 76, 53, 37, 60, 68, 54, 50, 53, 57, 60, 63, 67, 69, 88, 108, 108, 104, 105, 108, 100, 87, 84, 82, 73, 62, 51, 40, 0, 
    112, 88, 90, 85, 62, 30, 21, 43, 49, 45, 43, 41, 41, 46, 57, 68, 69, 85, 111, 117, 119, 120, 109, 96, 84, 81, 79, 70, 60, 48, 38, 0, 
    108, 86, 93, 97, 90, 54, 16, 34, 46, 48, 56, 55, 53, 58, 60, 65, 68, 77, 94, 104, 109, 117, 110, 89, 83, 82, 77, 68, 59, 52, 48, 0, 
    124, 114, 130, 143, 151, 101, 25, 23, 40, 49, 71, 78, 82, 84, 71, 68, 66, 64, 75, 87, 100, 109, 106, 91, 89, 88, 82, 77, 73, 69, 65, 0, 
    172, 165, 183, 197, 211, 134, 23, 20, 39, 42, 78, 101, 109, 109, 78, 68, 72, 66, 65, 71, 81, 90, 98, 94, 96, 101, 95, 88, 83, 80, 78, 0, 
    225, 210, 224, 234, 244, 143, 14, 26, 50, 43, 80, 117, 114, 113, 88, 71, 75, 71, 64, 65, 70, 73, 87, 91, 95, 106, 104, 99, 95, 90, 84, 0, 
    266, 236, 239, 239, 239, 150, 21, 30, 67, 64, 94, 131, 122, 108, 93, 78, 84, 80, 68, 66, 67, 61, 71, 91, 96, 107, 112, 106, 99, 90, 79, 0, 
    273, 231, 228, 226, 225, 170, 55, 21, 59, 76, 103, 133, 125, 101, 93, 82, 91, 91, 75, 71, 71, 57, 59, 88, 96, 100, 109, 104, 94, 82, 67, 0, 
    261, 218, 216, 213, 215, 196, 121, 60, 60, 60, 72, 104, 107, 87, 84, 86, 101, 107, 91, 81, 76, 60, 54, 82, 97, 88, 98, 98, 82, 67, 56, 0, 
    249, 208, 209, 213, 220, 214, 170, 124, 94, 55, 48, 96, 108, 84, 80, 94, 117, 123, 111, 94, 79, 63, 55, 73, 94, 81, 78, 80, 71, 64, 61, 0, 
    245, 213, 220, 226, 229, 210, 173, 168, 142, 90, 67, 107, 119, 88, 82, 97, 119, 129, 119, 100, 80, 66, 60, 63, 85, 80, 70, 81, 77, 69, 60, 0, 
    254, 222, 228, 239, 249, 237, 183, 214, 231, 150, 120, 123, 140, 114, 88, 99, 119, 130, 124, 105, 86, 74, 69, 60, 76, 83, 72, 81, 78, 56, 36, 0, 
    271, 245, 264, 290, 312, 309, 243, 222, 268, 226, 195, 139, 142, 140, 96, 93, 113, 125, 124, 111, 96, 85, 77, 63, 70, 85, 71, 68, 56, 29, 11, 0, 
    326, 307, 331, 352, 363, 367, 322, 252, 261, 244, 236, 151, 125, 157, 107, 89, 108, 121, 123, 117, 109, 99, 85, 68, 66, 79, 60, 42, 29, 5, 0, 0, 
    398, 367, 384, 393, 359, 347, 331, 238, 212, 228, 232, 152, 112, 149, 117, 92, 107, 120, 123, 121, 117, 107, 88, 69, 62, 71, 52, 21, 10, 1, 0, 0, 
    458, 411, 420, 403, 297, 243, 253, 194, 162, 185, 192, 133, 99, 127, 111, 93, 109, 119, 121, 122, 116, 101, 81, 63, 55, 61, 55, 28, 13, 9, 5, 0, 
    490, 418, 410, 369, 235, 170, 197, 158, 124, 132, 128, 102, 91, 95, 74, 80, 104, 110, 110, 109, 103, 94, 84, 70, 56, 54, 63, 52, 24, 11, 7, 0, 
    468, 366, 334, 290, 190, 141, 163, 135, 91, 78, 72, 69, 84, 92, 53, 46, 76, 84, 88, 99, 102, 97, 90, 72, 51, 48, 66, 72, 40, 12, 9, 0, 
    375, 278, 255, 226, 174, 147, 148, 126, 86, 50, 40, 52, 87, 98, 62, 42, 64, 79, 84, 99, 109, 110, 110, 90, 52, 39, 55, 75, 59, 26, 12, 0, 
    285, 201, 180, 164, 154, 147, 144, 131, 104, 76, 55, 62, 92, 106, 73, 39, 53, 76, 87, 116, 138, 130, 117, 101, 69, 42, 47, 62, 69, 47, 17, 0, 
    195, 141, 139, 140, 139, 135, 130, 128, 113, 82, 60, 53, 71, 88, 83, 62, 59, 78, 94, 130, 157, 140, 119, 104, 79, 53, 42, 47, 65, 64, 31, 0, 
    152, 122, 124, 125, 125, 124, 116, 103, 87, 74, 73, 64, 52, 59, 77, 70, 59, 72, 84, 114, 145, 132, 107, 99, 89, 60, 36, 34, 49, 63, 45, 0, 
    139, 109, 110, 111, 108, 95, 76, 60, 46, 50, 70, 64, 43, 58, 71, 56, 39, 47, 59, 77, 103, 106, 94, 88, 79, 54, 29, 24, 33, 45, 46, 0, 
    131, 98, 90, 79, 69, 55, 38, 26, 17, 35, 71, 72, 51, 53, 53, 37, 21, 22, 32, 40, 56, 69, 69, 64, 55, 34, 16, 15, 20, 24, 35, 0, 
    109, 65, 50, 39, 34, 28, 16, 12, 10, 33, 65, 67, 57, 51, 36, 20, 10, 11, 20, 19, 21, 34, 39, 36, 29, 14, 4, 8, 12, 10, 15, 0, 
    71, 29, 17, 13, 12, 11, 9, 8, 6, 26, 59, 56, 56, 45, 19, 10, 4, 2, 12, 12, 6, 14, 19, 15, 13, 5, 0, 0, 3, 2, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    43, 39, 41, 40, 41, 38, 40, 41, 40, 39, 40, 41, 43, 44, 46, 45, 44, 44, 44, 47, 49, 50, 52, 53, 54, 54, 54, 53, 57, 56, 55, 67, 
    24, 31, 35, 33, 30, 25, 32, 37, 34, 29, 27, 29, 28, 31, 35, 39, 40, 41, 39, 43, 44, 46, 49, 50, 51, 50, 48, 44, 46, 44, 42, 68, 
    23, 30, 33, 34, 26, 28, 44, 35, 30, 28, 23, 27, 31, 30, 29, 36, 42, 43, 41, 44, 44, 45, 45, 41, 39, 35, 33, 32, 36, 37, 37, 74, 
    25, 32, 33, 36, 27, 33, 49, 23, 31, 42, 34, 33, 40, 43, 35, 33, 38, 39, 39, 37, 33, 29, 29, 28, 29, 29, 30, 30, 34, 37, 38, 83, 
    26, 34, 33, 38, 31, 38, 51, 27, 32, 43, 37, 30, 29, 39, 42, 36, 36, 25, 23, 21, 24, 24, 25, 27, 30, 28, 31, 34, 39, 44, 46, 89, 
    27, 34, 33, 38, 39, 49, 58, 44, 36, 39, 38, 35, 34, 34, 31, 27, 31, 26, 25, 24, 26, 29, 26, 30, 34, 34, 39, 43, 44, 46, 46, 86, 
    28, 35, 32, 37, 48, 53, 46, 39, 44, 41, 41, 42, 42, 37, 33, 29, 26, 25, 30, 34, 26, 22, 27, 37, 39, 35, 35, 38, 39, 40, 41, 81, 
    27, 34, 29, 28, 29, 32, 34, 26, 38, 35, 29, 28, 27, 25, 28, 30, 32, 23, 21, 31, 33, 28, 30, 32, 32, 33, 34, 35, 37, 37, 36, 80, 
    19, 17, 9, 3, 0, 26, 51, 32, 38, 33, 27, 27, 19, 19, 26, 23, 30, 32, 25, 24, 27, 26, 28, 30, 25, 33, 34, 31, 29, 28, 29, 83, 
    0, 0, 0, 0, 0, 43, 69, 42, 39, 36, 29, 32, 24, 25, 36, 28, 26, 31, 32, 28, 26, 27, 28, 34, 28, 27, 27, 26, 28, 29, 31, 90, 
    0, 0, 0, 0, 0, 54, 69, 39, 39, 34, 15, 18, 25, 31, 43, 32, 27, 32, 32, 31, 28, 28, 25, 31, 30, 27, 28, 27, 28, 29, 31, 94, 
    0, 1, 2, 4, 6, 54, 68, 30, 34, 31, 6, 3, 20, 20, 36, 35, 24, 31, 33, 30, 30, 33, 26, 25, 24, 22, 27, 27, 29, 33, 37, 98, 
    0, 8, 11, 11, 11, 39, 67, 34, 33, 40, 25, 14, 27, 26, 27, 33, 22, 30, 34, 30, 30, 38, 31, 21, 26, 21, 25, 32, 35, 41, 45, 98, 
    0, 12, 13, 12, 10, 19, 47, 33, 11, 32, 45, 39, 43, 48, 34, 30, 18, 24, 30, 28, 28, 37, 35, 20, 27, 29, 26, 35, 41, 45, 45, 91, 
    0, 9, 9, 6, 2, 6, 28, 37, 16, 24, 26, 18, 24, 33, 30, 23, 13, 18, 25, 27, 29, 35, 35, 24, 23, 35, 28, 37, 44, 39, 34, 82, 
    0, 3, 0, 0, 0, 12, 28, 30, 42, 37, 9, 0, 15, 27, 24, 21, 17, 25, 29, 34, 34, 34, 33, 30, 22, 37, 31, 26, 30, 32, 36, 89, 
    0, 0, 1, 0, 0, 1, 9, 0, 0, 23, 20, 9, 13, 28, 22, 17, 16, 23, 28, 32, 33, 31, 30, 33, 23, 32, 33, 25, 35, 44, 53, 96, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 5, 29, 5, 32, 35, 20, 19, 21, 26, 30, 29, 29, 30, 35, 27, 27, 38, 36, 51, 58, 54, 82, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 23, 4, 48, 11, 24, 42, 26, 20, 22, 25, 27, 26, 27, 29, 33, 30, 27, 46, 45, 50, 53, 50, 78, 
    0, 0, 0, 0, 0, 0, 20, 58, 11, 9, 8, 63, 29, 11, 40, 30, 19, 22, 23, 23, 24, 27, 33, 35, 35, 31, 45, 45, 43, 48, 47, 77, 
    0, 0, 0, 0, 22, 21, 28, 71, 44, 16, 18, 53, 43, 18, 39, 37, 23, 22, 23, 23, 26, 32, 39, 41, 40, 34, 39, 42, 38, 44, 47, 77, 
    0, 0, 0, 0, 53, 19, 0, 26, 33, 34, 35, 43, 40, 35, 48, 43, 32, 30, 30, 31, 35, 35, 33, 33, 34, 32, 32, 40, 40, 41, 47, 79, 
    0, 0, 16, 39, 71, 35, 11, 27, 33, 39, 42, 42, 34, 32, 40, 35, 41, 45, 40, 33, 29, 27, 29, 37, 42, 37, 27, 34, 47, 42, 43, 81, 
    4, 37, 32, 28, 41, 40, 34, 47, 46, 34, 35, 36, 22, 26, 47, 30, 17, 26, 24, 20, 21, 24, 26, 31, 39, 37, 31, 31, 45, 45, 39, 79, 
    2, 27, 28, 30, 34, 35, 29, 28, 39, 37, 24, 17, 10, 22, 47, 50, 30, 26, 24, 12, 10, 18, 23, 32, 38, 31, 30, 29, 36, 47, 44, 78, 
    11, 33, 36, 32, 26, 22, 24, 25, 35, 54, 56, 42, 32, 33, 36, 45, 35, 28, 27, 11, 12, 26, 26, 28, 39, 42, 33, 32, 28, 42, 51, 78, 
    24, 32, 27, 23, 23, 24, 31, 37, 45, 49, 47, 44, 34, 32, 32, 41, 38, 29, 30, 20, 24, 41, 38, 31, 30, 43, 45, 40, 32, 34, 50, 85, 
    17, 26, 26, 28, 33, 40, 48, 51, 50, 38, 28, 41, 44, 28, 28, 43, 49, 41, 40, 31, 30, 42, 42, 33, 31, 42, 48, 44, 39, 35, 43, 93, 
    20, 31, 37, 45, 48, 50, 50, 48, 48, 37, 27, 35, 43, 34, 43, 47, 50, 46, 44, 40, 33, 37, 44, 45, 45, 48, 46, 43, 44, 42, 40, 92, 
    35, 50, 53, 52, 48, 44, 46, 44, 44, 33, 30, 38, 40, 40, 47, 46, 48, 45, 41, 45, 44, 41, 45, 48, 51, 51, 46, 42, 44, 47, 44, 86, 
    42, 54, 52, 48, 46, 47, 50, 46, 47, 35, 30, 39, 38, 45, 46, 47, 50, 47, 45, 49, 49, 43, 45, 45, 46, 50, 48, 45, 45, 50, 49, 80, 
    61, 79, 80, 78, 80, 80, 81, 82, 82, 73, 74, 88, 85, 95, 90, 82, 84, 83, 81, 85, 85, 81, 83, 82, 80, 84, 84, 80, 77, 80, 82, 97, 
    
    -- channel=124
    2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 4, 6, 7, 6, 7, 9, 11, 13, 16, 18, 20, 21, 20, 22, 24, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 8, 8, 6, 8, 10, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 8, 12, 12, 12, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 3, 10, 8, 13, 17, 18, 18, 20, 18, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 18, 17, 17, 18, 15, 15, 15, 16, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 17, 22, 20, 17, 8, 7, 5, 7, 13, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 18, 18, 18, 1, 0, 0, 0, 8, 10, 7, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 13, 11, 17, 1, 0, 0, 0, 2, 8, 7, 9, 10, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 11, 2, 7, 0, 0, 0, 0, 0, 5, 2, 5, 11, 9, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 3, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 8, 10, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 8, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 6, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 7, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 2, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 1, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 2, 5, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 9, 0, 0, 0, 13, 4, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 0, 8, 11, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 2, 0, 0, 0, 0, 1, 4, 3, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 4, 7, 3, 0, 0, 0, 5, 7, 2, 0, 0, 0, 
    16, 0, 0, 0, 2, 2, 0, 2, 3, 7, 0, 0, 0, 0, 0, 1, 1, 3, 3, 2, 3, 7, 5, 4, 3, 2, 4, 7, 5, 1, 1, 0, 
    34, 15, 18, 22, 21, 19, 17, 16, 18, 21, 18, 7, 8, 7, 12, 19, 18, 18, 20, 18, 17, 20, 19, 20, 20, 19, 19, 20, 21, 18, 17, 7, 
    
    -- channel=125
    12, 115, 108, 104, 101, 110, 122, 129, 125, 120, 113, 107, 99, 93, 91, 84, 72, 58, 52, 44, 38, 30, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    99, 233, 224, 216, 214, 225, 235, 243, 231, 223, 222, 220, 214, 203, 192, 179, 167, 152, 141, 127, 116, 100, 83, 66, 45, 31, 22, 21, 18, 14, 5, 0, 
    99, 233, 224, 212, 212, 214, 206, 212, 194, 202, 204, 207, 212, 201, 181, 163, 153, 143, 133, 119, 102, 86, 75, 66, 57, 55, 55, 61, 61, 59, 55, 0, 
    96, 227, 221, 208, 208, 203, 180, 173, 158, 175, 166, 163, 177, 174, 161, 148, 135, 131, 124, 124, 114, 110, 106, 105, 103, 107, 112, 121, 122, 117, 108, 15, 
    89, 217, 215, 204, 200, 187, 159, 143, 139, 143, 125, 120, 130, 132, 125, 120, 120, 140, 155, 169, 167, 164, 166, 166, 167, 170, 171, 173, 162, 145, 124, 22, 
    80, 202, 201, 196, 181, 149, 118, 109, 105, 105, 85, 78, 81, 88, 92, 99, 115, 151, 191, 221, 226, 221, 222, 217, 209, 197, 188, 180, 161, 137, 113, 11, 
    70, 186, 187, 182, 161, 118, 76, 63, 62, 66, 56, 53, 53, 56, 67, 89, 110, 148, 195, 235, 256, 253, 242, 229, 210, 196, 188, 174, 151, 126, 102, 3, 
    64, 178, 185, 190, 189, 145, 82, 55, 35, 54, 59, 66, 71, 73, 81, 97, 105, 127, 159, 197, 225, 238, 234, 217, 202, 191, 186, 169, 146, 126, 111, 10, 
    78, 212, 236, 262, 284, 241, 157, 76, 23, 47, 75, 101, 125, 128, 124, 117, 103, 106, 120, 146, 177, 202, 211, 202, 199, 196, 195, 182, 166, 154, 144, 32, 
    131, 305, 341, 378, 412, 352, 233, 97, 26, 48, 90, 134, 182, 191, 169, 139, 110, 106, 108, 113, 127, 150, 172, 184, 201, 211, 214, 205, 192, 184, 176, 54, 
    198, 414, 451, 483, 509, 420, 259, 109, 42, 62, 102, 150, 199, 221, 190, 155, 124, 115, 111, 104, 104, 116, 140, 159, 188, 211, 225, 229, 222, 214, 202, 68, 
    258, 496, 514, 525, 529, 439, 265, 129, 68, 94, 130, 176, 212, 222, 191, 159, 144, 133, 130, 114, 104, 101, 114, 137, 167, 207, 230, 243, 240, 227, 207, 71, 
    275, 508, 511, 510, 506, 448, 298, 158, 90, 107, 153, 202, 225, 216, 188, 158, 158, 156, 156, 134, 118, 104, 102, 123, 153, 194, 219, 234, 237, 218, 191, 59, 
    262, 485, 484, 482, 480, 458, 368, 242, 152, 117, 139, 171, 193, 192, 171, 152, 168, 183, 185, 162, 138, 113, 98, 114, 146, 175, 200, 210, 214, 192, 161, 38, 
    245, 458, 460, 466, 474, 472, 430, 349, 251, 169, 131, 137, 165, 182, 162, 154, 184, 210, 221, 194, 160, 122, 97, 103, 137, 155, 173, 172, 177, 166, 148, 33, 
    235, 449, 463, 479, 490, 481, 444, 407, 337, 271, 185, 168, 186, 191, 171, 161, 191, 226, 240, 216, 174, 131, 103, 96, 124, 137, 153, 156, 160, 163, 148, 38, 
    242, 464, 482, 503, 525, 524, 467, 465, 438, 400, 331, 260, 273, 241, 214, 187, 195, 231, 245, 225, 186, 144, 119, 101, 116, 129, 143, 153, 156, 155, 129, 17, 
    262, 504, 538, 582, 625, 647, 584, 532, 518, 498, 484, 368, 355, 282, 255, 206, 190, 219, 237, 226, 197, 165, 139, 114, 113, 127, 136, 149, 138, 121, 81, 0, 
    325, 609, 659, 710, 754, 789, 750, 654, 601, 538, 540, 421, 384, 304, 269, 224, 190, 209, 229, 227, 211, 190, 164, 133, 115, 121, 121, 121, 93, 63, 30, 0, 
    412, 751, 800, 838, 835, 834, 783, 672, 585, 497, 500, 425, 364, 293, 260, 229, 197, 209, 228, 230, 223, 209, 181, 144, 114, 113, 106, 88, 55, 29, 19, 0, 
    501, 882, 913, 913, 814, 717, 611, 533, 465, 396, 405, 361, 296, 247, 227, 214, 197, 211, 226, 231, 226, 210, 178, 137, 106, 101, 103, 87, 62, 38, 28, 0, 
    553, 935, 931, 889, 734, 568, 435, 378, 334, 284, 275, 244, 207, 185, 171, 171, 171, 197, 209, 211, 208, 195, 169, 138, 112, 100, 114, 114, 93, 63, 35, 0, 
    531, 878, 831, 759, 610, 456, 355, 307, 255, 196, 149, 126, 134, 152, 142, 130, 120, 139, 162, 176, 186, 187, 173, 148, 118, 101, 116, 137, 125, 88, 48, 0, 
    434, 716, 653, 587, 493, 410, 355, 312, 247, 161, 92, 66, 101, 145, 155, 127, 102, 110, 134, 155, 179, 200, 206, 184, 140, 107, 101, 135, 143, 113, 70, 0, 
    317, 518, 461, 415, 380, 356, 336, 311, 266, 204, 137, 105, 123, 166, 174, 130, 99, 97, 123, 167, 212, 244, 243, 212, 164, 118, 101, 115, 142, 132, 95, 0, 
    187, 349, 328, 321, 313, 305, 293, 287, 268, 231, 181, 137, 134, 151, 161, 142, 125, 118, 137, 192, 247, 280, 267, 222, 176, 134, 106, 100, 125, 139, 117, 6, 
    126, 272, 271, 272, 270, 269, 262, 250, 228, 205, 186, 161, 139, 124, 131, 134, 128, 119, 129, 181, 238, 269, 251, 207, 173, 138, 109, 88, 97, 123, 123, 17, 
    103, 235, 235, 240, 240, 229, 206, 176, 143, 130, 138, 141, 127, 116, 117, 126, 106, 93, 99, 133, 176, 204, 204, 180, 156, 126, 97, 71, 71, 93, 108, 14, 
    89, 217, 209, 199, 180, 156, 126, 95, 68, 73, 108, 140, 140, 123, 110, 105, 75, 63, 66, 78, 100, 122, 137, 137, 125, 99, 69, 49, 49, 62, 79, 0, 
    70, 176, 150, 124, 101, 83, 64, 49, 35, 56, 96, 135, 145, 126, 106, 77, 48, 41, 42, 45, 51, 61, 76, 89, 84, 63, 41, 29, 31, 37, 46, 0, 
    28, 101, 72, 53, 39, 38, 35, 32, 25, 45, 83, 116, 138, 116, 91, 56, 31, 25, 28, 33, 32, 35, 39, 47, 43, 33, 22, 12, 13, 17, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 66, 64, 66, 66, 66, 59, 59, 74, 97, 109, 110, 102, 85, 73, 64, 58, 55, 55, 52, 51, 48, 41, 39, 36, 34, 33, 33, 32, 33, 30, 6, 
    48, 70, 68, 68, 71, 65, 57, 76, 90, 106, 122, 121, 113, 109, 101, 83, 66, 57, 55, 55, 55, 52, 49, 51, 50, 49, 45, 40, 34, 31, 27, 0, 
    44, 67, 66, 63, 68, 62, 65, 91, 83, 98, 122, 132, 126, 121, 121, 113, 92, 73, 61, 63, 67, 67, 62, 57, 51, 45, 39, 36, 35, 34, 33, 3, 
    46, 67, 66, 63, 66, 63, 63, 78, 91, 120, 140, 155, 164, 155, 147, 137, 117, 101, 81, 72, 64, 62, 57, 54, 54, 54, 50, 46, 42, 40, 39, 9, 
    46, 68, 67, 64, 61, 55, 51, 68, 108, 132, 142, 150, 159, 170, 180, 172, 141, 108, 81, 70, 68, 68, 73, 69, 66, 61, 53, 51, 52, 53, 52, 18, 
    45, 68, 70, 66, 56, 57, 72, 87, 104, 132, 145, 150, 156, 169, 172, 170, 163, 139, 111, 95, 99, 100, 92, 80, 75, 69, 66, 63, 62, 60, 57, 18, 
    47, 68, 71, 73, 75, 70, 66, 90, 120, 152, 168, 170, 173, 172, 172, 171, 168, 173, 161, 134, 117, 112, 112, 109, 87, 67, 59, 58, 57, 57, 59, 19, 
    53, 82, 87, 88, 83, 48, 38, 88, 120, 147, 153, 149, 156, 159, 165, 179, 178, 175, 173, 167, 154, 150, 142, 121, 97, 69, 60, 65, 71, 72, 69, 17, 
    62, 85, 80, 78, 76, 50, 58, 92, 114, 134, 143, 138, 147, 151, 158, 172, 182, 185, 181, 182, 180, 174, 162, 137, 112, 91, 78, 74, 71, 69, 69, 19, 
    46, 75, 79, 88, 101, 84, 86, 93, 109, 136, 159, 154, 156, 157, 162, 175, 181, 186, 189, 190, 192, 192, 187, 166, 133, 103, 82, 77, 79, 79, 78, 24, 
    58, 97, 104, 108, 113, 92, 77, 90, 99, 123, 151, 159, 166, 182, 175, 175, 182, 179, 179, 187, 189, 189, 192, 181, 156, 123, 97, 88, 83, 78, 72, 21, 
    70, 104, 104, 108, 112, 97, 64, 76, 81, 93, 116, 143, 157, 172, 181, 176, 179, 168, 168, 176, 181, 181, 187, 185, 157, 135, 108, 87, 77, 70, 65, 21, 
    70, 106, 106, 107, 110, 104, 75, 76, 104, 97, 102, 129, 146, 153, 176, 180, 179, 171, 168, 170, 176, 179, 183, 185, 163, 138, 116, 89, 77, 69, 66, 24, 
    76, 109, 107, 107, 110, 104, 82, 61, 76, 92, 124, 149, 162, 172, 177, 179, 181, 177, 169, 169, 174, 180, 184, 185, 176, 146, 126, 95, 80, 75, 71, 22, 
    77, 111, 111, 110, 106, 99, 92, 82, 57, 75, 111, 124, 123, 145, 160, 170, 174, 171, 169, 167, 174, 182, 185, 182, 180, 152, 135, 116, 93, 71, 55, 9, 
    79, 110, 106, 107, 115, 128, 135, 157, 134, 102, 72, 81, 107, 126, 151, 169, 183, 185, 180, 176, 178, 183, 186, 181, 181, 160, 136, 112, 77, 56, 48, 17, 
    75, 118, 128, 140, 147, 142, 123, 140, 124, 106, 123, 95, 127, 111, 133, 167, 180, 187, 181, 178, 180, 181, 186, 182, 181, 167, 136, 107, 74, 64, 71, 35, 
    99, 143, 142, 131, 112, 105, 96, 114, 162, 136, 142, 100, 128, 122, 138, 168, 182, 184, 181, 179, 179, 183, 186, 187, 182, 170, 137, 114, 89, 70, 57, 16, 
    88, 117, 111, 113, 109, 120, 120, 99, 152, 170, 153, 111, 135, 152, 147, 171, 184, 185, 184, 183, 181, 181, 183, 186, 182, 170, 140, 108, 75, 48, 42, 11, 
    70, 126, 143, 148, 130, 151, 153, 137, 156, 170, 164, 151, 143, 155, 155, 166, 178, 183, 184, 181, 177, 175, 180, 184, 180, 164, 132, 90, 62, 43, 41, 12, 
    104, 154, 149, 135, 120, 169, 190, 187, 168, 155, 167, 175, 167, 159, 151, 152, 159, 173, 177, 173, 168, 174, 188, 188, 179, 154, 120, 81, 62, 52, 44, 10, 
    98, 131, 117, 115, 112, 117, 119, 124, 140, 153, 169, 177, 179, 166, 149, 138, 135, 157, 171, 177, 177, 176, 172, 164, 152, 134, 116, 87, 65, 63, 53, 12, 
    69, 127, 148, 157, 126, 81, 78, 88, 112, 143, 153, 164, 168, 138, 103, 121, 151, 167, 182, 180, 166, 157, 161, 166, 154, 131, 107, 91, 74, 67, 63, 18, 
    118, 157, 134, 106, 86, 86, 100, 108, 92, 97, 128, 145, 142, 123, 104, 91, 109, 134, 155, 168, 165, 162, 162, 157, 147, 133, 108, 97, 85, 68, 63, 23, 
    84, 95, 85, 90, 99, 99, 89, 81, 73, 58, 59, 77, 94, 120, 131, 118, 121, 138, 155, 166, 157, 151, 161, 166, 148, 123, 110, 94, 92, 78, 66, 30, 
    52, 89, 97, 97, 87, 79, 76, 76, 78, 84, 85, 86, 107, 123, 126, 121, 128, 145, 153, 155, 148, 149, 161, 172, 171, 140, 106, 88, 88, 87, 73, 26, 
    66, 88, 79, 74, 75, 79, 82, 84, 87, 92, 90, 75, 79, 105, 116, 112, 116, 126, 134, 143, 151, 154, 161, 168, 165, 142, 112, 90, 80, 84, 78, 21, 
    49, 69, 66, 69, 79, 89, 92, 87, 75, 69, 72, 77, 80, 86, 86, 101, 104, 107, 112, 118, 132, 139, 138, 134, 132, 124, 107, 83, 70, 71, 76, 25, 
    35, 62, 68, 78, 85, 84, 75, 67, 60, 65, 70, 76, 86, 86, 87, 87, 77, 81, 87, 86, 92, 105, 110, 109, 108, 100, 86, 73, 64, 61, 66, 26, 
    41, 72, 72, 69, 62, 54, 52, 57, 57, 65, 71, 77, 85, 83, 84, 70, 63, 65, 66, 69, 74, 81, 83, 86, 81, 72, 66, 64, 60, 56, 56, 24, 
    23, 28, 18, 16, 13, 18, 21, 19, 19, 23, 21, 19, 30, 23, 27, 28, 24, 23, 26, 26, 24, 24, 20, 21, 21, 19, 20, 22, 24, 20, 16, 0, 
    
    -- channel=127
    17, 1, 1, 4, 7, 9, 7, 4, 4, 6, 7, 12, 13, 14, 12, 10, 11, 12, 15, 16, 17, 18, 19, 21, 23, 26, 29, 32, 32, 34, 36, 36, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 7, 7, 10, 14, 18, 21, 24, 24, 23, 26, 26, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 3, 3, 3, 4, 6, 9, 12, 16, 17, 18, 20, 21, 22, 23, 21, 25, 22, 
    36, 0, 0, 0, 0, 0, 0, 1, 4, 1, 8, 16, 8, 1, 5, 12, 11, 10, 8, 9, 10, 15, 16, 15, 17, 18, 19, 19, 20, 18, 21, 19, 
    38, 0, 0, 0, 0, 0, 0, 0, 17, 12, 11, 20, 24, 16, 14, 20, 19, 16, 10, 5, 4, 9, 13, 13, 13, 15, 15, 14, 15, 17, 21, 20, 
    39, 0, 0, 0, 0, 1, 7, 4, 24, 15, 17, 25, 28, 32, 32, 33, 30, 21, 13, 2, 2, 1, 7, 7, 8, 10, 12, 11, 15, 19, 24, 23, 
    39, 0, 0, 0, 0, 4, 19, 23, 16, 18, 24, 29, 33, 39, 41, 41, 41, 32, 22, 5, 0, 0, 0, 5, 11, 12, 12, 11, 15, 22, 29, 27, 
    41, 0, 0, 0, 0, 0, 7, 27, 30, 21, 24, 26, 31, 33, 39, 44, 39, 38, 34, 17, 2, 0, 2, 12, 13, 13, 13, 16, 22, 29, 35, 30, 
    40, 0, 0, 0, 0, 0, 0, 24, 35, 27, 24, 21, 20, 23, 27, 38, 42, 36, 34, 32, 18, 14, 11, 8, 17, 17, 18, 24, 30, 35, 39, 27, 
    36, 0, 0, 0, 0, 0, 0, 7, 32, 27, 27, 19, 9, 7, 10, 21, 37, 37, 33, 33, 35, 28, 24, 16, 17, 24, 25, 30, 35, 37, 40, 27, 
    30, 0, 0, 0, 0, 0, 0, 0, 29, 23, 28, 19, 3, 0, 0, 10, 28, 32, 33, 34, 39, 37, 31, 26, 20, 29, 32, 35, 37, 36, 36, 22, 
    34, 0, 0, 0, 0, 0, 0, 2, 30, 15, 16, 20, 0, 0, 0, 2, 21, 25, 26, 36, 39, 36, 34, 30, 28, 34, 38, 36, 33, 31, 30, 18, 
    39, 0, 0, 0, 0, 0, 0, 0, 34, 19, 7, 15, 1, 0, 6, 8, 18, 20, 17, 26, 35, 33, 31, 35, 27, 36, 41, 32, 26, 23, 24, 16, 
    40, 0, 0, 0, 0, 0, 0, 0, 26, 28, 17, 15, 10, 0, 11, 19, 17, 15, 7, 13, 25, 28, 27, 36, 33, 27, 34, 30, 21, 18, 20, 17, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 26, 16, 9, 11, 23, 16, 10, 0, 1, 13, 23, 27, 32, 37, 21, 25, 28, 20, 20, 22, 17, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 27, 20, 16, 21, 28, 18, 3, 0, 0, 5, 19, 25, 28, 33, 22, 16, 27, 24, 22, 29, 24, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 7, 14, 23, 17, 2, 0, 0, 0, 12, 20, 23, 26, 26, 13, 24, 28, 35, 44, 41, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 17, 14, 2, 0, 0, 0, 5, 14, 18, 19, 25, 16, 25, 41, 48, 60, 50, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 2, 13, 0, 0, 0, 0, 1, 6, 13, 15, 23, 22, 33, 57, 62, 65, 50, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 10, 0, 0, 0, 0, 0, 3, 10, 14, 23, 31, 40, 64, 70, 73, 55, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 1, 9, 4, 0, 0, 0, 4, 8, 11, 17, 28, 39, 42, 63, 72, 73, 56, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 13, 14, 7, 1, 4, 6, 9, 13, 13, 20, 33, 46, 46, 53, 68, 72, 55, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 13, 14, 16, 21, 23, 17, 9, 10, 12, 10, 7, 13, 24, 41, 56, 56, 46, 59, 71, 54, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 20, 26, 20, 4, 15, 34, 18, 12, 11, 8, 2, 2, 10, 23, 44, 58, 64, 52, 47, 65, 52, 
    57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 24, 19, 12, 1, 19, 25, 13, 12, 4, 0, 0, 1, 16, 42, 59, 69, 63, 45, 52, 48, 
    54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 22, 30, 32, 18, 4, 7, 17, 11, 7, 0, 0, 0, 0, 13, 27, 58, 66, 71, 56, 43, 40, 
    46, 0, 0, 0, 0, 0, 0, 6, 14, 20, 21, 20, 33, 36, 24, 15, 11, 20, 17, 10, 1, 0, 0, 0, 13, 28, 44, 67, 72, 68, 50, 29, 
    52, 0, 0, 0, 5, 9, 17, 27, 38, 44, 45, 36, 29, 39, 40, 33, 31, 36, 35, 27, 22, 3, 0, 0, 13, 32, 49, 70, 75, 74, 65, 31, 
    50, 3, 11, 17, 25, 31, 40, 49, 58, 63, 62, 51, 34, 35, 44, 56, 57, 57, 56, 45, 42, 34, 22, 23, 31, 47, 62, 76, 82, 77, 73, 45, 
    56, 20, 31, 41, 49, 56, 60, 66, 73, 76, 71, 56, 43, 40, 57, 65, 72, 75, 73, 63, 57, 60, 57, 55, 58, 64, 72, 85, 89, 81, 74, 55, 
    71, 41, 51, 60, 69, 74, 76, 76, 76, 77, 75, 64, 51, 49, 63, 71, 84, 85, 82, 78, 73, 74, 74, 75, 77, 78, 82, 88, 89, 83, 75, 59, 
    73, 47, 53, 60, 65, 68, 67, 61, 62, 63, 65, 57, 52, 50, 52, 65, 70, 68, 69, 66, 63, 64, 66, 65, 69, 69, 68, 69, 71, 67, 62, 51, 
    
    -- channel=128
    120, 116, 97, 65, 108, 105, 94, 94, 91, 90, 98, 101, 99, 98, 95, 98, 105, 115, 112, 83, 95, 81, 87, 96, 88, 93, 91, 90, 92, 92, 93, 185, 
    103, 110, 81, 0, 12, 69, 57, 57, 58, 51, 48, 57, 62, 60, 54, 52, 66, 102, 125, 71, 43, 13, 15, 36, 45, 48, 46, 44, 49, 52, 53, 266, 
    103, 109, 101, 0, 0, 64, 60, 49, 49, 55, 40, 31, 52, 56, 47, 35, 34, 65, 118, 115, 40, 0, 2, 28, 35, 36, 39, 40, 46, 49, 50, 271, 
    104, 106, 111, 9, 0, 63, 66, 30, 27, 45, 56, 15, 22, 36, 31, 29, 20, 33, 94, 133, 41, 0, 0, 24, 29, 31, 35, 34, 37, 42, 43, 274, 
    105, 106, 112, 40, 0, 61, 79, 9, 0, 22, 62, 31, 6, 18, 15, 25, 27, 41, 86, 110, 13, 0, 0, 16, 24, 24, 25, 28, 30, 34, 37, 274, 
    105, 106, 108, 69, 0, 52, 88, 8, 0, 0, 50, 68, 41, 34, 20, 19, 29, 56, 69, 73, 0, 0, 0, 5, 12, 17, 12, 16, 21, 21, 28, 276, 
    122, 99, 105, 94, 12, 22, 63, 16, 0, 0, 35, 88, 84, 57, 40, 36, 31, 67, 45, 10, 0, 0, 0, 0, 1, 1, 0, 0, 0, 6, 8, 288, 
    160, 119, 106, 72, 0, 0, 37, 27, 0, 0, 18, 64, 89, 59, 47, 70, 46, 59, 36, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 296, 
    114, 133, 88, 1, 0, 0, 63, 56, 0, 0, 0, 22, 50, 54, 54, 73, 49, 47, 33, 0, 0, 23, 0, 0, 0, 0, 0, 21, 7, 0, 0, 303, 
    22, 81, 52, 0, 0, 19, 76, 80, 0, 0, 0, 5, 15, 38, 58, 74, 45, 48, 36, 0, 0, 1, 0, 0, 0, 0, 23, 38, 20, 0, 0, 306, 
    0, 35, 18, 0, 5, 23, 83, 75, 9, 0, 0, 0, 7, 29, 61, 82, 53, 44, 41, 0, 0, 0, 0, 0, 0, 0, 37, 48, 25, 1, 0, 293, 
    0, 25, 16, 0, 0, 28, 86, 55, 0, 0, 0, 0, 22, 52, 76, 67, 43, 50, 38, 0, 0, 0, 0, 0, 0, 0, 29, 55, 31, 17, 0, 281, 
    0, 18, 23, 4, 5, 27, 67, 52, 0, 0, 5, 6, 33, 66, 76, 48, 14, 43, 28, 0, 0, 0, 0, 0, 0, 0, 13, 51, 43, 23, 18, 280, 
    0, 20, 28, 12, 33, 30, 28, 63, 26, 20, 28, 16, 26, 50, 42, 16, 10, 35, 17, 11, 12, 0, 0, 0, 0, 0, 0, 27, 49, 20, 9, 284, 
    0, 21, 31, 10, 66, 58, 0, 49, 43, 41, 29, 0, 4, 57, 43, 0, 13, 49, 15, 9, 28, 0, 0, 0, 0, 0, 0, 0, 39, 12, 0, 288, 
    0, 18, 26, 8, 74, 90, 0, 6, 25, 9, 12, 5, 5, 48, 68, 0, 0, 52, 45, 0, 15, 13, 0, 0, 0, 0, 0, 0, 19, 1, 0, 295, 
    1, 29, 20, 10, 54, 106, 0, 0, 22, 18, 9, 33, 21, 6, 34, 58, 0, 16, 81, 0, 5, 58, 40, 0, 0, 0, 0, 15, 7, 0, 0, 302, 
    0, 55, 35, 15, 26, 76, 11, 0, 0, 26, 0, 17, 32, 4, 9, 91, 39, 0, 80, 36, 0, 61, 105, 69, 0, 0, 0, 34, 2, 0, 0, 310, 
    0, 64, 55, 14, 4, 20, 23, 0, 0, 0, 0, 0, 25, 14, 15, 75, 86, 0, 46, 50, 0, 42, 80, 100, 57, 0, 11, 40, 0, 0, 0, 315, 
    0, 47, 53, 1, 0, 0, 5, 15, 0, 0, 0, 0, 0, 13, 27, 44, 99, 38, 7, 31, 10, 47, 50, 68, 81, 37, 19, 43, 26, 0, 0, 293, 
    0, 27, 43, 0, 0, 8, 0, 11, 23, 2, 0, 0, 0, 0, 19, 9, 46, 71, 2, 10, 40, 69, 47, 48, 54, 27, 20, 48, 52, 40, 3, 250, 
    0, 14, 41, 17, 0, 5, 16, 0, 6, 6, 19, 33, 0, 0, 7, 0, 0, 55, 31, 36, 60, 66, 42, 29, 26, 27, 41, 59, 51, 41, 41, 233, 
    0, 2, 35, 41, 0, 0, 8, 1, 0, 0, 31, 60, 11, 0, 11, 0, 0, 27, 48, 77, 66, 40, 31, 25, 17, 40, 56, 54, 51, 48, 69, 230, 
    0, 0, 23, 58, 0, 0, 0, 0, 0, 0, 18, 38, 22, 5, 10, 6, 11, 22, 62, 91, 55, 19, 28, 30, 11, 38, 54, 47, 61, 73, 72, 222, 
    0, 3, 13, 55, 6, 0, 0, 0, 0, 16, 27, 7, 17, 18, 11, 7, 13, 35, 74, 81, 37, 21, 39, 37, 4, 28, 49, 53, 62, 68, 56, 221, 
    0, 9, 18, 42, 14, 0, 0, 0, 0, 52, 82, 3, 0, 20, 19, 14, 23, 49, 73, 69, 34, 33, 48, 41, 20, 26, 45, 61, 60, 58, 63, 227, 
    0, 15, 29, 41, 21, 0, 0, 2, 6, 81, 126, 10, 0, 12, 32, 27, 39, 55, 71, 65, 39, 39, 53, 42, 45, 49, 48, 46, 53, 63, 68, 226, 
    0, 20, 37, 50, 33, 0, 0, 0, 16, 62, 94, 11, 0, 22, 44, 44, 52, 60, 82, 62, 44, 44, 59, 49, 61, 70, 55, 34, 38, 51, 53, 231, 
    0, 23, 40, 59, 42, 0, 0, 0, 18, 32, 34, 14, 27, 49, 49, 56, 61, 67, 91, 58, 43, 45, 57, 55, 68, 72, 57, 38, 26, 37, 53, 236, 
    0, 29, 35, 67, 59, 0, 0, 0, 14, 20, 19, 28, 47, 55, 47, 58, 68, 85, 86, 51, 45, 50, 51, 55, 70, 73, 53, 34, 31, 44, 64, 235, 
    7, 32, 23, 56, 84, 0, 0, 0, 11, 12, 18, 43, 60, 63, 51, 59, 79, 95, 71, 49, 54, 54, 45, 53, 64, 61, 45, 45, 50, 53, 56, 232, 
    0, 29, 11, 29, 83, 28, 0, 0, 0, 0, 12, 64, 93, 83, 56, 45, 66, 72, 47, 41, 48, 35, 27, 41, 43, 44, 46, 48, 33, 25, 28, 223, 
    
    -- channel=129
    0, 0, 0, 19, 78, 140, 157, 146, 139, 138, 140, 143, 149, 149, 148, 148, 146, 129, 92, 61, 45, 74, 126, 176, 184, 178, 178, 179, 178, 174, 170, 72, 
    0, 0, 0, 25, 104, 202, 233, 217, 212, 214, 220, 220, 224, 231, 230, 234, 241, 231, 192, 139, 103, 135, 200, 267, 282, 275, 276, 276, 275, 271, 265, 149, 
    0, 0, 0, 10, 85, 180, 225, 212, 214, 230, 228, 228, 228, 245, 254, 258, 266, 260, 221, 155, 121, 158, 232, 297, 301, 291, 289, 289, 288, 285, 279, 159, 
    0, 0, 0, 0, 66, 146, 205, 201, 212, 247, 250, 235, 222, 225, 238, 251, 266, 261, 228, 182, 163, 190, 266, 321, 322, 316, 310, 304, 299, 291, 284, 162, 
    0, 0, 0, 0, 46, 115, 183, 194, 212, 257, 271, 247, 204, 188, 200, 216, 236, 232, 212, 189, 201, 230, 287, 321, 327, 327, 326, 321, 319, 316, 307, 182, 
    0, 0, 0, 0, 31, 104, 189, 212, 224, 265, 284, 256, 202, 165, 160, 177, 192, 182, 186, 194, 228, 269, 311, 329, 339, 345, 344, 344, 343, 338, 333, 204, 
    0, 7, 0, 0, 61, 163, 239, 235, 229, 258, 290, 275, 231, 191, 168, 156, 158, 150, 166, 197, 243, 284, 318, 325, 349, 367, 366, 362, 356, 344, 350, 223, 
    28, 115, 90, 100, 160, 225, 250, 239, 223, 234, 283, 294, 269, 233, 202, 174, 159, 149, 162, 192, 238, 286, 322, 332, 355, 368, 360, 344, 331, 332, 350, 234, 
    90, 219, 190, 200, 229, 265, 275, 242, 209, 221, 272, 290, 286, 266, 232, 193, 167, 139, 160, 186, 226, 287, 332, 349, 373, 382, 367, 348, 323, 319, 341, 226, 
    114, 293, 278, 264, 277, 307, 286, 242, 207, 220, 268, 288, 290, 276, 241, 193, 162, 153, 161, 186, 219, 280, 331, 354, 388, 398, 377, 352, 321, 306, 329, 218, 
    121, 312, 306, 301, 309, 317, 290, 255, 227, 238, 275, 290, 283, 263, 220, 180, 162, 157, 174, 190, 217, 272, 323, 357, 398, 405, 390, 363, 327, 303, 313, 201, 
    122, 317, 307, 304, 309, 312, 293, 266, 243, 248, 266, 273, 262, 244, 216, 188, 182, 183, 200, 202, 225, 267, 310, 356, 401, 412, 404, 380, 344, 314, 310, 193, 
    124, 323, 312, 307, 298, 299, 281, 259, 251, 235, 233, 234, 238, 241, 217, 200, 209, 217, 221, 215, 228, 257, 300, 351, 396, 412, 412, 398, 368, 338, 324, 206, 
    128, 328, 315, 311, 287, 274, 261, 251, 273, 253, 251, 259, 260, 249, 222, 205, 203, 229, 241, 226, 238, 272, 310, 347, 395, 411, 415, 409, 386, 360, 345, 224, 
    128, 331, 312, 309, 280, 256, 245, 244, 299, 285, 268, 263, 254, 239, 225, 221, 228, 237, 248, 244, 248, 274, 292, 328, 369, 402, 412, 407, 388, 369, 362, 237, 
    128, 329, 306, 294, 272, 245, 234, 234, 299, 301, 282, 261, 259, 257, 240, 217, 215, 220, 234, 246, 236, 249, 253, 258, 283, 336, 385, 389, 380, 372, 371, 249, 
    130, 324, 295, 272, 262, 248, 240, 248, 297, 314, 313, 305, 291, 267, 256, 226, 204, 209, 219, 238, 229, 251, 243, 211, 225, 266, 306, 329, 341, 354, 376, 258, 
    135, 329, 296, 269, 264, 270, 264, 259, 298, 321, 330, 325, 318, 303, 277, 246, 216, 196, 195, 229, 229, 243, 241, 200, 182, 211, 246, 275, 297, 313, 350, 244, 
    139, 341, 311, 285, 278, 290, 292, 284, 299, 311, 318, 324, 328, 314, 297, 275, 234, 209, 200, 226, 240, 239, 237, 205, 185, 184, 211, 245, 258, 267, 299, 198, 
    143, 353, 329, 303, 288, 300, 307, 301, 300, 306, 310, 310, 314, 309, 306, 302, 284, 260, 237, 238, 239, 220, 217, 202, 208, 213, 219, 227, 224, 218, 246, 163, 
    144, 359, 337, 313, 297, 303, 312, 316, 317, 314, 309, 296, 282, 281, 298, 305, 298, 287, 262, 237, 225, 204, 202, 209, 223, 229, 224, 216, 210, 205, 211, 124, 
    141, 359, 341, 317, 298, 300, 321, 329, 332, 330, 315, 291, 274, 267, 285, 295, 295, 297, 277, 230, 207, 191, 203, 217, 231, 232, 229, 220, 205, 194, 179, 91, 
    138, 356, 344, 319, 302, 295, 324, 340, 338, 338, 328, 302, 280, 274, 289, 290, 290, 295, 272, 225, 195, 191, 209, 223, 233, 238, 243, 225, 203, 186, 170, 91, 
    136, 350, 343, 321, 305, 294, 320, 341, 339, 327, 308, 282, 261, 277, 295, 291, 288, 282, 255, 217, 195, 192, 207, 220, 227, 233, 240, 225, 203, 185, 178, 94, 
    134, 347, 337, 320, 306, 296, 315, 333, 333, 306, 264, 223, 223, 272, 297, 288, 278, 267, 238, 209, 190, 187, 205, 212, 214, 218, 224, 211, 198, 192, 176, 85, 
    132, 343, 330, 314, 301, 292, 309, 330, 329, 294, 237, 200, 204, 264, 288, 271, 258, 245, 220, 193, 179, 184, 198, 201, 192, 192, 193, 188, 194, 193, 184, 100, 
    131, 339, 323, 306, 288, 288, 304, 329, 332, 298, 251, 217, 214, 257, 264, 246, 232, 216, 191, 173, 162, 174, 188, 187, 177, 171, 167, 174, 186, 195, 200, 109, 
    127, 331, 313, 296, 278, 275, 294, 328, 334, 312, 280, 249, 229, 240, 241, 222, 209, 196, 166, 154, 152, 172, 182, 182, 171, 165, 156, 159, 183, 204, 203, 110, 
    116, 310, 294, 282, 268, 261, 275, 316, 331, 318, 296, 274, 250, 241, 222, 203, 193, 169, 145, 141, 145, 165, 172, 176, 171, 164, 155, 165, 183, 193, 192, 106, 
    99, 282, 274, 274, 259, 248, 252, 293, 323, 319, 302, 281, 251, 208, 179, 171, 166, 150, 137, 135, 144, 159, 169, 175, 176, 169, 168, 170, 172, 178, 186, 107, 
    79, 248, 241, 251, 240, 223, 222, 262, 303, 305, 287, 251, 202, 155, 130, 125, 133, 132, 131, 134, 140, 154, 162, 171, 174, 169, 161, 153, 162, 179, 191, 108, 
    0, 68, 69, 76, 72, 57, 50, 68, 82, 81, 72, 57, 39, 17, 6, 9, 13, 13, 13, 7, 16, 21, 23, 26, 29, 24, 20, 24, 28, 30, 31, 0, 
    
    -- channel=130
    33, 17, 31, 84, 60, 2, 0, 0, 0, 0, 2, 3, 0, 0, 1, 4, 0, 0, 0, 0, 18, 47, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 15, 30, 119, 105, 13, 0, 0, 0, 0, 0, 10, 5, 0, 4, 7, 0, 0, 0, 0, 16, 81, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 17, 20, 105, 123, 23, 0, 9, 9, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 20, 100, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 18, 15, 83, 127, 34, 0, 27, 27, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 27, 91, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 19, 15, 58, 118, 50, 0, 40, 45, 0, 0, 0, 0, 0, 10, 9, 0, 0, 0, 0, 38, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 18, 18, 39, 111, 77, 6, 27, 49, 3, 0, 0, 0, 0, 19, 11, 0, 0, 0, 8, 43, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 0, 12, 48, 116, 72, 0, 0, 46, 14, 0, 0, 0, 0, 0, 0, 1, 0, 6, 41, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 0, 0, 51, 82, 31, 0, 0, 33, 26, 0, 0, 0, 0, 0, 0, 0, 0, 10, 54, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    68, 0, 0, 41, 42, 0, 0, 0, 29, 35, 0, 0, 0, 0, 0, 0, 0, 7, 4, 45, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    108, 0, 0, 11, 0, 0, 0, 0, 29, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    122, 0, 0, 0, 0, 0, 0, 0, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 26, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    122, 0, 0, 0, 0, 0, 0, 0, 14, 4, 0, 0, 0, 0, 0, 0, 10, 0, 0, 20, 9, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 1, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    123, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    119, 0, 0, 0, 0, 0, 42, 18, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    117, 0, 0, 0, 0, 0, 51, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 0, 0, 0, 0, 0, 0, 0, 
    115, 0, 0, 0, 0, 0, 30, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 16, 0, 0, 0, 38, 30, 0, 0, 0, 0, 0, 0, 
    118, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 26, 0, 0, 0, 31, 44, 11, 0, 0, 15, 0, 0, 
    123, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 12, 0, 0, 0, 0, 35, 25, 0, 0, 18, 6, 0, 
    129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 9, 0, 0, 16, 22, 0, 
    132, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 8, 0, 
    134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    134, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    131, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    129, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 5, 19, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    127, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 19, 69, 0, 0, 0, 0, 0, 0, 0, 10, 12, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    124, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 24, 54, 0, 0, 0, 0, 0, 0, 0, 19, 10, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 
    120, 0, 0, 0, 0, 13, 16, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 26, 5, 0, 0, 0, 0, 0, 23, 14, 0, 0, 0, 
    113, 0, 0, 0, 0, 15, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 23, 1, 0, 0, 0, 0, 6, 19, 11, 0, 0, 0, 
    104, 0, 0, 0, 0, 8, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 12, 2, 6, 0, 0, 0, 3, 5, 3, 0, 0, 0, 
    93, 0, 0, 0, 0, 0, 50, 5, 0, 0, 0, 0, 0, 0, 5, 15, 0, 0, 10, 18, 3, 6, 12, 0, 0, 0, 0, 2, 7, 5, 0, 0, 
    67, 11, 24, 12, 0, 15, 56, 26, 0, 0, 0, 0, 0, 2, 30, 37, 20, 14, 29, 28, 20, 27, 29, 17, 15, 17, 17, 19, 27, 27, 20, 0, 
    
    -- channel=131
    56, 38, 36, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71, 63, 75, 108, 124, 94, 79, 75, 70, 80, 102, 102, 85, 82, 85, 83, 69, 39, 15, 37, 88, 89, 63, 58, 64, 65, 68, 74, 76, 76, 77, 58, 
    71, 64, 71, 99, 133, 120, 98, 82, 56, 52, 71, 100, 95, 77, 74, 71, 67, 47, 14, 3, 31, 59, 63, 64, 73, 74, 79, 83, 82, 79, 78, 57, 
    70, 65, 69, 87, 131, 134, 106, 84, 48, 27, 36, 62, 94, 87, 75, 68, 66, 68, 61, 44, 29, 36, 57, 66, 70, 73, 78, 79, 79, 77, 75, 56, 
    69, 63, 64, 78, 123, 143, 107, 81, 57, 27, 21, 39, 89, 125, 131, 120, 104, 95, 87, 58, 38, 52, 82, 91, 78, 68, 69, 67, 68, 72, 72, 52, 
    69, 65, 62, 71, 110, 133, 92, 64, 58, 44, 29, 29, 61, 107, 125, 140, 143, 126, 107, 71, 30, 52, 94, 111, 94, 79, 69, 66, 61, 59, 57, 31, 
    41, 56, 69, 67, 58, 74, 70, 52, 52, 52, 43, 27, 20, 42, 67, 90, 117, 118, 95, 78, 47, 40, 72, 76, 55, 51, 50, 59, 78, 78, 68, 37, 
    0, 0, 10, 10, 0, 21, 55, 79, 88, 72, 51, 31, 1, 0, 15, 41, 56, 72, 64, 69, 77, 73, 80, 69, 42, 34, 48, 70, 98, 110, 88, 49, 
    25, 0, 0, 0, 0, 43, 86, 99, 99, 93, 71, 52, 29, 10, 11, 28, 46, 43, 53, 66, 83, 91, 80, 75, 69, 71, 87, 114, 128, 132, 115, 56, 
    100, 46, 16, 16, 44, 75, 87, 84, 66, 67, 71, 68, 59, 54, 50, 57, 61, 71, 65, 73, 81, 90, 87, 72, 68, 79, 87, 104, 123, 129, 134, 86, 
    117, 79, 76, 80, 81, 84, 89, 75, 52, 36, 46, 56, 59, 72, 83, 78, 61, 53, 60, 64, 75, 92, 114, 96, 76, 84, 94, 97, 115, 127, 136, 110, 
    122, 88, 81, 87, 99, 103, 91, 65, 55, 51, 50, 62, 70, 68, 77, 69, 51, 32, 39, 45, 60, 82, 107, 109, 92, 93, 97, 96, 106, 128, 138, 108, 
    128, 103, 99, 99, 107, 124, 106, 61, 64, 90, 102, 97, 81, 66, 48, 27, 18, 29, 28, 39, 56, 78, 91, 99, 95, 95, 89, 79, 80, 107, 116, 77, 
    130, 105, 104, 100, 100, 119, 121, 71, 49, 69, 85, 83, 67, 54, 57, 52, 25, 33, 53, 58, 55, 74, 96, 91, 95, 97, 91, 73, 68, 81, 90, 53, 
    133, 109, 103, 91, 85, 83, 102, 74, 28, 20, 5, 16, 39, 36, 36, 62, 84, 55, 63, 77, 52, 57, 97, 118, 100, 96, 93, 89, 89, 79, 85, 56, 
    133, 113, 116, 98, 78, 51, 66, 78, 43, 43, 50, 47, 61, 66, 23, 15, 81, 90, 58, 79, 90, 74, 122, 186, 176, 121, 100, 107, 116, 106, 94, 65, 
    132, 109, 125, 121, 91, 44, 30, 77, 69, 49, 53, 51, 45, 50, 47, 44, 77, 126, 84, 75, 101, 87, 106, 168, 233, 211, 157, 140, 134, 125, 108, 68, 
    132, 103, 108, 113, 85, 42, 12, 41, 78, 48, 18, 9, 1, 15, 35, 46, 59, 108, 109, 70, 73, 71, 55, 58, 106, 184, 202, 177, 161, 146, 126, 70, 
    133, 99, 83, 78, 63, 43, 32, 35, 75, 90, 68, 52, 32, 6, 15, 30, 29, 61, 111, 72, 63, 90, 84, 56, 39, 70, 115, 126, 134, 160, 169, 103, 
    133, 99, 81, 71, 67, 55, 59, 60, 63, 93, 100, 101, 98, 64, 37, 26, 10, 6, 52, 66, 63, 90, 104, 89, 62, 43, 53, 70, 90, 122, 161, 140, 
    132, 99, 87, 85, 92, 79, 69, 77, 67, 54, 62, 90, 109, 103, 76, 49, 25, 4, 10, 60, 88, 97, 89, 79, 59, 46, 58, 79, 88, 91, 107, 110, 
    133, 103, 90, 86, 97, 86, 62, 56, 63, 55, 50, 64, 87, 97, 88, 81, 81, 69, 52, 75, 105, 96, 72, 62, 62, 59, 70, 84, 81, 85, 97, 89, 
    132, 107, 99, 87, 92, 87, 62, 44, 46, 59, 64, 55, 51, 63, 70, 67, 74, 82, 83, 93, 96, 85, 69, 66, 70, 64, 64, 65, 70, 84, 98, 80, 
    131, 110, 111, 97, 86, 88, 74, 62, 56, 59, 70, 76, 50, 45, 58, 58, 59, 66, 81, 83, 78, 72, 73, 79, 78, 70, 59, 62, 71, 67, 66, 52, 
    131, 111, 119, 115, 95, 90, 80, 72, 76, 79, 103, 121, 100, 67, 68, 75, 75, 82, 83, 78, 77, 77, 84, 84, 87, 93, 85, 81, 75, 71, 66, 57, 
    129, 112, 123, 128, 120, 105, 85, 67, 70, 80, 87, 107, 108, 86, 84, 90, 94, 98, 92, 87, 85, 89, 87, 87, 85, 101, 113, 99, 79, 73, 74, 64, 
    129, 112, 124, 133, 136, 127, 98, 66, 62, 59, 27, 12, 49, 87, 98, 101, 104, 101, 98, 100, 93, 90, 89, 87, 89, 96, 107, 105, 85, 62, 54, 41, 
    132, 116, 125, 131, 139, 132, 103, 75, 67, 57, 18, 0, 28, 80, 106, 102, 100, 103, 104, 101, 94, 89, 85, 81, 81, 83, 87, 87, 84, 73, 63, 52, 
    141, 126, 130, 126, 135, 136, 105, 79, 72, 63, 51, 50, 66, 92, 99, 92, 89, 93, 101, 91, 87, 85, 83, 74, 71, 75, 74, 74, 77, 84, 85, 69, 
    153, 141, 138, 128, 126, 135, 119, 86, 74, 69, 67, 75, 94, 105, 103, 97, 88, 94, 93, 83, 85, 88, 87, 78, 75, 67, 63, 71, 84, 92, 89, 63, 
    156, 151, 149, 143, 130, 127, 126, 102, 80, 76, 78, 89, 109, 130, 139, 125, 106, 91, 76, 80, 82, 87, 81, 80, 76, 72, 75, 84, 90, 84, 74, 55, 
    221, 216, 227, 233, 226, 195, 195, 220, 215, 207, 208, 203, 187, 176, 175, 182, 177, 157, 149, 150, 157, 160, 165, 165, 163, 164, 165, 170, 167, 163, 161, 142, 
    
    -- channel=132
    0, 0, 0, 0, 0, 33, 45, 45, 46, 37, 30, 31, 36, 37, 34, 33, 43, 52, 43, 10, 0, 0, 13, 58, 69, 59, 58, 56, 58, 59, 56, 65, 
    0, 0, 0, 0, 0, 76, 111, 109, 117, 111, 96, 90, 96, 103, 98, 98, 114, 134, 135, 92, 38, 20, 57, 134, 148, 137, 135, 129, 129, 131, 127, 147, 
    0, 0, 0, 0, 0, 56, 115, 110, 124, 142, 125, 105, 105, 121, 120, 118, 130, 150, 165, 136, 57, 12, 78, 161, 163, 153, 149, 142, 141, 143, 139, 160, 
    0, 0, 0, 0, 0, 27, 104, 97, 120, 167, 168, 135, 111, 119, 121, 125, 138, 152, 169, 153, 76, 29, 107, 178, 176, 172, 166, 158, 156, 155, 152, 174, 
    0, 0, 0, 0, 0, 0, 84, 82, 111, 177, 205, 181, 127, 108, 105, 109, 130, 144, 152, 134, 84, 66, 134, 174, 178, 180, 178, 174, 175, 175, 170, 195, 
    0, 0, 0, 0, 0, 0, 71, 90, 110, 176, 226, 217, 155, 103, 80, 86, 108, 117, 124, 110, 96, 118, 162, 172, 185, 199, 197, 195, 197, 192, 187, 219, 
    0, 0, 0, 0, 0, 0, 91, 112, 113, 165, 229, 233, 189, 127, 88, 86, 90, 89, 96, 87, 110, 161, 183, 170, 200, 228, 224, 220, 215, 197, 195, 245, 
    0, 52, 17, 0, 0, 50, 118, 130, 112, 145, 212, 230, 213, 165, 127, 118, 97, 81, 88, 79, 111, 180, 190, 170, 216, 244, 233, 227, 203, 177, 186, 259, 
    0, 120, 76, 35, 52, 116, 157, 146, 102, 120, 190, 214, 215, 196, 169, 146, 112, 79, 92, 87, 108, 173, 181, 171, 226, 249, 235, 224, 180, 144, 163, 253, 
    0, 159, 137, 103, 120, 160, 171, 152, 97, 108, 176, 203, 207, 206, 190, 158, 114, 89, 99, 95, 105, 154, 164, 173, 226, 241, 229, 205, 152, 117, 134, 233, 
    0, 165, 160, 148, 154, 169, 178, 153, 102, 123, 181, 200, 202, 201, 181, 147, 106, 92, 110, 99, 109, 146, 149, 172, 227, 235, 227, 200, 144, 109, 111, 200, 
    0, 166, 164, 153, 152, 167, 177, 150, 112, 139, 182, 194, 195, 194, 173, 133, 104, 112, 132, 111, 124, 151, 141, 166, 225, 237, 229, 210, 158, 113, 105, 175, 
    0, 160, 161, 154, 146, 160, 156, 141, 134, 141, 165, 169, 171, 186, 168, 130, 116, 143, 149, 126, 141, 151, 138, 164, 218, 234, 233, 226, 189, 140, 115, 177, 
    0, 157, 156, 154, 153, 158, 126, 131, 169, 158, 165, 162, 166, 187, 170, 131, 124, 161, 159, 136, 152, 153, 143, 166, 214, 229, 234, 237, 224, 176, 135, 203, 
    0, 158, 153, 156, 168, 172, 109, 117, 193, 182, 173, 162, 167, 189, 180, 139, 137, 166, 158, 137, 147, 158, 139, 154, 195, 221, 229, 238, 239, 196, 158, 232, 
    0, 160, 149, 150, 175, 189, 115, 105, 197, 202, 192, 180, 182, 191, 188, 155, 129, 135, 150, 132, 127, 157, 137, 114, 130, 175, 211, 229, 226, 186, 170, 251, 
    0, 164, 143, 135, 161, 195, 146, 118, 194, 220, 209, 207, 207, 184, 185, 187, 137, 97, 134, 138, 111, 157, 159, 96, 68, 106, 158, 192, 184, 156, 173, 259, 
    0, 172, 148, 125, 144, 191, 180, 143, 182, 217, 216, 219, 232, 213, 196, 204, 159, 77, 103, 140, 104, 144, 171, 109, 52, 59, 105, 146, 141, 120, 155, 253, 
    0, 178, 160, 129, 138, 184, 198, 178, 178, 193, 207, 223, 242, 234, 220, 216, 179, 104, 92, 127, 117, 146, 158, 116, 92, 67, 79, 119, 117, 98, 123, 221, 
    0, 180, 171, 144, 144, 184, 197, 193, 185, 180, 193, 208, 220, 224, 232, 222, 206, 167, 119, 122, 139, 145, 128, 105, 120, 106, 100, 124, 119, 92, 96, 179, 
    0, 183, 181, 161, 151, 181, 195, 195, 195, 185, 190, 198, 181, 181, 212, 210, 205, 209, 161, 132, 150, 133, 105, 101, 123, 125, 127, 136, 124, 103, 94, 141, 
    0, 185, 187, 175, 153, 167, 200, 203, 201, 200, 206, 203, 165, 150, 184, 192, 197, 215, 190, 153, 140, 103, 94, 110, 128, 137, 147, 141, 118, 103, 98, 117, 
    0, 182, 185, 182, 156, 150, 199, 221, 216, 215, 226, 216, 170, 151, 176, 185, 189, 199, 190, 165, 117, 78, 96, 123, 132, 144, 160, 139, 117, 108, 98, 107, 
    0, 176, 174, 179, 156, 140, 193, 228, 229, 226, 227, 204, 162, 161, 181, 184, 185, 188, 182, 156, 100, 72, 103, 128, 125, 139, 160, 140, 123, 113, 97, 105, 
    0, 173, 163, 165, 148, 135, 184, 224, 229, 228, 223, 165, 125, 163, 188, 180, 178, 180, 171, 139, 92, 77, 109, 124, 115, 128, 148, 134, 120, 110, 96, 107, 
    0, 171, 154, 146, 131, 122, 169, 218, 224, 230, 222, 138, 86, 154, 186, 166, 162, 164, 150, 121, 85, 80, 108, 115, 104, 114, 121, 112, 109, 109, 106, 116, 
    0, 169, 149, 133, 111, 105, 148, 208, 223, 231, 223, 139, 90, 153, 171, 147, 142, 138, 123, 103, 70, 75, 103, 103, 100, 106, 94, 85, 94, 109, 114, 125, 
    0, 166, 144, 125, 99, 86, 127, 200, 225, 226, 212, 160, 130, 155, 149, 129, 125, 117, 104, 81, 54, 76, 98, 97, 96, 99, 79, 65, 82, 108, 117, 134, 
    0, 155, 131, 118, 96, 74, 109, 191, 225, 219, 198, 176, 164, 158, 130, 113, 115, 101, 87, 58, 44, 76, 88, 91, 96, 95, 73, 67, 81, 101, 114, 133, 
    0, 134, 110, 109, 98, 70, 91, 175, 218, 213, 195, 183, 171, 137, 100, 93, 99, 93, 72, 42, 51, 76, 79, 88, 99, 93, 77, 75, 84, 94, 105, 127, 
    0, 103, 77, 85, 91, 67, 69, 146, 203, 203, 189, 178, 153, 104, 65, 57, 74, 78, 56, 42, 59, 70, 69, 86, 96, 88, 79, 76, 80, 87, 99, 127, 
    0, 12, 0, 2, 17, 4, 0, 32, 77, 80, 75, 75, 60, 21, 0, 0, 0, 5, 0, 0, 0, 0, 0, 12, 18, 14, 13, 10, 5, 6, 16, 58, 
    
    -- channel=133
    0, 0, 2, 39, 85, 115, 108, 100, 99, 104, 108, 114, 110, 107, 108, 111, 106, 85, 58, 44, 46, 84, 105, 109, 121, 119, 122, 123, 123, 121, 119, 53, 
    1, 0, 19, 104, 166, 194, 191, 176, 169, 175, 177, 185, 191, 187, 189, 191, 184, 156, 109, 84, 85, 148, 197, 210, 214, 210, 213, 217, 214, 209, 204, 58, 
    0, 0, 7, 88, 163, 193, 188, 176, 170, 170, 180, 180, 192, 195, 196, 204, 204, 181, 131, 95, 107, 170, 211, 227, 227, 224, 225, 228, 225, 219, 214, 62, 
    1, 1, 1, 66, 149, 182, 179, 175, 180, 180, 177, 179, 181, 197, 213, 224, 227, 211, 160, 105, 130, 203, 236, 250, 244, 235, 231, 231, 228, 225, 219, 63, 
    1, 2, 0, 43, 129, 165, 170, 175, 187, 203, 184, 176, 174, 180, 198, 215, 222, 206, 166, 134, 166, 223, 254, 267, 264, 256, 248, 247, 241, 232, 227, 62, 
    2, 2, 2, 27, 111, 157, 168, 177, 195, 214, 197, 171, 150, 144, 165, 174, 183, 180, 155, 154, 206, 236, 256, 264, 264, 258, 260, 257, 255, 252, 246, 75, 
    22, 0, 1, 28, 115, 154, 166, 188, 212, 225, 211, 174, 141, 123, 130, 138, 146, 138, 145, 170, 220, 244, 256, 270, 269, 262, 269, 268, 267, 277, 274, 87, 
    67, 43, 17, 48, 124, 192, 213, 200, 210, 229, 224, 191, 160, 151, 136, 122, 127, 117, 138, 188, 231, 245, 263, 278, 277, 284, 284, 280, 283, 287, 296, 93, 
    128, 125, 119, 150, 206, 246, 217, 186, 201, 209, 222, 219, 197, 183, 164, 129, 125, 138, 142, 190, 231, 237, 274, 294, 291, 299, 289, 265, 268, 280, 298, 102, 
    209, 199, 198, 235, 256, 248, 209, 174, 191, 203, 217, 224, 218, 198, 174, 144, 140, 132, 144, 179, 218, 237, 286, 314, 307, 301, 288, 264, 259, 282, 300, 99, 
    232, 245, 240, 249, 261, 257, 212, 179, 190, 209, 217, 221, 218, 196, 167, 135, 139, 138, 137, 174, 205, 239, 289, 318, 319, 315, 293, 272, 262, 275, 299, 98, 
    239, 255, 253, 258, 265, 259, 217, 196, 202, 217, 224, 223, 215, 192, 149, 129, 139, 144, 143, 177, 194, 230, 288, 314, 322, 323, 303, 278, 270, 268, 286, 98, 
    247, 263, 254, 257, 259, 241, 223, 216, 210, 212, 210, 219, 204, 169, 146, 151, 162, 155, 169, 184, 195, 224, 282, 312, 323, 325, 314, 287, 273, 264, 277, 98, 
    249, 269, 254, 251, 239, 218, 219, 219, 212, 201, 182, 184, 185, 166, 148, 163, 202, 185, 185, 196, 205, 217, 268, 315, 322, 326, 321, 303, 278, 276, 284, 100, 
    249, 270, 257, 252, 216, 188, 207, 215, 213, 195, 192, 200, 200, 188, 170, 172, 179, 199, 196, 195, 208, 225, 269, 306, 331, 330, 330, 315, 288, 296, 303, 106, 
    249, 268, 251, 251, 205, 165, 199, 220, 239, 222, 216, 229, 211, 175, 166, 181, 182, 200, 206, 203, 211, 231, 243, 267, 314, 341, 338, 317, 295, 306, 318, 110, 
    250, 265, 244, 240, 208, 162, 197, 214, 240, 243, 227, 205, 197, 194, 178, 166, 186, 186, 192, 209, 210, 203, 196, 216, 229, 278, 318, 305, 301, 315, 323, 112, 
    253, 258, 236, 225, 213, 171, 194, 229, 235, 241, 245, 236, 220, 206, 197, 153, 156, 182, 175, 194, 206, 189, 163, 168, 193, 217, 249, 252, 266, 303, 323, 118, 
    260, 259, 236, 227, 227, 211, 209, 235, 245, 251, 267, 260, 244, 238, 214, 169, 154, 178, 160, 190, 208, 187, 172, 152, 161, 190, 202, 204, 227, 262, 293, 112, 
    265, 271, 245, 244, 246, 244, 232, 236, 256, 253, 255, 256, 249, 248, 230, 208, 169, 176, 170, 181, 200, 186, 180, 169, 155, 170, 182, 183, 199, 229, 251, 73, 
    266, 284, 260, 255, 251, 252, 251, 236, 241, 252, 243, 231, 243, 244, 231, 230, 214, 198, 209, 195, 186, 172, 175, 169, 170, 181, 189, 181, 177, 181, 204, 56, 
    267, 290, 268, 253, 251, 251, 251, 250, 243, 251, 244, 220, 223, 230, 232, 239, 238, 215, 215, 191, 168, 164, 173, 179, 186, 195, 186, 167, 164, 161, 169, 50, 
    266, 291, 273, 251, 248, 254, 254, 258, 262, 258, 236, 210, 217, 224, 224, 231, 233, 219, 200, 168, 158, 165, 179, 188, 198, 195, 176, 168, 163, 158, 146, 32, 
    262, 292, 279, 251, 254, 259, 263, 261, 264, 257, 228, 207, 229, 237, 229, 229, 227, 221, 189, 156, 155, 176, 187, 186, 198, 195, 185, 175, 160, 153, 136, 28, 
    258, 288, 282, 255, 260, 265, 266, 263, 259, 237, 198, 199, 225, 240, 235, 230, 227, 213, 180, 153, 162, 185, 182, 180, 193, 189, 186, 179, 165, 147, 145, 40, 
    256, 283, 280, 260, 260, 273, 269, 260, 254, 212, 153, 156, 196, 224, 231, 227, 218, 197, 170, 153, 167, 177, 172, 170, 182, 176, 172, 170, 166, 157, 151, 32, 
    254, 278, 272, 261, 259, 270, 270, 261, 252, 198, 135, 149, 185, 207, 219, 211, 196, 183, 159, 145, 164, 168, 164, 165, 160, 155, 153, 154, 164, 164, 150, 36, 
    249, 272, 264, 252, 248, 266, 272, 263, 252, 213, 164, 179, 201, 206, 198, 191, 177, 161, 140, 141, 153, 158, 156, 157, 146, 134, 137, 157, 165, 166, 165, 44, 
    241, 264, 257, 245, 237, 254, 269, 266, 252, 232, 212, 211, 203, 187, 181, 172, 158, 147, 123, 136, 145, 153, 155, 156, 143, 132, 138, 151, 165, 172, 169, 43, 
    226, 251, 250, 237, 228, 239, 254, 263, 251, 240, 234, 215, 184, 172, 173, 164, 153, 128, 116, 135, 141, 150, 153, 153, 143, 139, 140, 150, 165, 169, 160, 39, 
    204, 229, 240, 234, 220, 227, 237, 249, 249, 239, 228, 204, 175, 149, 144, 146, 137, 118, 121, 130, 139, 144, 153, 153, 147, 141, 146, 157, 159, 158, 152, 37, 
    126, 192, 196, 198, 180, 192, 202, 206, 225, 227, 216, 181, 141, 113, 107, 106, 104, 104, 113, 125, 128, 132, 141, 144, 143, 142, 140, 131, 135, 146, 157, 59, 
    
    -- channel=134
    36, 36, 22, 0, 38, 60, 53, 53, 49, 44, 48, 52, 52, 52, 48, 48, 56, 66, 63, 31, 31, 19, 39, 58, 54, 56, 52, 53, 56, 56, 55, 142, 
    29, 29, 20, 0, 0, 38, 36, 31, 27, 29, 22, 27, 35, 35, 31, 28, 36, 57, 76, 49, 1, 0, 12, 25, 30, 33, 32, 32, 35, 35, 35, 151, 
    29, 28, 28, 0, 0, 34, 36, 22, 22, 30, 29, 12, 26, 32, 30, 27, 25, 39, 69, 67, 3, 0, 10, 23, 27, 29, 30, 30, 33, 34, 34, 154, 
    29, 28, 30, 0, 0, 28, 36, 9, 12, 22, 40, 16, 10, 19, 20, 25, 23, 28, 48, 54, 3, 0, 8, 23, 28, 27, 28, 28, 28, 30, 30, 154, 
    29, 29, 30, 4, 0, 18, 40, 5, 0, 10, 40, 33, 9, 6, 0, 10, 19, 26, 33, 38, 2, 0, 1, 17, 25, 27, 23, 26, 27, 27, 29, 158, 
    30, 29, 31, 15, 0, 1, 44, 14, 0, 2, 31, 46, 27, 10, 2, 6, 6, 24, 18, 17, 10, 9, 1, 8, 17, 19, 15, 20, 25, 24, 26, 170, 
    52, 33, 29, 12, 0, 3, 42, 25, 0, 0, 17, 43, 47, 23, 20, 23, 4, 22, 11, 0, 3, 21, 5, 6, 20, 13, 15, 19, 12, 16, 17, 176, 
    74, 66, 36, 5, 2, 11, 41, 32, 0, 0, 8, 29, 45, 38, 32, 37, 19, 19, 14, 0, 0, 19, 0, 0, 15, 9, 14, 21, 6, 4, 11, 176, 
    46, 76, 50, 17, 7, 13, 46, 40, 0, 0, 1, 13, 24, 37, 37, 40, 18, 20, 15, 0, 0, 9, 1, 0, 4, 8, 19, 21, 11, 0, 1, 177, 
    11, 43, 36, 19, 11, 22, 53, 41, 3, 0, 0, 5, 12, 25, 35, 37, 14, 17, 15, 0, 0, 0, 0, 8, 7, 12, 34, 32, 21, 6, 0, 172, 
    3, 30, 23, 11, 14, 27, 54, 34, 9, 4, 4, 5, 16, 22, 31, 26, 17, 20, 16, 0, 0, 0, 0, 5, 11, 13, 35, 43, 26, 18, 0, 158, 
    0, 26, 25, 11, 12, 28, 47, 34, 6, 4, 10, 5, 16, 30, 33, 18, 10, 29, 14, 0, 1, 0, 0, 0, 9, 13, 30, 48, 33, 24, 14, 154, 
    0, 21, 25, 14, 21, 22, 27, 41, 12, 2, 5, 0, 12, 31, 29, 19, 11, 26, 12, 10, 3, 0, 0, 0, 6, 11, 25, 42, 45, 25, 19, 167, 
    3, 24, 28, 17, 40, 24, 0, 40, 25, 20, 10, 0, 15, 31, 18, 0, 17, 22, 9, 11, 12, 0, 0, 1, 6, 8, 13, 31, 49, 24, 19, 177, 
    5, 25, 30, 17, 50, 40, 0, 24, 29, 28, 25, 11, 10, 32, 30, 0, 0, 29, 17, 0, 21, 7, 0, 0, 9, 9, 6, 21, 34, 21, 17, 176, 
    7, 25, 24, 15, 41, 57, 0, 0, 26, 18, 13, 19, 9, 13, 33, 25, 0, 16, 40, 0, 8, 23, 1, 0, 0, 7, 9, 22, 16, 13, 18, 176, 
    8, 37, 22, 11, 22, 54, 0, 0, 17, 22, 8, 23, 21, 5, 15, 46, 0, 0, 50, 5, 0, 37, 38, 0, 0, 0, 4, 21, 8, 3, 19, 179, 
    6, 47, 31, 11, 11, 32, 25, 0, 0, 18, 12, 22, 32, 16, 13, 43, 30, 0, 34, 20, 0, 37, 48, 47, 5, 0, 0, 15, 0, 0, 12, 182, 
    2, 45, 43, 14, 12, 15, 21, 14, 0, 0, 1, 5, 21, 23, 23, 31, 53, 3, 7, 24, 9, 26, 27, 47, 43, 4, 5, 23, 7, 0, 0, 169, 
    0, 36, 43, 15, 10, 15, 11, 21, 15, 1, 0, 1, 0, 12, 23, 18, 49, 44, 0, 21, 23, 25, 15, 28, 35, 21, 19, 29, 21, 6, 0, 138, 
    0, 29, 40, 18, 3, 14, 14, 10, 20, 15, 16, 15, 0, 0, 12, 6, 24, 51, 20, 23, 24, 23, 18, 21, 24, 23, 22, 26, 22, 22, 14, 117, 
    0, 22, 38, 30, 0, 6, 20, 13, 11, 15, 29, 31, 0, 0, 9, 0, 3, 26, 32, 34, 19, 17, 22, 19, 16, 23, 27, 25, 25, 23, 25, 109, 
    0, 15, 31, 41, 0, 0, 12, 16, 11, 14, 26, 35, 14, 6, 15, 8, 8, 15, 35, 38, 19, 14, 21, 18, 8, 25, 31, 26, 32, 26, 25, 110, 
    0, 15, 23, 45, 9, 0, 5, 9, 9, 20, 25, 13, 14, 15, 15, 13, 14, 23, 37, 37, 20, 13, 21, 17, 4, 23, 29, 29, 30, 32, 31, 115, 
    0, 18, 21, 37, 18, 0, 5, 7, 5, 30, 30, 0, 0, 19, 16, 13, 16, 26, 35, 35, 16, 15, 23, 19, 6, 13, 24, 28, 26, 32, 29, 111, 
    0, 20, 25, 32, 20, 0, 7, 12, 10, 43, 47, 0, 0, 16, 18, 14, 19, 25, 34, 31, 13, 18, 25, 18, 17, 14, 14, 20, 28, 29, 29, 113, 
    0, 22, 29, 33, 22, 0, 4, 14, 17, 43, 57, 5, 0, 12, 20, 19, 22, 26, 36, 22, 14, 20, 26, 19, 25, 22, 15, 12, 21, 29, 32, 122, 
    1, 23, 31, 37, 27, 0, 0, 10, 20, 30, 38, 22, 15, 19, 21, 24, 25, 28, 37, 15, 18, 21, 25, 24, 29, 29, 20, 11, 13, 25, 29, 121, 
    1, 21, 26, 42, 33, 0, 0, 8, 19, 22, 21, 22, 27, 28, 21, 28, 29, 34, 32, 16, 22, 20, 23, 26, 33, 30, 21, 17, 15, 19, 27, 116, 
    1, 19, 19, 41, 46, 0, 0, 5, 15, 18, 19, 28, 30, 26, 20, 25, 32, 38, 25, 21, 22, 19, 19, 26, 31, 29, 25, 21, 16, 18, 26, 119, 
    4, 16, 15, 30, 55, 14, 0, 0, 13, 14, 20, 36, 34, 24, 13, 15, 31, 34, 24, 24, 22, 20, 19, 26, 26, 29, 24, 21, 17, 21, 25, 121, 
    0, 4, 0, 1, 25, 14, 0, 0, 0, 0, 0, 14, 22, 18, 6, 0, 10, 13, 9, 8, 8, 3, 1, 5, 7, 9, 7, 4, 0, 1, 4, 75, 
    
    -- channel=135
    70, 46, 45, 84, 104, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 46, 57, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 48, 50, 97, 152, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 84, 96, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 48, 48, 80, 155, 66, 0, 0, 14, 6, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 102, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 47, 47, 67, 142, 92, 0, 0, 45, 20, 0, 0, 13, 10, 4, 5, 0, 0, 0, 0, 0, 102, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    81, 47, 47, 59, 119, 112, 0, 3, 63, 42, 0, 0, 0, 15, 19, 25, 4, 0, 0, 0, 17, 84, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    81, 44, 48, 53, 100, 132, 19, 0, 55, 58, 3, 0, 0, 4, 28, 32, 15, 6, 0, 23, 49, 55, 12, 10, 3, 0, 0, 0, 0, 0, 0, 0, 
    97, 12, 39, 68, 114, 126, 20, 0, 38, 66, 12, 0, 0, 0, 19, 16, 8, 30, 15, 54, 76, 29, 0, 25, 17, 0, 0, 0, 0, 0, 0, 0, 
    162, 0, 5, 61, 106, 80, 0, 0, 21, 77, 27, 0, 0, 0, 0, 0, 0, 31, 24, 57, 87, 28, 0, 37, 23, 0, 0, 0, 0, 11, 16, 0, 
    218, 0, 0, 31, 71, 31, 0, 0, 8, 84, 43, 8, 0, 0, 0, 0, 0, 31, 24, 49, 83, 40, 4, 39, 18, 0, 0, 0, 0, 16, 34, 0, 
    260, 0, 0, 16, 29, 0, 0, 0, 9, 77, 44, 17, 5, 0, 0, 0, 0, 36, 24, 43, 76, 41, 26, 37, 3, 0, 0, 0, 0, 9, 32, 0, 
    275, 0, 0, 5, 12, 0, 0, 0, 21, 60, 27, 14, 4, 0, 0, 0, 13, 38, 18, 40, 72, 36, 39, 44, 0, 0, 0, 0, 0, 0, 16, 0, 
    278, 0, 0, 0, 10, 0, 0, 0, 16, 42, 16, 6, 9, 0, 0, 0, 36, 37, 5, 38, 57, 30, 43, 54, 6, 0, 0, 0, 0, 0, 2, 0, 
    278, 0, 0, 0, 2, 0, 0, 0, 0, 16, 14, 18, 24, 0, 0, 10, 39, 25, 0, 34, 33, 31, 52, 53, 9, 0, 0, 0, 0, 0, 0, 0, 
    278, 0, 0, 0, 0, 0, 0, 29, 0, 4, 9, 23, 35, 0, 0, 26, 57, 8, 0, 39, 27, 26, 55, 49, 6, 0, 0, 0, 0, 0, 2, 0, 
    280, 0, 0, 0, 0, 0, 0, 69, 0, 0, 0, 6, 21, 0, 0, 16, 61, 14, 0, 28, 36, 8, 31, 51, 17, 0, 0, 0, 0, 0, 8, 0, 
    282, 0, 0, 0, 0, 0, 0, 90, 0, 0, 0, 9, 2, 6, 2, 0, 20, 45, 0, 0, 50, 3, 0, 22, 55, 33, 5, 0, 0, 0, 12, 0, 
    285, 0, 0, 0, 9, 0, 0, 68, 32, 0, 0, 8, 0, 2, 16, 0, 0, 57, 23, 0, 51, 19, 0, 0, 48, 69, 34, 0, 0, 18, 16, 0, 
    289, 0, 0, 0, 24, 0, 0, 26, 37, 8, 2, 12, 0, 0, 8, 0, 0, 29, 53, 0, 36, 25, 0, 0, 7, 52, 55, 6, 0, 37, 32, 0, 
    293, 0, 0, 0, 28, 11, 0, 1, 12, 20, 16, 13, 0, 0, 0, 0, 0, 0, 48, 7, 21, 8, 0, 0, 0, 12, 48, 13, 0, 26, 39, 0, 
    298, 0, 0, 0, 27, 11, 0, 3, 0, 11, 19, 12, 8, 15, 0, 0, 0, 0, 1, 26, 1, 0, 0, 11, 0, 0, 24, 0, 0, 13, 29, 0, 
    300, 0, 0, 0, 17, 21, 0, 0, 0, 0, 2, 0, 3, 41, 10, 0, 7, 0, 0, 9, 0, 0, 3, 21, 2, 5, 4, 0, 0, 7, 10, 0, 
    301, 0, 0, 0, 2, 36, 10, 0, 0, 0, 0, 0, 0, 43, 18, 7, 17, 0, 0, 0, 0, 6, 25, 16, 10, 11, 0, 0, 0, 0, 0, 0, 
    299, 0, 0, 0, 0, 46, 24, 0, 0, 0, 0, 0, 0, 25, 12, 4, 13, 0, 0, 0, 0, 29, 30, 6, 14, 17, 0, 0, 0, 0, 0, 0, 
    296, 0, 0, 0, 0, 45, 32, 2, 0, 0, 0, 0, 6, 16, 0, 0, 3, 0, 0, 0, 0, 35, 22, 0, 15, 25, 0, 0, 0, 0, 0, 0, 
    294, 0, 0, 0, 0, 35, 36, 5, 0, 0, 0, 0, 57, 27, 0, 0, 0, 0, 0, 0, 0, 33, 13, 0, 16, 25, 0, 0, 0, 0, 0, 0, 
    292, 0, 0, 0, 0, 26, 40, 9, 0, 0, 0, 0, 89, 37, 0, 0, 0, 0, 0, 0, 5, 32, 6, 0, 15, 10, 1, 9, 6, 1, 0, 0, 
    291, 0, 0, 0, 0, 20, 48, 16, 0, 0, 0, 0, 66, 17, 0, 0, 0, 0, 0, 0, 18, 32, 4, 0, 13, 0, 4, 22, 26, 8, 0, 0, 
    286, 0, 0, 0, 0, 17, 57, 26, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 36, 27, 5, 4, 8, 0, 5, 30, 33, 15, 0, 0, 
    276, 0, 0, 0, 0, 11, 67, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 43, 16, 11, 11, 1, 0, 9, 28, 26, 15, 0, 0, 
    259, 0, 2, 0, 0, 0, 75, 53, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 24, 34, 12, 20, 15, 0, 0, 10, 17, 15, 15, 9, 0, 
    236, 0, 15, 8, 0, 0, 68, 74, 10, 0, 0, 0, 0, 0, 4, 25, 11, 0, 3, 31, 19, 15, 25, 16, 0, 0, 5, 12, 17, 22, 11, 0, 
    157, 5, 27, 20, 1, 0, 50, 70, 28, 13, 13, 0, 0, 0, 22, 37, 33, 15, 25, 34, 23, 25, 33, 25, 15, 21, 17, 20, 26, 32, 24, 0, 
    
    -- channel=136
    5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    
    -- channel=137
    3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 11, 0, 0, 0, 0, 0, 0, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 10, 2, 0, 0, 0, 0, 0, 36, 64, 42, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 9, 9, 0, 0, 0, 0, 0, 46, 91, 85, 48, 21, 0, 0, 0, 0, 0, 0, 0, 10, 28, 39, 22, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 8, 0, 0, 0, 0, 0, 45, 100, 110, 74, 35, 8, 0, 0, 0, 0, 3, 20, 38, 55, 57, 45, 39, 39, 35, 30, 23, 16, 8, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 43, 97, 118, 92, 51, 24, 4, 0, 3, 5, 13, 38, 61, 70, 67, 63, 66, 79, 77, 71, 64, 51, 48, 42, 
    0, 0, 0, 4, 5, 8, 0, 0, 40, 89, 113, 100, 72, 44, 29, 20, 13, 17, 19, 40, 70, 72, 69, 73, 85, 95, 89, 76, 63, 55, 60, 58, 
    14, 2, 0, 5, 25, 30, 8, 0, 31, 78, 103, 102, 87, 64, 48, 33, 24, 24, 28, 42, 67, 70, 62, 74, 90, 90, 77, 57, 36, 37, 54, 58, 
    20, 21, 14, 21, 40, 33, 8, 0, 21, 68, 97, 100, 89, 73, 55, 39, 33, 34, 37, 48, 62, 64, 57, 71, 83, 79, 58, 32, 11, 14, 38, 51, 
    23, 29, 29, 38, 42, 31, 10, 2, 23, 67, 94, 98, 86, 69, 51, 42, 36, 43, 47, 55, 64, 59, 58, 72, 81, 78, 56, 22, 3, 1, 14, 40, 
    23, 28, 30, 36, 35, 27, 11, 2, 28, 68, 88, 93, 83, 63, 48, 43, 49, 57, 61, 63, 73, 62, 60, 76, 87, 84, 65, 32, 6, 0, 0, 26, 
    16, 20, 22, 23, 16, 10, 5, 0, 27, 60, 75, 83, 79, 64, 54, 52, 65, 75, 74, 73, 81, 69, 62, 77, 88, 89, 78, 55, 23, 10, 6, 23, 
    12, 13, 13, 13, 0, 0, 0, 2, 33, 57, 72, 82, 83, 75, 64, 66, 72, 83, 77, 81, 83, 71, 65, 70, 78, 83, 86, 75, 49, 35, 30, 37, 
    13, 14, 13, 10, 0, 0, 0, 11, 47, 69, 75, 81, 92, 88, 73, 70, 75, 70, 65, 76, 73, 62, 54, 54, 59, 72, 84, 80, 70, 53, 51, 56, 
    17, 16, 16, 11, 0, 0, 0, 21, 59, 82, 87, 87, 95, 100, 85, 56, 58, 48, 38, 49, 55, 44, 22, 20, 30, 51, 70, 72, 68, 55, 58, 60, 
    20, 15, 14, 10, 7, 0, 0, 35, 74, 94, 100, 99, 97, 100, 92, 57, 29, 24, 14, 18, 37, 29, 1, 0, 0, 20, 41, 47, 42, 43, 52, 55, 
    25, 21, 13, 15, 18, 14, 6, 41, 83, 101, 105, 111, 109, 106, 99, 70, 14, 3, 2, 2, 17, 17, 0, 0, 0, 0, 11, 15, 13, 22, 38, 47, 
    29, 31, 18, 25, 34, 41, 41, 49, 77, 96, 102, 116, 119, 115, 108, 85, 29, 0, 5, 2, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 18, 35, 
    33, 41, 29, 35, 51, 57, 60, 58, 65, 82, 89, 101, 113, 113, 111, 99, 64, 19, 16, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    38, 49, 42, 43, 61, 66, 64, 64, 62, 72, 74, 78, 85, 88, 98, 93, 82, 50, 21, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    42, 55, 51, 47, 61, 70, 70, 66, 67, 71, 67, 62, 56, 61, 74, 77, 81, 66, 26, 4, 0, 0, 0, 0, 5, 8, 5, 0, 0, 0, 0, 0, 
    42, 56, 53, 46, 55, 70, 82, 79, 77, 75, 68, 52, 41, 47, 57, 62, 67, 58, 24, 0, 0, 0, 0, 6, 16, 17, 10, 0, 0, 0, 0, 0, 
    40, 51, 48, 41, 46, 68, 89, 94, 89, 75, 56, 41, 31, 39, 49, 51, 51, 42, 17, 0, 0, 0, 0, 6, 15, 17, 12, 0, 0, 0, 0, 0, 
    40, 46, 38, 33, 34, 61, 89, 99, 93, 66, 31, 15, 15, 31, 39, 35, 33, 25, 7, 0, 0, 0, 0, 3, 8, 15, 8, 0, 0, 0, 0, 0, 
    38, 41, 27, 18, 19, 48, 82, 96, 88, 56, 10, 0, 0, 20, 25, 17, 12, 8, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    36, 36, 18, 2, 2, 32, 73, 92, 83, 57, 7, 0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 29, 12, 0, 0, 22, 68, 95, 87, 65, 27, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    25, 20, 7, 0, 0, 18, 67, 100, 95, 72, 47, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    17, 11, 4, 0, 0, 12, 64, 98, 98, 76, 57, 34, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 1, 0, 0, 0, 1, 51, 87, 91, 74, 56, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 13, 41, 43, 33, 23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 79, 146, 138, 126, 116, 109, 115, 125, 126, 123, 120, 122, 129, 124, 91, 41, 30, 56, 118, 164, 161, 152, 150, 149, 151, 148, 142, 140, 0, 
    0, 0, 0, 129, 233, 213, 188, 184, 186, 186, 189, 197, 197, 194, 199, 210, 212, 183, 110, 65, 100, 209, 271, 255, 241, 237, 235, 238, 233, 225, 219, 0, 
    0, 0, 0, 96, 227, 216, 179, 194, 211, 210, 197, 208, 221, 221, 227, 238, 244, 218, 140, 70, 120, 255, 301, 272, 259, 252, 248, 249, 245, 238, 232, 0, 
    0, 0, 0, 61, 202, 206, 163, 200, 244, 245, 212, 200, 212, 217, 233, 247, 253, 234, 163, 92, 160, 291, 322, 296, 284, 274, 267, 262, 255, 247, 239, 0, 
    0, 0, 0, 31, 164, 195, 157, 200, 267, 284, 236, 190, 186, 187, 207, 227, 229, 207, 167, 141, 215, 302, 315, 305, 301, 292, 290, 290, 283, 275, 267, 0, 
    0, 0, 0, 10, 135, 207, 182, 210, 279, 307, 262, 189, 152, 156, 178, 187, 190, 171, 162, 198, 272, 310, 311, 318, 318, 314, 315, 315, 309, 303, 300, 9, 
    21, 0, 0, 43, 177, 248, 213, 211, 278, 313, 284, 219, 165, 156, 166, 153, 155, 153, 165, 237, 304, 297, 304, 340, 344, 344, 344, 328, 319, 324, 330, 20, 
    139, 63, 61, 132, 234, 279, 228, 188, 251, 305, 297, 257, 212, 192, 179, 146, 145, 155, 171, 250, 315, 294, 308, 356, 359, 351, 342, 311, 304, 332, 352, 26, 
    238, 148, 152, 223, 291, 291, 220, 168, 226, 290, 298, 282, 256, 229, 194, 138, 144, 160, 173, 243, 306, 303, 331, 377, 376, 366, 336, 287, 281, 319, 357, 30, 
    323, 225, 227, 279, 304, 284, 210, 162, 222, 287, 297, 292, 278, 243, 190, 146, 149, 167, 172, 231, 286, 301, 349, 386, 378, 368, 324, 271, 269, 302, 345, 30, 
    352, 272, 270, 291, 304, 286, 211, 177, 241, 290, 293, 292, 272, 226, 171, 139, 163, 177, 175, 229, 275, 295, 356, 387, 382, 373, 326, 270, 262, 282, 316, 24, 
    358, 283, 276, 289, 301, 280, 221, 202, 251, 282, 275, 273, 259, 214, 165, 158, 198, 195, 191, 237, 266, 286, 354, 392, 388, 379, 343, 288, 265, 271, 294, 17, 
    362, 287, 275, 285, 278, 251, 237, 225, 237, 244, 236, 252, 247, 203, 178, 201, 232, 215, 212, 240, 252, 281, 351, 390, 388, 384, 365, 321, 278, 275, 300, 19, 
    362, 287, 273, 279, 248, 209, 249, 255, 247, 247, 240, 261, 263, 208, 172, 222, 257, 225, 224, 254, 257, 283, 352, 387, 386, 385, 383, 352, 298, 292, 321, 26, 
    360, 283, 271, 279, 233, 172, 253, 285, 258, 255, 250, 260, 263, 228, 200, 230, 264, 235, 223, 257, 262, 272, 321, 369, 379, 383, 389, 363, 316, 317, 349, 31, 
    361, 272, 261, 271, 234, 160, 241, 309, 285, 266, 267, 269, 254, 236, 218, 206, 236, 245, 212, 236, 264, 243, 233, 275, 333, 368, 381, 350, 319, 342, 363, 30, 
    364, 258, 241, 254, 245, 193, 237, 312, 311, 298, 301, 283, 258, 257, 245, 189, 190, 244, 208, 218, 269, 237, 191, 193, 250, 308, 328, 304, 307, 355, 368, 28, 
    373, 256, 228, 251, 266, 238, 250, 300, 317, 310, 324, 323, 287, 277, 268, 193, 154, 224, 208, 200, 258, 230, 167, 158, 195, 249, 273, 251, 270, 336, 361, 25, 
    381, 269, 236, 262, 289, 282, 280, 290, 305, 315, 327, 327, 310, 300, 275, 224, 172, 197, 217, 219, 251, 217, 175, 158, 158, 206, 242, 227, 234, 280, 320, 16, 
    392, 290, 253, 271, 303, 299, 293, 293, 297, 308, 315, 308, 310, 310, 292, 273, 234, 208, 229, 236, 227, 188, 186, 190, 176, 202, 226, 203, 200, 232, 266, 5, 
    396, 310, 274, 272, 301, 308, 301, 297, 299, 308, 296, 269, 285, 304, 289, 291, 279, 235, 236, 230, 191, 173, 192, 208, 207, 219, 218, 191, 183, 197, 210, 0, 
    397, 321, 287, 261, 291, 317, 314, 310, 312, 312, 289, 244, 260, 293, 287, 295, 296, 258, 232, 192, 162, 180, 208, 217, 228, 231, 207, 185, 177, 173, 163, 0, 
    394, 324, 300, 255, 279, 324, 328, 325, 330, 321, 287, 244, 259, 287, 283, 289, 291, 268, 218, 160, 157, 200, 218, 219, 241, 236, 204, 190, 178, 163, 149, 0, 
    388, 320, 304, 256, 273, 327, 336, 329, 328, 306, 254, 239, 268, 286, 281, 280, 279, 255, 200, 148, 167, 212, 214, 207, 235, 237, 208, 189, 176, 159, 151, 0, 
    383, 311, 299, 261, 270, 322, 336, 326, 321, 266, 188, 211, 276, 287, 274, 272, 264, 234, 183, 149, 178, 210, 202, 197, 222, 223, 199, 188, 174, 159, 151, 0, 
    378, 303, 288, 256, 261, 312, 333, 324, 313, 242, 142, 188, 280, 277, 255, 252, 240, 209, 167, 149, 177, 200, 185, 185, 197, 187, 179, 182, 181, 175, 164, 0, 
    374, 294, 274, 246, 248, 298, 332, 326, 305, 238, 157, 207, 274, 256, 230, 222, 207, 184, 146, 138, 171, 187, 174, 175, 172, 157, 157, 175, 192, 186, 172, 0, 
    366, 282, 263, 232, 229, 285, 332, 332, 304, 254, 211, 234, 255, 224, 206, 200, 182, 159, 124, 134, 170, 179, 168, 170, 158, 135, 145, 178, 198, 195, 180, 0, 
    344, 262, 255, 224, 207, 265, 326, 332, 305, 276, 260, 256, 229, 195, 191, 180, 160, 133, 108, 134, 165, 165, 166, 170, 151, 136, 151, 177, 193, 192, 176, 0, 
    313, 240, 251, 228, 191, 236, 311, 328, 306, 288, 279, 241, 187, 159, 163, 164, 144, 112, 108, 141, 157, 158, 171, 169, 154, 148, 158, 169, 178, 181, 176, 0, 
    270, 209, 231, 221, 173, 197, 282, 315, 298, 278, 254, 200, 139, 109, 121, 135, 124, 107, 118, 143, 143, 153, 170, 168, 155, 147, 150, 157, 170, 181, 178, 0, 
    114, 69, 86, 82, 50, 57, 112, 134, 118, 108, 97, 59, 21, 12, 23, 35, 29, 17, 31, 41, 36, 44, 55, 50, 45, 46, 42, 40, 49, 60, 60, 0, 
    
    -- channel=139
    59, 61, 49, 17, 29, 27, 27, 34, 35, 33, 34, 32, 30, 31, 29, 28, 31, 40, 49, 44, 52, 20, 9, 21, 19, 22, 21, 21, 25, 26, 26, 103, 
    53, 58, 44, 0, 0, 10, 10, 14, 12, 7, 5, 8, 9, 7, 2, 0, 3, 14, 29, 26, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 120, 
    53, 56, 52, 0, 0, 13, 15, 9, 6, 5, 0, 0, 2, 0, 0, 0, 0, 10, 45, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 121, 
    53, 55, 56, 10, 0, 16, 20, 2, 0, 1, 5, 0, 8, 15, 7, 2, 0, 8, 40, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 
    53, 53, 54, 27, 0, 14, 18, 0, 0, 0, 12, 12, 11, 20, 17, 17, 16, 25, 37, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 123, 
    53, 55, 56, 41, 0, 0, 5, 0, 0, 0, 15, 25, 18, 15, 6, 16, 24, 34, 28, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 
    35, 42, 50, 24, 0, 0, 0, 0, 0, 0, 7, 20, 15, 1, 2, 17, 13, 26, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 139, 
    8, 0, 0, 0, 0, 0, 7, 12, 0, 0, 0, 11, 15, 0, 4, 19, 6, 13, 5, 0, 0, 6, 0, 0, 0, 0, 0, 4, 0, 0, 0, 144, 
    10, 22, 0, 0, 0, 0, 16, 19, 0, 0, 0, 4, 10, 11, 15, 32, 22, 17, 12, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 150, 
    0, 14, 2, 0, 0, 0, 25, 22, 0, 0, 0, 0, 0, 15, 29, 37, 15, 17, 14, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 153, 
    0, 0, 0, 0, 0, 0, 26, 10, 0, 0, 0, 0, 2, 21, 37, 37, 13, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 147, 
    0, 0, 0, 0, 0, 4, 21, 2, 0, 0, 3, 3, 12, 19, 24, 13, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 131, 
    0, 0, 0, 0, 0, 12, 13, 4, 0, 9, 23, 10, 10, 25, 21, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 123, 
    0, 0, 0, 0, 12, 15, 0, 6, 0, 0, 0, 0, 0, 17, 22, 6, 0, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 132, 
    0, 0, 0, 0, 20, 18, 0, 0, 0, 0, 0, 0, 4, 18, 5, 0, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 139, 
    0, 0, 4, 0, 22, 28, 0, 0, 0, 2, 6, 1, 0, 14, 16, 2, 0, 17, 15, 0, 9, 12, 7, 9, 10, 0, 0, 0, 0, 0, 0, 143, 
    0, 3, 5, 0, 11, 24, 0, 0, 0, 0, 0, 0, 0, 0, 7, 32, 0, 0, 31, 0, 0, 12, 12, 0, 0, 9, 12, 18, 0, 0, 0, 144, 
    0, 8, 1, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 12, 0, 31, 5, 0, 23, 30, 6, 0, 0, 4, 19, 1, 0, 0, 150, 
    0, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 15, 18, 0, 7, 0, 0, 23, 27, 29, 16, 0, 0, 3, 0, 0, 0, 161, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 5, 0, 0, 0, 8, 24, 12, 15, 16, 0, 0, 15, 10, 0, 0, 146, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 7, 0, 9, 16, 0, 6, 25, 22, 1, 3, 4, 0, 8, 21, 15, 7, 2, 124, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 0, 0, 0, 0, 16, 9, 26, 26, 11, 0, 0, 0, 4, 11, 15, 13, 19, 28, 117, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 4, 9, 0, 0, 0, 0, 0, 0, 20, 34, 13, 0, 2, 4, 0, 4, 12, 9, 15, 18, 21, 104, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 18, 18, 0, 0, 0, 0, 0, 5, 27, 30, 6, 0, 8, 10, 0, 11, 15, 14, 21, 18, 15, 104, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 18, 42, 14, 0, 0, 0, 0, 5, 17, 29, 27, 7, 2, 13, 10, 0, 15, 22, 21, 18, 22, 24, 112, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 23, 38, 0, 0, 3, 5, 3, 11, 21, 30, 28, 7, 8, 18, 14, 10, 20, 25, 20, 15, 15, 13, 103, 
    0, 0, 1, 7, 0, 0, 0, 0, 0, 21, 26, 0, 0, 7, 12, 11, 20, 24, 35, 29, 10, 12, 20, 13, 21, 23, 17, 13, 13, 12, 13, 107, 
    0, 0, 4, 10, 2, 0, 0, 0, 0, 9, 13, 0, 0, 14, 14, 14, 19, 25, 40, 19, 8, 13, 17, 12, 22, 26, 17, 4, 4, 12, 18, 116, 
    0, 7, 7, 14, 8, 0, 0, 0, 0, 0, 0, 0, 12, 19, 13, 18, 25, 33, 39, 13, 13, 18, 18, 15, 24, 24, 11, 3, 6, 15, 22, 116, 
    0, 9, 3, 15, 14, 0, 0, 0, 0, 0, 0, 8, 29, 35, 25, 27, 30, 38, 27, 11, 17, 16, 12, 16, 23, 17, 10, 12, 15, 15, 16, 109, 
    1, 14, 8, 21, 32, 0, 0, 0, 0, 3, 12, 35, 46, 44, 35, 34, 40, 38, 19, 17, 21, 16, 12, 19, 21, 23, 24, 22, 13, 8, 12, 113, 
    72, 96, 92, 103, 119, 91, 73, 99, 116, 117, 116, 122, 112, 93, 77, 80, 94, 95, 90, 91, 93, 90, 93, 101, 100, 100, 96, 94, 93, 98, 103, 159, 
    
    -- channel=140
    26, 26, 37, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 18, 26, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 18, 22, 35, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 17, 19, 32, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 16, 16, 26, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 16, 15, 21, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 9, 14, 17, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=141
    0, 0, 0, 32, 144, 246, 264, 252, 242, 233, 234, 242, 247, 246, 246, 250, 249, 218, 153, 100, 88, 158, 230, 298, 316, 305, 306, 306, 304, 300, 293, 132, 
    0, 0, 0, 104, 274, 414, 452, 438, 434, 421, 417, 421, 431, 439, 440, 450, 464, 441, 353, 257, 224, 308, 435, 539, 548, 534, 532, 530, 526, 518, 506, 259, 
    0, 0, 0, 69, 245, 389, 448, 446, 463, 473, 452, 450, 459, 480, 492, 506, 528, 516, 434, 313, 265, 354, 503, 598, 590, 575, 567, 562, 556, 548, 537, 279, 
    0, 0, 0, 34, 204, 338, 412, 437, 490, 539, 510, 475, 459, 476, 503, 527, 553, 550, 480, 362, 330, 426, 578, 651, 638, 622, 606, 593, 584, 572, 557, 293, 
    0, 0, 0, 7, 158, 281, 369, 420, 510, 596, 580, 513, 451, 430, 456, 485, 515, 507, 460, 388, 407, 502, 623, 665, 665, 657, 649, 639, 632, 621, 604, 323, 
    0, 0, 0, 0, 123, 255, 364, 435, 530, 626, 636, 548, 436, 376, 376, 402, 436, 422, 411, 415, 488, 583, 656, 676, 690, 699, 698, 692, 687, 676, 664, 366, 
    0, 6, 0, 21, 162, 322, 429, 470, 538, 628, 667, 592, 474, 389, 354, 350, 363, 347, 371, 438, 547, 627, 670, 689, 729, 761, 759, 746, 735, 716, 719, 411, 
    78, 176, 125, 160, 291, 455, 506, 483, 517, 595, 663, 633, 553, 473, 417, 371, 344, 330, 360, 451, 571, 645, 683, 710, 769, 800, 782, 751, 719, 710, 740, 441, 
    211, 375, 324, 358, 477, 576, 549, 478, 478, 548, 639, 654, 620, 563, 496, 405, 361, 335, 368, 451, 557, 640, 695, 744, 811, 828, 788, 728, 666, 666, 725, 439, 
    325, 549, 516, 539, 598, 626, 555, 471, 452, 528, 625, 655, 645, 603, 525, 430, 373, 353, 377, 443, 528, 621, 696, 763, 825, 828, 772, 692, 622, 622, 691, 417, 
    362, 624, 611, 621, 643, 643, 568, 487, 474, 550, 628, 650, 634, 587, 496, 407, 369, 367, 391, 443, 516, 607, 693, 767, 835, 836, 778, 688, 613, 592, 640, 379, 
    370, 642, 630, 634, 645, 640, 576, 511, 512, 572, 618, 629, 609, 555, 469, 403, 399, 409, 436, 463, 522, 596, 677, 764, 841, 848, 801, 717, 636, 589, 607, 344, 
    372, 649, 630, 630, 616, 605, 568, 525, 537, 547, 560, 573, 560, 525, 467, 436, 459, 479, 488, 490, 534, 585, 661, 761, 836, 853, 828, 767, 680, 623, 613, 341, 
    371, 647, 622, 622, 581, 551, 542, 535, 577, 554, 548, 559, 563, 534, 473, 468, 501, 528, 524, 524, 551, 590, 670, 758, 831, 851, 851, 816, 740, 682, 656, 378, 
    371, 647, 617, 620, 568, 507, 517, 545, 614, 587, 566, 568, 579, 554, 505, 498, 531, 543, 533, 540, 551, 593, 646, 725, 797, 839, 856, 837, 782, 730, 718, 426, 
    373, 640, 605, 603, 565, 488, 505, 558, 650, 642, 621, 605, 595, 568, 526, 490, 513, 516, 510, 531, 541, 564, 558, 593, 667, 760, 824, 817, 777, 746, 755, 452, 
    377, 629, 581, 565, 558, 514, 522, 583, 668, 690, 676, 644, 620, 592, 564, 506, 474, 476, 477, 517, 528, 540, 510, 463, 500, 606, 699, 720, 713, 727, 765, 461, 
    387, 631, 567, 543, 558, 559, 566, 605, 668, 697, 711, 708, 681, 647, 612, 530, 442, 437, 437, 485, 505, 517, 481, 393, 392, 475, 557, 589, 611, 663, 735, 449, 
    398, 650, 583, 560, 582, 619, 629, 634, 665, 690, 721, 735, 727, 700, 655, 582, 471, 435, 435, 476, 515, 516, 480, 397, 375, 409, 462, 503, 527, 570, 651, 393, 
    409, 680, 617, 597, 615, 652, 663, 656, 661, 674, 693, 705, 716, 706, 689, 652, 568, 507, 486, 490, 517, 486, 454, 421, 421, 431, 457, 472, 471, 485, 544, 320, 
    417, 706, 655, 626, 633, 661, 676, 672, 666, 672, 666, 649, 649, 654, 672, 672, 640, 590, 549, 512, 497, 444, 421, 434, 458, 475, 487, 472, 445, 432, 454, 251, 
    420, 720, 677, 633, 630, 654, 687, 695, 693, 695, 674, 622, 595, 603, 640, 663, 666, 637, 581, 503, 448, 404, 421, 459, 493, 507, 499, 464, 424, 407, 395, 195, 
    416, 721, 691, 633, 623, 647, 702, 727, 730, 725, 693, 627, 590, 595, 624, 643, 649, 635, 570, 475, 404, 395, 442, 483, 514, 518, 507, 465, 423, 401, 368, 167, 
    409, 711, 689, 633, 619, 645, 711, 744, 744, 719, 664, 612, 586, 609, 633, 634, 632, 611, 541, 444, 388, 407, 454, 479, 502, 515, 512, 468, 430, 392, 359, 168, 
    403, 698, 675, 628, 610, 641, 704, 740, 738, 675, 586, 535, 542, 610, 638, 625, 611, 581, 507, 420, 393, 415, 449, 459, 476, 493, 491, 459, 425, 390, 366, 175, 
    398, 686, 654, 609, 589, 624, 686, 728, 721, 639, 511, 453, 491, 588, 616, 590, 567, 533, 463, 400, 387, 405, 427, 433, 433, 440, 435, 420, 413, 407, 389, 185, 
    394, 675, 631, 585, 557, 594, 665, 719, 712, 627, 501, 453, 492, 570, 569, 531, 505, 469, 406, 367, 358, 384, 406, 405, 394, 388, 372, 378, 403, 416, 406, 199, 
    384, 658, 610, 557, 522, 559, 642, 716, 714, 646, 556, 518, 529, 540, 511, 476, 450, 412, 353, 330, 330, 374, 389, 387, 372, 349, 333, 354, 399, 428, 427, 217, 
    361, 622, 582, 533, 493, 523, 612, 705, 713, 668, 616, 586, 551, 505, 463, 429, 406, 359, 308, 294, 313, 360, 372, 377, 363, 342, 329, 352, 396, 424, 420, 212, 
    323, 567, 545, 519, 473, 488, 573, 675, 705, 679, 643, 591, 519, 441, 395, 382, 366, 320, 283, 279, 315, 348, 364, 374, 371, 351, 343, 360, 386, 401, 402, 202, 
    271, 492, 483, 486, 440, 438, 514, 621, 676, 660, 617, 544, 445, 344, 302, 303, 304, 286, 269, 282, 310, 331, 351, 371, 369, 349, 346, 351, 366, 383, 396, 204, 
    108, 220, 222, 232, 204, 191, 236, 314, 355, 348, 324, 269, 190, 118, 91, 100, 111, 104, 105, 118, 129, 138, 155, 166, 167, 160, 155, 147, 152, 170, 187, 81, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 15, 71, 99, 115, 127, 120, 117, 124, 130, 130, 131, 134, 138, 137, 127, 110, 87, 77, 84, 101, 105, 130, 141, 140, 144, 148, 148, 146, 144, 43, 
    0, 2, 7, 60, 103, 115, 129, 121, 108, 107, 123, 133, 132, 138, 140, 141, 134, 104, 58, 48, 86, 109, 117, 142, 146, 147, 150, 155, 155, 153, 151, 48, 
    0, 3, 4, 45, 97, 109, 125, 116, 95, 95, 98, 115, 106, 103, 112, 123, 129, 118, 92, 69, 84, 104, 128, 153, 159, 159, 158, 157, 154, 149, 145, 41, 
    1, 4, 4, 29, 86, 105, 122, 116, 94, 92, 85, 94, 105, 106, 113, 116, 117, 112, 101, 92, 101, 109, 134, 149, 152, 153, 155, 158, 160, 158, 157, 49, 
    1, 1, 0, 17, 81, 114, 126, 121, 110, 94, 83, 85, 94, 103, 118, 114, 114, 108, 103, 96, 110, 131, 163, 170, 165, 156, 157, 152, 149, 152, 151, 42, 
    24, 20, 12, 40, 106, 126, 112, 108, 110, 99, 96, 89, 89, 96, 91, 95, 110, 98, 100, 99, 96, 116, 148, 163, 160, 158, 158, 151, 151, 156, 157, 40, 
    35, 75, 75, 82, 72, 91, 116, 116, 110, 101, 102, 89, 77, 78, 75, 79, 91, 81, 83, 100, 107, 123, 152, 148, 131, 132, 128, 134, 158, 166, 169, 48, 
    19, 45, 63, 68, 83, 134, 139, 128, 131, 109, 99, 98, 88, 75, 75, 62, 58, 65, 69, 95, 118, 135, 163, 162, 158, 161, 161, 167, 174, 175, 170, 50, 
    89, 115, 97, 107, 140, 151, 131, 124, 124, 111, 111, 115, 108, 92, 79, 72, 84, 71, 75, 96, 109, 131, 152, 167, 176, 170, 171, 180, 178, 185, 188, 53, 
    106, 155, 149, 149, 152, 152, 139, 132, 111, 104, 109, 110, 104, 97, 85, 80, 78, 75, 78, 95, 104, 135, 163, 172, 177, 179, 179, 181, 182, 183, 192, 66, 
    107, 154, 149, 154, 155, 155, 146, 129, 108, 97, 96, 99, 101, 107, 100, 93, 83, 72, 82, 92, 98, 129, 170, 179, 185, 190, 192, 187, 192, 190, 199, 83, 
    116, 168, 158, 160, 158, 152, 146, 124, 117, 104, 95, 108, 106, 86, 81, 85, 80, 67, 86, 81, 91, 121, 155, 175, 186, 189, 190, 186, 185, 192, 201, 80, 
    118, 177, 167, 165, 148, 150, 151, 121, 136, 141, 141, 133, 109, 91, 73, 63, 71, 86, 92, 94, 114, 130, 148, 174, 187, 190, 188, 180, 169, 189, 188, 58, 
    118, 177, 166, 162, 136, 135, 147, 117, 118, 98, 91, 84, 80, 87, 100, 107, 87, 98, 108, 111, 100, 112, 141, 159, 182, 192, 192, 175, 168, 185, 182, 61, 
    119, 176, 159, 150, 123, 102, 124, 112, 116, 106, 94, 103, 112, 90, 69, 70, 92, 97, 105, 117, 98, 114, 128, 141, 153, 176, 185, 179, 184, 184, 186, 68, 
    119, 175, 167, 151, 128, 97, 118, 121, 122, 138, 146, 122, 111, 109, 84, 67, 115, 116, 96, 129, 137, 126, 144, 186, 177, 155, 156, 166, 186, 193, 194, 72, 
    122, 173, 172, 160, 138, 99, 91, 123, 124, 115, 111, 108, 110, 108, 102, 89, 96, 121, 98, 117, 122, 96, 105, 122, 159, 176, 173, 170, 171, 179, 186, 68, 
    125, 173, 164, 155, 133, 113, 101, 118, 134, 121, 116, 108, 96, 100, 98, 92, 89, 123, 114, 118, 119, 107, 109, 83, 91, 136, 152, 152, 162, 168, 171, 55, 
    127, 178, 157, 146, 132, 127, 119, 118, 144, 152, 145, 133, 123, 107, 102, 114, 98, 107, 127, 102, 101, 115, 123, 110, 104, 108, 106, 106, 124, 153, 176, 60, 
    124, 180, 164, 156, 146, 138, 139, 138, 134, 143, 137, 127, 139, 124, 110, 104, 87, 81, 109, 99, 106, 117, 120, 112, 107, 97, 98, 107, 117, 119, 132, 55, 
    123, 179, 165, 155, 154, 142, 137, 146, 138, 129, 124, 128, 139, 133, 128, 126, 121, 109, 103, 103, 115, 115, 106, 107, 105, 105, 111, 113, 106, 94, 97, 41, 
    123, 179, 168, 154, 157, 142, 130, 131, 139, 139, 131, 122, 129, 133, 127, 129, 134, 129, 111, 110, 122, 111, 102, 106, 115, 112, 108, 108, 98, 105, 112, 40, 
    120, 181, 175, 156, 160, 147, 135, 129, 127, 124, 112, 101, 109, 121, 123, 121, 119, 117, 110, 112, 107, 103, 104, 108, 112, 100, 104, 99, 96, 103, 96, 20, 
    120, 180, 179, 165, 161, 153, 141, 138, 134, 114, 97, 113, 112, 120, 129, 124, 119, 114, 112, 101, 99, 106, 109, 112, 111, 102, 101, 101, 106, 89, 79, 18, 
    118, 179, 182, 177, 165, 161, 146, 139, 138, 119, 114, 127, 116, 119, 129, 129, 124, 119, 107, 96, 106, 106, 106, 104, 102, 103, 103, 106, 103, 100, 107, 37, 
    117, 178, 180, 181, 178, 173, 152, 137, 132, 116, 98, 104, 104, 116, 130, 126, 118, 115, 99, 98, 104, 102, 103, 104, 95, 102, 109, 103, 98, 101, 95, 20, 
    114, 175, 177, 179, 177, 176, 159, 139, 134, 122, 87, 70, 87, 121, 126, 122, 119, 108, 94, 107, 101, 101, 104, 102, 95, 91, 92, 103, 106, 96, 91, 21, 
    108, 170, 173, 173, 172, 170, 153, 138, 133, 129, 111, 100, 113, 121, 120, 111, 102, 94, 93, 100, 88, 95, 96, 94, 90, 89, 95, 97, 97, 98, 99, 32, 
    108, 170, 172, 168, 167, 165, 147, 133, 131, 132, 131, 122, 107, 100, 100, 96, 96, 90, 96, 91, 90, 100, 101, 94, 92, 95, 90, 86, 95, 107, 107, 33, 
    104, 160, 159, 158, 150, 154, 145, 123, 124, 124, 113, 100, 103, 100, 93, 91, 83, 84, 88, 79, 89, 94, 94, 92, 95, 82, 78, 91, 107, 107, 98, 21, 
    22, 64, 63, 65, 56, 58, 48, 17, 13, 20, 26, 35, 42, 44, 47, 39, 25, 18, 7, 13, 19, 17, 13, 15, 15, 15, 26, 25, 14, 4, 7, 0, 
    
    -- channel=143
    43, 40, 47, 55, 34, 25, 28, 24, 20, 22, 26, 31, 30, 30, 29, 25, 20, 17, 22, 33, 29, 32, 21, 8, 19, 23, 25, 23, 22, 25, 27, 4, 
    46, 35, 39, 66, 67, 20, 13, 8, 0, 0, 9, 12, 13, 12, 12, 9, 0, 0, 0, 0, 27, 20, 10, 1, 0, 5, 4, 6, 7, 8, 12, 0, 
    47, 35, 38, 57, 73, 27, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 22, 4, 0, 0, 0, 0, 0, 0, 2, 6, 0, 
    48, 35, 37, 48, 73, 39, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 36, 37, 40, 68, 52, 16, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    51, 37, 38, 38, 59, 56, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 31, 38, 40, 44, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 5, 20, 27, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 14, 2, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 3, 0, 0, 0, 0, 1, 8, 3, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 11, 6, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 10, 8, 14, 5, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 
    55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 6, 6, 9, 9, 13, 3, 4, 0, 0, 0, 0, 5, 3, 0, 0, 0, 
    65, 0, 1, 1, 0, 0, 14, 0, 0, 0, 0, 0, 0, 14, 32, 34, 26, 24, 19, 30, 23, 22, 21, 20, 14, 15, 21, 20, 18, 18, 16, 8, 
    
    -- channel=144
    114, 57, 62, 46, 55, 58, 63, 56, 73, 77, 67, 78, 74, 85, 78, 68, 60, 47, 50, 52, 53, 43, 50, 54, 70, 68, 60, 58, 81, 67, 76, 174, 
    0, 0, 1, 0, 0, 1, 26, 6, 11, 25, 8, 6, 2, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 22, 3, 0, 31, 27, 17, 262, 
    0, 0, 0, 0, 0, 0, 45, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 0, 271, 
    0, 0, 0, 0, 0, 0, 52, 11, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 0, 0, 0, 281, 
    0, 0, 0, 0, 0, 0, 80, 34, 0, 35, 0, 6, 27, 0, 5, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 0, 12, 22, 0, 0, 0, 297, 
    0, 0, 0, 0, 0, 0, 119, 83, 0, 31, 6, 7, 20, 5, 19, 18, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 14, 39, 0, 0, 0, 305, 
    0, 0, 0, 0, 0, 0, 91, 108, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 8, 22, 52, 18, 0, 0, 306, 
    0, 0, 0, 0, 0, 0, 47, 88, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 24, 31, 31, 0, 0, 296, 
    0, 0, 0, 0, 9, 0, 41, 79, 0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 29, 46, 36, 0, 273, 
    0, 0, 0, 0, 5, 0, 56, 75, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 41, 42, 14, 0, 266, 
    0, 0, 0, 0, 44, 13, 59, 45, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 290, 
    0, 0, 0, 0, 63, 33, 57, 44, 0, 0, 16, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 307, 
    0, 0, 0, 5, 29, 8, 75, 92, 62, 2, 0, 0, 16, 12, 5, 11, 19, 22, 4, 8, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 307, 
    0, 0, 0, 25, 36, 1, 73, 85, 56, 0, 0, 0, 0, 27, 23, 14, 6, 0, 0, 0, 37, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 307, 
    0, 0, 11, 20, 52, 33, 65, 39, 0, 0, 4, 0, 0, 17, 37, 18, 0, 0, 0, 7, 50, 41, 16, 0, 0, 0, 0, 0, 0, 0, 0, 306, 
    0, 5, 70, 35, 34, 24, 26, 45, 13, 12, 47, 58, 47, 37, 51, 45, 26, 33, 39, 46, 58, 40, 27, 15, 3, 0, 9, 0, 0, 0, 0, 306, 
    0, 27, 126, 67, 7, 0, 0, 68, 64, 34, 65, 69, 72, 36, 51, 77, 74, 87, 96, 72, 92, 87, 61, 82, 51, 16, 13, 0, 0, 0, 0, 307, 
    0, 12, 105, 57, 0, 0, 55, 62, 60, 27, 17, 0, 38, 25, 56, 90, 97, 72, 73, 15, 35, 103, 77, 81, 36, 0, 0, 0, 0, 0, 0, 312, 
    0, 4, 99, 49, 0, 34, 143, 70, 5, 12, 30, 0, 15, 8, 49, 39, 26, 0, 1, 0, 0, 40, 30, 16, 0, 0, 0, 0, 0, 0, 0, 314, 
    0, 19, 115, 60, 0, 50, 165, 83, 0, 9, 75, 67, 35, 13, 30, 0, 0, 23, 10, 0, 2, 13, 8, 15, 0, 17, 71, 36, 0, 0, 0, 311, 
    0, 9, 122, 100, 8, 41, 127, 86, 47, 28, 59, 75, 70, 50, 32, 0, 0, 58, 27, 0, 12, 28, 20, 27, 0, 3, 100, 63, 0, 0, 0, 309, 
    0, 0, 110, 109, 71, 45, 73, 91, 94, 58, 47, 54, 70, 47, 72, 24, 0, 40, 60, 40, 40, 55, 24, 48, 53, 8, 48, 53, 3, 0, 0, 308, 
    0, 0, 102, 78, 59, 88, 58, 88, 109, 81, 74, 29, 21, 0, 87, 99, 25, 12, 70, 56, 38, 57, 0, 12, 119, 21, 0, 12, 37, 0, 0, 302, 
    0, 0, 114, 94, 11, 76, 72, 64, 99, 90, 90, 48, 19, 0, 83, 146, 37, 0, 25, 54, 15, 38, 0, 0, 130, 96, 0, 26, 66, 0, 0, 292, 
    0, 0, 126, 145, 41, 14, 18, 51, 94, 109, 96, 86, 78, 49, 80, 111, 58, 0, 21, 69, 22, 34, 9, 34, 107, 105, 58, 67, 47, 0, 0, 285, 
    0, 0, 95, 136, 62, 0, 0, 55, 90, 110, 107, 96, 93, 94, 88, 82, 91, 47, 0, 0, 0, 1, 2, 104, 101, 70, 76, 69, 30, 0, 0, 275, 
    0, 0, 13, 54, 45, 15, 0, 70, 64, 80, 108, 107, 95, 98, 93, 85, 103, 49, 0, 0, 0, 3, 1, 116, 146, 100, 71, 42, 15, 0, 0, 266, 
    0, 0, 0, 6, 48, 50, 0, 72, 54, 54, 98, 123, 105, 95, 91, 72, 65, 41, 0, 0, 0, 3, 12, 127, 142, 111, 64, 22, 11, 0, 0, 260, 
    0, 0, 0, 13, 33, 57, 0, 61, 62, 52, 87, 117, 103, 87, 84, 69, 48, 41, 31, 23, 7, 0, 0, 136, 134, 92, 61, 27, 13, 0, 0, 254, 
    0, 0, 3, 8, 17, 54, 48, 53, 57, 59, 78, 100, 100, 83, 81, 78, 70, 57, 48, 35, 16, 0, 0, 117, 149, 86, 61, 44, 12, 0, 0, 249, 
    0, 0, 0, 0, 5, 49, 90, 53, 47, 62, 82, 87, 93, 79, 74, 73, 71, 63, 59, 51, 37, 30, 24, 80, 139, 103, 60, 45, 0, 0, 0, 250, 
    0, 0, 0, 0, 0, 20, 106, 71, 47, 59, 70, 65, 62, 56, 51, 53, 50, 36, 30, 33, 26, 22, 22, 49, 92, 85, 45, 0, 0, 0, 0, 244, 
    
    -- channel=145
    122, 253, 250, 253, 251, 241, 228, 208, 188, 188, 191, 189, 198, 215, 224, 240, 261, 278, 282, 278, 273, 270, 268, 266, 257, 247, 237, 243, 229, 224, 207, 111, 
    148, 381, 376, 373, 369, 367, 339, 305, 274, 272, 270, 268, 285, 295, 311, 330, 351, 362, 378, 383, 380, 374, 369, 372, 373, 372, 358, 349, 336, 331, 321, 199, 
    159, 400, 399, 399, 395, 384, 347, 304, 254, 245, 255, 244, 258, 266, 277, 300, 320, 337, 362, 360, 369, 360, 358, 367, 378, 381, 369, 355, 344, 346, 343, 218, 
    162, 406, 405, 406, 406, 389, 330, 258, 188, 172, 188, 180, 187, 192, 191, 208, 230, 241, 272, 289, 313, 337, 348, 358, 377, 376, 368, 359, 346, 347, 352, 230, 
    162, 411, 410, 411, 407, 390, 317, 238, 151, 122, 146, 143, 156, 154, 152, 163, 166, 168, 190, 219, 258, 295, 346, 363, 373, 369, 358, 340, 329, 327, 353, 240, 
    162, 411, 409, 409, 400, 383, 317, 234, 153, 118, 160, 163, 179, 175, 168, 175, 164, 160, 167, 178, 229, 275, 320, 365, 377, 362, 343, 315, 303, 306, 340, 235, 
    161, 409, 410, 404, 386, 365, 308, 241, 165, 139, 212, 239, 236, 227, 202, 188, 183, 171, 175, 183, 205, 262, 298, 330, 363, 356, 336, 324, 305, 300, 317, 208, 
    161, 410, 410, 401, 378, 360, 298, 237, 171, 152, 213, 236, 230, 227, 200, 193, 203, 199, 196, 209, 213, 232, 275, 314, 346, 357, 358, 339, 306, 268, 282, 184, 
    160, 408, 408, 399, 374, 343, 261, 199, 161, 140, 198, 229, 226, 220, 193, 182, 193, 203, 203, 216, 219, 245, 264, 288, 349, 384, 383, 358, 331, 304, 309, 202, 
    157, 402, 406, 397, 354, 299, 201, 171, 137, 124, 163, 174, 169, 179, 165, 162, 173, 184, 186, 196, 205, 230, 258, 281, 329, 368, 385, 391, 375, 363, 359, 228, 
    146, 382, 399, 392, 340, 284, 206, 159, 99, 86, 118, 133, 133, 143, 139, 141, 146, 148, 146, 158, 170, 192, 218, 240, 286, 344, 392, 408, 401, 387, 386, 252, 
    130, 358, 381, 370, 327, 276, 192, 145, 80, 61, 98, 127, 131, 133, 118, 108, 107, 111, 121, 135, 148, 157, 166, 201, 264, 345, 392, 411, 410, 410, 410, 268, 
    116, 329, 338, 326, 288, 251, 180, 152, 98, 106, 118, 136, 138, 135, 127, 110, 109, 125, 150, 163, 164, 153, 155, 189, 234, 285, 335, 370, 387, 407, 411, 267, 
    110, 309, 309, 288, 244, 217, 178, 170, 137, 120, 103, 119, 116, 113, 101, 88, 90, 97, 108, 114, 116, 112, 116, 144, 180, 228, 270, 307, 336, 377, 410, 267, 
    113, 302, 273, 231, 182, 183, 200, 205, 156, 104, 82, 71, 46, 48, 54, 52, 52, 53, 62, 66, 71, 67, 62, 83, 105, 136, 163, 207, 275, 339, 399, 269, 
    105, 277, 225, 186, 150, 182, 210, 197, 131, 96, 81, 94, 89, 90, 78, 58, 35, 6, 0, 6, 11, 21, 13, 0, 15, 46, 96, 151, 219, 305, 387, 269, 
    103, 290, 240, 196, 148, 176, 184, 155, 94, 85, 105, 128, 118, 126, 101, 90, 65, 57, 71, 95, 102, 108, 94, 66, 79, 102, 129, 165, 217, 290, 363, 266, 
    110, 298, 231, 187, 140, 152, 145, 110, 66, 84, 109, 118, 105, 117, 114, 130, 127, 152, 159, 165, 176, 177, 167, 152, 159, 158, 170, 173, 178, 240, 323, 258, 
    117, 308, 238, 192, 138, 132, 119, 85, 36, 65, 78, 81, 78, 97, 90, 130, 159, 172, 150, 150, 156, 178, 171, 142, 162, 159, 165, 142, 129, 213, 300, 250, 
    119, 317, 246, 183, 107, 89, 91, 71, 16, 29, 48, 58, 50, 51, 63, 114, 117, 145, 162, 157, 155, 153, 148, 145, 166, 167, 144, 118, 110, 186, 274, 241, 
    115, 315, 254, 190, 100, 78, 76, 58, 14, 7, 13, 27, 31, 48, 53, 64, 68, 93, 88, 77, 73, 74, 81, 82, 98, 89, 96, 108, 114, 184, 261, 232, 
    112, 314, 255, 199, 101, 70, 80, 51, 27, 13, 0, 18, 40, 84, 85, 83, 47, 63, 110, 129, 111, 101, 127, 140, 137, 131, 94, 113, 133, 176, 244, 225, 
    110, 304, 241, 180, 96, 62, 83, 83, 63, 36, 0, 0, 17, 53, 54, 45, 30, 67, 116, 147, 134, 127, 156, 165, 146, 103, 53, 68, 81, 143, 230, 221, 
    99, 283, 222, 155, 65, 59, 97, 112, 106, 52, 6, 0, 0, 12, 18, 26, 15, 33, 74, 111, 132, 137, 161, 151, 120, 75, 26, 33, 68, 138, 218, 209, 
    83, 262, 220, 172, 106, 87, 138, 131, 119, 70, 24, 0, 0, 0, 0, 2, 0, 0, 62, 163, 237, 248, 249, 186, 147, 76, 5, 14, 46, 121, 207, 195, 
    70, 244, 237, 221, 172, 132, 132, 130, 140, 86, 46, 16, 0, 0, 0, 0, 0, 3, 75, 160, 237, 245, 240, 185, 115, 23, 0, 12, 46, 122, 199, 185, 
    71, 243, 251, 239, 191, 146, 148, 128, 142, 86, 62, 26, 0, 0, 0, 0, 1, 31, 84, 137, 198, 218, 227, 179, 118, 15, 0, 15, 50, 124, 195, 176, 
    78, 250, 244, 227, 205, 172, 160, 119, 118, 78, 65, 38, 6, 0, 0, 0, 9, 27, 45, 79, 139, 173, 192, 156, 108, 12, 0, 10, 47, 124, 194, 175, 
    72, 233, 225, 221, 205, 174, 145, 103, 95, 68, 62, 43, 16, 0, 0, 3, 9, 23, 41, 57, 81, 104, 129, 114, 78, 13, 0, 5, 47, 124, 198, 176, 
    61, 220, 214, 210, 203, 183, 144, 89, 67, 57, 54, 40, 22, 16, 15, 19, 22, 28, 35, 49, 64, 79, 99, 97, 74, 17, 0, 12, 63, 142, 219, 179, 
    58, 222, 222, 227, 221, 197, 145, 97, 46, 41, 42, 41, 43, 40, 39, 43, 43, 49, 62, 77, 88, 95, 105, 101, 86, 49, 30, 51, 105, 182, 238, 180, 
    0, 27, 27, 27, 23, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 35, 9, 
    
    -- channel=146
    85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    147, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    158, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    161, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    161, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 2, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    161, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    161, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 26, 0, 
    160, 0, 0, 0, 0, 0, 0, 0, 9, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 11, 0, 
    161, 0, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    162, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    163, 0, 0, 0, 0, 0, 0, 0, 0, 24, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 
    158, 0, 0, 0, 0, 0, 0, 0, 0, 24, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 30, 9, 0, 0, 0, 0, 0, 0, 
    151, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 38, 17, 0, 0, 0, 0, 0, 0, 
    144, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 13, 12, 6, 25, 40, 0, 0, 0, 
    139, 0, 0, 0, 8, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 42, 17, 16, 68, 20, 0, 0, 
    138, 0, 0, 0, 28, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 17, 10, 0, 0, 0, 19, 43, 13, 0, 45, 35, 0, 0, 
    124, 0, 0, 0, 35, 29, 0, 0, 27, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 3, 18, 0, 0, 20, 62, 4, 0, 
    128, 0, 0, 0, 33, 2, 0, 0, 53, 24, 0, 0, 0, 0, 0, 12, 2, 0, 0, 14, 0, 0, 0, 0, 9, 0, 0, 0, 18, 83, 29, 0, 
    132, 0, 0, 0, 24, 3, 0, 0, 35, 21, 0, 0, 0, 18, 7, 40, 21, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 20, 99, 53, 0, 
    136, 0, 0, 0, 0, 4, 0, 0, 0, 14, 7, 0, 4, 11, 3, 23, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 89, 66, 0, 
    140, 0, 0, 0, 0, 0, 0, 0, 0, 3, 21, 25, 25, 22, 0, 0, 22, 41, 0, 0, 0, 0, 5, 5, 0, 0, 20, 0, 0, 79, 83, 0, 
    143, 0, 0, 0, 0, 1, 0, 0, 0, 0, 9, 36, 34, 38, 0, 0, 30, 80, 0, 0, 0, 0, 12, 9, 0, 0, 54, 4, 0, 99, 97, 0, 
    141, 0, 0, 0, 9, 21, 22, 0, 0, 0, 0, 23, 35, 44, 0, 0, 31, 84, 19, 0, 3, 0, 2, 0, 0, 0, 44, 9, 0, 118, 101, 0, 
    138, 0, 0, 0, 0, 39, 30, 0, 0, 0, 0, 0, 14, 30, 10, 0, 20, 67, 78, 32, 0, 0, 0, 0, 0, 0, 17, 16, 35, 128, 91, 0, 
    129, 0, 0, 0, 0, 2, 36, 0, 0, 0, 0, 0, 0, 15, 19, 24, 13, 41, 109, 60, 0, 0, 0, 0, 0, 0, 20, 37, 49, 110, 79, 0, 
    133, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 15, 19, 26, 21, 44, 105, 58, 0, 0, 0, 0, 0, 0, 33, 54, 46, 90, 69, 0, 
    138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 18, 25, 25, 32, 65, 42, 6, 1, 0, 0, 0, 0, 40, 58, 42, 86, 64, 0, 
    131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 16, 20, 26, 24, 22, 17, 17, 18, 0, 0, 0, 0, 39, 51, 44, 96, 57, 0, 
    126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 11, 11, 16, 19, 16, 17, 16, 6, 0, 0, 0, 36, 46, 61, 99, 31, 0, 
    124, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 5, 8, 2, 3, 13, 13, 5, 6, 5, 0, 0, 0, 0, 24, 46, 72, 70, 0, 0, 
    68, 0, 0, 0, 0, 0, 0, 0, 12, 5, 1, 6, 7, 9, 8, 4, 6, 13, 12, 4, 4, 4, 2, 0, 0, 0, 19, 40, 54, 41, 0, 0, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84, 45, 43, 40, 39, 40, 44, 73, 82, 53, 26, 18, 18, 7, 0, 0, 0, 15, 43, 60, 64, 68, 78, 75, 54, 32, 34, 54, 74, 56, 44, 17, 
    80, 36, 36, 33, 28, 29, 27, 54, 75, 77, 70, 59, 77, 88, 87, 90, 90, 87, 90, 100, 110, 103, 92, 84, 69, 54, 55, 78, 95, 68, 44, 30, 
    84, 38, 39, 39, 41, 43, 49, 59, 74, 74, 73, 84, 80, 103, 124, 134, 142, 135, 125, 138, 131, 123, 95, 72, 76, 79, 83, 107, 114, 95, 63, 34, 
    91, 51, 52, 52, 50, 55, 53, 63, 86, 62, 43, 47, 40, 41, 55, 69, 99, 117, 128, 159, 160, 108, 80, 64, 65, 83, 97, 111, 131, 128, 96, 40, 
    90, 52, 52, 52, 54, 55, 23, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 49, 111, 114, 62, 54, 53, 68, 100, 114, 131, 147, 124, 56, 
    91, 53, 53, 51, 61, 67, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86, 124, 77, 62, 68, 75, 87, 89, 123, 137, 77, 
    91, 52, 52, 53, 53, 56, 39, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 115, 126, 87, 63, 48, 43, 66, 89, 123, 96, 
    91, 52, 52, 51, 40, 42, 42, 2, 3, 17, 46, 71, 63, 4, 0, 0, 0, 0, 0, 0, 0, 0, 37, 78, 63, 47, 40, 42, 63, 66, 64, 57, 
    96, 55, 53, 49, 49, 76, 62, 20, 0, 0, 0, 11, 39, 13, 0, 0, 0, 0, 0, 0, 0, 0, 2, 51, 49, 35, 30, 25, 0, 0, 0, 0, 
    107, 62, 53, 50, 50, 40, 33, 9, 21, 42, 15, 2, 16, 15, 0, 0, 2, 13, 18, 13, 15, 7, 11, 64, 98, 75, 51, 29, 6, 0, 0, 0, 
    110, 73, 62, 59, 41, 0, 0, 0, 27, 61, 45, 4, 0, 0, 4, 8, 16, 24, 20, 15, 31, 53, 55, 67, 83, 81, 60, 49, 51, 51, 52, 31, 
    95, 75, 75, 80, 71, 55, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 61, 56, 61, 79, 87, 76, 56, 51, 52, 31, 
    83, 54, 77, 85, 78, 77, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 46, 70, 96, 128, 139, 135, 100, 56, 51, 31, 
    70, 31, 56, 87, 84, 45, 8, 0, 0, 0, 3, 30, 50, 55, 37, 24, 28, 41, 63, 87, 95, 79, 66, 79, 99, 115, 116, 119, 131, 87, 51, 30, 
    79, 52, 57, 92, 106, 62, 2, 0, 0, 6, 16, 26, 31, 44, 44, 41, 63, 78, 79, 81, 65, 63, 80, 83, 99, 87, 64, 59, 82, 96, 60, 29, 
    81, 56, 44, 34, 48, 54, 70, 90, 34, 0, 0, 0, 0, 0, 0, 0, 12, 28, 24, 15, 0, 0, 18, 49, 45, 26, 0, 0, 12, 74, 66, 29, 
    55, 8, 4, 0, 19, 31, 84, 117, 75, 0, 2, 16, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 69, 78, 31, 
    65, 20, 24, 38, 64, 64, 58, 59, 56, 36, 42, 77, 107, 100, 68, 4, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 54, 84, 97, 92, 36, 
    75, 26, 11, 24, 77, 105, 59, 22, 31, 60, 61, 43, 51, 79, 84, 78, 62, 43, 67, 84, 86, 84, 88, 86, 79, 82, 53, 56, 66, 65, 70, 36, 
    80, 32, 10, 2, 44, 98, 72, 23, 31, 60, 66, 36, 3, 0, 7, 55, 102, 68, 15, 18, 34, 39, 37, 19, 34, 70, 48, 0, 0, 37, 65, 35, 
    77, 37, 21, 5, 4, 12, 47, 26, 23, 48, 69, 69, 24, 0, 0, 11, 78, 73, 29, 29, 39, 33, 29, 7, 0, 61, 58, 0, 0, 27, 68, 39, 
    65, 27, 27, 34, 52, 13, 0, 3, 0, 21, 48, 58, 61, 32, 11, 4, 36, 36, 0, 0, 0, 0, 0, 0, 0, 0, 47, 53, 32, 50, 68, 37, 
    62, 21, 24, 44, 83, 88, 0, 0, 0, 1, 36, 57, 84, 122, 139, 92, 54, 75, 92, 39, 13, 1, 1, 50, 82, 47, 70, 110, 105, 74, 55, 28, 
    56, 21, 9, 0, 19, 46, 34, 0, 0, 4, 25, 47, 62, 82, 98, 89, 66, 93, 114, 57, 1, 0, 1, 25, 80, 91, 57, 55, 42, 32, 43, 26, 
    52, 15, 0, 0, 0, 0, 0, 18, 16, 8, 1, 27, 51, 54, 53, 53, 51, 49, 34, 0, 0, 0, 0, 0, 0, 41, 65, 42, 10, 7, 24, 19, 
    45, 4, 0, 0, 0, 0, 7, 20, 15, 9, 1, 15, 44, 58, 54, 47, 31, 11, 37, 94, 105, 87, 63, 49, 49, 54, 61, 42, 13, 9, 16, 8, 
    31, 1, 10, 18, 12, 0, 21, 42, 18, 22, 22, 24, 34, 40, 37, 33, 29, 23, 38, 93, 124, 104, 70, 44, 53, 56, 44, 35, 24, 20, 15, 6, 
    32, 7, 14, 17, 10, 0, 19, 63, 45, 32, 32, 32, 31, 36, 36, 37, 48, 62, 67, 63, 56, 48, 42, 28, 16, 47, 49, 40, 34, 19, 5, 1, 
    46, 13, 11, 3, 0, 0, 15, 50, 53, 36, 36, 40, 32, 30, 32, 29, 31, 34, 37, 39, 46, 54, 63, 55, 28, 30, 49, 41, 23, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 29, 54, 51, 43, 35, 30, 15, 9, 10, 11, 10, 6, 2, 8, 19, 30, 33, 23, 6, 19, 17, 0, 0, 0, 0, 
    144, 121, 116, 113, 114, 110, 98, 74, 98, 109, 105, 95, 83, 78, 74, 74, 76, 78, 79, 76, 74, 82, 89, 94, 83, 67, 59, 68, 89, 107, 134, 136, 
    
    -- channel=148
    0, 137, 131, 125, 131, 144, 144, 118, 96, 106, 112, 108, 102, 106, 107, 100, 107, 121, 137, 149, 147, 137, 134, 141, 145, 137, 107, 96, 102, 105, 86, 103, 
    0, 247, 241, 234, 235, 257, 260, 216, 171, 183, 197, 190, 188, 191, 194, 194, 205, 218, 236, 245, 241, 231, 225, 233, 247, 246, 213, 188, 190, 193, 175, 220, 
    0, 269, 267, 266, 262, 273, 283, 240, 174, 181, 204, 195, 204, 201, 200, 220, 225, 236, 249, 231, 224, 220, 217, 222, 242, 250, 235, 208, 191, 193, 198, 255, 
    0, 286, 284, 283, 282, 288, 297, 247, 170, 177, 193, 189, 208, 190, 181, 201, 194, 204, 218, 192, 184, 194, 203, 218, 241, 242, 237, 214, 172, 170, 205, 272, 
    0, 294, 293, 293, 292, 300, 304, 255, 168, 174, 197, 194, 220, 200, 195, 206, 185, 191, 197, 166, 155, 160, 191, 230, 250, 237, 228, 200, 152, 139, 189, 275, 
    0, 294, 293, 293, 296, 301, 302, 266, 179, 170, 212, 218, 240, 229, 228, 239, 221, 218, 214, 183, 157, 149, 177, 235, 263, 244, 226, 193, 147, 119, 155, 264, 
    0, 294, 292, 292, 299, 289, 285, 289, 202, 162, 228, 255, 267, 265, 261, 263, 259, 249, 244, 232, 195, 167, 171, 211, 256, 253, 222, 198, 163, 124, 131, 237, 
    0, 294, 291, 296, 303, 277, 272, 303, 213, 157, 229, 254, 271, 287, 271, 269, 271, 267, 263, 258, 250, 217, 174, 186, 238, 250, 234, 216, 187, 138, 118, 211, 
    0, 292, 289, 297, 302, 271, 266, 289, 206, 163, 240, 247, 263, 296, 271, 258, 261, 260, 267, 261, 262, 275, 209, 175, 230, 253, 253, 252, 227, 183, 155, 223, 
    0, 287, 289, 297, 301, 273, 248, 265, 188, 170, 239, 228, 229, 264, 250, 242, 248, 247, 257, 254, 250, 282, 246, 196, 221, 251, 269, 290, 268, 230, 216, 270, 
    0, 271, 284, 298, 311, 279, 242, 246, 168, 143, 201, 213, 214, 228, 227, 228, 231, 231, 232, 230, 229, 258, 255, 211, 210, 242, 277, 298, 288, 267, 266, 322, 
    0, 253, 274, 294, 302, 260, 233, 244, 161, 111, 154, 199, 213, 218, 208, 201, 200, 202, 200, 202, 206, 210, 213, 195, 184, 221, 271, 296, 293, 293, 293, 345, 
    0, 236, 258, 281, 266, 224, 224, 245, 169, 131, 156, 199, 221, 235, 222, 195, 189, 193, 200, 211, 214, 179, 160, 156, 147, 179, 235, 266, 277, 291, 294, 344, 
    0, 231, 253, 262, 229, 191, 195, 213, 180, 174, 186, 204, 213, 236, 221, 183, 172, 175, 182, 198, 201, 157, 124, 125, 135, 170, 208, 227, 240, 272, 293, 344, 
    0, 237, 245, 222, 176, 159, 170, 194, 196, 199, 202, 180, 150, 163, 169, 148, 138, 141, 153, 163, 164, 134, 109, 113, 121, 142, 169, 184, 195, 240, 287, 345, 
    0, 231, 236, 196, 127, 125, 155, 201, 204, 190, 183, 167, 141, 138, 135, 125, 103, 79, 78, 81, 81, 84, 73, 61, 69, 91, 143, 176, 162, 203, 276, 346, 
    0, 240, 247, 204, 105, 98, 152, 201, 173, 152, 155, 147, 147, 154, 137, 140, 105, 72, 79, 84, 90, 120, 100, 67, 72, 90, 146, 189, 173, 187, 253, 345, 
    0, 246, 241, 205, 103, 101, 161, 158, 99, 118, 139, 129, 145, 164, 164, 178, 133, 120, 133, 122, 134, 184, 158, 119, 119, 121, 172, 196, 173, 167, 219, 339, 
    0, 260, 254, 214, 103, 108, 171, 120, 36, 92, 130, 117, 112, 125, 138, 153, 147, 178, 174, 157, 169, 213, 194, 160, 162, 168, 210, 193, 154, 147, 188, 330, 
    0, 267, 263, 218, 90, 83, 146, 103, 28, 69, 110, 112, 91, 83, 97, 111, 132, 204, 203, 180, 192, 202, 188, 183, 175, 191, 223, 180, 126, 117, 160, 320, 
    0, 261, 269, 237, 105, 70, 106, 95, 52, 46, 56, 79, 83, 87, 90, 86, 100, 158, 158, 140, 145, 150, 141, 137, 142, 144, 172, 159, 127, 116, 146, 311, 
    0, 257, 271, 246, 122, 74, 91, 88, 72, 40, 17, 41, 66, 103, 124, 127, 72, 82, 137, 160, 144, 138, 137, 139, 168, 156, 110, 137, 163, 126, 128, 304, 
    0, 264, 274, 235, 110, 81, 101, 103, 103, 63, 13, 5, 24, 64, 111, 132, 49, 27, 106, 162, 135, 138, 139, 129, 193, 153, 45, 94, 152, 108, 114, 303, 
    0, 272, 282, 231, 73, 55, 106, 125, 149, 97, 29, 4, 0, 21, 64, 98, 30, 0, 73, 138, 132, 149, 153, 139, 195, 148, 34, 61, 110, 77, 110, 307, 
    0, 278, 289, 246, 106, 52, 104, 152, 184, 124, 53, 17, 0, 0, 9, 32, 12, 0, 40, 119, 174, 204, 213, 191, 200, 117, 28, 38, 56, 53, 122, 311, 
    0, 262, 278, 267, 181, 117, 110, 160, 200, 134, 83, 43, 3, 0, 0, 0, 2, 5, 3, 73, 179, 214, 218, 223, 192, 66, 11, 22, 47, 72, 140, 311, 
    0, 246, 257, 269, 239, 188, 147, 157, 189, 129, 109, 70, 12, 0, 0, 0, 9, 17, 8, 72, 181, 215, 222, 237, 204, 57, 0, 9, 54, 96, 152, 306, 
    0, 244, 251, 260, 256, 222, 164, 150, 168, 118, 117, 89, 27, 0, 0, 0, 8, 25, 34, 76, 147, 174, 198, 226, 187, 43, 0, 3, 58, 101, 154, 306, 
    0, 250, 254, 253, 238, 219, 172, 141, 138, 106, 111, 88, 38, 5, 3, 10, 17, 34, 56, 78, 103, 123, 157, 200, 163, 37, 0, 6, 55, 91, 159, 311, 
    0, 255, 254, 246, 232, 226, 198, 136, 98, 91, 97, 76, 44, 25, 22, 31, 36, 41, 50, 68, 85, 102, 126, 163, 149, 46, 0, 12, 54, 92, 185, 320, 
    1, 252, 250, 253, 247, 243, 219, 146, 68, 71, 78, 65, 54, 49, 49, 57, 60, 60, 69, 86, 99, 108, 119, 135, 137, 76, 23, 34, 68, 125, 221, 321, 
    0, 109, 109, 112, 112, 116, 115, 59, 0, 3, 6, 0, 0, 0, 1, 7, 7, 3, 7, 21, 28, 29, 34, 41, 43, 18, 0, 0, 0, 38, 102, 183, 
    
    -- channel=149
    108, 162, 158, 156, 149, 155, 139, 137, 137, 127, 111, 108, 122, 113, 119, 122, 130, 147, 160, 171, 171, 171, 169, 175, 163, 154, 148, 147, 147, 142, 134, 58, 
    256, 273, 272, 283, 279, 259, 230, 220, 220, 209, 206, 208, 216, 228, 243, 262, 285, 307, 307, 303, 299, 300, 297, 295, 275, 263, 265, 279, 258, 253, 239, 73, 
    269, 293, 290, 289, 294, 274, 227, 199, 211, 205, 199, 215, 217, 236, 255, 270, 298, 297, 301, 313, 303, 298, 299, 298, 288, 285, 284, 294, 278, 271, 266, 79, 
    277, 304, 304, 306, 307, 285, 215, 179, 179, 172, 170, 166, 172, 183, 195, 208, 231, 240, 258, 286, 302, 282, 286, 293, 293, 295, 289, 283, 291, 291, 288, 89, 
    284, 309, 307, 309, 307, 284, 208, 139, 113, 108, 120, 105, 101, 117, 111, 116, 138, 147, 171, 198, 251, 285, 280, 280, 291, 287, 276, 274, 289, 306, 300, 94, 
    284, 308, 309, 309, 298, 269, 189, 120, 81, 73, 92, 90, 74, 87, 87, 83, 92, 84, 97, 134, 178, 249, 301, 285, 281, 277, 258, 252, 266, 292, 306, 98, 
    284, 309, 308, 306, 284, 268, 191, 106, 106, 114, 130, 132, 127, 110, 109, 113, 108, 102, 93, 111, 169, 212, 275, 305, 282, 268, 262, 233, 239, 258, 296, 100, 
    283, 307, 309, 299, 272, 261, 195, 102, 119, 135, 165, 194, 190, 163, 144, 135, 132, 129, 129, 123, 147, 208, 247, 271, 277, 265, 252, 231, 222, 248, 278, 84, 
    282, 308, 311, 293, 257, 244, 186, 109, 119, 151, 162, 180, 165, 148, 131, 124, 135, 139, 138, 155, 145, 152, 217, 260, 268, 267, 267, 256, 226, 218, 244, 61, 
    279, 308, 309, 291, 243, 218, 163, 86, 106, 120, 124, 143, 137, 124, 119, 119, 129, 138, 131, 155, 157, 146, 193, 236, 274, 300, 296, 257, 239, 227, 248, 75, 
    268, 308, 308, 288, 231, 191, 105, 54, 92, 107, 116, 119, 110, 102, 102, 107, 113, 121, 119, 134, 149, 145, 174, 223, 268, 304, 300, 280, 276, 288, 295, 90, 
    255, 290, 300, 274, 208, 182, 117, 62, 66, 85, 84, 86, 86, 78, 81, 91, 97, 98, 101, 112, 126, 133, 156, 202, 244, 279, 302, 310, 308, 308, 308, 88, 
    235, 268, 279, 250, 210, 187, 131, 69, 53, 54, 60, 74, 77, 79, 66, 64, 68, 71, 81, 91, 105, 118, 122, 160, 225, 284, 307, 316, 318, 310, 308, 89, 
    221, 251, 235, 207, 187, 175, 129, 80, 46, 72, 90, 96, 83, 72, 73, 65, 64, 77, 103, 109, 109, 113, 116, 153, 204, 239, 253, 270, 305, 320, 309, 88, 
    213, 229, 197, 169, 157, 170, 139, 111, 77, 89, 75, 88, 97, 74, 68, 69, 76, 87, 96, 84, 67, 75, 92, 112, 137, 161, 183, 217, 258, 303, 314, 88, 
    210, 216, 175, 137, 127, 150, 161, 138, 111, 68, 61, 52, 39, 23, 26, 31, 36, 46, 50, 45, 44, 35, 39, 69, 83, 106, 104, 136, 219, 276, 309, 88, 
    213, 196, 121, 93, 118, 161, 164, 116, 99, 67, 52, 59, 61, 56, 53, 32, 34, 25, 11, 16, 24, 20, 17, 18, 27, 44, 66, 105, 183, 255, 306, 90, 
    199, 195, 124, 101, 134, 173, 126, 84, 58, 75, 86, 102, 102, 120, 86, 59, 65, 50, 51, 92, 88, 78, 79, 53, 78, 106, 102, 120, 183, 264, 304, 91, 
    213, 218, 137, 101, 129, 146, 74, 57, 52, 67, 98, 111, 91, 98, 94, 113, 113, 122, 134, 166, 172, 134, 130, 135, 157, 172, 141, 131, 154, 229, 281, 88, 
    219, 219, 136, 88, 115, 114, 55, 41, 60, 60, 57, 55, 54, 70, 67, 104, 144, 153, 123, 120, 122, 125, 123, 119, 141, 126, 112, 92, 93, 194, 276, 86, 
    218, 223, 142, 82, 89, 73, 43, 37, 41, 44, 33, 38, 42, 41, 49, 94, 92, 83, 92, 96, 91, 84, 88, 92, 110, 105, 75, 71, 84, 177, 272, 86, 
    217, 222, 143, 77, 74, 76, 36, 37, 22, 26, 31, 36, 45, 61, 53, 45, 69, 89, 83, 60, 59, 57, 71, 88, 77, 46, 62, 83, 89, 186, 271, 82, 
    208, 217, 141, 86, 68, 82, 72, 35, 13, 11, 20, 42, 49, 90, 74, 57, 60, 80, 94, 90, 84, 71, 104, 121, 78, 82, 89, 94, 107, 191, 261, 75, 
    196, 208, 122, 73, 79, 61, 92, 72, 25, 25, 12, 34, 55, 82, 49, 24, 49, 98, 113, 137, 129, 116, 150, 152, 78, 78, 88, 77, 63, 153, 243, 70, 
    180, 185, 108, 52, 55, 66, 82, 94, 59, 33, 14, 11, 17, 36, 21, 0, 27, 84, 112, 127, 131, 113, 131, 124, 30, 9, 43, 42, 52, 148, 228, 61, 
    170, 175, 118, 69, 59, 82, 130, 105, 60, 36, 21, 3, 0, 6, 8, 13, 14, 34, 91, 146, 193, 190, 182, 110, 56, 29, 24, 36, 60, 150, 219, 46, 
    164, 175, 150, 120, 116, 112, 135, 101, 68, 49, 28, 16, 8, 3, 5, 10, 10, 42, 124, 176, 214, 209, 198, 111, 40, 22, 21, 42, 68, 148, 208, 40, 
    162, 174, 180, 164, 128, 101, 119, 91, 85, 63, 37, 16, 8, 6, 9, 19, 25, 53, 125, 149, 146, 149, 150, 84, 17, 5, 25, 53, 72, 147, 202, 35, 
    161, 175, 170, 148, 125, 100, 114, 78, 78, 63, 39, 20, 17, 16, 20, 29, 44, 53, 66, 77, 93, 116, 126, 66, 30, 3, 27, 54, 72, 147, 195, 32, 
    157, 159, 145, 139, 134, 104, 84, 64, 64, 59, 42, 27, 25, 24, 23, 26, 30, 39, 49, 58, 74, 94, 107, 50, 19, 15, 26, 46, 78, 153, 185, 32, 
    145, 150, 145, 139, 132, 107, 71, 48, 51, 53, 48, 40, 27, 32, 31, 30, 34, 43, 50, 55, 62, 72, 81, 53, 18, 20, 26, 46, 98, 160, 192, 34, 
    101, 164, 167, 173, 170, 141, 87, 83, 60, 52, 44, 48, 54, 55, 56, 58, 58, 64, 73, 81, 88, 91, 96, 84, 56, 47, 59, 79, 126, 187, 210, 65, 
    
    -- channel=150
    56, 57, 59, 49, 51, 62, 67, 48, 52, 59, 51, 50, 50, 59, 54, 46, 47, 47, 53, 59, 61, 53, 54, 58, 71, 62, 52, 47, 73, 57, 56, 156, 
    0, 10, 14, 12, 1, 19, 32, 8, 3, 16, 11, 5, 11, 9, 13, 13, 3, 7, 2, 4, 14, 11, 1, 5, 19, 24, 24, 9, 27, 26, 20, 158, 
    0, 7, 8, 8, 4, 16, 44, 13, 0, 7, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 7, 11, 2, 2, 5, 13, 20, 16, 12, 21, 18, 159, 
    0, 1, 2, 1, 2, 16, 51, 9, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 7, 0, 4, 19, 19, 5, 10, 17, 166, 
    0, 0, 0, 0, 1, 17, 62, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 10, 6, 3, 19, 25, 4, 0, 9, 177, 
    0, 0, 0, 0, 5, 8, 63, 57, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 4, 13, 15, 14, 31, 8, 0, 0, 179, 
    0, 0, 0, 3, 9, 0, 45, 68, 0, 0, 0, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 17, 19, 33, 26, 0, 0, 169, 
    0, 0, 0, 8, 15, 0, 40, 44, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 5, 8, 25, 34, 33, 12, 0, 153, 
    0, 0, 0, 8, 19, 0, 34, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 4, 17, 37, 27, 20, 0, 152, 
    0, 0, 0, 10, 31, 0, 22, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 28, 29, 20, 11, 171, 
    0, 0, 0, 15, 43, 6, 28, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 14, 9, 6, 179, 
    0, 0, 0, 17, 30, 18, 43, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 0, 0, 15, 13, 1, 39, 24, 11, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 0, 9, 8, 19, 0, 24, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 13, 27, 0, 8, 5, 19, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 11, 46, 4, 0, 0, 18, 45, 8, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 7, 62, 22, 0, 0, 20, 14, 16, 0, 1, 9, 39, 13, 25, 30, 14, 11, 20, 0, 22, 40, 5, 13, 0, 0, 0, 0, 0, 0, 0, 175, 
    3, 15, 64, 22, 0, 7, 44, 0, 0, 0, 0, 0, 5, 1, 25, 16, 27, 31, 33, 9, 21, 51, 38, 38, 21, 8, 0, 0, 0, 0, 0, 177, 
    0, 16, 58, 16, 0, 20, 63, 13, 0, 0, 9, 0, 0, 0, 0, 0, 15, 11, 0, 0, 0, 5, 9, 8, 0, 14, 13, 0, 0, 0, 0, 177, 
    0, 15, 68, 32, 0, 6, 56, 30, 0, 0, 8, 18, 3, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 175, 
    0, 8, 70, 47, 1, 0, 34, 31, 17, 0, 0, 10, 16, 7, 12, 0, 0, 2, 7, 0, 0, 0, 0, 2, 0, 0, 13, 16, 0, 0, 0, 175, 
    0, 1, 64, 39, 23, 21, 13, 28, 30, 10, 2, 0, 6, 0, 40, 17, 0, 0, 18, 4, 0, 8, 0, 4, 42, 0, 0, 18, 9, 0, 0, 173, 
    0, 0, 61, 29, 0, 37, 16, 24, 42, 23, 19, 0, 0, 0, 37, 42, 0, 0, 30, 22, 5, 23, 0, 0, 79, 8, 0, 0, 2, 0, 0, 168, 
    0, 0, 62, 40, 0, 0, 15, 32, 43, 32, 24, 13, 0, 0, 3, 31, 3, 0, 0, 12, 0, 14, 0, 0, 41, 29, 0, 0, 0, 0, 0, 160, 
    0, 0, 49, 55, 9, 0, 0, 30, 33, 38, 31, 23, 18, 9, 5, 17, 16, 0, 0, 9, 8, 13, 5, 38, 25, 18, 12, 5, 0, 0, 0, 151, 
    0, 0, 22, 55, 37, 5, 0, 24, 21, 32, 41, 31, 21, 23, 20, 17, 24, 0, 0, 0, 13, 17, 10, 70, 51, 14, 8, 4, 0, 0, 0, 142, 
    0, 0, 0, 22, 30, 14, 0, 32, 12, 18, 41, 39, 24, 22, 22, 15, 21, 10, 0, 0, 0, 0, 0, 55, 49, 25, 6, 0, 0, 0, 0, 137, 
    0, 0, 0, 0, 11, 18, 0, 27, 11, 10, 29, 39, 30, 24, 24, 15, 10, 9, 0, 0, 0, 0, 0, 58, 39, 25, 10, 0, 0, 0, 0, 133, 
    0, 0, 0, 0, 4, 20, 1, 8, 11, 10, 20, 33, 30, 22, 22, 17, 9, 2, 0, 0, 0, 0, 0, 51, 50, 19, 8, 1, 0, 0, 0, 128, 
    0, 0, 0, 0, 0, 23, 25, 0, 7, 13, 18, 21, 30, 22, 20, 20, 16, 9, 6, 1, 0, 0, 0, 23, 55, 22, 7, 3, 0, 0, 0, 125, 
    0, 0, 0, 0, 0, 18, 47, 8, 3, 10, 16, 19, 24, 21, 20, 20, 16, 11, 12, 13, 4, 1, 0, 14, 41, 31, 12, 0, 0, 0, 0, 126, 
    0, 0, 0, 0, 0, 0, 29, 22, 8, 7, 9, 13, 14, 12, 11, 12, 10, 4, 3, 6, 4, 2, 3, 9, 22, 27, 15, 0, 0, 0, 0, 69, 
    
    -- channel=151
    235, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 9, 1, 14, 18, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    325, 0, 0, 0, 9, 1, 0, 0, 12, 15, 7, 17, 15, 15, 13, 15, 15, 14, 3, 0, 0, 0, 1, 9, 0, 0, 0, 0, 0, 0, 3, 0, 
    340, 0, 0, 0, 2, 0, 0, 0, 16, 26, 15, 37, 19, 25, 42, 27, 26, 29, 1, 8, 0, 0, 4, 17, 6, 0, 0, 0, 0, 0, 4, 0, 
    352, 0, 0, 0, 1, 0, 0, 0, 24, 43, 24, 67, 26, 36, 65, 38, 51, 58, 19, 40, 18, 4, 22, 25, 1, 2, 0, 0, 0, 22, 10, 0, 
    357, 2, 4, 3, 2, 0, 0, 0, 32, 77, 53, 86, 49, 57, 73, 47, 65, 73, 45, 60, 61, 45, 36, 27, 0, 0, 0, 0, 0, 33, 27, 0, 
    357, 1, 4, 3, 0, 0, 0, 0, 10, 110, 79, 81, 53, 64, 72, 52, 58, 63, 63, 64, 64, 85, 61, 26, 0, 0, 0, 0, 0, 31, 46, 0, 
    357, 2, 5, 1, 0, 0, 0, 0, 0, 138, 90, 70, 36, 31, 58, 55, 57, 60, 57, 73, 60, 60, 76, 46, 1, 0, 0, 0, 0, 4, 48, 0, 
    356, 2, 5, 1, 0, 0, 0, 0, 0, 133, 74, 66, 50, 9, 49, 72, 65, 70, 57, 66, 76, 34, 59, 72, 18, 0, 0, 0, 0, 0, 35, 0, 
    355, 3, 5, 0, 0, 0, 0, 0, 31, 141, 67, 69, 80, 14, 46, 81, 73, 78, 62, 62, 91, 32, 38, 89, 36, 6, 1, 0, 0, 0, 24, 0, 
    352, 6, 7, 0, 0, 0, 9, 0, 50, 131, 58, 67, 88, 44, 60, 80, 79, 75, 67, 61, 96, 57, 33, 80, 56, 25, 9, 0, 0, 0, 11, 0, 
    339, 19, 12, 0, 0, 0, 12, 0, 48, 118, 79, 70, 77, 67, 75, 77, 79, 73, 72, 75, 96, 79, 51, 67, 83, 63, 26, 0, 0, 0, 4, 0, 
    322, 33, 17, 0, 0, 0, 11, 0, 28, 102, 109, 82, 72, 62, 69, 75, 78, 76, 82, 89, 79, 80, 79, 76, 100, 87, 36, 0, 4, 4, 4, 0, 
    303, 35, 19, 0, 0, 0, 14, 0, 27, 78, 100, 79, 82, 55, 46, 67, 79, 82, 87, 83, 43, 46, 74, 73, 95, 85, 41, 21, 21, 7, 3, 0, 
    299, 28, 8, 0, 0, 4, 26, 0, 34, 58, 80, 62, 84, 67, 39, 57, 74, 80, 81, 73, 30, 27, 59, 72, 86, 76, 47, 44, 67, 35, 2, 0, 
    298, 16, 0, 0, 16, 35, 43, 0, 12, 53, 70, 48, 76, 86, 69, 69, 79, 87, 84, 77, 57, 57, 73, 75, 80, 76, 69, 63, 106, 90, 13, 0, 
    285, 6, 0, 0, 42, 73, 52, 0, 0, 59, 77, 53, 60, 63, 73, 54, 47, 71, 71, 75, 81, 60, 64, 78, 87, 109, 107, 84, 118, 132, 35, 0, 
    287, 0, 0, 0, 47, 85, 35, 0, 7, 74, 72, 54, 51, 27, 51, 20, 24, 68, 61, 65, 94, 34, 20, 67, 66, 109, 111, 79, 97, 127, 65, 0, 
    293, 0, 0, 0, 53, 77, 0, 0, 75, 97, 57, 46, 68, 43, 53, 18, 45, 47, 30, 35, 68, 12, 0, 33, 37, 70, 55, 37, 69, 112, 108, 0, 
    308, 0, 0, 0, 53, 81, 0, 0, 99, 105, 54, 37, 65, 65, 78, 56, 80, 20, 15, 50, 63, 17, 9, 31, 44, 69, 7, 11, 77, 120, 144, 0, 
    311, 0, 0, 0, 31, 90, 0, 0, 76, 89, 73, 40, 51, 73, 78, 83, 124, 39, 29, 66, 67, 45, 51, 61, 61, 79, 5, 2, 83, 135, 165, 0, 
    307, 0, 0, 0, 4, 68, 30, 5, 43, 57, 83, 66, 62, 65, 69, 63, 99, 66, 45, 55, 61, 55, 63, 75, 56, 67, 51, 38, 70, 118, 173, 0, 
    305, 7, 0, 0, 10, 41, 31, 33, 26, 33, 71, 79, 96, 85, 62, 0, 62, 127, 84, 34, 54, 67, 67, 105, 27, 0, 96, 90, 36, 82, 182, 0, 
    304, 9, 0, 0, 21, 69, 22, 45, 18, 5, 48, 63, 96, 90, 74, 0, 30, 135, 99, 3, 35, 52, 39, 89, 0, 0, 83, 106, 36, 91, 197, 0, 
    303, 15, 0, 0, 15, 102, 64, 54, 0, 0, 29, 51, 78, 86, 85, 12, 40, 112, 112, 35, 50, 60, 32, 59, 0, 0, 73, 90, 53, 121, 205, 0, 
    297, 30, 0, 0, 4, 87, 91, 65, 0, 0, 17, 34, 52, 66, 69, 49, 58, 93, 142, 125, 67, 42, 26, 24, 0, 0, 63, 67, 74, 136, 196, 0, 
    289, 43, 26, 0, 0, 33, 78, 68, 0, 12, 14, 10, 34, 53, 57, 63, 63, 65, 133, 158, 49, 14, 5, 0, 0, 0, 65, 77, 92, 128, 180, 0, 
    280, 52, 39, 8, 0, 5, 52, 65, 0, 35, 21, 0, 22, 53, 58, 64, 71, 67, 110, 141, 60, 38, 33, 0, 0, 0, 65, 92, 103, 118, 169, 0, 
    277, 45, 37, 25, 14, 5, 26, 58, 0, 50, 31, 0, 16, 49, 56, 58, 66, 70, 87, 104, 74, 70, 65, 0, 0, 8, 66, 94, 103, 119, 169, 0, 
    280, 42, 33, 26, 25, 16, 8, 38, 17, 56, 34, 15, 20, 44, 55, 57, 65, 71, 74, 76, 77, 84, 77, 22, 0, 9, 69, 90, 99, 130, 166, 0, 
    278, 40, 43, 41, 38, 19, 0, 10, 49, 59, 34, 29, 34, 42, 55, 54, 54, 60, 68, 69, 73, 80, 77, 44, 0, 0, 68, 90, 102, 145, 147, 0, 
    274, 49, 56, 45, 41, 24, 0, 0, 57, 59, 45, 44, 46, 45, 54, 50, 50, 59, 68, 60, 57, 63, 61, 44, 4, 3, 55, 90, 114, 138, 111, 0, 
    197, 59, 61, 54, 51, 41, 19, 1, 58, 60, 53, 53, 52, 52, 58, 55, 53, 58, 64, 58, 54, 58, 56, 51, 32, 28, 51, 69, 97, 106, 79, 8, 
    
    -- channel=152
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=153
    55, 83, 77, 78, 84, 83, 73, 61, 57, 60, 65, 71, 76, 82, 85, 87, 91, 95, 99, 94, 88, 84, 82, 87, 81, 74, 65, 63, 58, 58, 57, 22, 
    96, 126, 121, 120, 132, 127, 109, 89, 86, 100, 101, 110, 112, 120, 124, 125, 132, 134, 137, 129, 117, 109, 112, 117, 120, 111, 96, 86, 86, 82, 88, 65, 
    106, 147, 146, 145, 146, 144, 129, 111, 110, 129, 138, 139, 139, 142, 144, 147, 151, 149, 138, 122, 107, 100, 103, 112, 122, 117, 100, 80, 82, 83, 95, 79, 
    118, 163, 161, 161, 160, 155, 143, 136, 147, 169, 184, 187, 184, 180, 175, 178, 173, 168, 150, 120, 98, 94, 103, 109, 116, 113, 93, 68, 62, 75, 95, 80, 
    123, 170, 169, 169, 167, 160, 150, 150, 179, 216, 235, 248, 242, 236, 233, 226, 217, 214, 186, 145, 114, 100, 108, 115, 112, 101, 80, 54, 42, 61, 90, 75, 
    123, 170, 169, 169, 167, 165, 157, 158, 206, 251, 276, 287, 285, 289, 291, 284, 276, 272, 248, 204, 161, 129, 117, 122, 115, 97, 77, 46, 34, 47, 79, 73, 
    123, 169, 170, 168, 165, 162, 170, 180, 224, 263, 281, 283, 289, 306, 325, 328, 321, 315, 305, 276, 215, 163, 136, 120, 117, 100, 78, 56, 37, 39, 68, 68, 
    123, 168, 169, 167, 164, 159, 184, 208, 236, 263, 274, 270, 279, 297, 328, 340, 336, 330, 323, 318, 274, 195, 157, 121, 118, 111, 90, 72, 46, 33, 52, 61, 
    122, 167, 167, 169, 166, 159, 201, 220, 238, 261, 280, 275, 290, 301, 324, 338, 331, 325, 322, 319, 320, 246, 181, 144, 128, 125, 117, 94, 73, 58, 61, 65, 
    119, 163, 165, 166, 165, 171, 217, 228, 249, 276, 293, 283, 298, 306, 317, 328, 323, 315, 320, 313, 327, 292, 223, 181, 149, 148, 148, 135, 113, 105, 105, 84, 
    112, 154, 162, 164, 169, 180, 222, 227, 235, 257, 273, 277, 288, 297, 306, 313, 312, 304, 309, 304, 318, 312, 256, 215, 181, 169, 166, 163, 150, 147, 151, 109, 
    100, 142, 156, 156, 163, 163, 210, 209, 212, 221, 242, 273, 280, 284, 286, 283, 282, 279, 281, 276, 277, 274, 240, 209, 182, 172, 171, 170, 170, 169, 169, 123, 
    87, 130, 140, 137, 131, 134, 184, 194, 207, 217, 248, 283, 297, 294, 285, 271, 267, 271, 278, 267, 244, 220, 195, 174, 151, 151, 154, 159, 165, 168, 169, 122, 
    86, 121, 125, 118, 95, 101, 141, 170, 210, 243, 278, 287, 303, 294, 278, 260, 256, 263, 272, 261, 226, 186, 166, 162, 157, 158, 155, 161, 165, 167, 169, 122, 
    84, 103, 100, 89, 75, 83, 104, 139, 218, 253, 272, 242, 243, 242, 232, 221, 224, 232, 237, 230, 201, 177, 167, 170, 169, 176, 176, 179, 181, 175, 169, 122, 
    68, 86, 75, 64, 69, 77, 84, 127, 202, 232, 242, 202, 192, 195, 189, 172, 162, 153, 149, 156, 148, 146, 144, 136, 151, 177, 197, 204, 192, 186, 172, 123, 
    64, 90, 82, 72, 70, 74, 76, 129, 172, 196, 196, 171, 171, 182, 173, 152, 126, 113, 111, 130, 132, 129, 121, 106, 129, 169, 211, 224, 192, 187, 172, 122, 
    77, 107, 108, 89, 76, 71, 70, 111, 153, 167, 171, 160, 177, 191, 182, 168, 137, 131, 133, 147, 160, 155, 134, 123, 139, 174, 207, 209, 183, 177, 171, 121, 
    95, 128, 126, 99, 85, 79, 76, 82, 132, 151, 155, 143, 155, 164, 170, 173, 164, 169, 171, 177, 190, 191, 171, 166, 182, 187, 192, 186, 176, 169, 176, 123, 
    102, 134, 129, 100, 84, 86, 84, 74, 115, 143, 147, 140, 136, 144, 154, 163, 183, 194, 197, 203, 208, 204, 200, 195, 198, 202, 188, 174, 172, 165, 177, 126, 
    102, 135, 136, 111, 84, 89, 92, 86, 99, 111, 120, 134, 135, 148, 141, 147, 174, 180, 183, 190, 195, 188, 189, 184, 174, 189, 184, 173, 174, 169, 172, 125, 
    104, 143, 143, 121, 93, 86, 101, 97, 89, 83, 85, 115, 132, 162, 149, 132, 136, 151, 160, 168, 170, 166, 174, 172, 152, 156, 165, 172, 175, 167, 167, 125, 
    117, 164, 151, 118, 100, 88, 110, 118, 98, 79, 63, 81, 110, 142, 138, 110, 98, 116, 131, 143, 150, 153, 159, 158, 132, 113, 128, 154, 161, 151, 166, 132, 
    139, 195, 169, 114, 86, 99, 120, 139, 126, 91, 65, 62, 80, 95, 111, 90, 71, 92, 122, 131, 146, 156, 153, 146, 140, 98, 97, 124, 136, 143, 181, 146, 
    161, 223, 200, 140, 96, 110, 142, 158, 150, 104, 74, 58, 56, 58, 73, 70, 63, 82, 125, 141, 167, 177, 171, 151, 137, 94, 82, 96, 115, 149, 204, 159, 
    161, 229, 225, 181, 146, 137, 157, 168, 159, 124, 92, 64, 49, 44, 49, 55, 61, 76, 110, 142, 168, 176, 176, 156, 112, 76, 70, 90, 122, 171, 225, 169, 
    156, 221, 224, 212, 194, 173, 165, 163, 155, 141, 111, 73, 49, 42, 47, 57, 67, 75, 101, 145, 170, 182, 179, 160, 107, 58, 60, 94, 137, 189, 235, 173, 
    154, 221, 221, 221, 214, 184, 161, 158, 147, 146, 124, 83, 51, 43, 49, 58, 70, 82, 101, 139, 162, 179, 189, 158, 105, 52, 57, 97, 143, 195, 238, 176, 
    161, 233, 233, 225, 215, 185, 151, 152, 138, 141, 124, 88, 59, 51, 56, 64, 75, 92, 108, 129, 147, 165, 184, 156, 99, 56, 59, 94, 142, 194, 241, 180, 
    171, 247, 246, 237, 226, 201, 158, 144, 127, 131, 115, 92, 69, 67, 72, 78, 84, 93, 105, 119, 133, 147, 160, 147, 94, 60, 63, 92, 145, 199, 254, 186, 
    178, 256, 257, 252, 241, 221, 172, 137, 113, 116, 106, 92, 84, 87, 94, 100, 103, 108, 116, 126, 135, 142, 147, 141, 110, 79, 81, 109, 157, 213, 265, 183, 
    124, 164, 163, 159, 155, 147, 114, 78, 64, 65, 60, 53, 54, 58, 66, 69, 70, 71, 76, 82, 86, 88, 89, 86, 75, 55, 53, 70, 101, 140, 168, 125, 
    
    -- channel=154
    268, 234, 229, 231, 240, 224, 189, 178, 187, 180, 176, 188, 200, 205, 211, 232, 250, 261, 264, 256, 247, 246, 251, 251, 229, 212, 212, 227, 202, 185, 193, 10, 
    430, 360, 353, 361, 372, 346, 280, 255, 270, 268, 266, 278, 286, 298, 319, 339, 366, 380, 378, 373, 359, 354, 361, 367, 348, 328, 325, 330, 305, 286, 298, 20, 
    454, 386, 382, 382, 390, 366, 273, 234, 264, 257, 264, 275, 271, 293, 313, 325, 354, 358, 357, 361, 348, 339, 354, 371, 367, 355, 336, 324, 320, 323, 329, 24, 
    469, 399, 399, 400, 401, 359, 238, 181, 213, 206, 223, 232, 212, 234, 245, 245, 280, 284, 291, 321, 324, 324, 354, 368, 367, 365, 334, 307, 320, 347, 349, 24, 
    479, 407, 406, 408, 401, 363, 227, 143, 176, 181, 203, 212, 192, 210, 210, 199, 223, 224, 225, 254, 298, 333, 366, 369, 357, 350, 318, 278, 300, 347, 363, 28, 
    478, 406, 407, 406, 385, 349, 234, 129, 171, 208, 233, 237, 218, 232, 232, 219, 220, 213, 217, 229, 267, 340, 383, 375, 354, 329, 299, 258, 268, 325, 368, 33, 
    477, 406, 409, 397, 358, 342, 254, 124, 185, 274, 299, 303, 273, 254, 254, 244, 243, 237, 232, 254, 270, 306, 367, 374, 348, 324, 302, 273, 256, 288, 352, 34, 
    477, 406, 409, 390, 343, 342, 267, 134, 195, 279, 288, 315, 295, 258, 262, 264, 265, 267, 258, 271, 279, 280, 335, 362, 349, 337, 323, 277, 241, 255, 317, 29, 
    475, 405, 407, 383, 327, 310, 242, 133, 215, 284, 269, 296, 282, 236, 245, 261, 269, 278, 265, 291, 297, 256, 311, 376, 371, 369, 359, 306, 265, 274, 325, 30, 
    470, 404, 407, 377, 288, 259, 200, 126, 205, 249, 226, 253, 248, 219, 230, 245, 256, 261, 250, 273, 302, 272, 293, 357, 377, 395, 387, 347, 321, 333, 361, 37, 
    452, 399, 405, 371, 284, 242, 184, 113, 163, 205, 198, 213, 212, 206, 214, 221, 225, 226, 220, 240, 272, 267, 270, 316, 371, 407, 405, 379, 372, 385, 392, 39, 
    426, 388, 390, 339, 258, 246, 193, 99, 122, 173, 190, 205, 197, 189, 186, 186, 187, 190, 206, 221, 227, 233, 241, 290, 364, 414, 415, 406, 408, 408, 408, 41, 
    393, 362, 352, 294, 238, 241, 180, 116, 131, 175, 199, 211, 215, 189, 174, 175, 185, 201, 231, 230, 204, 204, 214, 254, 326, 374, 379, 394, 407, 408, 407, 41, 
    381, 337, 303, 251, 216, 221, 185, 149, 148, 176, 196, 195, 202, 170, 149, 150, 160, 176, 197, 187, 152, 149, 172, 218, 274, 306, 308, 346, 401, 411, 408, 41, 
    380, 310, 229, 178, 188, 228, 228, 184, 167, 161, 151, 131, 139, 133, 121, 121, 136, 148, 154, 138, 107, 110, 129, 154, 182, 210, 229, 279, 376, 418, 410, 40, 
    356, 278, 173, 131, 177, 239, 241, 175, 133, 154, 157, 141, 134, 130, 121, 88, 74, 71, 65, 80, 78, 62, 66, 74, 112, 165, 188, 235, 350, 422, 413, 40, 
    361, 276, 160, 117, 190, 251, 197, 118, 110, 150, 158, 164, 151, 152, 136, 93, 87, 105, 98, 136, 155, 109, 97, 101, 126, 182, 216, 243, 326, 414, 419, 40, 
    360, 272, 158, 110, 201, 234, 118, 62, 123, 159, 159, 163, 163, 177, 158, 141, 159, 170, 165, 201, 220, 172, 155, 160, 192, 229, 220, 214, 269, 381, 423, 42, 
    380, 290, 167, 105, 191, 196, 58, 34, 123, 148, 131, 131, 130, 145, 153, 190, 213, 189, 178, 222, 231, 183, 174, 177, 227, 243, 182, 170, 217, 348, 428, 47, 
    388, 296, 166, 78, 145, 156, 46, 32, 94, 118, 99, 85, 93, 122, 120, 189, 236, 196, 189, 209, 205, 189, 191, 194, 222, 216, 138, 124, 183, 334, 433, 51, 
    385, 305, 181, 81, 108, 122, 66, 44, 51, 66, 73, 78, 85, 105, 107, 141, 157, 133, 131, 140, 137, 125, 146, 151, 157, 160, 130, 138, 179, 323, 432, 54, 
    382, 313, 179, 81, 109, 104, 83, 63, 33, 38, 53, 85, 114, 162, 122, 72, 120, 182, 171, 145, 150, 144, 184, 222, 138, 111, 167, 177, 163, 300, 428, 55, 
    375, 310, 173, 63, 106, 118, 110, 100, 46, 24, 27, 56, 92, 141, 104, 26, 76, 187, 185, 151, 168, 158, 202, 237, 110, 61, 141, 153, 130, 280, 424, 56, 
    364, 298, 153, 42, 85, 128, 156, 144, 71, 25, 15, 34, 61, 96, 67, 7, 50, 146, 165, 150, 185, 184, 205, 203, 77, 33, 108, 112, 103, 273, 417, 53, 
    349, 289, 179, 71, 107, 155, 198, 170, 89, 39, 19, 11, 17, 38, 30, 12, 32, 111, 207, 253, 278, 254, 258, 188, 48, 21, 57, 71, 109, 279, 403, 48, 
    331, 287, 233, 157, 136, 164, 225, 176, 97, 72, 35, 3, 0, 0, 6, 19, 21, 63, 201, 285, 286, 268, 254, 141, 21, 13, 40, 76, 128, 278, 388, 47, 
    324, 296, 272, 221, 179, 162, 216, 167, 106, 98, 52, 7, 0, 3, 10, 30, 47, 88, 205, 269, 260, 258, 255, 125, 1, 0, 40, 94, 141, 270, 373, 46, 
    324, 290, 282, 251, 209, 163, 188, 149, 106, 113, 67, 14, 3, 12, 19, 35, 52, 84, 156, 197, 205, 227, 240, 105, 0, 0, 42, 100, 144, 269, 367, 45, 
    320, 278, 261, 239, 216, 172, 156, 122, 102, 109, 71, 30, 16, 24, 32, 45, 65, 83, 103, 124, 151, 186, 203, 97, 0, 1, 44, 90, 143, 277, 360, 42, 
    310, 261, 251, 244, 234, 180, 117, 94, 100, 98, 67, 46, 35, 40, 49, 53, 59, 74, 92, 108, 131, 157, 172, 100, 8, 7, 48, 91, 169, 299, 358, 36, 
    301, 270, 272, 265, 249, 202, 101, 70, 86, 83, 71, 66, 62, 66, 73, 72, 77, 96, 115, 123, 134, 147, 156, 117, 52, 37, 70, 128, 220, 322, 351, 33, 
    142, 106, 108, 106, 101, 72, 12, 0, 14, 11, 3, 4, 4, 6, 11, 10, 10, 20, 30, 31, 34, 39, 41, 28, 0, 0, 4, 37, 97, 146, 148, 0, 
    
    -- channel=155
    17, 5, 5, 1, 10, 15, 26, 22, 22, 19, 11, 7, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 7, 6, 13, 5, 0, 0, 17, 11, 6, 97, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 8, 5, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 129, 
    0, 0, 0, 0, 0, 0, 16, 8, 0, 12, 9, 8, 14, 6, 8, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 137, 
    0, 0, 0, 0, 0, 0, 46, 37, 24, 36, 18, 31, 31, 15, 27, 28, 16, 32, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 140, 
    0, 0, 0, 0, 0, 0, 39, 31, 20, 31, 6, 16, 20, 0, 9, 8, 3, 19, 19, 15, 4, 0, 0, 0, 0, 0, 3, 5, 0, 0, 0, 148, 
    0, 0, 0, 0, 0, 0, 40, 35, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 0, 0, 156, 
    0, 0, 0, 0, 0, 0, 36, 61, 0, 0, 0, 0, 0, 0, 11, 16, 12, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 158, 
    0, 0, 0, 0, 0, 0, 26, 64, 0, 0, 17, 15, 25, 19, 11, 12, 7, 8, 6, 2, 12, 0, 0, 0, 0, 0, 0, 2, 15, 0, 0, 150, 
    0, 0, 0, 0, 0, 0, 45, 63, 0, 0, 0, 0, 22, 30, 11, 8, 3, 1, 9, 0, 5, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 125, 
    0, 0, 0, 0, 20, 21, 50, 59, 0, 13, 19, 0, 18, 30, 18, 12, 10, 8, 21, 1, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 131, 
    0, 0, 0, 0, 21, 0, 25, 48, 17, 29, 35, 19, 19, 23, 22, 18, 20, 23, 25, 16, 9, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 155, 
    0, 0, 0, 6, 30, 9, 34, 51, 22, 10, 21, 15, 14, 18, 25, 28, 27, 24, 12, 8, 8, 18, 22, 0, 0, 0, 0, 0, 0, 0, 0, 159, 
    0, 0, 0, 21, 26, 18, 56, 54, 7, 0, 3, 8, 16, 18, 16, 19, 14, 4, 0, 2, 8, 2, 12, 0, 0, 0, 0, 0, 0, 0, 0, 159, 
    0, 0, 5, 22, 22, 7, 33, 31, 25, 15, 19, 14, 31, 50, 36, 29, 29, 30, 30, 51, 55, 34, 27, 13, 2, 2, 11, 1, 0, 0, 0, 159, 
    0, 0, 28, 38, 37, 1, 0, 10, 28, 38, 48, 47, 44, 59, 53, 42, 34, 33, 34, 48, 57, 45, 35, 24, 23, 21, 22, 0, 0, 0, 0, 159, 
    0, 18, 51, 32, 15, 0, 12, 44, 36, 36, 21, 10, 2, 9, 25, 42, 48, 57, 58, 49, 45, 47, 54, 56, 42, 21, 20, 0, 0, 0, 0, 160, 
    0, 0, 45, 22, 0, 0, 38, 72, 49, 28, 19, 10, 17, 2, 12, 28, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 160, 
    0, 0, 57, 38, 0, 0, 61, 48, 35, 25, 23, 32, 56, 31, 40, 28, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 14, 2, 0, 0, 161, 
    0, 0, 52, 37, 1, 29, 81, 31, 16, 38, 39, 28, 39, 40, 57, 13, 17, 38, 45, 26, 34, 56, 52, 49, 19, 24, 43, 36, 16, 0, 0, 161, 
    0, 0, 54, 47, 10, 44, 82, 42, 21, 37, 47, 37, 28, 18, 27, 8, 29, 28, 9, 5, 21, 23, 17, 18, 0, 35, 57, 25, 5, 0, 0, 158, 
    0, 0, 55, 48, 10, 25, 61, 51, 41, 37, 51, 49, 37, 19, 24, 7, 33, 59, 46, 39, 45, 48, 33, 34, 28, 38, 50, 16, 0, 0, 0, 158, 
    0, 0, 60, 59, 28, 17, 36, 49, 48, 33, 40, 33, 31, 4, 27, 29, 12, 5, 6, 6, 4, 11, 0, 0, 13, 10, 15, 20, 19, 0, 0, 160, 
    0, 0, 64, 62, 41, 43, 17, 28, 47, 40, 43, 28, 43, 34, 82, 74, 16, 0, 29, 23, 7, 21, 0, 3, 79, 34, 14, 57, 58, 0, 0, 158, 
    0, 2, 72, 65, 22, 43, 19, 20, 51, 46, 49, 38, 35, 29, 74, 79, 30, 12, 56, 47, 21, 31, 1, 28, 105, 60, 17, 38, 36, 0, 0, 159, 
    0, 6, 56, 43, 0, 0, 1, 40, 57, 51, 48, 47, 44, 36, 46, 56, 45, 11, 0, 0, 0, 0, 0, 7, 51, 55, 41, 35, 14, 0, 0, 159, 
    0, 0, 25, 27, 4, 0, 0, 40, 49, 47, 47, 50, 53, 54, 51, 47, 48, 18, 0, 0, 5, 17, 11, 70, 72, 50, 45, 30, 13, 0, 0, 155, 
    0, 0, 8, 36, 36, 22, 0, 41, 40, 42, 57, 56, 47, 47, 45, 37, 34, 8, 0, 7, 31, 29, 22, 83, 86, 54, 34, 20, 17, 0, 0, 154, 
    0, 0, 6, 19, 29, 30, 2, 52, 41, 39, 57, 60, 48, 44, 43, 37, 40, 38, 11, 11, 14, 8, 13, 75, 72, 54, 32, 18, 20, 0, 0, 150, 
    0, 5, 9, 13, 19, 37, 21, 47, 41, 38, 53, 58, 48, 43, 43, 38, 32, 30, 29, 28, 23, 18, 25, 83, 66, 48, 34, 24, 15, 0, 0, 150, 
    0, 9, 12, 10, 7, 30, 43, 39, 37, 41, 50, 51, 46, 38, 37, 36, 35, 30, 26, 24, 20, 19, 20, 68, 73, 43, 30, 23, 0, 0, 0, 147, 
    0, 0, 0, 0, 4, 25, 50, 33, 38, 46, 46, 38, 38, 31, 29, 32, 30, 21, 16, 14, 11, 10, 11, 38, 58, 33, 16, 4, 0, 0, 0, 145, 
    79, 105, 110, 112, 112, 120, 135, 89, 74, 78, 82, 83, 85, 84, 86, 86, 83, 81, 86, 93, 91, 90, 90, 98, 105, 94, 78, 68, 71, 86, 106, 205, 
    
    -- channel=156
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 
    
    -- channel=157
    238, 483, 468, 464, 474, 472, 438, 403, 374, 370, 369, 369, 378, 387, 400, 414, 447, 486, 514, 523, 512, 502, 502, 508, 487, 458, 423, 428, 409, 400, 370, 187, 
    471, 803, 789, 789, 802, 791, 725, 651, 601, 599, 612, 612, 626, 650, 674, 708, 762, 798, 829, 831, 814, 801, 800, 807, 796, 768, 730, 720, 693, 670, 646, 369, 
    504, 861, 854, 850, 854, 837, 741, 647, 582, 578, 611, 605, 628, 653, 677, 726, 770, 786, 817, 801, 792, 777, 780, 799, 817, 812, 781, 747, 718, 710, 718, 422, 
    529, 898, 895, 895, 896, 858, 725, 599, 509, 496, 529, 523, 534, 540, 551, 586, 619, 642, 683, 692, 702, 720, 752, 783, 818, 819, 786, 737, 706, 722, 758, 448, 
    543, 918, 914, 916, 908, 871, 712, 548, 446, 426, 467, 471, 480, 477, 476, 483, 495, 512, 533, 552, 600, 658, 745, 793, 814, 796, 757, 693, 664, 696, 757, 457, 
    542, 917, 915, 914, 895, 855, 698, 517, 428, 414, 489, 506, 515, 514, 508, 508, 495, 487, 491, 493, 542, 625, 733, 811, 817, 779, 727, 646, 616, 644, 726, 452, 
    542, 915, 915, 904, 869, 832, 696, 538, 467, 476, 594, 641, 632, 617, 594, 575, 562, 541, 535, 544, 556, 614, 698, 774, 804, 777, 717, 652, 604, 607, 684, 420, 
    541, 914, 915, 898, 851, 811, 695, 570, 493, 501, 620, 679, 668, 664, 633, 614, 618, 608, 601, 612, 606, 621, 662, 717, 780, 777, 737, 678, 609, 572, 625, 376, 
    539, 912, 913, 892, 827, 769, 659, 537, 490, 515, 617, 660, 649, 638, 603, 593, 611, 622, 616, 649, 646, 631, 647, 693, 776, 811, 804, 750, 672, 613, 644, 382, 
    534, 905, 911, 885, 788, 717, 576, 479, 453, 477, 544, 568, 569, 568, 553, 560, 577, 593, 591, 617, 640, 646, 655, 686, 765, 839, 856, 825, 762, 724, 745, 442, 
    514, 878, 899, 877, 781, 680, 531, 444, 391, 414, 467, 493, 498, 502, 503, 516, 523, 531, 531, 548, 588, 614, 626, 660, 737, 826, 881, 882, 855, 848, 859, 512, 
    481, 836, 870, 839, 739, 643, 527, 431, 335, 334, 393, 453, 462, 460, 449, 447, 450, 453, 468, 488, 518, 540, 553, 605, 690, 807, 890, 919, 916, 916, 916, 544, 
    437, 780, 803, 769, 676, 609, 516, 441, 333, 334, 387, 454, 477, 470, 440, 411, 412, 430, 470, 491, 489, 470, 462, 511, 608, 729, 818, 870, 893, 913, 917, 543, 
    420, 738, 732, 684, 589, 548, 491, 443, 379, 401, 421, 457, 467, 456, 417, 373, 370, 394, 437, 453, 423, 376, 367, 428, 521, 617, 679, 750, 821, 881, 917, 543, 
    417, 707, 648, 561, 477, 487, 494, 474, 455, 433, 403, 377, 357, 355, 339, 318, 326, 347, 374, 370, 332, 298, 296, 339, 391, 456, 510, 592, 717, 824, 905, 544, 
    394, 669, 562, 459, 394, 452, 504, 498, 440, 394, 372, 343, 305, 300, 280, 247, 221, 194, 186, 198, 190, 184, 184, 185, 238, 312, 389, 486, 631, 774, 886, 546, 
    396, 665, 527, 423, 368, 448, 481, 448, 357, 340, 346, 354, 334, 351, 311, 271, 222, 191, 192, 235, 253, 257, 233, 188, 223, 298, 399, 491, 601, 750, 858, 544, 
    394, 668, 526, 423, 377, 430, 405, 328, 263, 317, 353, 373, 380, 409, 377, 368, 317, 324, 342, 377, 412, 413, 366, 318, 354, 412, 473, 503, 548, 691, 808, 533, 
    425, 712, 558, 435, 377, 390, 323, 222, 190, 286, 322, 322, 314, 342, 356, 404, 418, 462, 449, 470, 503, 497, 457, 424, 476, 496, 501, 467, 459, 612, 763, 521, 
    438, 726, 562, 410, 321, 314, 260, 182, 159, 233, 251, 237, 225, 250, 268, 362, 444, 495, 479, 471, 483, 479, 464, 457, 489, 496, 451, 376, 364, 543, 731, 512, 
    434, 729, 582, 424, 283, 256, 223, 180, 140, 150, 161, 187, 193, 216, 229, 289, 330, 355, 351, 348, 348, 334, 345, 342, 373, 387, 358, 337, 354, 530, 711, 502, 
    429, 731, 588, 435, 283, 232, 228, 187, 135, 107, 99, 155, 201, 290, 279, 259, 248, 302, 356, 371, 349, 326, 371, 404, 374, 352, 320, 354, 396, 527, 682, 491, 
    424, 725, 580, 414, 277, 238, 267, 237, 177, 118, 65, 94, 155, 262, 265, 214, 167, 246, 338, 384, 362, 346, 407, 436, 377, 302, 244, 309, 356, 477, 652, 486, 
    421, 712, 554, 371, 226, 227, 305, 315, 269, 162, 68, 65, 99, 175, 187, 142, 111, 200, 313, 369, 394, 411, 453, 452, 371, 244, 191, 233, 266, 417, 632, 481, 
    408, 692, 566, 384, 253, 253, 357, 386, 342, 203, 99, 52, 36, 58, 69, 63, 64, 154, 297, 422, 534, 554, 569, 479, 344, 183, 116, 141, 193, 392, 628, 471, 
    384, 669, 607, 487, 370, 339, 409, 411, 374, 244, 146, 71, 18, 0, 6, 25, 37, 91, 243, 423, 583, 612, 598, 464, 299, 125, 73, 118, 200, 411, 627, 459, 
    369, 651, 642, 590, 506, 432, 443, 395, 377, 271, 195, 107, 32, 2, 10, 36, 64, 123, 276, 449, 581, 609, 605, 472, 285, 90, 52, 124, 230, 431, 619, 447, 
    366, 648, 656, 628, 562, 471, 441, 373, 350, 278, 227, 134, 52, 17, 26, 51, 84, 142, 250, 360, 448, 499, 535, 420, 247, 63, 46, 130, 242, 435, 613, 444, 
    366, 647, 631, 597, 545, 469, 415, 340, 302, 261, 226, 149, 78, 50, 54, 78, 112, 155, 204, 255, 314, 381, 442, 366, 213, 65, 51, 125, 238, 428, 610, 444, 
    359, 624, 603, 584, 557, 488, 392, 298, 246, 234, 209, 156, 105, 90, 92, 106, 120, 143, 175, 215, 264, 318, 370, 323, 199, 83, 60, 128, 259, 450, 640, 450, 
    348, 617, 615, 612, 590, 532, 394, 278, 197, 198, 189, 162, 144, 143, 147, 156, 164, 183, 212, 245, 276, 301, 329, 305, 224, 136, 112, 186, 324, 520, 685, 452, 
    178, 336, 340, 342, 334, 297, 207, 116, 63, 63, 57, 50, 47, 52, 60, 66, 67, 76, 96, 115, 128, 138, 147, 137, 95, 48, 34, 76, 177, 306, 396, 253, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    99, 143, 143, 148, 152, 130, 118, 125, 115, 88, 80, 78, 72, 79, 81, 85, 105, 124, 140, 144, 148, 152, 158, 153, 143, 140, 139, 152, 144, 153, 134, 22, 
    100, 147, 146, 142, 139, 129, 106, 106, 104, 85, 83, 74, 80, 93, 87, 95, 125, 125, 147, 159, 160, 162, 167, 160, 149, 139, 141, 157, 167, 154, 139, 32, 
    94, 139, 140, 143, 142, 127, 77, 69, 57, 43, 55, 36, 52, 65, 63, 80, 87, 78, 102, 128, 159, 166, 160, 151, 152, 154, 158, 168, 180, 161, 150, 45, 
    101, 147, 146, 146, 144, 137, 105, 80, 48, 25, 32, 22, 26, 38, 45, 53, 59, 63, 80, 101, 133, 162, 160, 144, 155, 156, 153, 164, 176, 177, 167, 45, 
    101, 146, 146, 146, 134, 125, 80, 47, 31, 0, 0, 0, 0, 0, 0, 0, 4, 15, 29, 68, 102, 115, 138, 143, 143, 146, 151, 156, 176, 187, 177, 44, 
    101, 147, 147, 141, 128, 130, 71, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 96, 112, 137, 131, 142, 164, 160, 167, 172, 172, 46, 
    101, 146, 147, 138, 134, 137, 67, 15, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 139, 138, 140, 149, 136, 121, 115, 143, 170, 47, 
    100, 146, 146, 138, 116, 96, 38, 18, 9, 12, 44, 60, 17, 8, 0, 0, 0, 0, 0, 6, 0, 21, 90, 131, 152, 144, 136, 142, 156, 158, 167, 52, 
    98, 145, 147, 136, 94, 83, 44, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 48, 78, 101, 124, 139, 136, 139, 123, 120, 22, 
    93, 141, 144, 131, 110, 121, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 59, 104, 133, 135, 127, 106, 105, 115, 12, 
    97, 134, 133, 114, 84, 52, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 21, 79, 128, 132, 138, 147, 145, 146, 146, 30, 
    84, 119, 116, 108, 91, 54, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 31, 39, 60, 89, 117, 134, 143, 146, 146, 30, 
    78, 120, 107, 104, 91, 85, 50, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 31, 67, 99, 110, 115, 123, 138, 146, 30, 
    74, 93, 75, 71, 56, 76, 72, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 25, 39, 53, 67, 95, 115, 121, 144, 30, 
    54, 74, 71, 87, 78, 60, 31, 0, 6, 0, 0, 22, 23, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 25, 39, 97, 114, 137, 30, 
    85, 120, 71, 70, 71, 64, 36, 24, 7, 0, 0, 0, 0, 0, 0, 0, 30, 47, 45, 51, 34, 29, 55, 53, 57, 30, 2, 11, 56, 100, 129, 31, 
    57, 77, 25, 28, 36, 51, 50, 63, 6, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 2, 0, 3, 0, 0, 0, 7, 90, 120, 27, 
    59, 91, 52, 46, 45, 32, 34, 45, 0, 0, 0, 31, 30, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 42, 103, 115, 23, 
    68, 94, 47, 36, 42, 29, 18, 6, 0, 0, 0, 6, 15, 28, 27, 4, 0, 49, 64, 51, 44, 49, 50, 53, 55, 17, 21, 39, 28, 73, 105, 19, 
    67, 93, 43, 40, 49, 44, 12, 0, 0, 0, 0, 0, 0, 0, 0, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 1, 3, 58, 97, 16, 
    71, 94, 40, 19, 13, 28, 9, 0, 0, 0, 1, 0, 0, 0, 0, 0, 28, 43, 36, 35, 36, 27, 42, 42, 30, 35, 11, 0, 0, 58, 97, 13, 
    59, 81, 36, 24, 2, 0, 23, 6, 0, 0, 0, 2, 0, 0, 0, 0, 15, 6, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 65, 94, 10, 
    45, 63, 24, 26, 35, 3, 10, 0, 0, 0, 0, 0, 16, 26, 10, 0, 0, 0, 0, 8, 6, 0, 21, 9, 0, 14, 22, 35, 34, 60, 73, 0, 
    37, 46, 26, 34, 48, 52, 12, 0, 0, 0, 0, 0, 3, 18, 26, 2, 0, 38, 102, 103, 100, 80, 75, 75, 60, 3, 0, 13, 12, 43, 61, 0, 
    32, 42, 26, 0, 0, 0, 24, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 15, 21, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 28, 54, 0, 
    34, 40, 17, 0, 0, 0, 28, 5, 9, 0, 0, 0, 1, 1, 0, 1, 1, 10, 30, 32, 52, 62, 54, 16, 5, 6, 7, 0, 0, 23, 40, 0, 
    36, 31, 30, 32, 20, 10, 21, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 63, 79, 69, 52, 21, 10, 0, 0, 0, 0, 27, 39, 0, 
    15, 27, 37, 33, 16, 0, 15, 11, 10, 0, 0, 0, 0, 0, 0, 0, 6, 14, 13, 12, 9, 6, 5, 0, 0, 0, 0, 0, 3, 29, 31, 0, 
    20, 28, 19, 19, 21, 9, 3, 13, 5, 0, 0, 0, 0, 2, 0, 0, 0, 2, 4, 6, 7, 12, 18, 0, 0, 0, 2, 3, 20, 34, 28, 0, 
    24, 27, 25, 22, 13, 3, 0, 7, 0, 0, 1, 7, 0, 2, 0, 0, 0, 3, 7, 8, 13, 17, 20, 11, 0, 6, 8, 16, 24, 19, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 7, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 2, 0, 0, 0, 0, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 5, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 21, 5, 1, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 11, 17, 15, 26, 0, 0, 21, 18, 0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 24, 24, 22, 17, 18, 12, 0, 0, 0, 0, 0, 0, 0, 16, 10, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 24, 22, 21, 16, 4, 4, 0, 0, 0, 0, 0, 0, 0, 23, 12, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 21, 20, 18, 1, 0, 2, 0, 0, 0, 0, 0, 0, 22, 14, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 17, 12, 12, 8, 0, 0, 0, 0, 0, 0, 0, 3, 21, 13, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 22, 10, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 0, 0, 0, 0, 
    46, 0, 0, 0, 0, 0, 0, 0, 16, 17, 13, 12, 20, 17, 18, 16, 16, 15, 13, 9, 8, 6, 5, 5, 5, 3, 23, 28, 6, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
