LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias
					-- layer=0
					-11382, -1814, 11868, -522, -1631, 597, -2891, -200, -289, 3459, 357, 335, 5731, 485, 1682, 3401, 655, -9010, -399, 242, -552, 1885, 599, -186, 5308, 1070, 1584, 2367, 12, -2715, -663, 2588, 259, -520, -3099, -2342, -1295, 943, 1284, -6732, 1739, 921, 11797, 213, -153, 225, 1431, 851, -1680, 6007, -802, 1214, 1143, -1664, 2406, 6352, -899, 1682, 149, -2412, -997, -1864, -23, -274, -6222, -3625, -3480, -4305, -140, 2587, -211, 3618, 321, -961, -1340, 1594, -8848, 375, -2659, 911, -299, 2603, 1284, -5804, 147, 454, 134, 1805, 1723, 689, -192, 1228, 4832, 1343, -11189, -672, 2040, -4837, 241, 324, -762, 337, -16063, 237, 353, -4997, 2135, -1574, 540, -882, -4819, -706, -538, 6619, 520, -1021, -800, -326, 291, 30, 1830, 2243, -516, 3881, -86, 701, -1373, 195,

					-- weights
					-- layer=0 filter=0 channel=0
					-10, 5, -5, -10, -2, 5, 0, -23, -10,
					-- layer=0 filter=0 channel=1
					10, -5, 8, 4, 22, 14, -7, 12, 13,
					-- layer=0 filter=0 channel=2
					0, 21, 2, -3, 24, 11, -3, 9, -5,
					-- layer=0 filter=1 channel=0
					-4, -38, 0, -9, 17, 9, 24, 16, -8,
					-- layer=0 filter=1 channel=1
					-33, -11, 4, -17, 3, 15, 26, 26, -20,
					-- layer=0 filter=1 channel=2
					-44, -47, -15, -5, 7, 11, 36, 19, 14,
					-- layer=0 filter=2 channel=0
					-3, -13, 14, 5, -16, -15, -15, -15, -22,
					-- layer=0 filter=2 channel=1
					0, -21, -13, -19, -7, -29, 7, 0, 0,
					-- layer=0 filter=2 channel=2
					27, -10, 16, -17, -8, -22, -14, -19, -14,
					-- layer=0 filter=3 channel=0
					5, -9, -18, 12, -15, 0, -3, -8, -21,
					-- layer=0 filter=3 channel=1
					-22, 0, -11, 6, 3, -20, -9, 8, 6,
					-- layer=0 filter=3 channel=2
					-8, 9, -10, -16, 0, -22, -17, -19, -21,
					-- layer=0 filter=4 channel=0
					3, 10, -11, -14, 10, -9, -14, 0, -16,
					-- layer=0 filter=4 channel=1
					2, -18, 10, -3, -1, -4, 4, -20, 10,
					-- layer=0 filter=4 channel=2
					13, -4, 8, -18, -11, -18, -5, 9, 0,
					-- layer=0 filter=5 channel=0
					-3, -23, 13, -19, 12, -17, 18, 4, 1,
					-- layer=0 filter=5 channel=1
					-20, -20, -11, -12, -23, 0, 38, 17, 14,
					-- layer=0 filter=5 channel=2
					-32, -37, -20, -8, 3, -14, 32, 45, 36,
					-- layer=0 filter=6 channel=0
					19, 35, 23, 28, 32, 0, 12, 20, 22,
					-- layer=0 filter=6 channel=1
					-12, 9, 11, -1, -14, -12, -8, -30, -21,
					-- layer=0 filter=6 channel=2
					4, -11, 6, -24, -26, -29, -7, -36, -17,
					-- layer=0 filter=7 channel=0
					-24, -2, 34, -27, 3, 33, -12, -4, 12,
					-- layer=0 filter=7 channel=1
					-28, -13, 30, -22, -11, 37, -26, -2, 32,
					-- layer=0 filter=7 channel=2
					-13, -10, 30, -36, -8, 28, -26, 5, 18,
					-- layer=0 filter=8 channel=0
					-38, -44, -18, 13, 10, 28, 21, 10, 21,
					-- layer=0 filter=8 channel=1
					-16, -12, -26, -14, -5, -1, 28, 23, 14,
					-- layer=0 filter=8 channel=2
					-5, -24, -33, -20, 11, 16, 27, 28, 4,
					-- layer=0 filter=9 channel=0
					31, 2, -34, -10, -8, -33, -10, -4, 8,
					-- layer=0 filter=9 channel=1
					40, 38, 1, 26, -7, -12, -26, -21, 10,
					-- layer=0 filter=9 channel=2
					43, 14, -38, -8, -33, -29, -32, -25, -23,
					-- layer=0 filter=10 channel=0
					-17, 4, 32, -29, 9, 30, -35, -6, 28,
					-- layer=0 filter=10 channel=1
					-15, 15, 1, -38, -5, 41, -42, 2, 38,
					-- layer=0 filter=10 channel=2
					-30, 4, 14, -25, 0, 8, -24, 11, 35,
					-- layer=0 filter=11 channel=0
					-7, -8, -12, -13, -6, 2, -19, -1, -29,
					-- layer=0 filter=11 channel=1
					-6, -6, -10, 9, -2, -19, -2, -6, -13,
					-- layer=0 filter=11 channel=2
					31, 31, 14, 26, 2, 18, 3, 19, 7,
					-- layer=0 filter=12 channel=0
					21, 22, 58, 17, 11, 1, -42, -43, -59,
					-- layer=0 filter=12 channel=1
					14, 27, 64, -15, -5, 3, -42, -95, -76,
					-- layer=0 filter=12 channel=2
					10, 5, 40, -18, -20, 15, -53, -96, -69,
					-- layer=0 filter=13 channel=0
					8, 8, 0, 41, 20, -8, 38, 30, 15,
					-- layer=0 filter=13 channel=1
					1, 5, -23, -15, -10, -20, -23, -28, -6,
					-- layer=0 filter=13 channel=2
					13, -13, -24, 9, -2, -18, 13, -19, -4,
					-- layer=0 filter=14 channel=0
					-33, 26, 49, -44, -20, 24, -15, -20, -14,
					-- layer=0 filter=14 channel=1
					-30, 21, 44, -26, -9, 47, -31, -11, -6,
					-- layer=0 filter=14 channel=2
					-31, 36, 34, -54, 18, 20, -31, 7, 0,
					-- layer=0 filter=15 channel=0
					-5, -33, 22, 30, -6, -10, 40, 25, -4,
					-- layer=0 filter=15 channel=1
					-22, -47, -21, 11, -43, -41, 6, 21, -7,
					-- layer=0 filter=15 channel=2
					9, -48, -8, 36, -33, -21, 47, 19, -23,
					-- layer=0 filter=16 channel=0
					-23, -10, -17, -18, -15, -8, 34, 19, 40,
					-- layer=0 filter=16 channel=1
					-23, -11, -27, 1, -27, 8, 22, 28, 23,
					-- layer=0 filter=16 channel=2
					-2, -13, -12, -26, -1, 6, 2, 31, 10,
					-- layer=0 filter=17 channel=0
					12, 0, 4, 10, 14, 13, 23, 18, 8,
					-- layer=0 filter=17 channel=1
					-7, -26, -35, -11, 0, -3, -24, -25, 3,
					-- layer=0 filter=17 channel=2
					21, 12, -15, 14, 14, 14, 18, 6, 11,
					-- layer=0 filter=18 channel=0
					25, 18, 4, 6, -4, -2, -30, -19, -13,
					-- layer=0 filter=18 channel=1
					-2, 0, 22, -2, 0, -9, -31, -26, -10,
					-- layer=0 filter=18 channel=2
					22, 21, 29, 14, 12, 12, -13, -13, -22,
					-- layer=0 filter=19 channel=0
					28, 0, 6, -16, -37, -34, -8, 19, 32,
					-- layer=0 filter=19 channel=1
					32, 16, 4, -33, -32, -40, -8, 24, 32,
					-- layer=0 filter=19 channel=2
					35, 8, -5, -16, -39, -17, -14, 12, 29,
					-- layer=0 filter=20 channel=0
					10, 14, 16, 30, 20, 35, 36, 40, 26,
					-- layer=0 filter=20 channel=1
					-11, -21, -29, -29, -31, -19, 4, -3, -13,
					-- layer=0 filter=20 channel=2
					15, -11, 0, -18, -14, -7, 6, -10, -7,
					-- layer=0 filter=21 channel=0
					-23, 5, -3, -12, 11, 1, 15, 7, -16,
					-- layer=0 filter=21 channel=1
					-5, 24, 15, 5, 26, 13, 21, 7, 21,
					-- layer=0 filter=21 channel=2
					-21, -25, -8, -16, -16, 0, -15, -17, -12,
					-- layer=0 filter=22 channel=0
					-13, 4, 0, 32, 35, 14, 30, 27, 34,
					-- layer=0 filter=22 channel=1
					-31, -33, -31, -27, -3, -17, -6, -8, -30,
					-- layer=0 filter=22 channel=2
					5, -2, 12, 20, -8, 18, -11, 7, -10,
					-- layer=0 filter=23 channel=0
					15, -43, 20, 22, -47, 22, -2, -16, 20,
					-- layer=0 filter=23 channel=1
					10, -51, 32, 21, -50, 16, 22, -22, 17,
					-- layer=0 filter=23 channel=2
					17, -39, 31, 25, -47, 31, 23, -35, -5,
					-- layer=0 filter=24 channel=0
					13, -19, -28, -1, -8, -24, -17, -5, 12,
					-- layer=0 filter=24 channel=1
					23, 19, -17, 19, 23, 0, 15, 23, 25,
					-- layer=0 filter=24 channel=2
					12, -12, -21, -17, 0, -26, 10, -16, -3,
					-- layer=0 filter=25 channel=0
					1, -30, 10, -31, -14, 36, 7, 5, 32,
					-- layer=0 filter=25 channel=1
					-16, -32, 11, -43, -16, 35, -15, 30, 26,
					-- layer=0 filter=25 channel=2
					-19, -10, -4, -43, -9, 34, -28, 21, 42,
					-- layer=0 filter=26 channel=0
					26, -10, -27, 27, -6, -15, 27, 27, -1,
					-- layer=0 filter=26 channel=1
					17, -19, -34, 18, -19, -37, -4, 4, -12,
					-- layer=0 filter=26 channel=2
					43, 9, -12, 47, -6, -31, 7, 0, -31,
					-- layer=0 filter=27 channel=0
					-43, -36, -45, -46, -32, -41, -30, -16, -36,
					-- layer=0 filter=27 channel=1
					15, 3, 25, 16, 23, -5, 11, 3, 4,
					-- layer=0 filter=27 channel=2
					11, 15, 20, 14, 13, 25, 22, 11, 9,
					-- layer=0 filter=28 channel=0
					-35, 3, 15, -27, 26, -1, 0, 14, 17,
					-- layer=0 filter=28 channel=1
					-33, 25, 27, -29, 15, 23, -28, 7, 12,
					-- layer=0 filter=28 channel=2
					-46, 14, 8, -47, 0, 37, -31, 14, 28,
					-- layer=0 filter=29 channel=0
					-33, -6, -25, -22, -31, -25, -36, -25, -39,
					-- layer=0 filter=29 channel=1
					13, 17, 26, -2, 2, 27, 11, 17, 16,
					-- layer=0 filter=29 channel=2
					7, 0, -8, -2, 9, -1, 15, 20, -5,
					-- layer=0 filter=30 channel=0
					28, 32, 13, -8, -22, -3, -23, -25, -8,
					-- layer=0 filter=30 channel=1
					29, 9, 22, 14, -25, -1, -28, -2, 12,
					-- layer=0 filter=30 channel=2
					29, 33, -3, -13, -15, -14, -26, -1, -9,
					-- layer=0 filter=31 channel=0
					14, 25, 28, 5, 8, 0, 11, -18, -18,
					-- layer=0 filter=31 channel=1
					-4, -23, 11, -39, -18, -16, -39, -32, -23,
					-- layer=0 filter=31 channel=2
					-2, 22, 1, 7, -14, 17, -2, 8, 0,
					-- layer=0 filter=32 channel=0
					26, -5, -4, 31, -28, -14, 26, -13, -18,
					-- layer=0 filter=32 channel=1
					29, -25, -3, 31, -8, -29, 18, -4, -21,
					-- layer=0 filter=32 channel=2
					36, -1, -28, 21, -15, -4, 19, -18, -11,
					-- layer=0 filter=33 channel=0
					-16, -1, -2, 5, 10, 17, -14, 12, 16,
					-- layer=0 filter=33 channel=1
					12, -9, -9, -6, -22, -15, -15, -8, -21,
					-- layer=0 filter=33 channel=2
					-13, 14, 1, 1, -20, -12, 12, -8, -9,
					-- layer=0 filter=34 channel=0
					-6, 26, 20, 24, 2, 1, 28, 20, 17,
					-- layer=0 filter=34 channel=1
					7, -1, -27, -8, -19, -27, -28, -24, -5,
					-- layer=0 filter=34 channel=2
					1, -16, -18, -33, -11, -6, -8, -32, -18,
					-- layer=0 filter=35 channel=0
					-13, -17, 0, 7, -23, -28, -17, 8, -4,
					-- layer=0 filter=35 channel=1
					-5, -21, -4, -5, -24, -15, 9, 1, -7,
					-- layer=0 filter=35 channel=2
					-17, -2, -20, 6, -15, -4, 14, -7, -14,
					-- layer=0 filter=36 channel=0
					0, -18, -14, -11, -7, -16, -20, -26, -5,
					-- layer=0 filter=36 channel=1
					12, 15, -13, -15, -11, -8, 0, 14, -19,
					-- layer=0 filter=36 channel=2
					18, 28, 26, 21, 34, 15, 14, 23, 20,
					-- layer=0 filter=37 channel=0
					13, 2, 0, 2, -20, -15, -5, 7, 8,
					-- layer=0 filter=37 channel=1
					-21, -23, -18, -22, -3, -20, 19, 37, 41,
					-- layer=0 filter=37 channel=2
					-12, -15, -19, -25, -20, 6, 26, 21, 42,
					-- layer=0 filter=38 channel=0
					26, 25, 9, -2, 31, 13, 15, 29, 25,
					-- layer=0 filter=38 channel=1
					-21, 7, 1, -4, 4, -7, -3, -12, -16,
					-- layer=0 filter=38 channel=2
					10, -16, -20, -21, -27, -23, -7, -12, -3,
					-- layer=0 filter=39 channel=0
					-33, -26, -22, 4, -18, -11, 0, 16, 15,
					-- layer=0 filter=39 channel=1
					-8, 5, 0, 7, -16, -18, 11, 5, 3,
					-- layer=0 filter=39 channel=2
					8, 3, -1, 20, 13, 24, 6, 13, 28,
					-- layer=0 filter=40 channel=0
					1, 21, 26, 22, 33, 20, -10, 8, 21,
					-- layer=0 filter=40 channel=1
					0, -1, -10, -22, -22, -22, -26, -28, -32,
					-- layer=0 filter=40 channel=2
					-2, 29, 32, -13, 0, 0, -22, -24, -6,
					-- layer=0 filter=41 channel=0
					46, 9, -28, 20, -47, -38, -11, -49, 30,
					-- layer=0 filter=41 channel=1
					30, 17, -25, 41, -11, -31, 8, -45, 31,
					-- layer=0 filter=41 channel=2
					42, -3, -19, 39, -23, -11, 8, -35, 13,
					-- layer=0 filter=42 channel=0
					-15, 2, 0, -2, -5, -15, -19, 2, 5,
					-- layer=0 filter=42 channel=1
					-7, -21, 8, -29, -39, 2, -21, -15, -9,
					-- layer=0 filter=42 channel=2
					-6, -3, 29, -13, -29, -17, -11, -12, 10,
					-- layer=0 filter=43 channel=0
					-37, -39, -7, -4, -13, 3, 2, 47, 35,
					-- layer=0 filter=43 channel=1
					-36, -47, 1, -8, 7, 14, 26, 29, 28,
					-- layer=0 filter=43 channel=2
					-21, -36, 0, -6, 11, 6, -10, 28, 10,
					-- layer=0 filter=44 channel=0
					13, -10, -18, 23, 0, -11, 28, 10, -27,
					-- layer=0 filter=44 channel=1
					22, -5, -16, 8, 7, -38, 29, 0, -32,
					-- layer=0 filter=44 channel=2
					25, -8, -17, 33, 17, -42, 33, -2, -35,
					-- layer=0 filter=45 channel=0
					10, -8, -5, -7, 2, -8, 25, 9, 1,
					-- layer=0 filter=45 channel=1
					-10, -7, -26, 23, 15, -23, 11, 25, 1,
					-- layer=0 filter=45 channel=2
					-15, -27, -27, 13, -15, -40, -5, 19, -19,
					-- layer=0 filter=46 channel=0
					21, 12, 24, -33, -20, -29, 4, 14, 21,
					-- layer=0 filter=46 channel=1
					12, 12, 18, -33, -40, -49, 7, 19, 15,
					-- layer=0 filter=46 channel=2
					3, 7, 28, -34, -41, -42, 42, 13, 25,
					-- layer=0 filter=47 channel=0
					18, -9, 2, 35, -20, -1, 23, -47, -6,
					-- layer=0 filter=47 channel=1
					4, -19, -3, 17, -53, 12, 32, -31, 19,
					-- layer=0 filter=47 channel=2
					6, -28, 11, 6, -51, 39, 1, -49, 46,
					-- layer=0 filter=48 channel=0
					3, -16, 7, 0, -1, 13, 4, -11, 11,
					-- layer=0 filter=48 channel=1
					25, 25, 18, 19, 17, 25, -13, 3, 14,
					-- layer=0 filter=48 channel=2
					-29, -22, -19, -7, -9, -32, -30, -30, 6,
					-- layer=0 filter=49 channel=0
					1, 16, 21, 18, 8, -5, 8, -14, 6,
					-- layer=0 filter=49 channel=1
					20, -4, -18, 20, -6, 12, 5, -16, -6,
					-- layer=0 filter=49 channel=2
					-2, -15, -33, -25, -22, -29, -10, -40, 6,
					-- layer=0 filter=50 channel=0
					3, -16, -21, 1, -9, 10, 7, 6, 1,
					-- layer=0 filter=50 channel=1
					6, -3, -8, -20, -24, -9, -34, -18, -25,
					-- layer=0 filter=50 channel=2
					13, 13, -10, 0, 2, -10, -23, -18, -4,
					-- layer=0 filter=51 channel=0
					2, -1, 26, -10, 14, 29, -18, -1, 14,
					-- layer=0 filter=51 channel=1
					0, -12, 29, -12, -2, 31, -22, 18, 15,
					-- layer=0 filter=51 channel=2
					-32, -4, -11, -42, 5, -16, -35, 0, -14,
					-- layer=0 filter=52 channel=0
					-18, -19, -11, 12, -5, 6, 0, -13, -13,
					-- layer=0 filter=52 channel=1
					12, -4, -7, 6, 20, 18, -17, -4, -10,
					-- layer=0 filter=52 channel=2
					-22, -15, -23, 8, 15, 11, -3, -17, 4,
					-- layer=0 filter=53 channel=0
					-12, -9, 15, -9, -7, 12, 10, 3, -12,
					-- layer=0 filter=53 channel=1
					-2, 0, -8, -8, -21, -18, -25, -4, -4,
					-- layer=0 filter=53 channel=2
					-12, -27, -6, -5, 2, -13, -19, -6, 3,
					-- layer=0 filter=54 channel=0
					24, -17, -5, -29, -29, 6, -27, 25, 38,
					-- layer=0 filter=54 channel=1
					-14, -26, 6, -51, -30, 32, -6, 40, 48,
					-- layer=0 filter=54 channel=2
					5, -16, -20, -41, -34, 29, -29, 39, 47,
					-- layer=0 filter=55 channel=0
					-22, -22, -15, 0, -29, -24, -3, -26, -23,
					-- layer=0 filter=55 channel=1
					-11, 14, -16, 5, -9, 6, 0, 1, 1,
					-- layer=0 filter=55 channel=2
					18, 7, -5, 21, 30, 22, 15, 9, 24,
					-- layer=0 filter=56 channel=0
					-19, -4, -1, -2, 12, -6, -11, 1, -3,
					-- layer=0 filter=56 channel=1
					-3, 3, 12, -5, -14, 13, -7, -12, -8,
					-- layer=0 filter=56 channel=2
					-17, -1, -7, 0, 9, -11, -19, 5, 9,
					-- layer=0 filter=57 channel=0
					3, 15, 21, -19, 5, 28, -20, 1, 36,
					-- layer=0 filter=57 channel=1
					-25, -17, -1, -31, -9, 17, -42, -20, 20,
					-- layer=0 filter=57 channel=2
					-26, 19, 11, -21, 5, 14, -26, 15, 25,
					-- layer=0 filter=58 channel=0
					21, -25, 4, 8, -25, 26, -13, -22, 32,
					-- layer=0 filter=58 channel=1
					11, -38, 23, 13, -46, 36, 4, -44, 37,
					-- layer=0 filter=58 channel=2
					7, -3, -1, 3, -35, 7, 19, -40, 34,
					-- layer=0 filter=59 channel=0
					-23, -28, 0, -13, 2, 8, -1, 7, -12,
					-- layer=0 filter=59 channel=1
					-9, -15, -7, 0, -17, 5, 8, 6, -20,
					-- layer=0 filter=59 channel=2
					-14, -3, 5, -15, -11, 11, 0, 2, -6,
					-- layer=0 filter=60 channel=0
					-16, 3, -25, -25, 0, -20, 3, -19, -12,
					-- layer=0 filter=60 channel=1
					-9, 13, -5, -18, 2, -17, -8, -10, -25,
					-- layer=0 filter=60 channel=2
					-5, 9, -14, -15, -7, -2, -27, 9, -5,
					-- layer=0 filter=61 channel=0
					9, -23, -8, 3, -22, -3, 12, 2, -9,
					-- layer=0 filter=61 channel=1
					-17, -22, -18, 10, -15, -8, -17, 2, 0,
					-- layer=0 filter=61 channel=2
					-25, -18, -13, 5, -3, 8, -19, -5, -8,
					-- layer=0 filter=62 channel=0
					-1, -32, -29, -17, -14, 10, 4, 42, 38,
					-- layer=0 filter=62 channel=1
					-18, -19, -16, 0, -12, 4, -1, 31, 30,
					-- layer=0 filter=62 channel=2
					-1, -35, -25, -7, -4, -7, 24, 27, 26,
					-- layer=0 filter=63 channel=0
					8, -5, -21, -19, -25, -29, -5, -14, -29,
					-- layer=0 filter=63 channel=1
					-4, 25, 23, 19, 18, 4, -2, -12, -18,
					-- layer=0 filter=63 channel=2
					13, 20, 24, 25, 5, 20, 4, 5, 9,
					-- layer=0 filter=64 channel=0
					3, -8, 8, 14, 16, 14, 15, 6, 4,
					-- layer=0 filter=64 channel=1
					-32, -4, 1, -10, 9, 7, 4, -22, -4,
					-- layer=0 filter=64 channel=2
					-29, -24, -4, -25, -1, 0, 12, 14, -22,
					-- layer=0 filter=65 channel=0
					-13, 4, -9, -9, -1, 3, 7, 17, 9,
					-- layer=0 filter=65 channel=1
					9, 21, 8, -7, 18, 25, 16, 19, 17,
					-- layer=0 filter=65 channel=2
					-22, -8, 3, -7, -25, -26, -24, -25, -35,
					-- layer=0 filter=66 channel=0
					-12, -7, 9, -20, -20, -2, -15, -19, -24,
					-- layer=0 filter=66 channel=1
					10, 21, -1, 20, 0, -2, 9, 23, 0,
					-- layer=0 filter=66 channel=2
					-7, -10, 17, -3, 21, 24, 16, 6, 21,
					-- layer=0 filter=67 channel=0
					19, 25, 19, -11, 18, -8, 4, -6, -12,
					-- layer=0 filter=67 channel=1
					37, 16, 26, 5, 15, 33, 7, 6, 0,
					-- layer=0 filter=67 channel=2
					-41, -31, -40, -33, -50, -32, 1, -15, -13,
					-- layer=0 filter=68 channel=0
					14, -4, -12, 20, 15, -35, 10, 18, -23,
					-- layer=0 filter=68 channel=1
					5, 21, -33, 25, 16, -34, 18, 13, -36,
					-- layer=0 filter=68 channel=2
					13, 23, -28, 29, 21, -46, 9, 1, -24,
					-- layer=0 filter=69 channel=0
					0, -25, -29, 18, -21, -38, 26, 41, 24,
					-- layer=0 filter=69 channel=1
					-20, -40, -23, 8, -13, -11, 37, 33, 8,
					-- layer=0 filter=69 channel=2
					15, -31, -4, 15, -10, -36, 33, 22, 6,
					-- layer=0 filter=70 channel=0
					33, 32, 33, -1, 20, 25, -24, -15, -11,
					-- layer=0 filter=70 channel=1
					-6, -17, -14, 1, -16, 3, 6, -22, -9,
					-- layer=0 filter=70 channel=2
					-26, -5, -2, -16, -40, -20, 10, -2, -13,
					-- layer=0 filter=71 channel=0
					-25, -24, 4, -30, -9, -22, -6, 7, -5,
					-- layer=0 filter=71 channel=1
					23, 20, 28, -4, 13, 18, 2, 30, 29,
					-- layer=0 filter=71 channel=2
					-12, -23, -5, -5, -12, -20, 7, -11, -11,
					-- layer=0 filter=72 channel=0
					1, 28, -3, 5, -38, -13, -13, 13, 12,
					-- layer=0 filter=72 channel=1
					31, 6, 16, -14, -30, -21, -20, 14, 12,
					-- layer=0 filter=72 channel=2
					30, 11, 16, 8, -27, -40, -15, -15, 12,
					-- layer=0 filter=73 channel=0
					-14, -11, -16, -23, -5, 7, 11, 5, -20,
					-- layer=0 filter=73 channel=1
					-4, 12, 15, -17, 4, 8, -16, 11, -17,
					-- layer=0 filter=73 channel=2
					10, -20, 2, 3, -3, -19, 10, 9, -19,
					-- layer=0 filter=74 channel=0
					14, 32, -7, 11, 17, -2, -10, 1, -27,
					-- layer=0 filter=74 channel=1
					10, 35, -11, -10, 25, -39, -3, 3, -41,
					-- layer=0 filter=74 channel=2
					-12, 24, 10, 6, 14, -40, -3, 7, -35,
					-- layer=0 filter=75 channel=0
					-7, 14, 45, -28, -38, -16, -4, -9, -40,
					-- layer=0 filter=75 channel=1
					24, 12, 53, -6, -3, 14, -2, -20, -23,
					-- layer=0 filter=75 channel=2
					8, 14, 60, -15, -27, 2, -3, -38, -29,
					-- layer=0 filter=76 channel=0
					22, 0, -23, 8, 1, -11, 9, -14, -21,
					-- layer=0 filter=76 channel=1
					33, 22, 5, 25, 14, -24, 14, -27, -8,
					-- layer=0 filter=76 channel=2
					34, 30, -5, 35, -2, -20, -6, -3, -31,
					-- layer=0 filter=77 channel=0
					-7, 4, -16, -19, 8, -14, 10, 6, -18,
					-- layer=0 filter=77 channel=1
					28, 24, -4, 25, 25, 22, -6, 28, 21,
					-- layer=0 filter=77 channel=2
					-30, -26, -8, -21, -4, -5, -13, -26, 3,
					-- layer=0 filter=78 channel=0
					7, -1, 5, -20, 6, 0, 2, -7, -18,
					-- layer=0 filter=78 channel=1
					-15, -7, -17, -37, 0, 18, -36, 1, 17,
					-- layer=0 filter=78 channel=2
					-15, 16, 5, -10, 7, 8, -21, 18, 19,
					-- layer=0 filter=79 channel=0
					-8, -38, -26, -5, -15, 6, 18, 39, 42,
					-- layer=0 filter=79 channel=1
					-13, -28, -31, -17, -24, 12, 25, 19, 36,
					-- layer=0 filter=79 channel=2
					-18, 6, -20, 10, -18, -12, 16, 5, 32,
					-- layer=0 filter=80 channel=0
					-20, -12, -6, -12, 1, 10, -1, -11, -16,
					-- layer=0 filter=80 channel=1
					0, 0, -17, -11, -14, 10, 8, -8, 0,
					-- layer=0 filter=80 channel=2
					-4, -11, 2, -3, -11, 7, 2, 9, -18,
					-- layer=0 filter=81 channel=0
					-33, -30, -34, 0, 10, -22, -4, -6, 12,
					-- layer=0 filter=81 channel=1
					29, 20, 14, 23, 23, 23, 27, 13, 35,
					-- layer=0 filter=81 channel=2
					-32, 0, -6, 3, -23, -8, -27, -7, 9,
					-- layer=0 filter=82 channel=0
					11, -19, 3, 19, -2, -2, 1, -1, 8,
					-- layer=0 filter=82 channel=1
					4, 28, 27, 11, 20, 25, 7, 22, 7,
					-- layer=0 filter=82 channel=2
					-28, -33, -23, -14, -4, -24, -8, -25, -14,
					-- layer=0 filter=83 channel=0
					11, -15, -27, 30, 21, -27, 31, 11, 6,
					-- layer=0 filter=83 channel=1
					-7, -44, -27, 35, 19, -25, 23, 6, 14,
					-- layer=0 filter=83 channel=2
					-20, -49, -30, 32, 6, -26, 29, 25, -4,
					-- layer=0 filter=84 channel=0
					-1, 1, 0, 30, 4, 4, -13, -12, -10,
					-- layer=0 filter=84 channel=1
					25, 15, 0, 34, 25, -19, -17, -43, -27,
					-- layer=0 filter=84 channel=2
					25, 31, 21, 24, 7, -15, -17, -45, -40,
					-- layer=0 filter=85 channel=0
					31, -36, 20, 5, -18, 2, -7, -13, 24,
					-- layer=0 filter=85 channel=1
					17, -37, 18, 23, -33, 4, 3, -35, 33,
					-- layer=0 filter=85 channel=2
					26, -39, 0, 8, -31, 21, -2, -29, 42,
					-- layer=0 filter=86 channel=0
					0, 14, 13, -18, -5, -11, 1, 3, 12,
					-- layer=0 filter=86 channel=1
					-16, -10, -14, -16, -21, -20, 0, -19, -19,
					-- layer=0 filter=86 channel=2
					-4, 14, 12, 21, 19, 29, 29, 23, 21,
					-- layer=0 filter=87 channel=0
					34, 34, 6, -12, -21, -28, -25, -14, 28,
					-- layer=0 filter=87 channel=1
					27, 14, -19, -15, -40, -45, 4, 13, 15,
					-- layer=0 filter=87 channel=2
					30, 7, -12, -26, -54, -9, 0, 10, 44,
					-- layer=0 filter=88 channel=0
					13, -13, 5, -15, -5, 2, -4, -15, 15,
					-- layer=0 filter=88 channel=1
					4, 18, -2, 23, 0, 0, 11, 19, -8,
					-- layer=0 filter=88 channel=2
					-26, -14, -31, 0, -11, -32, -30, -36, -12,
					-- layer=0 filter=89 channel=0
					-10, -8, 13, 21, 11, -15, 7, -11, 3,
					-- layer=0 filter=89 channel=1
					12, 24, 26, 33, 31, 12, 29, 21, -10,
					-- layer=0 filter=89 channel=2
					-11, -9, -11, -14, -28, -18, -12, -23, -33,
					-- layer=0 filter=90 channel=0
					21, -5, -37, 26, 13, -30, 27, 22, -26,
					-- layer=0 filter=90 channel=1
					17, -7, -28, 9, 20, -25, 8, 2, -11,
					-- layer=0 filter=90 channel=2
					32, -1, -37, 16, -8, -28, 24, 29, -26,
					-- layer=0 filter=91 channel=0
					32, 36, 34, 33, 11, 12, 16, 17, 18,
					-- layer=0 filter=91 channel=1
					-17, -20, -2, 1, -20, 3, -22, -18, -5,
					-- layer=0 filter=91 channel=2
					-20, -1, -4, -30, -6, 4, -21, -15, 0,
					-- layer=0 filter=92 channel=0
					30, -17, -64, 40, -16, -52, 40, 13, -53,
					-- layer=0 filter=92 channel=1
					27, -11, -44, 28, -11, -54, 47, 10, -40,
					-- layer=0 filter=92 channel=2
					1, 8, -32, 36, 14, -38, 31, 0, -47,
					-- layer=0 filter=93 channel=0
					2, -19, -4, -7, -2, -5, 2, -14, 17,
					-- layer=0 filter=93 channel=1
					0, 17, 21, 21, 21, 25, 25, 30, 17,
					-- layer=0 filter=93 channel=2
					-17, -10, -20, -10, -1, -11, -4, -7, -20,
					-- layer=0 filter=94 channel=0
					-12, 19, 19, -15, -4, 13, 7, 6, -14,
					-- layer=0 filter=94 channel=1
					-9, 2, 14, -1, -18, -2, -20, -4, -7,
					-- layer=0 filter=94 channel=2
					12, 27, 16, 10, 26, 21, -12, 15, 17,
					-- layer=0 filter=95 channel=0
					-4, 19, 31, -11, 1, -14, 10, -26, -32,
					-- layer=0 filter=95 channel=1
					27, 33, 10, 18, 20, -3, -4, -26, -39,
					-- layer=0 filter=95 channel=2
					24, 31, 9, 5, -11, 11, -13, -38, -30,
					-- layer=0 filter=96 channel=0
					-15, -16, -2, 7, 5, -30, -25, -17, -34,
					-- layer=0 filter=96 channel=1
					-3, 5, 6, 4, 10, -13, 10, 0, -20,
					-- layer=0 filter=96 channel=2
					-10, -16, -14, -4, 2, 6, -7, -22, 2,
					-- layer=0 filter=97 channel=0
					-8, -25, -27, 0, 8, -3, -1, 15, 2,
					-- layer=0 filter=97 channel=1
					13, 12, 19, 2, 4, 23, 17, 11, 14,
					-- layer=0 filter=97 channel=2
					-11, -5, 13, 7, 9, 14, -2, 19, -18,
					-- layer=0 filter=98 channel=0
					-31, -47, -22, 19, 28, 19, 1, 32, 32,
					-- layer=0 filter=98 channel=1
					-38, -22, -36, -4, 3, 18, 0, 24, 27,
					-- layer=0 filter=98 channel=2
					-17, -27, -21, 15, 13, 13, -3, 2, 16,
					-- layer=0 filter=99 channel=0
					-21, 27, -3, -32, 37, 2, -37, 32, -17,
					-- layer=0 filter=99 channel=1
					-16, 42, -22, -13, 40, -5, -39, 33, 2,
					-- layer=0 filter=99 channel=2
					-18, 45, -29, -37, 44, -12, -35, 16, 12,
					-- layer=0 filter=100 channel=0
					-1, 10, 4, -2, -17, -33, -10, -33, -37,
					-- layer=0 filter=100 channel=1
					-12, 6, 14, -1, -15, -1, 4, -9, 6,
					-- layer=0 filter=100 channel=2
					20, 19, 1, 25, 22, -4, 23, 19, -5,
					-- layer=0 filter=101 channel=0
					14, 19, 30, 27, 31, 25, 15, 4, 7,
					-- layer=0 filter=101 channel=1
					2, 0, 11, -21, 0, -5, 12, -19, -4,
					-- layer=0 filter=101 channel=2
					-24, -12, -21, -3, -4, -27, -7, -18, -23,
					-- layer=0 filter=102 channel=0
					26, 28, 24, 13, 13, 2, -12, 17, 12,
					-- layer=0 filter=102 channel=1
					11, 2, 14, -21, 7, 3, 3, -28, -4,
					-- layer=0 filter=102 channel=2
					-7, 8, 12, 4, -5, 12, 0, 10, -12,
					-- layer=0 filter=103 channel=0
					2, -14, -10, -18, 0, 6, -23, -36, -26,
					-- layer=0 filter=103 channel=1
					8, -13, 8, 5, 9, -20, -13, -9, -23,
					-- layer=0 filter=103 channel=2
					27, 7, 5, 19, 16, 3, 2, 15, 17,
					-- layer=0 filter=104 channel=0
					20, -18, 8, -1, -27, 20, 10, -23, 3,
					-- layer=0 filter=104 channel=1
					24, -31, 2, 8, -44, 9, 1, -25, 17,
					-- layer=0 filter=104 channel=2
					24, -36, 13, 15, -29, 21, 19, -20, 7,
					-- layer=0 filter=105 channel=0
					-21, 0, -13, -27, 6, 14, -30, 6, -6,
					-- layer=0 filter=105 channel=1
					8, 24, 15, 16, 15, 17, -6, -1, 21,
					-- layer=0 filter=105 channel=2
					-6, 7, 10, 0, 26, 18, -1, 1, 13,
					-- layer=0 filter=106 channel=0
					22, 25, 6, 33, 27, 20, 23, 12, -14,
					-- layer=0 filter=106 channel=1
					14, -10, -12, 23, -10, -28, 11, -14, -35,
					-- layer=0 filter=106 channel=2
					10, -5, -29, 1, -24, -11, 14, -20, -31,
					-- layer=0 filter=107 channel=0
					-24, -11, 9, 8, -3, -7, -2, -11, 1,
					-- layer=0 filter=107 channel=1
					-10, -24, -26, 5, 11, -1, 11, 2, -15,
					-- layer=0 filter=107 channel=2
					-23, -23, -7, -21, 4, -14, -21, -16, 1,
					-- layer=0 filter=108 channel=0
					12, -10, -22, 14, -8, -8, 20, -6, 4,
					-- layer=0 filter=108 channel=1
					32, -15, -24, 42, -6, -15, 41, -18, -25,
					-- layer=0 filter=108 channel=2
					35, -4, -33, 28, -22, -33, 39, -6, -12,
					-- layer=0 filter=109 channel=0
					8, -10, -3, -5, 8, -11, -17, 4, 1,
					-- layer=0 filter=109 channel=1
					-2, 8, 8, 0, -18, 9, -19, -4, 0,
					-- layer=0 filter=109 channel=2
					2, -19, -15, -10, -13, -3, 10, -5, -9,
					-- layer=0 filter=110 channel=0
					-25, -3, 10, 6, 5, 6, -12, -5, -14,
					-- layer=0 filter=110 channel=1
					-2, 4, 20, -1, -5, -5, -28, 8, 8,
					-- layer=0 filter=110 channel=2
					-4, 0, 0, -3, 6, 2, -17, -23, 8,
					-- layer=0 filter=111 channel=0
					5, 26, 4, -2, 7, 9, -19, -40, -4,
					-- layer=0 filter=111 channel=1
					18, 31, 17, 14, 25, 0, -34, -31, -12,
					-- layer=0 filter=111 channel=2
					28, 9, 8, 14, 10, -9, -30, -37, -10,
					-- layer=0 filter=112 channel=0
					-22, 8, 0, 12, 32, 22, -14, -24, -39,
					-- layer=0 filter=112 channel=1
					8, 13, 3, 35, 3, 16, -5, -36, -21,
					-- layer=0 filter=112 channel=2
					3, -16, 0, 14, 32, 30, -7, -25, -34,
					-- layer=0 filter=113 channel=0
					3, 15, 29, 5, 26, 2, 8, 24, 24,
					-- layer=0 filter=113 channel=1
					-33, -37, 5, -48, -38, -11, -20, -28, 14,
					-- layer=0 filter=113 channel=2
					-10, -11, -5, -7, -31, -8, -16, -6, 5,
					-- layer=0 filter=114 channel=0
					-33, -38, -14, -18, -32, -28, 33, 16, 13,
					-- layer=0 filter=114 channel=1
					-29, -2, -24, 8, -9, -23, 33, 19, 3,
					-- layer=0 filter=114 channel=2
					-10, -4, 12, 8, 9, -19, 20, 38, 31,
					-- layer=0 filter=115 channel=0
					-17, 0, 26, -14, 15, 31, -24, 5, 28,
					-- layer=0 filter=115 channel=1
					-30, -25, 11, -32, -26, -4, -17, -15, 12,
					-- layer=0 filter=115 channel=2
					12, 25, 19, 10, 25, 1, 5, 9, 30,
					-- layer=0 filter=116 channel=0
					0, -6, 4, -3, 10, -16, -14, -9, -4,
					-- layer=0 filter=116 channel=1
					2, -8, -7, -13, -10, -9, -14, 2, -11,
					-- layer=0 filter=116 channel=2
					-21, 10, 9, 13, -5, -10, 4, -15, 0,
					-- layer=0 filter=117 channel=0
					3, -1, -3, -4, 27, 29, -27, -23, -7,
					-- layer=0 filter=117 channel=1
					-3, -6, -3, 11, 30, 44, -25, -32, -20,
					-- layer=0 filter=117 channel=2
					0, 5, -20, 27, 22, 36, -11, -31, -29,
					-- layer=0 filter=118 channel=0
					35, 19, 15, 2, 15, -22, -26, -18, -9,
					-- layer=0 filter=118 channel=1
					33, 17, 4, 20, 15, -14, -23, -13, -29,
					-- layer=0 filter=118 channel=2
					34, 14, 12, -9, 0, -14, -12, -22, -25,
					-- layer=0 filter=119 channel=0
					34, -15, -16, 38, -21, -17, 2, 1, -14,
					-- layer=0 filter=119 channel=1
					35, -1, -39, 35, 2, -36, 27, -19, 0,
					-- layer=0 filter=119 channel=2
					40, -6, -35, 13, -5, -15, 17, -9, -8,
					-- layer=0 filter=120 channel=0
					7, -13, -7, -5, 1, 18, -6, 12, 12,
					-- layer=0 filter=120 channel=1
					-6, 2, 0, 1, 9, 31, 11, 5, 16,
					-- layer=0 filter=120 channel=2
					-33, -27, -6, -35, -26, 14, -22, -19, 25,
					-- layer=0 filter=121 channel=0
					15, 11, 9, -42, -35, -22, 7, -21, -8,
					-- layer=0 filter=121 channel=1
					10, 31, 30, -33, -13, 7, -4, 2, -14,
					-- layer=0 filter=121 channel=2
					11, 2, -10, -29, 2, -12, 25, 5, 14,
					-- layer=0 filter=122 channel=0
					-8, -4, -11, -16, -9, -5, -18, -1, -3,
					-- layer=0 filter=122 channel=1
					-3, 3, -9, 0, 10, 13, 11, -15, -1,
					-- layer=0 filter=122 channel=2
					-8, -6, -5, 15, -6, 0, -1, -10, -9,
					-- layer=0 filter=123 channel=0
					-14, -7, 10, -33, -36, 0, -17, -33, -18,
					-- layer=0 filter=123 channel=1
					18, 16, 9, -14, -18, 5, 18, 0, 16,
					-- layer=0 filter=123 channel=2
					15, 14, 19, -5, 14, -11, 9, 9, 5,
					-- layer=0 filter=124 channel=0
					-8, -23, -9, 10, 11, -18, 0, -18, -6,
					-- layer=0 filter=124 channel=1
					-20, 6, 9, 3, 10, -13, -19, 15, 13,
					-- layer=0 filter=124 channel=2
					-16, -26, 3, 1, -14, -24, -16, 6, -11,
					-- layer=0 filter=125 channel=0
					42, 23, 32, 18, 23, 28, -17, -16, -8,
					-- layer=0 filter=125 channel=1
					-15, 0, -13, -25, 10, 17, -20, -14, 1,
					-- layer=0 filter=125 channel=2
					-31, -14, -27, -34, -28, -23, 1, 4, 14,
					-- layer=0 filter=126 channel=0
					-1, -23, -32, 31, 19, 18, -9, 8, -15,
					-- layer=0 filter=126 channel=1
					-24, -27, -2, 27, 26, 27, -12, 13, 6,
					-- layer=0 filter=126 channel=2
					-30, -34, -37, 30, 9, 19, -10, 17, 15,
					-- layer=0 filter=127 channel=0
					35, 21, 19, 8, -4, -18, -28, -16, -19,
					-- layer=0 filter=127 channel=1
					-1, 31, 32, -3, 0, -18, -9, -1, -27,
					-- layer=0 filter=127 channel=2
					22, 2, 12, 21, 0, 2, -25, -21, -24,

					-- test image
					-- image=0 channel=0 column=0
					158,159,165,166,160,156,162,159,158,159,161,160,161,166,169,170,167,162,160,160,156,149,150,148,149,143,140,141,143,137,126,116,
					-- image=0 channel=0 column=1
					152,151,159,166,162,160,164,162,163,156,155,159,163,170,171,171,169,160,154,151,145,139,140,141,149,147,145,142,143,136,125,119,
					-- image=0 channel=0 column=2
					151,151,158,167,160,163,165,165,163,162,158,157,161,166,167,169,170,159,145,121,110,98,101,114,120,134,143,140,142,139,130,120,
					-- image=0 channel=0 column=3
					155,155,160,174,167,167,169,169,165,165,167,191,177,157,162,164,158,149,104,103,98,92,80,74,86,83,113,132,140,140,136,127,
					-- image=0 channel=0 column=4
					155,156,161,170,169,163,169,166,164,164,173,246,195,151,146,142,111,78,85,113,112,106,97,93,74,84,85,105,128,138,133,129,
					-- image=0 channel=0 column=5
					148,133,130,147,161,165,167,167,163,165,163,180,157,128,97,66,69,66,89,118,122,119,114,94,99,91,58,67,108,140,138,134,
					-- image=0 channel=0 column=6
					127,109,47,88,153,170,168,170,169,166,164,147,129,127,100,68,78,72,83,132,146,124,105,107,115,85,63,46,79,132,141,134,
					-- image=0 channel=0 column=7
					131,99,42,70,143,167,165,168,171,161,140,120,130,144,116,88,91,85,77,124,163,136,102,106,100,85,54,49,57,107,138,136,
					-- image=0 channel=0 column=8
					170,103,54,124,153,161,163,166,165,174,113,125,157,156,121,86,82,84,80,81,138,146,113,87,83,86,71,56,40,74,133,137,
					-- image=0 channel=0 column=9
					180,134,94,154,174,158,156,153,207,237,207,156,174,148,125,93,86,74,59,76,137,143,133,106,86,87,84,75,50,40,95,132,
					-- image=0 channel=0 column=10
					183,108,142,165,177,155,159,122,213,237,220,164,183,156,125,120,78,80,45,91,175,157,155,107,87,103,88,78,59,41,59,104,
					-- image=0 channel=0 column=11
					188,100,135,170,187,166,173,134,117,194,199,170,185,189,134,117,102,84,38,125,210,160,146,93,83,94,104,85,73,55,62,76,
					-- image=0 channel=0 column=12
					189,90,127,175,174,166,178,159,97,168,168,137,186,216,160,123,120,115,50,150,194,155,123,91,84,84,95,86,84,73,79,73,
					-- image=0 channel=0 column=13
					189,93,152,185,119,136,173,167,103,147,145,167,189,226,180,141,126,117,71,154,186,149,114,87,80,72,80,99,100,90,97,94,
					-- image=0 channel=0 column=14
					194,108,168,186,105,99,156,167,100,115,138,198,190,172,145,154,146,103,71,152,179,137,130,110,85,91,95,109,115,100,97,117,
					-- image=0 channel=0 column=15
					197,132,172,184,130,78,140,155,115,130,143,230,242,145,135,131,121,108,95,144,168,152,112,87,71,87,105,112,120,103,121,136,
					-- image=0 channel=0 column=16
					203,146,168,191,168,78,126,138,138,96,154,173,162,140,113,113,101,105,112,171,156,148,135,109,78,79,94,101,107,125,151,144,
					-- image=0 channel=0 column=17
					214,163,164,183,176,94,96,156,148,106,129,118,114,116,102,115,86,101,144,118,68,128,133,75,60,58,71,102,116,143,150,140,
					-- image=0 channel=0 column=18
					212,178,167,173,176,124,86,141,153,135,104,77,134,124,129,147,85,92,150,132,117,107,75,64,44,65,86,133,155,160,154,151,
					-- image=0 channel=0 column=19
					199,187,171,174,177,144,86,119,122,137,144,70,129,108,145,184,116,73,131,137,134,89,51,52,47,90,121,163,171,164,158,149,
					-- image=0 channel=0 column=20
					165,195,179,177,181,152,99,131,171,103,93,80,93,122,178,191,150,100,89,87,60,46,38,24,46,60,108,144,144,128,127,120,
					-- image=0 channel=0 column=21
					117,195,177,178,181,138,83,150,245,219,133,134,149,176,190,194,168,125,110,61,35,34,49,58,61,58,69,72,78,69,59,55,
					-- image=0 channel=0 column=22
					79,175,174,176,177,140,109,211,253,252,208,124,114,124,116,122,104,68,68,60,52,50,51,56,56,51,43,51,59,48,43,42,
					-- image=0 channel=0 column=23
					41,96,144,168,178,165,165,246,253,227,110,60,53,49,49,48,45,42,46,42,38,46,46,43,42,46,46,50,55,53,51,45,
					-- image=0 channel=0 column=24
					29,29,59,131,166,132,194,254,241,141,61,50,50,51,49,50,47,42,39,34,35,39,38,42,45,56,62,59,56,50,46,51,
					-- image=0 channel=0 column=25
					48,30,34,73,128,128,215,256,187,66,54,50,52,52,46,45,43,41,36,39,40,40,43,46,59,62,64,59,54,50,70,83,
					-- image=0 channel=0 column=26
					52,35,31,41,66,128,224,240,124,58,49,56,54,44,44,47,46,43,43,44,44,45,54,58,54,46,43,36,51,73,85,76,
					-- image=0 channel=0 column=27
					50,35,29,35,44,78,202,211,97,65,54,48,58,48,40,45,47,48,47,46,51,39,39,48,47,39,28,40,67,67,46,51,
					-- image=0 channel=0 column=28
					50,35,32,33,41,46,104,170,64,54,52,53,61,58,54,45,42,41,46,49,46,42,40,39,37,40,44,63,47,31,15,51,
					-- image=0 channel=0 column=29
					68,42,31,38,37,43,42,71,49,31,27,38,49,56,58,53,56,60,57,53,50,45,39,33,42,62,79,73,56,38,13,40,
					-- image=0 channel=0 column=30
					61,49,35,43,39,42,44,40,42,27,23,30,27,29,36,47,56,62,66,75,69,49,43,43,60,85,109,93,60,26,29,20,
					-- image=0 channel=0 column=31
					54,56,45,43,40,40,40,38,36,26,22,29,25,29,19,18,32,47,61,74,66,53,52,45,67,89,105,89,48,24,34,21,
					-- image=0 channel=1 column=0
					112,111,116,118,112,109,115,113,111,113,116,111,111,117,117,119,117,113,111,112,109,107,107,106,107,101,98,97,97,95,91,85,
					-- image=0 channel=1 column=1
					112,110,114,116,112,113,117,114,116,110,111,110,113,119,117,115,115,111,112,115,110,104,102,100,105,102,102,97,98,95,91,88,
					-- image=0 channel=1 column=2
					110,109,111,111,106,115,117,117,115,115,114,109,111,115,114,113,116,114,111,96,90,78,77,85,86,96,103,99,99,98,95,89,
					-- image=0 channel=1 column=3
					107,110,109,112,110,117,120,119,115,117,123,146,130,111,115,114,112,111,80,87,90,90,75,63,70,62,85,98,102,101,99,94,
					-- image=0 channel=1 column=4
					107,114,115,114,114,113,120,116,113,116,128,214,156,114,111,108,80,53,69,103,110,114,102,94,72,78,73,83,96,101,94,93,
					-- image=0 channel=1 column=5
					109,104,100,112,115,113,116,115,111,116,118,138,122,102,75,50,58,56,83,113,121,122,116,96,100,91,58,58,84,105,98,95,
					-- image=0 channel=1 column=6
					100,95,37,74,117,118,115,118,117,116,120,107,98,108,87,67,83,75,84,130,142,118,99,102,111,83,71,47,61,98,99,93,
					-- image=0 channel=1 column=7
					115,96,43,64,111,117,114,116,119,113,109,94,110,131,106,87,95,88,77,118,153,124,93,98,93,81,60,53,47,83,103,97,
					-- image=0 channel=1 column=8
					161,105,58,121,124,113,117,122,121,135,89,105,141,143,111,80,81,85,78,71,125,135,103,79,77,82,73,57,35,59,106,103,
					-- image=0 channel=1 column=9
					176,139,100,154,149,116,116,118,180,214,180,131,153,131,110,85,84,74,57,68,125,133,124,98,81,85,85,76,49,30,75,103,
					-- image=0 channel=1 column=10
					183,116,151,169,156,112,118,89,197,224,191,135,159,137,108,111,76,80,44,85,165,147,147,100,83,102,88,79,59,36,46,81,
					-- image=0 channel=1 column=11
					191,108,144,175,167,120,123,93,95,182,171,142,161,171,119,107,98,84,38,121,201,152,139,89,80,93,104,87,75,53,55,56,
					-- image=0 channel=1 column=12
					194,96,134,180,156,123,123,109,68,154,144,114,166,202,149,113,114,114,50,147,187,149,118,88,83,84,95,87,87,73,74,55,
					-- image=0 channel=1 column=13
					192,95,154,188,110,106,124,116,72,132,125,149,174,216,172,131,117,114,71,152,181,144,110,85,80,73,80,100,101,88,89,73,
					-- image=0 channel=1 column=14
					196,107,167,186,109,89,119,122,74,106,123,185,180,165,140,143,136,100,71,152,175,133,128,109,86,93,96,110,116,96,85,95,
					-- image=0 channel=1 column=15
					197,129,167,178,137,83,120,125,94,120,131,221,236,138,130,121,112,104,88,134,159,147,108,85,72,88,104,109,110,86,96,104,
					-- image=0 channel=1 column=16
					203,146,164,182,170,86,125,126,121,80,143,163,152,132,106,106,101,101,90,143,138,141,130,105,76,79,93,91,83,88,108,104,
					-- image=0 channel=1 column=17
					215,166,167,184,182,102,96,149,137,93,116,105,102,105,91,110,91,103,128,96,56,120,126,69,56,56,70,93,94,112,116,110,
					-- image=0 channel=1 column=18
					211,184,175,181,184,131,88,139,148,128,90,64,121,111,117,143,92,96,139,117,109,99,68,59,41,62,69,105,119,120,115,111,
					-- image=0 channel=1 column=19
					192,189,176,179,182,149,90,121,124,136,134,59,118,97,134,176,118,75,119,124,129,86,49,51,49,90,91,118,121,113,111,107,
					-- image=0 channel=1 column=20
					156,193,178,173,181,157,103,135,175,105,90,77,90,118,173,182,148,100,78,77,61,52,46,33,57,71,100,125,123,109,113,105,
					-- image=0 channel=1 column=21
					120,200,178,169,179,144,87,153,247,222,140,141,156,182,196,192,172,133,109,62,49,54,70,81,85,84,99,101,104,96,92,90,
					-- image=0 channel=1 column=22
					105,197,183,172,177,146,112,211,252,253,224,143,132,141,133,133,124,93,87,82,84,84,85,93,94,91,96,104,108,97,97,95,
					-- image=0 channel=1 column=23
					89,137,168,174,182,170,166,245,251,231,136,88,80,76,75,72,79,81,81,82,86,90,89,87,89,93,94,96,96,94,95,90,
					-- image=0 channel=1 column=24
					91,87,102,153,179,136,189,250,245,159,94,84,84,85,83,84,86,84,82,79,83,86,85,89,92,103,103,101,102,99,94,103,
					-- image=0 channel=1 column=25
					111,94,85,106,148,136,213,253,198,93,91,88,90,90,83,82,82,81,80,83,86,89,92,95,108,110,109,108,108,105,123,137,
					-- image=0 channel=1 column=26
					114,99,86,83,95,145,229,245,143,92,87,94,92,82,82,83,84,83,86,88,90,97,106,110,105,97,95,91,108,130,138,125,
					-- image=0 channel=1 column=27
					110,98,89,86,83,106,219,228,126,104,94,87,97,87,80,82,84,87,89,89,97,92,93,102,101,93,85,101,129,126,98,96,
					-- image=0 channel=1 column=28
					108,97,92,88,88,84,133,197,100,97,94,95,103,100,96,83,79,80,88,92,92,95,93,92,90,93,102,125,110,90,60,93,
					-- image=0 channel=1 column=29
					124,100,88,91,87,89,79,107,89,77,71,82,93,100,102,92,94,99,99,97,95,94,88,83,91,112,132,131,116,97,64,85,
					-- image=0 channel=1 column=30
					116,102,85,91,90,92,88,81,85,72,67,74,71,73,80,86,95,101,109,119,113,95,88,88,105,130,156,145,115,82,82,64,
					-- image=0 channel=1 column=31
					107,105,89,86,89,92,87,81,79,69,66,73,69,73,63,58,70,87,104,119,111,96,95,87,109,131,146,135,99,77,84,67,
					-- image=0 channel=2 column=0
					49,47,51,53,46,41,47,45,44,41,41,52,49,41,45,44,40,38,39,43,44,45,45,43,44,39,43,41,38,36,36,33,
					-- image=0 channel=2 column=1
					51,40,45,56,49,43,47,45,46,38,41,54,52,41,40,33,30,33,41,50,53,55,52,48,50,46,45,38,34,31,32,34,
					-- image=0 channel=2 column=2
					47,33,36,48,42,44,45,45,43,43,48,57,51,38,37,35,39,47,54,49,52,50,47,50,48,55,51,39,35,34,34,33,
					-- image=0 channel=2 column=3
					40,32,31,44,43,46,48,48,44,45,57,95,75,41,47,54,58,67,47,65,76,84,66,50,52,39,45,46,43,39,39,36,
					-- image=0 channel=2 column=4
					41,48,49,47,43,40,47,44,41,42,59,164,107,56,60,71,50,31,56,98,111,118,105,93,67,70,47,45,48,46,36,36,
					-- image=0 channel=2 column=5
					54,64,57,53,44,39,41,41,37,39,42,85,78,58,43,31,43,45,76,110,120,122,116,96,97,86,47,37,49,58,44,40,
					-- image=0 channel=2 column=6
					57,80,17,28,48,43,40,43,42,37,39,52,59,75,70,57,72,64,74,121,132,108,90,94,103,77,69,39,36,58,48,39,
					-- image=0 channel=2 column=7
					90,92,38,41,56,42,36,39,49,51,51,49,77,107,93,79,88,82,69,107,140,112,81,88,84,74,58,49,32,50,51,39,
					-- image=0 channel=2 column=8
					144,105,59,113,82,43,41,50,66,95,59,78,121,128,101,74,77,82,73,61,112,123,93,70,69,76,67,53,27,35,59,45,
					-- image=0 channel=2 column=9
					163,143,105,149,112,51,47,60,146,198,166,119,145,125,107,79,79,71,53,58,112,122,114,89,74,78,78,71,43,15,44,57,
					-- image=0 channel=2 column=10
					175,122,158,168,122,50,51,47,179,226,188,131,155,132,104,104,69,77,40,77,154,137,138,92,77,96,79,73,59,33,31,46,
					-- image=0 channel=2 column=11
					189,116,153,178,136,59,55,44,80,188,164,133,151,159,106,95,89,79,34,113,192,142,130,82,75,88,94,81,78,55,48,26,
					-- image=0 channel=2 column=12
					194,105,144,185,133,68,53,47,44,152,126,94,148,183,129,98,105,109,47,140,178,140,111,83,79,80,85,81,89,73,64,24,
					-- image=0 channel=2 column=13
					193,103,163,192,98,66,58,50,39,120,103,127,155,200,157,117,107,109,68,147,174,136,104,80,76,70,72,94,99,81,69,34,
					-- image=0 channel=2 column=14
					196,112,172,188,109,67,62,55,34,88,103,169,169,159,140,134,125,95,70,149,170,127,122,105,83,91,90,104,111,80,53,47,
					-- image=0 channel=2 column=15
					197,136,174,181,142,77,88,77,52,93,116,211,230,137,130,112,101,95,75,118,146,138,101,80,68,87,99,99,93,54,48,48,
					-- image=0 channel=2 column=16
					204,160,178,188,172,90,126,113,82,37,133,155,141,117,88,90,92,87,58,104,109,126,118,97,72,77,94,82,55,45,55,46,
					-- image=0 channel=2 column=17
					215,180,184,194,186,105,102,145,111,61,105,95,89,89,73,98,88,95,102,64,32,105,115,61,51,53,65,78,64,68,64,54,
					-- image=0 channel=2 column=18
					205,192,189,193,188,133,96,143,141,111,80,55,108,96,100,133,93,93,120,93,92,86,58,52,39,60,40,59,62,54,45,46,
					-- image=0 channel=2 column=19
					180,187,181,185,184,152,99,132,130,135,126,51,108,86,123,168,118,73,103,105,118,78,44,50,52,93,60,68,64,52,50,46,
					-- image=0 channel=2 column=20
					146,187,175,172,180,160,111,146,185,111,87,73,86,116,173,177,148,101,66,63,57,54,51,41,69,83,75,82,76,61,69,63,
					-- image=0 channel=2 column=21
					124,200,176,168,179,147,91,159,250,225,144,147,164,192,208,197,181,143,109,62,58,68,87,102,110,111,122,119,120,112,112,115,
					-- image=0 channel=2 column=22
					133,213,192,177,182,150,113,209,247,252,232,157,149,162,156,152,148,119,104,101,111,110,115,125,131,130,135,141,142,132,137,132,
					-- image=0 channel=2 column=23
					135,168,188,188,192,174,164,237,241,228,153,111,105,105,107,101,115,120,113,116,125,125,126,128,132,139,137,137,135,134,139,133,
					-- image=0 channel=2 column=24
					141,130,134,176,191,137,181,242,245,175,127,118,119,121,120,116,117,117,115,113,120,125,125,130,134,145,142,142,146,144,140,149,
					-- image=0 channel=2 column=25
					162,140,124,136,167,143,209,249,205,118,128,125,127,127,121,115,113,112,113,117,123,131,134,138,150,152,147,149,154,152,167,182,
					-- image=0 channel=2 column=26
					165,147,130,122,126,164,234,247,153,114,123,131,129,119,119,119,119,119,123,127,131,141,150,154,150,141,140,138,158,178,182,169,
					-- image=0 channel=2 column=27
					162,149,138,133,126,138,233,234,140,126,129,124,133,123,116,119,122,126,130,132,140,138,139,148,147,139,133,153,182,176,142,139,
					-- image=0 channel=2 column=28
					161,147,143,141,138,125,159,211,119,121,128,130,139,135,131,120,118,120,130,135,136,139,138,136,135,138,151,178,164,140,103,136,
					-- image=0 channel=2 column=29
					177,148,137,146,139,132,113,133,114,105,105,117,128,135,137,128,131,137,139,138,137,136,131,125,133,154,179,181,168,146,108,127,
					-- image=0 channel=2 column=30
					168,148,132,143,139,134,125,112,115,104,102,109,106,108,115,120,128,135,144,156,152,134,127,127,144,170,197,190,164,130,126,107,
					-- image=0 channel=2 column=31
					160,149,132,134,134,132,123,115,114,105,101,108,104,108,98,89,100,118,137,152,145,131,130,123,145,167,182,175,145,124,129,110,

					others=>0 );
END inmem_package;
