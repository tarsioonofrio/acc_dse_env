library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -23047, -94993, -94140, 53301, 113833, -542, 21988, 596, -23155, 2651,

    -- weights
    -- filter=0 channel=0
    6, -16, 240, 90, -217, -159, -22, 26, -79, -7, -24, -245, -239, 111, 0, -29, 35, 109, 111, -53, 80, 2, 2, -293, 39, 64, -69, -73, -39, 33, -188, -112, -31, -82, 84, -11, -19, -93, 31, -104, 8, 58, -5, -37, -164, -110, 152, -1, 24, -175, -226, 174, -134, 51, -26, 45, 36, -34, -49, 31, -31, -109, 9, -35, -20, 50, -43, 56, -201, 16, 23, -20, 18, 51, 84, -46, -92, 135, -28, -84, 204, 31, 45, 42, -1, 18, -67, 122, 63, 16, 65, -109, -58, 151, -7, 83, 115, -15, 2, -4, -6, -15, -112, 44, -3, -47, -25, -7, -49, -34, -12, -87, 65, -18, 31, 31, -43, -32, -17, 8, -129, -40, -6, -85, 62, -116, -193, 15, -11, 57, 194, 52, 275, -20, -26, -41, 84, -41, -145, -23, 32, 46, -23, 47, 39, 22, 49, 120, -85, 22, 27, -152, -124, -54, -32, -104, 2, -9, 72, 140, 59, 166, 82, 15, -5, -47, -16, -48, -14, -74, -101, 36, 3, -83, 2, -458, -20, -175, -51, 64, -152, -95, 9, -105, -18, -53, 58, 44, -145, -98, -203, -20, 2, -116, 11, 15, -50, -69, -4, 104, -58, -64, -342, -85, -59, -306, 22, 15, 68, 18, 93, 17, -38, 23, -81, 12, 4, -52, 56, 5, -187, -166, 13, -101, 82, -67, -16, -22, 79, 2, -76, -148, 66, 5, -36, 35, 32, -57, -3, 123, -30, 105, 18, 45, 17, -119, 3, 130, 53, 17, -75, -295, 87, 77, -101, 80, -7, -140, -174, -67, 193, 36, -24, 79, 35, 58, -318, 10, -62, -201, -4, -59, 80, -87, 143, 35, 159, 16, -156, 156, 67, -40, -159, 76, -193, -13, -86, -23, 77, 20, -50, -3, 75, -1, -245, -45, -76, 87, -2, 142, 101, -133, -12, 127, 31, -112, -60, -33, -12, -37, -14, -142, 147, -18, -4, -108, 71, 77, 11, -28, -2, -128, 79, 21, 69, -67, 12, -73, 228, -68, -157, -38, 41, -51, 3, 138, 36, -119, 5, -6, -65, 4, -29, -448, -89, -209, -94, -103, -236, 7, -10, 76, -55, -61, -5, -1, -107, 49, -182, -127, 42, -156, -109, 111, -37, -137, -82, -237, -6, -13, 146, 14, -57, -38, -6, -202, 57, -128, 113, -113, -3, -15, -185, 55, 8, 25, -100, -112, 62, -110, 18, -11, 38, -5, -171, -33, 33, -13, 7, -48, 77, -1, 201, -86, 20, 10, -64, -57, -148, 45, 41, -142, 14, -6, -61, -232, 253, 102, -5, -6, 40, 3, 5, -234, 73, 20, -112, 53, -91, -109, 67, 112, -122, -5, 71, -155, 48, -75, 9, 151, -88, 126, -79, -128, 5, -107, -122, 29, -7, 36, 43, -92, 147, -72, 20, 27, 56, -61, -99, -21, -56, -44, -21, 21, -52, 43, 172, -88, 9, 6, -31, 49, -92, 27, -23, -6, -212, 11, -171, 50, 241, 12, -67, 7, 51, -12, -132, 42, 30, -43, 71, -48, -39, 20, 34, -242, -51, 50, -87, 6, 45, 43, -32, -35, -90, 74, 118, -225, -58, -151, -33, -31, -12, -41, 12, 61, 151, -58, 18, 144, 48, -132, -59, -13, 92, 54, 9, -14, -74, 39, 121, -31, -39, -10, -30, -84, 3, -17, -189, -63, -32, -40, 104, 58, 73, -51, -33, -17, -156, 16, 167, -268, 13, -108, -66, 87, -100, -158, -163, 74, -57, -126, -218, -107, 94, -21, 6, -10, 31, -158, 178, -97, 192, 13, 63, 17,
    -- filter=0 channel=1
    -10, -60, -195, -117, 130, 19, -21, 16, -110, -53, -16, 94, -1, 136, -12, -67, 37, -90, 70, -6, 90, -17, -8, -112, 24, 35, -115, 15, -34, 87, 182, 120, -32, -5, -53, -3, 94, 0, -69, -56, -98, -39, 46, -30, -12, -102, 34, -282, -18, -5, 28, -112, -40, -17, 21, -125, -12, 11, -116, -132, -130, 123, 44, -108, -18, 82, 132, -52, -247, 60, 17, 93, -18, -56, -216, -206, -126, 32, 13, 56, -15, -93, -2, -196, 130, -26, -80, -84, -127, 22, -42, 4, -122, 53, -10, -10, -177, 96, 10, -10, -39, -33, -100, -153, -43, -80, -87, 52, 87, 116, -12, -54, 16, 40, 91, -171, -21, -122, -25, 8, -18, 114, 56, 24, 114, 63, -6, -12, 24, 65, 334, 42, 125, 81, -27, 87, -75, 8, -84, 62, -64, -65, 19, -7, 10, 104, -30, 14, 28, -12, -3, -87, 21, 70, -152, 139, -221, 166, 35, 53, 107, -160, -110, -17, -60, 27, 141, 0, -23, -26, 7, -83, -54, 56, -1, -193, -182, -21, 32, -94, -10, -8, 25, 49, -73, 131, -5, -302, 34, -65, -35, -5, 0, 0, 115, 49, -137, 1, -35, 64, -129, 48, -176, -32, -57, 146, -19, 40, -57, -184, -27, -21, 95, -20, -24, 60, 55, -6, -9, 58, -48, -137, -303, -46, -152, 35, -226, -10, -175, 79, 181, 111, -37, -82, 26, 8, -237, -48, -80, -48, -8, -76, 19, -55, 92, 80, -8, 34, 86, -22, -3, -347, 45, -156, -47, -36, -26, -165, 26, 99, -261, 54, -17, 58, -16, 17, 138, -113, -162, 76, 12, -44, 202, -292, 88, 101, -37, 9, 96, -94, -33, -27, -74, 7, -282, -196, -36, -415, -211, -10, -33, 23, -145, -64, -65, 10, 67, -172, 54, 6, -196, -46, -136, 30, 32, -14, -44, -25, -5, 151, -1, 104, 66, 16, 224, -8, 101, 16, -99, 0, -20, -109, -362, 52, -213, 64, -8, 39, -12, 97, -158, 0, -12, 9, -5, 37, 49, -109, -41, -190, -26, -23, -1, 105, 107, 13, -110, 46, -106, -120, 13, -297, -126, 129, -28, 11, -39, 27, 156, 192, -86, -20, -188, -60, -36, 49, -147, -46, -371, -154, 22, -39, -88, 117, 3, -642, -15, 72, 18, 25, -19, -219, -223, -87, -19, -264, -81, 29, -25, 53, -13, 109, -91, 152, -270, -30, -202, 105, -20, 5, -98, 0, 13, -228, 82, -18, -145, 142, -91, -65, -5, 184, -57, -185, 100, -171, -130, -192, 80, -13, -250, 42, -199, -19, -125, 90, -234, -1, -97, -39, 222, -46, 159, 64, -171, 49, 86, 0, 10, 10, 146, -3, -191, -116, 198, 12, -36, -30, 8, -73, -56, 25, -485, 43, 22, -37, 106, 63, -457, 59, -60, 147, -6, -86, 113, 49, -103, -204, 183, -12, -30, -120, 111, 73, -4, 147, 43, 28, -104, 21, -10, 0, 65, -14, -150, 0, 1, -99, 0, -26, -196, 80, -64, -115, 7, 104, 134, -118, 149, 6, -83, 81, 0, -119, 120, -20, -31, 30, 74, -94, -130, 60, -20, -230, -219, -131, 109, 6, 4, -19, 101, 219, -519, 8, 78, 83, -25, 56, 61, -171, -35, -130, 119, 16, -12, 7, 19, -23, -33, 47, -97, 51, -139, -79, -81, 60, 155, 3, 60, 0, -310, -19, -158, -137, -200, -104, -19, -50, -213, 60, 2, 69, 80, 65, -66, 31, 7, -306, 105, -25, -107, 21, -158, 3, -152, -37,
    -- filter=0 channel=2
    24, 76, -344, -29, -85, 24, -6, -34, 18, -47, -14, 51, 4, -206, 27, 65, -26, -70, -48, 52, -54, 3, -65, 18, -47, -50, 7, -11, 74, 31, -123, -33, 140, -21, -79, 20, -142, -12, 20, -93, -35, 5, -25, -31, -5, -15, -40, 261, -14, 30, 2, -41, 30, -73, -24, -18, -67, -56, -36, -68, -64, 16, -83, 32, 3, -135, -124, -11, -163, -41, 0, 29, -17, -36, -41, 84, 30, -105, -22, -91, -7, 49, 23, 84, -77, 14, 50, -32, 106, -60, 96, -24, 39, 92, -99, -25, 86, 5, -24, 12, -23, 14, -104, -80, 4, 34, 55, 8, -1, 20, -6, -67, -47, -96, -45, -7, -78, -31, 2, -111, -106, 49, -46, -117, -88, 107, -21, -71, -22, -34, -69, -68, -154, -123, 19, 120, -48, -46, -101, 4, -143, 15, -10, -5, -24, 13, 37, -87, 62, -20, -130, -135, -113, 17, -11, -41, 12, 138, -116, -32, 95, -4, 39, -6, -14, -71, 52, -83, 50, -20, 98, -97, 7, 75, -45, 67, 16, -41, 78, -68, -33, -34, -34, 27, -2, 5, 44, -105, -7, 39, 22, -107, 0, 69, -49, 109, -346, -13, -20, -175, 105, -98, -170, 79, 0, -53, 18, -72, 189, 13, -26, 11, -91, 2, -51, -177, -16, -8, 49, -20, 20, 60, 1, 70, 68, 6, -24, -23, 2, -11, 0, -20, -142, 34, -11, -32, -5, -27, 77, -61, -32, -3, -20, -11, 12, -63, -20, 104, 43, 27, -19, -142, -56, 7, -50, 25, -24, -187, -38, 102, -144, -77, -1, -64, 42, -101, -122, -32, 15, -5, 5, 45, -132, -56, -10, -86, -28, -3, -22, 47, -16, 68, 67, -10, 26, -20, -78, -46, 77, 83, -8, -27, -1, -49, 48, -57, -77, 40, 30, 74, 41, 127, -15, -107, -54, 60, 4, 0, -53, 59, -14, -96, -164, 46, -131, 38, -152, -65, -132, -77, -21, 0, 198, 45, -34, -156, 13, 23, 58, -39, -147, -58, 50, -59, 16, -37, -34, 58, 7, 5, 27, 25, -187, -153, -38, 65, 13, 1, 15, -52, 114, 64, 80, 70, 52, 11, -36, -24, 104, -183, 94, -22, 53, -37, 59, 25, -32, 0, 0, -36, -71, -25, -27, -84, 4, -155, -99, 28, 91, -107, -28, -7, 54, -73, 10, -33, -167, 53, -426, -147, 17, -33, 63, -70, -3, 14, 11, -79, 6, 47, 129, 31, 84, -17, -177, -5, -88, -171, 14, -13, -55, -87, 111, 16, -196, 11, 61, 78, -31, 18, 161, -93, -350, 88, 167, 10, 22, 8, 7, -79, 20, -279, -123, 15, 46, -121, -6, 53, 17, 13, -147, 76, 61, -54, -132, 26, 61, -6, 10, -133, 57, -51, 39, -111, -26, 95, 2, -78, 174, 0, 22, 133, -24, 20, -57, 13, -3, 30, -129, -7, -98, -12, -50, 26, -1, -141, 21, -50, -125, -80, 14, -51, -32, 24, 26, -85, -262, -7, 22, -126, 0, 5, 74, -47, 83, -83, -52, -13, 3, -82, -44, 67, 19, -3, -87, 63, 24, -163, -88, -28, 7, -62, -20, 34, 211, 76, 161, -103, 9, 53, -4, -69, 22, 28, 12, -199, 16, -87, -86, -21, 30, 14, -53, 6, -86, -131, -46, -19, 27, 0, 36, -31, -79, -89, 165, 26, -84, 5, -36, 90, -244, -31, 81, 1, 70, 73, 42, -68, 60, -307, -67, -133, -71, -113, -36, -36, -3, 4, -18, 65, 21, -227, 2, 13, 63, -125,
    -- filter=0 channel=3
    -10, -16, -193, -28, -260, -56, -1, -27, -22, -59, -20, -79, 47, -98, 14, -6, -27, 55, 0, -75, -57, -8, -32, -20, -65, 83, 84, 7, -29, -6, -117, -75, 70, -12, -89, -14, 11, -47, -35, -25, -67, 64, 36, -80, 15, 30, -6, -145, -22, 14, -21, 86, -24, -77, 4, -13, 88, -39, -53, -10, -33, -22, -20, 59, -23, -50, -90, -86, -144, -61, 0, -20, 7, 1, 8, 83, -32, -25, -5, -5, -13, -15, -18, -37, -61, -26, -23, 43, -122, 32, 22, 20, 64, -9, -138, -11, 30, -81, -38, -19, -26, -67, 90, 5, -161, 33, 14, -23, 15, 45, -79, 4, 57, 0, -79, 38, 50, -28, -4, 53, -35, -59, 102, -81, -72, -49, 29, 13, 8, -16, -212, -70, -85, -46, -18, -12, 23, -108, -117, 0, 1, 46, -11, 66, -28, -34, 21, 34, 49, -31, -50, -44, -51, 27, -2, 10, 37, -40, -111, -9, -126, -50, 20, -23, -71, -42, -145, -47, -47, 13, 47, -47, 14, 0, 16, -154, -39, -1, 82, -33, 13, -121, -27, 28, -28, -36, -109, 20, -116, 25, 6, 62, 4, -34, 45, -6, 148, 75, -12, -73, -25, 24, 64, 69, -9, -144, 14, -14, -109, 6, 82, 21, 22, 14, -79, -31, -70, 36, -40, -70, 17, 43, -44, 116, 80, -30, -22, 1, -86, -15, -334, -73, 29, -33, 37, -118, -14, 52, -51, -47, -70, -83, -60, 16, -198, -40, -10, 51, -98, -123, -134, 49, -21, 37, 20, -60, 14, -37, 57, -102, -108, 4, 3, 43, 8, -104, 122, 88, 32, 15, 0, -48, -128, -34, -48, 58, -81, -13, -87, -2, -144, -11, -18, -63, 66, 0, 0, -5, -23, -105, -118, -20, 40, 63, -10, 16, 6, -22, 24, -113, 7, 38, 61, -122, -175, 1, 46, -35, -31, -93, -22, 59, -237, -83, -88, -82, 47, 34, 17, 54, 15, 0, -24, -69, -78, -39, 1, 26, 0, -54, 26, 30, 0, 11, 21, -49, -102, -18, -28, 37, -18, 20, -88, 114, -73, 2, -33, -42, 83, -55, -94, -101, -47, -38, -27, -18, 55, 5, -45, -2, 0, 46, -4, -161, -43, 51, 18, -103, 91, 31, -18, -10, -25, -85, 1, 112, -18, -45, -29, -153, -11, 5, -5, 37, 22, -55, 122, 16, 117, 40, 23, -83, 32, -34, 15, -9, -1, -107, -7, 2, 4, 93, -107, 19, -40, 20, 5, 24, 89, 5, 56, -117, -80, 52, -109, 10, 7, -9, 19, -12, 17, 58, -57, -35, -75, -38, 89, -77, 16, 61, -99, -76, 75, 2, 0, -42, -96, -4, -10, -39, -46, -26, 48, 41, -153, 0, 1, -89, 25, 81, -115, -106, -103, -6, 30, -5, -43, -48, 102, -19, 26, -120, 21, -54, 37, 13, -124, 59, -10, -12, -97, -10, 15, 11, -69, -67, 23, -15, 38, -18, -136, -56, -28, 0, -92, -2, -137, -15, -27, 70, 2, 0, -54, -2, -67, 36, -30, -4, 0, -12, -28, -84, -2, -31, -40, 66, 11, -21, 9, 93, 19, -16, -4, 71, 1, -18, -169, -59, -11, -23, -33, -73, 3, -54, 68, 64, -14, 49, -23, -17, -48, 83, -21, -3, -27, 27, -21, -34, 11, -18, 53, -60, 91, 66, -66, -25, -62, 6, -13, -42, -24, -40, 30, 54, 23, 34, -38, 35, 23, -48, -32, 33, -22, -122, -94, -118, -38, 5, -6, -27, -14, -227, -22, -9, -58, -16,
    -- filter=0 channel=4
    -12, -71, 5, 15, -41, -78, -2, -64, -94, 66, -26, 53, 57, 38, -9, -8, 85, 45, -105, -25, -44, 4, -26, 79, -108, -35, -119, -45, 83, 36, 55, -125, -268, -127, 58, -2, 41, 4, 0, 7, -28, -81, -34, -33, -94, 48, -71, -98, -38, 7, -108, -18, 63, 32, 17, 90, -95, -30, 130, -149, 100, -107, -25, -75, 18, 3, -350, -86, 64, -131, 7, -24, -13, 0, -68, 118, 25, -51, 21, -214, -35, -36, -142, -17, -45, -22, -76, -46, -132, 47, -124, -72, 43, 32, 51, -30, -243, 119, 52, 10, 66, -23, 29, 92, 27, 33, -92, -52, -116, -62, 25, -259, -42, -162, 34, 133, 26, -17, 18, 130, 85, -117, -47, 52, -18, -74, -20, -95, -1, -42, -46, -71, -9, -58, 5, -81, 50, -99, 43, -3, -5, -124, -4, -105, -77, -42, -34, 63, 20, -14, 44, 100, -69, -32, -66, -86, 88, 29, 77, -19, -116, 53, 72, -26, -70, 92, -121, 4, -37, -136, -122, 34, -4, -152, -52, -119, -9, -88, 40, 60, 0, 29, -18, -21, -117, -70, -8, -145, 89, 10, 74, 20, -1, 46, -16, -113, -84, -33, -6, -60, 49, 41, -147, -27, -27, -116, 6, -29, -11, 39, -84, 40, -43, -19, 161, 9, 81, -14, -124, -79, 3, 68, 163, -6, 30, -82, 41, -5, 25, 27, 112, 63, 100, 46, -64, 67, 42, 77, -80, -227, -64, 31, -76, -98, 7, 55, 2, 25, -130, 56, 30, 17, -33, -200, -34, 64, -3, -4, 8, -86, -213, -106, -15, -103, -30, -1, -36, 52, -91, 44, 18, -105, -209, 50, -193, -32, -43, 13, 171, -134, 14, -83, 67, -187, 32, -46, -35, -58, 0, -25, 59, 22, 22, -7, -103, 63, 4, 11, -60, -123, 75, 40, -108, -246, -26, 40, -42, 104, -80, 63, -6, -31, -60, -140, -53, -81, -131, -148, 53, 39, -13, -12, 62, -47, 14, -77, -21, -31, -67, 22, -31, 13, -118, -53, 13, -155, -27, 86, -110, 25, -29, 6, 174, -37, 6, 55, 62, -50, 80, -57, -71, 9, -55, 17, 58, 23, -46, 57, -49, 60, 56, -10, 2, -38, 83, 12, -14, 54, -30, 15, -59, 138, -18, 67, 5, -56, -4, -13, 76, -279, -121, -82, 100, 36, 22, -22, -2, -110, -210, -82, 1, -185, -178, -58, 58, 4, 8, 18, -7, -61, -18, -101, -43, 49, -44, 22, 124, 23, 100, -11, -120, -80, 13, 44, -144, 16, -16, -20, -7, 18, 105, -45, 56, 59, 1, -35, -54, 60, 26, -70, 38, 175, -96, -90, 29, -164, 39, 35, -18, -164, -16, -201, -2, -29, 77, -94, 66, 48, -6, 102, -83, -86, -76, -51, -26, -138, -118, -64, 189, -23, -91, -193, -15, -41, -60, 38, -143, 13, -3, -18, -74, -48, 13, 27, 11, -177, 14, 1, -201, -46, -100, -80, 24, 4, -44, -139, -166, 98, -77, -69, 35, -81, 24, -91, 16, -62, -25, -51, -77, 34, 4, 91, 1, -30, -117, -166, -27, -153, -111, -36, 42, 36, 11, 37, -39, -69, -96, -13, 1, 7, -205, 58, 156, -28, -33, 56, -9, -168, -64, 22, -98, -46, -18, 24, 154, -48, -43, 83, 7, -94, 43, 40, -414, 29, 112, -80, -42, -11, 16, 49, -64, 34, 88, -70, 20, -56, -63, 32, 0, 27, -151, -19, -32, -58, 37, 17, 2, 38, -161, -34, 24, -345, -25, -45, 42, -16,
    -- filter=0 channel=5
    -16, -70, -126, -78, -113, 57, 15, -64, -17, -79, -59, -44, 65, 10, -5, 104, -89, -52, -24, 8, -9, 4, -46, -57, -33, -10, 26, -32, -50, 19, 28, -103, -1, -17, -37, -1, -110, -63, -64, -24, 69, 75, 43, 1, 29, 82, -92, -34, -172, -4, -68, 45, -5, -31, -24, -81, -8, -33, 88, -98, 101, 4, -6, 73, -20, 51, -98, -98, -335, 69, 3, -98, -72, -45, -56, 52, 35, -29, -5, 3, -9, -30, -113, 39, 21, -6, -6, -76, -108, 14, 61, 13, -4, -16, -96, -71, 33, -112, -87, -8, 24, -98, -179, -31, -101, 26, 58, 95, 100, 113, -33, 47, -64, -63, -97, 9, 20, 31, -28, 4, 42, -36, -32, -80, -13, -56, 33, -24, -23, -109, -172, -68, -234, 28, -18, -2, -51, -12, 71, -40, -121, -63, 2, -6, -131, 27, -38, -14, 66, -10, 29, 35, 16, 45, -22, -14, -8, -55, 53, 5, -61, -96, -61, -18, 46, -95, -119, -62, -13, 80, 33, 67, -5, 53, 21, 46, -98, -29, -116, -35, 13, 73, 5, -1, -101, 18, -31, 186, -8, 11, 39, 55, 16, -1, -135, -45, 30, 64, 18, -134, -30, -101, 7, 24, 45, -114, -13, 29, -137, -1, 24, -21, 43, -4, 65, -27, -76, -35, 53, -57, 35, 114, 47, -15, 45, -66, 0, 0, -55, -87, -168, 6, -57, -39, 19, -53, 53, -5, -13, 104, -72, -58, -59, 23, -76, -15, -38, -87, -139, -158, -124, 88, -98, 74, -52, 25, -14, 97, -168, -128, -137, 103, -9, -112, -7, -81, -76, 124, 26, -52, 18, -10, 8, -49, -66, -28, 62, 5, 64, -22, -60, -63, 91, -72, 1, 4, -45, -15, -13, -133, -63, 3, 29, -117, 141, -3, -187, -37, 48, -60, 56, -30, -28, 54, -116, 8, -1, 0, -81, -7, 3, 40, -55, -65, -126, -533, -53, 40, 33, 57, -17, 59, -57, -99, -109, 18, 5, -41, 35, -112, 111, -12, -6, -28, -5, -41, -108, -21, -68, 2, 43, 9, -62, -29, -68, 19, 81, -15, 60, -99, -13, -22, -10, -113, -28, -26, 8, -50, -146, 4, -72, 37, 29, -10, -47, -4, 0, -27, 37, 5, -169, -121, -32, 2, -43, 99, -67, -3, -94, -98, -88, 14, 24, 62, 23, 56, -38, -31, -74, 51, 6, -32, 58, -85, -57, -4, 55, 34, 8, 13, -79, 7, -27, 53, -74, 25, 52, -28, -44, 44, 0, -131, -11, 55, -49, 87, -49, -7, 6, -24, 7, -38, 92, -15, -45, -131, 93, -20, 17, 17, -73, -47, 26, 48, -80, -32, -40, 26, -8, -59, -138, -81, 96, 33, -126, 101, -85, -52, -14, -58, -160, -95, -44, 91, 8, -63, -30, -111, -281, -18, 0, -18, -9, -45, -14, -31, 47, 19, 5, 19, 38, 0, 62, -29, 4, -141, -90, 8, -14, 41, -108, -116, 3, 1, -57, -14, 213, -17, -177, 6, 17, -85, -20, 27, -49, 45, 37, 11, -55, -10, -17, -31, -20, -23, 62, 67, -78, -87, 50, -15, -26, 0, -17, 118, -175, 0, -304, -48, -10, -24, -97, -86, -138, -11, 5, -102, -15, 12, -87, 18, -139, 65, -73, -10, -11, 25, -20, 9, 63, -78, 45, -63, 12, 94, -14, 8, -49, -25, 10, -80, -67, 14, -22, 58, 54, -46, -3, 70, -10, -5, 6, 30, -67, -145, -23, -162, 0, 39, -68, 76, -54, -11, 45, -133, -47, 9,
    -- filter=0 channel=6
    17, -69, 0, 84, -169, 0, 9, -308, 19, -110, 65, 29, 46, -149, 7, -75, -199, -38, 29, 53, -98, -2, -79, -166, 86, -10, 176, -27, -37, -47, 161, 42, -108, 84, -243, 1, 13, 13, -122, -241, -17, 14, -55, -52, 46, 10, -66, -134, -52, -152, 70, -97, -31, -46, 15, -193, 22, -98, 195, -17, -272, -232, 97, -126, 14, -34, 118, 249, 137, -142, -19, -135, -22, -57, -85, -15, -11, -65, -16, -25, -86, -96, 112, 29, -117, 0, -98, -156, 240, 57, -168, 4, 19, -124, 3, 47, -121, 27, -66, -8, -23, 85, 168, 104, 143, -105, -13, 52, -240, -111, -9, -320, -188, 1, 44, -113, 129, -7, 27, -84, -119, -254, -1, -56, 38, -63, -45, -46, 20, -17, -234, 49, -5, 24, 14, -12, -39, -5, -10, 59, -8, 105, -22, -13, 29, 2, -198, -96, -118, -20, -81, 116, 44, 76, 20, -14, 78, -6, -86, -227, 15, 53, -124, -11, 89, 57, 114, -20, 14, 150, 75, -45, -122, 17, 20, -274, -94, 63, -58, 37, 100, -87, 9, -75, -28, -23, -162, -157, -267, 17, 64, -158, 20, -46, -138, 31, -179, 17, 3, 104, -33, 66, 86, 32, -45, -69, 18, -74, -145, -7, 87, 76, -22, 24, -131, -26, -9, -78, 115, -16, 11, -4, 19, -53, -223, -3, -108, 3, 81, -109, 55, -155, -44, 162, -53, -109, -6, 104, 31, -175, 82, -10, -70, -89, 22, -12, 6, -132, -19, 41, -18, -125, -142, 49, 51, -102, 2, 1, -257, 131, 182, -9, -14, -125, -134, 47, -36, -55, -106, 99, 0, 0, -266, 161, -33, 75, -89, 26, -208, -38, -128, 117, -99, -46, 192, 54, 69, 212, -162, 104, -201, 22, -55, -62, 47, -183, 174, 144, 114, -79, -153, 10, -16, -533, -208, 22, -41, 20, 23, -262, 2, -40, -71, -39, -1, -43, -189, -42, 47, -129, -10, -101, -104, 55, -137, -19, -23, -46, -42, -65, -492, 62, -11, -155, 19, 29, 48, -9, 9, 2, -83, 6, -238, -107, 96, 45, 30, -5, 91, 57, -204, -53, -87, 27, -117, 23, 67, -218, 102, -176, -78, 91, 117, -65, 79, 16, -14, -39, -121, 42, 11, 63, 119, -64, -5, -125, -90, 55, 104, 54, -85, 15, 69, -100, -19, 91, -36, 77, 51, 46, -26, -112, -114, -72, -76, -22, 35, -42, 19, -133, -23, -27, -195, 41, -23, -17, -231, -11, -10, -144, -25, -62, 69, 48, 118, 32, -67, -23, -171, 10, 22, -184, -77, 14, -79, 15, -23, -313, 2, 51, -178, -70, 0, 28, 37, 19, -67, -95, -21, 48, 100, 44, 57, 65, -41, -30, 39, 19, 11, -29, -111, -78, 72, -14, 9, -114, -4, -36, -45, 40, 79, -118, 0, 10, -128, -15, -25, -4, -35, 15, -79, 16, -13, -148, 4, -114, 46, 17, -70, 74, 92, -89, -74, -22, 37, -47, -165, -91, -76, 7, 29, -45, 49, 36, -292, 142, -46, 62, -13, 104, 27, -314, -9, 59, 30, 23, 123, -76, -14, 50, 46, -32, -2, -6, -335, 55, -114, 77, 19, -197, -21, -208, -4, 15, -16, -193, -21, -12, -102, -21, -48, 59, 1, -7, 6, -12, 16, -7, -25, -40, 87, -73, -63, -150, -215, -18, -182, 9, 39, -33, 14, -102, -54, -85, -36, -107, 95, -79, -72, -86, -125, 26, 116, 101, -92, -42, 2, -184, -35, -61, 93, -129, -3, -79, 128, -8,
    -- filter=0 channel=7
    -20, 15, 35, -119, 39, 9, -2, 10, 41, -20, -128, -10, -7, -61, -8, -71, -33, 3, -99, 5, -85, 11, 14, 137, 61, -133, -56, 126, -17, -82, -539, 38, 80, 28, -38, -15, 18, 49, 4, 133, 24, 28, 50, 82, -42, -55, -94, 116, 0, 118, 60, -190, -85, 77, 2, 63, -70, -13, -57, -114, -19, -26, -147, 49, -19, -149, 1, 6, 203, 42, -22, -91, 8, -10, 8, -97, 63, -114, 4, -19, -11, -31, -56, 80, -8, -27, 73, 107, -188, -87, -6, 20, -16, -162, 15, -58, 129, -58, 32, 9, -35, 79, -103, -52, -103, -24, -13, -286, 77, -118, -128, 122, 7, 72, -147, 9, -111, -6, -8, -14, -120, -75, -94, 12, -61, -157, -23, 135, 5, -135, -71, 15, 68, 61, -11, -21, 18, 77, 13, -43, 61, -24, -22, -108, -85, -164, 66, -86, -42, 11, 85, 67, 2, -141, 15, -25, -1, -86, -71, -14, 29, -141, 28, 1, -148, -27, -42, 41, 23, 51, -21, -30, -63, -14, -87, 159, 73, 80, -181, 38, -83, 64, -5, 6, 46, -117, -75, -219, -140, -45, -1, 62, 11, -55, -81, -207, -74, -31, -34, -257, 7, 34, 140, 28, -51, 167, -8, -94, 6, 31, -80, 50, -112, -4, 115, 13, 106, 181, 28, -122, 80, -47, -96, -3, -466, 18, 19, 10, 6, -66, 50, 51, 14, -18, 58, 0, 61, -72, -94, 104, 33, 87, 58, -71, 53, 120, -8, -241, -224, -61, -29, 73, 43, -154, 32, 30, 2, 274, 148, -94, -154, -46, -21, -60, -181, 63, -37, -128, 16, -177, 22, -16, -137, 58, -120, -9, 85, 18, 145, -125, 114, -1, -13, -127, -192, -40, -217, -105, 51, -12, 91, -21, -90, -78, -58, 97, -174, -155, -94, -47, -85, 3, 0, -1, 55, -21, 13, -65, 124, 29, -17, 65, -44, -161, -195, -387, -16, -182, 17, 80, -26, 40, 33, -27, -259, 102, 22, -123, -141, 22, 146, 28, -4, -15, 24, -124, -98, -19, -200, -107, 7, -17, 69, -47, -20, -30, 6, -43, -179, 43, 35, -11, 125, -98, 113, 4, 26, -68, -142, 89, 28, -152, -21, 21, -17, 60, -53, 35, 141, -2, -71, -121, 29, 60, -7, 182, -49, -36, -101, -267, 3, -33, 68, -50, -23, 125, -67, -345, -186, -40, -14, 49, -95, 21, -130, 107, 53, -121, 17, -38, 91, 11, -57, 99, 21, 3, 56, -72, 133, 157, -87, -124, -64, -124, -151, 6, -145, 19, 79, 20, -14, -35, -263, -8, 59, 25, -66, 127, 111, -59, 120, 217, 63, -76, 18, -71, 132, 65, -12, -46, -101, -36, -15, -30, -64, -151, 94, 5, 13, -148, 48, -163, 73, -114, 0, 15, -109, 160, -15, 13, -70, -208, -19, -25, -157, -23, 41, -51, -117, 3, -30, 15, 11, 46, -66, -130, 29, 52, -22, 41, -198, -28, -1, 17, 33, -164, 105, 60, 11, -15, -44, -161, -9, -37, 12, -22, -14, 23, -265, -222, 149, -14, -29, 96, 56, 36, -185, 15, -10, -140, 131, -6, -1, -86, 19, -126, -182, 86, 10, 15, -60, -35, -100, 25, -80, 79, -19, -94, -61, 99, -103, -99, -27, 6, -8, 14, 83, 69, -1, -125, -89, 55, -255, 81, 63, -167, -31, 3, 90, -46, 32, 8, 151, -43, 42, -93, 7, 79, -18, -41, 105, -91, -143, -56, 82, -1, -32, 104, -199, -88, -73, -42, -24, -14, 10, 37,
    -- filter=0 channel=8
    3, 151, 245, -25, 289, -9, -34, 63, 97, -17, -105, 137, -113, -61, -7, -299, 21, -63, 9, 46, -54, -6, 32, -28, -101, -11, 4, -84, -191, -28, -14, 128, -8, 40, 123, 3, -41, 121, -193, 32, -96, -202, -75, 9, -154, -149, 87, -342, 43, -66, 8, -75, 221, 187, 3, 0, -40, 63, 52, 195, -56, -98, -112, -157, 8, -10, -15, -89, 95, 28, 9, -8, 73, -46, -65, -172, 38, -76, -10, 50, -144, 41, 27, -72, -56, 19, -15, 24, 25, -92, -141, -14, -135, -42, -347, 109, -51, -77, -38, 15, 0, 9, 58, -40, 65, -125, -104, 25, -18, -77, 143, -133, 57, 212, 11, -20, -91, -89, -26, -35, -222, -98, -4, -134, -83, -41, 34, -14, -15, 104, 51, -35, -192, -13, 4, -171, -81, -52, -29, -76, 123, -202, 18, -21, 29, -79, 17, -36, -40, -20, -26, -129, 55, -108, -36, -106, -118, -56, -151, -1, -59, -77, -141, 2, -10, 20, -72, 109, -15, -325, -113, 11, 117, -48, 155, 61, 80, -70, -77, 66, -55, 88, -12, -57, -33, -11, 79, 220, 79, -189, -101, -22, 23, 25, -120, 72, -284, -94, -4, 13, 25, -57, -20, -104, -65, -94, 1, -83, -54, -4, -197, -100, -46, -4, -32, 63, -14, -86, -276, -12, -285, -37, 43, -14, 4, 96, 175, 22, 117, 29, 14, -65, -108, -136, -39, 111, -148, -74, 32, -182, 18, -100, 62, 109, -59, -2, 17, -121, -153, -9, 94, 79, -10, -6, 75, -19, 6, -93, -167, 39, 396, 26, -4, 108, 7, -35, 31, -160, 87, -89, -19, 144, 80, 38, 26, -31, -76, -7, -146, 126, -36, 20, -79, 98, -268, 5, -36, -46, -75, -3, 64, -23, -72, 233, -7, -99, 93, -40, -40, -48, -65, 18, 221, 9, -29, 35, 8, 0, 10, -162, -19, -160, -24, 56, -49, 155, -8, 193, 89, -21, -7, 43, -397, 31, 189, -63, 9, -37, -127, -106, 147, -43, 64, -115, -3, 47, -25, 10, 65, -25, -54, 15, 18, 132, -17, -44, -66, -10, -78, -89, -38, -43, 2, 88, -72, -21, 32, 76, 94, 85, -98, 5, 24, 53, -190, -169, 218, -11, 11, 85, -22, 64, 0, -16, 12, -31, 12, -33, -97, 90, 25, 65, -14, 43, -16, -45, 30, 41, 269, -152, 0, 77, 50, -188, 73, -312, -272, -164, -9, -25, -169, 34, -51, -119, -43, 23, -40, 18, 33, 82, -109, -88, -302, -169, 47, -95, -286, -177, -19, 2, -131, 40, 187, -287, -136, 20, 139, -28, -93, 113, -61, -299, -92, -98, 35, 153, -196, -157, -27, 34, 39, 38, 31, -26, 4, 225, -164, 5, -14, -69, -193, 261, -243, -66, 6, 63, 21, -82, -10, -42, -47, 14, -13, 60, 81, -195, 14, -134, -225, 14, 16, -17, 4, -169, -71, -2, -106, -155, 143, -143, 6, 140, -42, 3, 107, 170, -212, -112, 199, 115, 37, 69, -154, -115, 152, -626, -165, 38, 159, 116, 17, -171, 13, 70, 122, -1, -30, 237, -81, 349, -171, -102, 20, -91, -69, -187, 120, -197, -25, 25, -77, -238, 49, -47, -119, -123, -8, 113, 19, -158, 11, -24, -225, 5, -186, -26, -67, -34, 40, -63, -62, 33, 192, -110, -260, 93, 148, 6, -108, -30, 170, 77, -150, 137, -8, 81, -84, -68, -120, -247, 5, 114, 45, 151, -56, 131, 7, -39, 157, 20, -28, 171, -91, 226, -94, 47,
    -- filter=0 channel=9
    -10, -130, 49, -76, 112, 7, -18, 113, 107, 78, -96, -152, -8, -55, 4, -34, -47, -65, -29, -16, 0, 8, 17, -43, 55, 64, -24, -68, -118, -24, -100, 134, -11, -19, 79, -5, -8, -24, 116, 43, 123, -68, -51, 76, 60, 73, 16, -32, 100, -65, 40, -36, -121, -134, -24, 49, -172, 101, -59, -288, 35, 77, 65, 15, -12, -8, 5, -67, -177, 6, -21, 43, 44, 51, -23, -76, -60, 15, -7, 166, -100, 54, -11, -186, 32, 22, -14, -197, -9, -88, 15, 44, -187, -111, 0, -102, -76, -20, 54, -6, -39, 32, -24, -149, 41, 4, 57, 69, -106, 14, -86, -61, 35, -18, 47, -111, -90, 70, 15, -59, 55, 222, -2, -26, -11, 120, 134, 3, -2, -53, -116, -56, -51, -82, -18, -33, -42, 82, -117, -4, 71, -71, -1, -35, 41, 109, -18, -53, -68, -7, -91, -250, 163, -6, 128, 79, -173, -185, -206, -19, -72, -86, 20, 0, 73, -18, 65, -34, -16, -66, -1, 19, 45, -59, 14, 47, 29, 54, -85, -85, 76, -37, -15, 80, 59, 74, -40, -70, 143, -143, -199, 5, -23, -70, -70, -126, -101, -44, -13, 35, 63, 21, -41, -214, 74, 166, -10, 148, -72, -121, -41, -185, 90, -15, 8, -164, -137, -23, -91, 106, -81, -220, -113, -153, -7, -86, 38, 23, -14, -53, 71, -77, -5, -184, -114, -36, -10, -32, 58, -444, 48, -46, 68, -3, 9, -82, 11, -96, 79, 125, 97, -190, 8, -88, 0, -72, -18, 99, -26, -115, 31, -58, -14, -104, 117, -25, -25, -123, -104, -146, -28, -58, -27, 1, 36, -196, -100, -22, 20, -235, 50, 20, 34, 167, -119, 158, 23, 82, -128, -64, 40, 6, -52, -135, 66, -152, -66, -40, -226, 62, -35, -54, -97, 61, 175, -153, -40, 15, 51, 17, 6, 63, 96, 149, 123, 98, 65, 34, -7, -99, -17, 39, -189, -61, 29, 31, 21, -68, -60, 91, -57, -3, -82, 52, -5, -19, -14, 60, 82, -47, 38, -25, 47, 138, 92, -150, -124, 88, -95, 230, -295, 62, -56, -172, -56, 23, -90, -127, -47, -117, -155, -72, -234, -17, 39, -3, 78, -144, 13, -132, 46, -67, 81, -29, 3, 263, 55, 0, -104, 122, 51, 27, -97, 15, 22, -92, -229, -34, -270, 126, -10, -28, -28, 43, 43, 38, -81, 10, 7, 41, 28, -202, -81, -176, 87, -9, 28, 11, -141, -147, 82, 229, -76, -81, 20, -110, -22, -134, -50, -24, -89, -23, 90, 102, -104, 0, -282, -20, -2, -73, 10, -257, -55, -59, -66, 98, 92, -17, -12, -135, -20, -268, -129, -112, 53, -64, 10, 29, -14, 130, 19, 52, -297, 57, 17, -102, -2, 32, -108, -21, -22, -85, 16, 55, -23, -129, 58, -2, 115, 11, 53, 16, -97, -167, 33, 214, 62, -8, -10, -137, 14, 102, -73, 4, -38, -61, 96, -55, 92, 17, -190, 30, -74, 80, 8, -158, -65, -32, 69, -21, -110, -26, 1, -204, -112, -233, -58, -130, 9, -174, -63, -4, 15, -75, -107, 11, -170, 67, 9, -173, 137, 133, 100, 6, -122, 35, 16, -10, 65, -67, 62, -135, 121, -24, 8, 8, -119, -114, -67, 159, -52, -11, -98, -229, -205, -30, 47, -17, -119, 8, -119, 42, -212, 49, -153, 13, 0, -57, -22, -125, 23, -14, 131, 41, 49, 121, -28, -88, -95, 68, -224, 75, -21, -14, -91, -5,

    others => 0);
end iwght_package;
