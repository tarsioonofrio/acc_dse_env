library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    80, 312, 318, 
    543, 209, 307, 
    0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=2
    106, 16, 0, 
    280, 0, 0, 
    0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 
    563, 168, 0, 
    100, 0, 0, 
    
    -- channel=4
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=6
    218, 181, 200, 
    84, 0, 0, 
    0, 268, 604, 
    
    -- channel=7
    114, 0, 0, 
    98, 0, 0, 
    0, 0, 0, 
    
    -- channel=8
    318, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=12
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 
    0, 137, 0, 
    0, 0, 0, 
    
    -- channel=14
    221, 0, 473, 
    50, 0, 0, 
    0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 
    0, 0, 507, 
    0, 114, 116, 
    
    -- channel=17
    58, 214, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=22
    478, 201, 693, 
    299, 0, 283, 
    486, 0, 124, 
    
    -- channel=23
    281, 0, 250, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=24
    52, 164, 319, 
    0, 183, 213, 
    0, 60, 671, 
    
    -- channel=25
    0, 0, 0, 
    0, 45, 0, 
    0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=28
    589, 186, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=29
    12, 0, 0, 
    467, 0, 191, 
    0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 
    0, 142, 125, 
    0, 0, 0, 
    
    -- channel=31
    47, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=33
    207, 45, 0, 
    114, 0, 0, 
    0, 0, 0, 
    
    -- channel=34
    195, 578, 0, 
    368, 165, 0, 
    889, 0, 0, 
    
    -- channel=35
    0, 0, 0, 
    0, 0, 0, 
    0, 168, 108, 
    
    -- channel=36
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 
    334, 308, 0, 
    176, 0, 42, 
    
    -- channel=40
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=41
    40, 0, 308, 
    381, 0, 0, 
    104, 0, 0, 
    
    -- channel=42
    0, 736, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=44
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 
    0, 0, 0, 
    326, 0, 0, 
    
    -- channel=47
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=48
    156, 0, 304, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=50
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=51
    0, 150, 0, 
    0, 95, 0, 
    0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=54
    313, 154, 0, 
    251, 265, 0, 
    0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 
    0, 464, 0, 
    0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=59
    61, 20, 0, 
    187, 0, 392, 
    0, 0, 0, 
    
    -- channel=60
    117, 114, 0, 
    328, 28, 0, 
    54, 0, 0, 
    
    -- channel=61
    0, 274, 0, 
    0, 563, 469, 
    199, 0, 0, 
    
    -- channel=62
    0, 0, 0, 
    0, 62, 0, 
    0, 0, 0, 
    
    -- channel=63
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=64
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=65
    396, 0, 0, 
    326, 343, 753, 
    0, 352, 0, 
    
    -- channel=66
    614, 0, 604, 
    496, 0, 0, 
    360, 10, 0, 
    
    -- channel=67
    301, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=68
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=69
    0, 0, 260, 
    137, 0, 146, 
    0, 0, 166, 
    
    -- channel=70
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=71
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=72
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=73
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=75
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=77
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=78
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=79
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=80
    0, 0, 303, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 
    102, 192, 0, 
    8, 0, 0, 
    
    -- channel=83
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=85
    125, 325, 14, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=88
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=89
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=90
    13, 0, 338, 
    217, 0, 0, 
    386, 378, 0, 
    
    -- channel=91
    0, 0, 298, 
    350, 406, 250, 
    0, 0, 0, 
    
    -- channel=92
    0, 0, 310, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=93
    0, 0, 0, 
    278, 0, 0, 
    0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 
    46, 0, 0, 
    0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=96
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 
    286, 0, 180, 
    0, 0, 0, 
    
    -- channel=99
    307, 97, 120, 
    182, 0, 0, 
    0, 0, 0, 
    
    -- channel=100
    0, 475, 0, 
    0, 233, 0, 
    0, 311, 0, 
    
    -- channel=101
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=102
    0, 0, 268, 
    0, 75, 0, 
    0, 0, 0, 
    
    -- channel=103
    157, 59, 127, 
    641, 0, 0, 
    0, 0, 302, 
    
    -- channel=104
    0, 0, 0, 
    0, 0, 0, 
    0, 251, 0, 
    
    -- channel=105
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 
    0, 0, 0, 
    0, 293, 0, 
    
    -- channel=109
    0, 0, 66, 
    0, 0, 0, 
    399, 0, 29, 
    
    -- channel=110
    0, 0, 0, 
    205, 205, 0, 
    155, 0, 0, 
    
    -- channel=111
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=112
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=113
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=114
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=115
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=116
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=117
    0, 210, 0, 
    0, 386, 0, 
    0, 0, 0, 
    
    -- channel=118
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=119
    0, 134, 8, 
    0, 0, 0, 
    0, 0, 55, 
    
    -- channel=120
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=121
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 
    0, 0, 115, 
    146, 0, 0, 
    
    -- channel=124
    0, 30, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=125
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=128
    0, 0, 0, 
    0, 0, 69, 
    0, 0, 0, 
    
    -- channel=129
    0, 0, 0, 
    0, 0, 0, 
    163, 0, 0, 
    
    -- channel=130
    0, 0, 21, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=131
    0, 0, 0, 
    0, 0, 0, 
    0, 11, 250, 
    
    -- channel=132
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=133
    0, 0, 0, 
    0, 0, 0, 
    0, 110, 0, 
    
    -- channel=134
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=135
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=136
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=137
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=138
    0, 40, 258, 
    0, 188, 304, 
    0, 106, 173, 
    
    -- channel=139
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=140
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=141
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=142
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=143
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=144
    0, 0, 0, 
    0, 13, 0, 
    0, 0, 0, 
    
    -- channel=145
    0, 0, 577, 
    600, 313, 290, 
    191, 0, 0, 
    
    -- channel=146
    0, 0, 0, 
    54, 380, 5, 
    489, 340, 801, 
    
    -- channel=147
    288, 50, 58, 
    0, 0, 33, 
    0, 156, 176, 
    
    -- channel=148
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=149
    0, 0, 0, 
    200, 0, 0, 
    0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=152
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=153
    0, 0, 0, 
    0, 0, 0, 
    0, 432, 465, 
    
    -- channel=154
    0, 0, 0, 
    304, 0, 0, 
    0, 0, 0, 
    
    -- channel=155
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=156
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=157
    193, 202, 272, 
    0, 235, 0, 
    80, 0, 0, 
    
    -- channel=158
    473, 528, 0, 
    654, 256, 0, 
    0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=160
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=161
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=162
    142, 108, 0, 
    340, 0, 19, 
    0, 0, 0, 
    
    -- channel=163
    0, 0, 0, 
    0, 371, 120, 
    0, 0, 0, 
    
    -- channel=164
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=165
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=166
    0, 361, 0, 
    0, 0, 0, 
    136, 0, 0, 
    
    -- channel=167
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=168
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=169
    0, 0, 0, 
    0, 217, 16, 
    0, 0, 0, 
    
    -- channel=170
    0, 0, 0, 
    0, 0, 112, 
    0, 0, 0, 
    
    -- channel=171
    0, 0, 0, 
    0, 0, 84, 
    0, 0, 0, 
    
    -- channel=172
    10, 35, 0, 
    0, 287, 383, 
    0, 0, 0, 
    
    -- channel=173
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=174
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=176
    0, 0, 434, 
    0, 0, 0, 
    0, 153, 0, 
    
    -- channel=177
    0, 0, 0, 
    0, 0, 161, 
    0, 0, 0, 
    
    -- channel=178
    0, 30, 470, 
    161, 103, 40, 
    0, 0, 0, 
    
    -- channel=179
    289, 0, 0, 
    0, 0, 97, 
    687, 795, 110, 
    
    -- channel=180
    16, 0, 0, 
    14, 0, 0, 
    0, 0, 0, 
    
    -- channel=181
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=182
    0, 112, 0, 
    0, 22, 289, 
    0, 0, 0, 
    
    -- channel=183
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=184
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=185
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=186
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=187
    0, 0, 0, 
    123, 0, 116, 
    0, 0, 0, 
    
    -- channel=188
    0, 0, 0, 
    0, 0, 0, 
    0, 170, 219, 
    
    -- channel=189
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=190
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=191
    0, 0, 93, 
    165, 312, 0, 
    0, 0, 0, 
    
    -- channel=192
    0, 0, 0, 
    0, 0, 141, 
    492, 0, 0, 
    
    -- channel=193
    0, 0, 0, 
    0, 0, 0, 
    0, 496, 0, 
    
    -- channel=194
    0, 0, 0, 
    0, 131, 0, 
    0, 0, 0, 
    
    -- channel=195
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=196
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=197
    0, 0, 0, 
    176, 0, 0, 
    0, 0, 0, 
    
    -- channel=198
    0, 0, 419, 
    0, 846, 0, 
    404, 0, 15, 
    
    -- channel=199
    532, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=200
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=201
    257, 10, 295, 
    0, 287, 0, 
    0, 0, 0, 
    
    -- channel=202
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=203
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=204
    0, 0, 293, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=205
    592, 0, 0, 
    267, 0, 0, 
    0, 0, 0, 
    
    -- channel=206
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=207
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=208
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=209
    245, 81, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=210
    773, 0, 442, 
    0, 0, 0, 
    170, 0, 0, 
    
    -- channel=211
    0, 16, 0, 
    0, 122, 0, 
    233, 128, 162, 
    
    -- channel=212
    187, 462, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=213
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=214
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=215
    81, 0, 272, 
    0, 95, 130, 
    0, 0, 0, 
    
    -- channel=216
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=217
    117, 0, 303, 
    510, 0, 0, 
    631, 0, 0, 
    
    -- channel=218
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=219
    0, 0, 145, 
    0, 0, 109, 
    0, 0, 0, 
    
    -- channel=220
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=221
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=222
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=223
    0, 9, 0, 
    53, 0, 0, 
    24, 0, 0, 
    
    -- channel=224
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=225
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=226
    0, 0, 49, 
    0, 465, 0, 
    0, 0, 0, 
    
    -- channel=227
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=228
    0, 514, 0, 
    0, 0, 0, 
    315, 88, 98, 
    
    -- channel=229
    0, 258, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=230
    345, 0, 0, 
    117, 0, 0, 
    746, 0, 0, 
    
    -- channel=231
    0, 13, 0, 
    0, 0, 229, 
    0, 0, 0, 
    
    -- channel=232
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=233
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=234
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=235
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=236
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=237
    167, 84, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=238
    0, 0, 0, 
    35, 0, 58, 
    0, 0, 0, 
    
    -- channel=239
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=240
    0, 0, 0, 
    0, 0, 0, 
    0, 760, 62, 
    
    -- channel=241
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=242
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=243
    0, 0, 45, 
    481, 81, 281, 
    0, 0, 0, 
    
    -- channel=244
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=245
    0, 347, 0, 
    513, 0, 75, 
    0, 0, 0, 
    
    -- channel=246
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=247
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 53, 
    
    -- channel=248
    623, 0, 21, 
    283, 0, 0, 
    0, 0, 0, 
    
    -- channel=249
    163, 236, 395, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=250
    0, 0, 68, 
    0, 117, 0, 
    666, 0, 0, 
    
    -- channel=251
    0, 18, 0, 
    0, 27, 205, 
    0, 0, 0, 
    
    -- channel=252
    345, 147, 0, 
    0, 0, 430, 
    0, 0, 0, 
    
    -- channel=253
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=254
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=255
    361, 0, 0, 
    0, 0, 0, 
    0, 120, 253, 
    
    -- channel=256
    118, 0, 58, 
    0, 218, 387, 
    422, 0, 0, 
    
    -- channel=257
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=258
    0, 0, 0, 
    0, 0, 219, 
    393, 222, 63, 
    
    -- channel=259
    0, 0, 166, 
    278, 0, 0, 
    158, 0, 353, 
    
    -- channel=260
    0, 0, 68, 
    608, 0, 0, 
    0, 0, 0, 
    
    -- channel=261
    193, 0, 88, 
    149, 0, 0, 
    0, 0, 0, 
    
    -- channel=262
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=263
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=264
    0, 0, 0, 
    0, 0, 323, 
    0, 144, 0, 
    
    -- channel=265
    0, 0, 0, 
    204, 0, 255, 
    0, 0, 0, 
    
    -- channel=266
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=267
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=268
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=269
    0, 0, 91, 
    0, 48, 0, 
    0, 0, 0, 
    
    -- channel=270
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=271
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=272
    0, 0, 401, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=273
    96, 186, 0, 
    81, 131, 184, 
    302, 0, 0, 
    
    -- channel=274
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=275
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=276
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=277
    0, 0, 0, 
    0, 0, 0, 
    0, 59, 546, 
    
    -- channel=278
    497, 0, 286, 
    454, 0, 0, 
    0, 32, 359, 
    
    -- channel=279
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=280
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=281
    0, 0, 0, 
    0, 0, 0, 
    0, 258, 0, 
    
    -- channel=282
    0, 0, 0, 
    0, 0, 0, 
    0, 655, 0, 
    
    -- channel=283
    106, 21, 40, 
    287, 76, 157, 
    77, 0, 0, 
    
    -- channel=284
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 141, 
    
    -- channel=285
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=286
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=287
    0, 0, 0, 
    0, 105, 0, 
    0, 0, 0, 
    
    -- channel=288
    0, 97, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=289
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=290
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=291
    369, 386, 446, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=292
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=293
    154, 29, 30, 
    633, 373, 76, 
    0, 0, 0, 
    
    -- channel=294
    0, 0, 35, 
    401, 718, 0, 
    0, 0, 0, 
    
    -- channel=295
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=296
    0, 0, 0, 
    177, 0, 896, 
    0, 0, 42, 
    
    -- channel=297
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=298
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=299
    0, 320, 0, 
    0, 220, 21, 
    158, 0, 0, 
    
    -- channel=300
    0, 0, 318, 
    0, 0, 0, 
    0, 90, 0, 
    
    -- channel=301
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=302
    186, 208, 204, 
    0, 0, 329, 
    0, 0, 0, 
    
    -- channel=303
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=304
    0, 86, 0, 
    153, 0, 0, 
    0, 205, 0, 
    
    -- channel=305
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=306
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=307
    0, 0, 0, 
    0, 0, 0, 
    0, 194, 137, 
    
    -- channel=308
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 74, 
    
    -- channel=309
    0, 0, 0, 
    0, 0, 127, 
    3, 0, 0, 
    
    -- channel=310
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=311
    0, 181, 229, 
    781, 105, 0, 
    141, 0, 0, 
    
    -- channel=312
    0, 0, 0, 
    130, 0, 0, 
    0, 0, 0, 
    
    -- channel=313
    383, 0, 0, 
    0, 0, 167, 
    27, 0, 0, 
    
    -- channel=314
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=315
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=316
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=317
    0, 0, 0, 
    0, 0, 31, 
    0, 0, 0, 
    
    -- channel=318
    0, 0, 0, 
    0, 1, 0, 
    0, 0, 0, 
    
    -- channel=319
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=320
    0, 0, 0, 
    67, 57, 0, 
    0, 0, 0, 
    
    -- channel=321
    99, 319, 229, 
    240, 0, 53, 
    0, 0, 0, 
    
    -- channel=322
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=323
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=324
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=325
    443, 86, 0, 
    478, 451, 582, 
    0, 0, 0, 
    
    -- channel=326
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=327
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=328
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=329
    0, 0, 0, 
    0, 0, 0, 
    0, 115, 0, 
    
    -- channel=330
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=331
    0, 0, 444, 
    604, 0, 0, 
    238, 0, 0, 
    
    -- channel=332
    0, 164, 0, 
    349, 0, 0, 
    0, 0, 0, 
    
    -- channel=333
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=334
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=335
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=336
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=337
    0, 0, 218, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=338
    353, 3, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=339
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=340
    0, 190, 0, 
    58, 71, 122, 
    0, 0, 83, 
    
    -- channel=341
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=342
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=343
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=344
    0, 0, 479, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=345
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=346
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=347
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=348
    158, 0, 0, 
    489, 334, 333, 
    183, 0, 0, 
    
    -- channel=349
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=350
    0, 127, 370, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=351
    0, 0, 0, 
    0, 0, 0, 
    148, 560, 0, 
    
    -- channel=352
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=353
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=354
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=355
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=356
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=357
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=358
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=359
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=360
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=361
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=362
    225, 216, 517, 
    45, 0, 482, 
    0, 0, 0, 
    
    -- channel=363
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=364
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=365
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=366
    0, 0, 0, 
    210, 0, 0, 
    0, 0, 0, 
    
    -- channel=367
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=368
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=369
    0, 0, 0, 
    0, 0, 0, 
    0, 165, 232, 
    
    -- channel=370
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=371
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=372
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=373
    0, 108, 51, 
    132, 0, 0, 
    0, 0, 0, 
    
    -- channel=374
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=375
    0, 0, 32, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=376
    0, 0, 0, 
    400, 0, 268, 
    316, 0, 192, 
    
    -- channel=377
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=378
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=379
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=380
    0, 432, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=381
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=382
    77, 0, 0, 
    0, 0, 446, 
    0, 0, 0, 
    
    -- channel=383
    0, 0, 0, 
    0, 0, 12, 
    186, 0, 466, 
    
    -- channel=384
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=385
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=386
    129, 530, 213, 
    0, 190, 0, 
    0, 0, 0, 
    
    -- channel=387
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=388
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=389
    0, 118, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=390
    0, 0, 439, 
    0, 0, 605, 
    0, 473, 0, 
    
    -- channel=391
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=392
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=393
    0, 0, 11, 
    114, 0, 0, 
    104, 0, 0, 
    
    -- channel=394
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=395
    0, 0, 0, 
    0, 0, 0, 
    0, 505, 355, 
    
    -- channel=396
    0, 0, 0, 
    0, 0, 0, 
    0, 414, 315, 
    
    -- channel=397
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=398
    34, 437, 660, 
    0, 0, 0, 
    0, 33, 0, 
    
    -- channel=399
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=400
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=401
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=402
    0, 258, 136, 
    149, 0, 76, 
    0, 296, 0, 
    
    -- channel=403
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=404
    190, 140, 151, 
    245, 0, 231, 
    0, 0, 0, 
    
    -- channel=405
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=406
    0, 0, 0, 
    0, 0, 47, 
    711, 0, 0, 
    
    -- channel=407
    214, 290, 564, 
    152, 0, 0, 
    0, 0, 0, 
    
    -- channel=408
    0, 0, 371, 
    314, 0, 66, 
    0, 0, 0, 
    
    -- channel=409
    0, 0, 0, 
    0, 201, 0, 
    121, 0, 0, 
    
    -- channel=410
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=411
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=412
    0, 0, 0, 
    47, 104, 390, 
    700, 0, 0, 
    
    -- channel=413
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=414
    0, 0, 364, 
    286, 0, 0, 
    0, 0, 0, 
    
    -- channel=415
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=416
    407, 0, 0, 
    2, 0, 0, 
    0, 0, 0, 
    
    -- channel=417
    0, 137, 0, 
    258, 0, 0, 
    0, 49, 457, 
    
    -- channel=418
    0, 0, 381, 
    566, 580, 0, 
    0, 0, 0, 
    
    -- channel=419
    0, 340, 0, 
    0, 277, 0, 
    0, 0, 0, 
    
    -- channel=420
    0, 0, 0, 
    0, 112, 0, 
    0, 0, 0, 
    
    -- channel=421
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=422
    238, 291, 53, 
    704, 0, 0, 
    0, 0, 21, 
    
    -- channel=423
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=424
    0, 476, 0, 
    0, 0, 457, 
    0, 0, 0, 
    
    -- channel=425
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=426
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=427
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=428
    671, 0, 561, 
    0, 24, 0, 
    0, 0, 0, 
    
    -- channel=429
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=430
    0, 527, 0, 
    0, 140, 119, 
    0, 0, 0, 
    
    -- channel=431
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=432
    0, 0, 0, 
    4, 0, 0, 
    0, 506, 179, 
    
    -- channel=433
    681, 0, 302, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=434
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=435
    0, 0, 0, 
    117, 67, 0, 
    124, 0, 0, 
    
    -- channel=436
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 159, 
    
    -- channel=437
    0, 0, 0, 
    196, 0, 783, 
    754, 539, 114, 
    
    -- channel=438
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=439
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=440
    0, 0, 0, 
    0, 0, 0, 
    0, 178, 98, 
    
    -- channel=441
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=442
    165, 0, 0, 
    0, 4, 0, 
    0, 0, 0, 
    
    -- channel=443
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=444
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=445
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=446
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=447
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=448
    107, 0, 382, 
    0, 640, 135, 
    0, 0, 0, 
    
    -- channel=449
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=450
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=451
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=452
    0, 0, 40, 
    0, 285, 44, 
    377, 0, 0, 
    
    -- channel=453
    260, 0, 0, 
    0, 0, 0, 
    49, 0, 0, 
    
    -- channel=454
    687, 0, 0, 
    0, 0, 139, 
    0, 0, 0, 
    
    -- channel=455
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=456
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=457
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=458
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=459
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=460
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=461
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=462
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=463
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=464
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=465
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=466
    0, 0, 0, 
    0, 0, 114, 
    0, 0, 0, 
    
    -- channel=467
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=468
    0, 0, 0, 
    102, 0, 498, 
    509, 825, 319, 
    
    -- channel=469
    0, 0, 9, 
    35, 0, 0, 
    0, 0, 0, 
    
    -- channel=470
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=471
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=472
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=473
    0, 19, 374, 
    0, 0, 44, 
    0, 0, 19, 
    
    -- channel=474
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=475
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=476
    0, 189, 0, 
    416, 0, 244, 
    0, 0, 0, 
    
    -- channel=477
    0, 136, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=478
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=479
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=480
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=481
    0, 0, 0, 
    0, 29, 70, 
    0, 0, 0, 
    
    -- channel=482
    0, 287, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=483
    0, 0, 0, 
    361, 2, 384, 
    0, 0, 64, 
    
    -- channel=484
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=485
    0, 0, 0, 
    0, 0, 18, 
    0, 0, 0, 
    
    -- channel=486
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=487
    0, 0, 120, 
    208, 0, 197, 
    0, 0, 0, 
    
    -- channel=488
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=489
    159, 659, 139, 
    0, 86, 0, 
    0, 344, 0, 
    
    -- channel=490
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=491
    0, 63, 0, 
    0, 220, 0, 
    0, 0, 0, 
    
    -- channel=492
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=493
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=494
    269, 0, 142, 
    0, 0, 215, 
    0, 0, 0, 
    
    -- channel=495
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 652, 
    
    -- channel=496
    0, 0, 0, 
    0, 0, 256, 
    650, 0, 0, 
    
    -- channel=497
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=498
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=499
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=500
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=501
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=502
    133, 379, 0, 
    131, 0, 554, 
    1038, 0, 0, 
    
    -- channel=503
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=504
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=505
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=506
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=507
    0, 0, 0, 
    0, 224, 308, 
    33, 0, 0, 
    
    -- channel=508
    0, 0, 378, 
    0, 0, 0, 
    0, 608, 154, 
    
    -- channel=509
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=510
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=511
    0, 0, 100, 
    655, 0, 199, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
