library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    47, 47, 52, 47, 47, 45, 54, 54, 41, 24, 23, 39, 43, 41, 35, 
    52, 52, 53, 46, 53, 64, 27, 29, 5, 24, 2, 6, 26, 43, 38, 
    2, 65, 53, 50, 51, 22, 2, 0, 12, 41, 0, 5, 0, 21, 54, 
    0, 80, 48, 53, 26, 38, 4, 0, 1, 41, 0, 0, 0, 0, 66, 
    0, 44, 26, 67, 28, 14, 0, 0, 0, 71, 2, 0, 8, 0, 26, 
    0, 26, 25, 11, 41, 12, 0, 0, 0, 107, 0, 0, 11, 0, 2, 
    0, 0, 33, 4, 46, 50, 0, 0, 0, 80, 0, 0, 9, 13, 0, 
    0, 0, 0, 12, 32, 34, 0, 0, 0, 59, 0, 0, 14, 10, 32, 
    0, 1, 0, 37, 0, 7, 0, 0, 34, 0, 0, 0, 17, 48, 48, 
    0, 0, 0, 37, 0, 13, 42, 0, 0, 0, 0, 0, 38, 59, 29, 
    34, 0, 0, 96, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    26, 31, 30, 31, 31, 31, 32, 33, 35, 27, 15, 14, 20, 29, 30, 
    28, 39, 33, 34, 28, 40, 39, 35, 15, 1, 12, 16, 7, 8, 26, 
    30, 0, 32, 33, 34, 19, 8, 4, 5, 0, 3, 0, 11, 1, 10, 
    32, 4, 31, 32, 41, 4, 27, 6, 0, 0, 0, 3, 0, 6, 0, 
    0, 15, 27, 0, 31, 28, 13, 8, 3, 0, 9, 17, 1, 6, 7, 
    0, 0, 16, 44, 0, 0, 13, 9, 22, 0, 2, 0, 0, 0, 7, 
    0, 10, 0, 41, 1, 0, 1, 0, 10, 0, 0, 4, 0, 0, 5, 
    0, 0, 0, 17, 6, 1, 0, 0, 0, 1, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 16, 0, 21, 5, 0, 0, 0, 30, 
    0, 0, 0, 0, 5, 0, 0, 19, 10, 0, 0, 0, 0, 20, 20, 
    0, 0, 0, 0, 9, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    9, 6, 8, 5, 7, 10, 5, 6, 8, 7, 7, 13, 10, 5, 8, 
    12, 9, 8, 3, 12, 17, 0, 1, 2, 34, 14, 16, 26, 25, 9, 
    0, 36, 10, 6, 12, 23, 0, 22, 27, 47, 0, 2, 0, 31, 27, 
    0, 67, 9, 15, 0, 31, 3, 0, 10, 53, 0, 8, 3, 8, 59, 
    0, 30, 0, 48, 0, 0, 0, 0, 3, 76, 3, 0, 17, 0, 32, 
    0, 13, 0, 0, 55, 0, 0, 0, 0, 106, 0, 0, 25, 3, 5, 
    0, 0, 12, 0, 56, 32, 0, 0, 0, 89, 0, 0, 25, 29, 0, 
    0, 0, 0, 1, 39, 27, 0, 2, 0, 54, 0, 0, 32, 8, 4, 
    0, 4, 0, 37, 0, 24, 10, 13, 34, 6, 31, 0, 35, 33, 13, 
    0, 1, 0, 59, 0, 0, 36, 0, 0, 0, 0, 28, 41, 29, 3, 
    55, 0, 0, 90, 0, 0, 9, 0, 0, 3, 35, 28, 28, 40, 26, 
    59, 28, 0, 49, 0, 0, 36, 35, 22, 27, 27, 29, 29, 26, 19, 
    12, 55, 54, 0, 0, 20, 17, 23, 26, 29, 33, 27, 17, 24, 31, 
    11, 29, 72, 0, 2, 26, 15, 22, 25, 24, 24, 27, 25, 38, 2, 
    0, 26, 30, 37, 21, 36, 25, 19, 24, 23, 14, 31, 47, 2, 0, 
    
    -- channel=3
    5, 6, 0, 0, 0, 2, 1, 2, 2, 16, 27, 20, 5, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 17, 35, 0, 0, 0, 18, 16, 1, 
    36, 36, 1, 0, 0, 34, 23, 15, 0, 0, 0, 0, 0, 20, 6, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 14, 0, 9, 5, 6, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 13, 
    12, 0, 0, 15, 52, 22, 0, 0, 0, 0, 5, 14, 1, 0, 0, 
    0, 0, 28, 0, 10, 0, 9, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 30, 25, 6, 0, 6, 0, 4, 8, 0, 
    0, 0, 0, 0, 0, 34, 2, 0, 0, 0, 28, 36, 12, 0, 0, 
    7, 0, 0, 0, 6, 13, 0, 0, 0, 45, 33, 9, 0, 0, 7, 
    2, 0, 0, 0, 0, 0, 4, 36, 23, 0, 0, 0, 0, 18, 20, 
    49, 27, 0, 0, 52, 57, 27, 25, 16, 4, 0, 0, 0, 0, 0, 
    0, 36, 10, 7, 52, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 40, 46, 13, 0, 0, 0, 0, 0, 0, 7, 0, 0, 24, 
    0, 0, 3, 31, 11, 16, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    14, 17, 20, 18, 16, 19, 19, 18, 16, 12, 6, 10, 14, 8, 5, 
    16, 21, 23, 18, 25, 51, 14, 16, 0, 11, 3, 0, 0, 10, 10, 
    0, 24, 20, 18, 19, 8, 0, 0, 0, 31, 0, 0, 0, 0, 15, 
    0, 29, 16, 25, 14, 25, 17, 0, 0, 23, 0, 0, 0, 0, 16, 
    0, 45, 7, 63, 82, 42, 0, 0, 0, 30, 14, 0, 0, 0, 0, 
    0, 28, 4, 0, 25, 16, 16, 0, 0, 78, 0, 0, 0, 0, 0, 
    0, 1, 1, 0, 29, 47, 28, 8, 0, 67, 0, 0, 0, 4, 0, 
    8, 18, 0, 14, 30, 66, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    15, 33, 0, 27, 0, 0, 0, 0, 18, 0, 0, 0, 0, 3, 18, 
    22, 24, 0, 31, 0, 0, 28, 25, 0, 0, 0, 0, 12, 29, 12, 
    49, 26, 0, 91, 43, 25, 53, 19, 0, 0, 0, 5, 1, 9, 0, 
    4, 33, 23, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 50, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 10, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 9, 14, 0, 0, 
    19, 19, 0, 0, 0, 0, 26, 13, 4, 0, 0, 0, 0, 0, 0, 
    33, 53, 9, 18, 89, 53, 0, 0, 0, 0, 16, 15, 6, 15, 0, 
    0, 0, 3, 0, 0, 0, 14, 11, 11, 27, 0, 0, 0, 9, 21, 
    0, 0, 0, 0, 0, 6, 4, 7, 6, 10, 0, 0, 0, 8, 11, 
    1, 9, 20, 17, 14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 2, 0, 9, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 2, 7, 0, 0, 40, 0, 0, 0, 0, 27, 18, 0, 
    0, 0, 0, 31, 94, 73, 33, 0, 8, 4, 17, 42, 20, 0, 0, 
    0, 0, 21, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 10, 2, 0, 13, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 23, 16, 3, 
    
    -- channel=6
    22, 21, 25, 26, 26, 21, 28, 26, 24, 17, 5, 4, 11, 20, 18, 
    24, 26, 30, 28, 26, 32, 34, 17, 4, 0, 5, 0, 0, 0, 17, 
    9, 0, 26, 25, 32, 12, 0, 0, 0, 12, 15, 0, 15, 0, 1, 
    10, 12, 26, 23, 23, 0, 24, 13, 5, 7, 4, 7, 0, 0, 0, 
    4, 46, 33, 14, 46, 64, 14, 1, 0, 0, 15, 18, 0, 0, 5, 
    9, 6, 22, 48, 0, 0, 17, 9, 8, 22, 25, 0, 0, 0, 3, 
    2, 30, 0, 15, 14, 15, 21, 12, 0, 31, 0, 0, 0, 1, 12, 
    16, 1, 19, 6, 32, 35, 6, 0, 0, 32, 1, 0, 0, 9, 0, 
    17, 12, 12, 0, 30, 0, 0, 9, 0, 29, 0, 0, 0, 0, 35, 
    1, 17, 1, 8, 3, 8, 0, 30, 25, 0, 0, 0, 3, 33, 19, 
    0, 16, 0, 16, 54, 49, 44, 0, 0, 0, 0, 5, 3, 0, 0, 
    0, 0, 4, 73, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    
    -- channel=7
    38, 41, 37, 39, 38, 35, 44, 41, 37, 45, 45, 41, 34, 33, 32, 
    35, 38, 40, 43, 35, 34, 40, 51, 49, 10, 11, 14, 22, 34, 37, 
    61, 46, 40, 39, 39, 60, 29, 4, 0, 10, 24, 11, 24, 18, 36, 
    29, 3, 42, 37, 46, 9, 29, 14, 16, 20, 30, 21, 11, 11, 22, 
    11, 33, 42, 5, 52, 21, 32, 14, 22, 0, 15, 18, 12, 15, 8, 
    1, 41, 38, 23, 41, 15, 34, 14, 23, 0, 43, 16, 16, 12, 0, 
    0, 61, 29, 46, 33, 9, 68, 22, 32, 22, 28, 8, 1, 3, 16, 
    0, 33, 4, 37, 13, 67, 53, 32, 20, 27, 25, 11, 8, 29, 13, 
    15, 30, 11, 26, 14, 15, 8, 19, 8, 24, 29, 26, 3, 9, 31, 
    29, 24, 31, 0, 34, 8, 0, 34, 13, 48, 37, 2, 16, 39, 43, 
    38, 23, 30, 0, 27, 18, 52, 66, 42, 7, 0, 0, 9, 27, 22, 
    39, 30, 19, 44, 82, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 
    1, 17, 0, 85, 9, 0, 1, 0, 0, 0, 0, 0, 9, 1, 0, 
    0, 0, 7, 92, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 30, 
    1, 0, 0, 22, 1, 0, 9, 0, 0, 0, 0, 0, 0, 7, 0, 
    
    -- channel=8
    0, 2, 0, 2, 1, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 4, 0, 22, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 4, 0, 0, 7, 0, 0, 0, 7, 6, 3, 0, 0, 
    29, 0, 5, 0, 8, 0, 8, 0, 0, 0, 30, 0, 0, 0, 0, 
    36, 8, 24, 0, 45, 23, 34, 12, 0, 0, 18, 16, 0, 3, 0, 
    14, 22, 38, 0, 0, 10, 48, 15, 23, 0, 37, 18, 0, 0, 0, 
    22, 38, 5, 17, 0, 0, 24, 29, 23, 0, 38, 11, 0, 0, 6, 
    26, 45, 11, 18, 0, 0, 46, 0, 12, 0, 22, 13, 0, 0, 10, 
    39, 18, 38, 0, 1, 0, 8, 1, 0, 10, 0, 7, 0, 0, 0, 
    25, 16, 55, 0, 16, 0, 0, 30, 1, 0, 3, 0, 0, 0, 2, 
    0, 19, 50, 0, 88, 14, 0, 17, 26, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 46, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 34, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 48, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 5, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 0, 4, 0, 8, 0, 0, 0, 0, 0, 
    0, 8, 0, 13, 0, 0, 0, 0, 0, 0, 11, 0, 1, 0, 0, 
    15, 6, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    38, 1, 0, 23, 0, 0, 27, 27, 3, 0, 0, 1, 4, 6, 0, 
    53, 44, 0, 16, 7, 27, 20, 20, 21, 17, 22, 21, 23, 20, 22, 
    21, 44, 33, 21, 1, 19, 17, 17, 15, 18, 18, 21, 27, 28, 24, 
    26, 25, 54, 42, 18, 16, 11, 16, 21, 23, 25, 34, 26, 37, 42, 
    23, 31, 29, 21, 16, 33, 35, 23, 18, 15, 16, 20, 23, 16, 15, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 3, 7, 6, 3, 6, 2, 0, 2, 0, 0, 0, 2, 0, 0, 
    5, 8, 6, 3, 11, 72, 5, 0, 0, 12, 21, 0, 0, 0, 0, 
    0, 0, 3, 4, 0, 0, 0, 0, 3, 41, 25, 31, 0, 0, 0, 
    0, 30, 0, 8, 5, 19, 35, 14, 6, 5, 27, 0, 0, 0, 0, 
    52, 63, 8, 42, 116, 72, 30, 20, 0, 39, 48, 18, 17, 6, 0, 
    30, 52, 21, 0, 8, 37, 66, 28, 8, 78, 32, 3, 7, 16, 16, 
    62, 24, 0, 0, 0, 74, 31, 47, 6, 49, 24, 17, 10, 29, 17, 
    71, 64, 25, 15, 16, 47, 16, 0, 11, 29, 28, 3, 7, 2, 16, 
    76, 62, 30, 40, 22, 0, 9, 23, 31, 0, 0, 0, 0, 20, 18, 
    63, 60, 38, 45, 15, 16, 52, 63, 11, 0, 0, 0, 13, 20, 0, 
    52, 59, 23, 129, 146, 72, 50, 22, 16, 3, 18, 36, 18, 0, 0, 
    0, 45, 67, 105, 0, 0, 0, 0, 0, 4, 11, 13, 27, 24, 23, 
    17, 0, 79, 39, 0, 23, 13, 12, 13, 20, 29, 36, 20, 21, 57, 
    21, 16, 9, 2, 15, 24, 25, 13, 17, 24, 17, 10, 18, 44, 0, 
    24, 23, 5, 0, 0, 0, 1, 23, 35, 40, 19, 24, 69, 49, 15, 
    
    -- channel=12
    1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 4, 0, 4, 4, 0, 0, 0, 1, 0, 0, 7, 4, 0, 
    0, 11, 1, 0, 6, 0, 0, 0, 10, 35, 0, 0, 0, 16, 7, 
    0, 64, 0, 1, 0, 3, 0, 0, 0, 55, 0, 0, 0, 0, 43, 
    0, 35, 0, 44, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 31, 
    0, 0, 0, 14, 32, 0, 0, 0, 0, 134, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 46, 34, 0, 0, 0, 101, 0, 0, 2, 9, 0, 
    0, 0, 0, 0, 37, 51, 0, 0, 0, 66, 0, 0, 16, 3, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 15, 0, 18, 0, 17, 14, 16, 
    0, 0, 0, 38, 0, 1, 14, 0, 3, 0, 0, 0, 29, 25, 0, 
    28, 0, 0, 113, 0, 0, 32, 0, 0, 0, 3, 9, 9, 0, 0, 
    42, 2, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 45, 47, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 4, 0, 0, 6, 0, 0, 0, 0, 0, 0, 24, 0, 0, 
    
    -- channel=13
    36, 42, 41, 39, 38, 41, 44, 46, 40, 28, 23, 30, 36, 34, 33, 
    41, 49, 44, 41, 43, 50, 25, 32, 24, 21, 4, 2, 13, 31, 31, 
    11, 41, 43, 44, 43, 33, 17, 7, 7, 20, 0, 0, 0, 5, 37, 
    0, 26, 38, 45, 30, 30, 13, 0, 0, 17, 0, 0, 0, 0, 35, 
    0, 14, 18, 43, 27, 3, 0, 0, 0, 29, 6, 0, 1, 0, 1, 
    0, 5, 16, 23, 39, 13, 12, 0, 0, 43, 0, 0, 2, 0, 0, 
    0, 0, 19, 29, 34, 29, 5, 0, 0, 35, 0, 0, 0, 6, 0, 
    0, 0, 0, 21, 22, 20, 0, 0, 0, 26, 0, 0, 3, 1, 13, 
    0, 0, 0, 21, 0, 10, 7, 4, 8, 9, 10, 0, 6, 24, 30, 
    0, 0, 0, 17, 0, 0, 16, 9, 0, 0, 0, 0, 13, 33, 25, 
    21, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    70, 70, 71, 70, 71, 67, 74, 80, 75, 66, 59, 60, 60, 60, 61, 
    72, 72, 73, 72, 72, 57, 59, 68, 59, 37, 13, 20, 40, 58, 59, 
    55, 77, 74, 76, 76, 70, 53, 36, 19, 10, 0, 0, 0, 30, 55, 
    0, 31, 68, 77, 64, 53, 18, 2, 4, 20, 8, 11, 6, 5, 47, 
    0, 0, 49, 66, 14, 2, 6, 3, 4, 23, 5, 0, 4, 0, 20, 
    0, 8, 45, 54, 48, 26, 9, 2, 0, 21, 3, 6, 7, 0, 0, 
    0, 0, 50, 55, 36, 29, 16, 8, 0, 18, 3, 0, 4, 4, 0, 
    0, 0, 3, 36, 28, 21, 5, 18, 9, 22, 13, 1, 7, 9, 26, 
    0, 0, 0, 17, 17, 27, 19, 9, 14, 24, 28, 13, 12, 25, 45, 
    7, 0, 0, 1, 0, 10, 18, 0, 0, 26, 12, 6, 8, 42, 58, 
    14, 0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 4, 6, 
    0, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 6, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 
    22, 10, 0, 0, 10, 0, 0, 0, 1, 0, 5, 7, 4, 8, 0, 
    16, 17, 0, 0, 0, 0, 14, 1, 11, 1, 15, 2, 0, 4, 0, 
    14, 32, 0, 0, 0, 7, 16, 5, 1, 0, 6, 3, 6, 0, 0, 
    27, 32, 13, 6, 0, 4, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    26, 25, 28, 17, 12, 0, 1, 12, 0, 3, 17, 13, 0, 0, 0, 
    37, 20, 29, 7, 25, 13, 29, 50, 39, 24, 30, 38, 42, 44, 43, 
    74, 53, 32, 8, 55, 65, 58, 58, 62, 64, 70, 73, 76, 73, 77, 
    83, 59, 32, 30, 72, 65, 66, 62, 65, 68, 76, 77, 80, 86, 86, 
    96, 79, 46, 77, 65, 66, 65, 64, 70, 74, 81, 87, 88, 89, 95, 
    92, 87, 67, 78, 65, 68, 74, 70, 67, 71, 76, 77, 78, 90, 92, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 4, 14, 16, 0, 0, 
    5, 0, 0, 0, 0, 16, 30, 35, 0, 0, 0, 0, 0, 6, 0, 
    7, 0, 0, 0, 6, 6, 0, 0, 0, 0, 2, 0, 10, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 
    2, 0, 0, 11, 15, 0, 0, 0, 4, 0, 0, 13, 0, 0, 0, 
    0, 2, 12, 2, 0, 0, 0, 0, 0, 0, 12, 8, 5, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 9, 0, 0, 8, 18, 0, 0, 0, 
    0, 0, 10, 0, 0, 25, 22, 4, 0, 30, 7, 21, 7, 0, 0, 
    0, 0, 8, 1, 0, 0, 0, 0, 0, 0, 11, 5, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 17, 23, 
    0, 0, 0, 0, 30, 57, 41, 39, 16, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 2, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 8, 33, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=17
    39, 39, 38, 36, 37, 34, 44, 49, 35, 25, 27, 34, 33, 35, 32, 
    39, 42, 41, 39, 35, 3, 23, 28, 30, 0, 0, 0, 19, 30, 29, 
    18, 50, 42, 42, 42, 51, 15, 9, 0, 0, 0, 0, 0, 15, 31, 
    0, 9, 36, 38, 20, 10, 0, 0, 0, 7, 0, 0, 0, 0, 35, 
    0, 0, 21, 11, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 19, 
    0, 0, 19, 33, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 18, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 1, 0, 11, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 25, 0, 0, 0, 14, 0, 7, 10, 10, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 22, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 32, 10, 0, 0, 0, 25, 13, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 4, 29, 24, 31, 0, 3, 
    57, 0, 8, 0, 7, 0, 32, 10, 14, 0, 41, 4, 17, 12, 0, 
    60, 45, 22, 0, 72, 24, 42, 24, 15, 0, 38, 34, 15, 30, 0, 
    16, 47, 31, 0, 0, 4, 65, 32, 49, 0, 43, 26, 5, 21, 20, 
    17, 71, 10, 19, 0, 5, 48, 38, 48, 0, 50, 28, 8, 12, 27, 
    26, 68, 21, 37, 0, 6, 38, 12, 28, 0, 37, 30, 0, 10, 14, 
    47, 41, 44, 27, 3, 0, 23, 25, 11, 23, 0, 12, 0, 12, 8, 
    36, 34, 75, 11, 39, 0, 0, 66, 8, 0, 17, 0, 11, 5, 3, 
    27, 32, 68, 0, 119, 47, 9, 35, 45, 21, 13, 18, 14, 15, 16, 
    0, 20, 47, 25, 64, 18, 7, 6, 20, 13, 21, 19, 28, 28, 27, 
    40, 0, 0, 60, 36, 24, 25, 22, 21, 21, 25, 28, 29, 22, 35, 
    41, 30, 0, 84, 23, 21, 33, 23, 18, 22, 22, 24, 29, 22, 36, 
    44, 30, 21, 27, 15, 7, 14, 24, 25, 34, 32, 22, 25, 56, 55, 
    
    -- channel=20
    40, 33, 39, 36, 37, 36, 39, 40, 36, 28, 23, 28, 28, 32, 29, 
    38, 38, 41, 36, 42, 21, 31, 26, 13, 14, 2, 13, 25, 29, 28, 
    13, 35, 41, 37, 45, 29, 0, 10, 22, 26, 1, 0, 0, 33, 25, 
    0, 55, 36, 41, 20, 30, 3, 10, 5, 48, 0, 13, 0, 5, 43, 
    0, 25, 24, 68, 0, 32, 0, 0, 0, 59, 2, 0, 4, 0, 45, 
    10, 2, 17, 56, 16, 17, 0, 0, 0, 85, 0, 0, 13, 0, 5, 
    15, 0, 23, 0, 36, 34, 0, 0, 0, 62, 0, 0, 13, 13, 5, 
    14, 0, 24, 0, 50, 33, 0, 2, 0, 53, 0, 0, 19, 16, 16, 
    0, 0, 0, 4, 31, 18, 0, 0, 23, 9, 19, 0, 22, 22, 38, 
    0, 7, 0, 26, 0, 33, 26, 0, 31, 2, 0, 2, 21, 38, 24, 
    4, 9, 0, 69, 0, 6, 26, 0, 0, 0, 1, 2, 6, 0, 0, 
    19, 2, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=21
    9, 14, 12, 10, 10, 13, 12, 11, 9, 9, 11, 13, 14, 13, 12, 
    9, 15, 14, 11, 12, 12, 8, 13, 17, 7, 6, 8, 9, 8, 10, 
    10, 10, 9, 10, 10, 20, 0, 5, 8, 21, 5, 8, 11, 8, 13, 
    3, 12, 5, 12, 8, 9, 10, 8, 9, 20, 2, 11, 3, 5, 20, 
    0, 14, 2, 18, 16, 25, 8, 4, 10, 17, 5, 5, 11, 9, 18, 
    0, 0, 0, 19, 8, 4, 1, 7, 8, 27, 0, 0, 11, 10, 10, 
    0, 4, 0, 12, 32, 4, 4, 0, 4, 32, 0, 0, 8, 7, 4, 
    0, 0, 0, 2, 23, 18, 1, 6, 0, 27, 0, 0, 11, 11, 3, 
    0, 1, 0, 3, 1, 11, 0, 4, 4, 17, 0, 4, 13, 8, 13, 
    0, 0, 0, 19, 0, 14, 9, 8, 5, 4, 10, 13, 17, 19, 8, 
    2, 0, 0, 13, 0, 3, 21, 4, 0, 11, 3, 11, 7, 0, 0, 
    5, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 2, 0, 2, 4, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 1, 3, 0, 0, 2, 4, 0, 0, 0, 0, 1, 3, 
    6, 4, 0, 0, 1, 31, 0, 0, 0, 9, 13, 11, 0, 0, 0, 
    0, 0, 3, 4, 3, 0, 1, 12, 8, 9, 0, 0, 0, 0, 0, 
    5, 27, 1, 5, 2, 9, 9, 0, 0, 0, 0, 0, 1, 1, 0, 
    0, 10, 0, 0, 0, 0, 0, 3, 0, 20, 15, 0, 5, 1, 0, 
    0, 0, 0, 3, 0, 0, 15, 7, 12, 15, 0, 0, 0, 0, 9, 
    2, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 11, 12, 12, 0, 
    1, 4, 0, 0, 0, 0, 0, 0, 0, 3, 0, 11, 0, 0, 4, 
    0, 0, 2, 0, 4, 0, 17, 17, 0, 16, 0, 0, 1, 14, 5, 
    0, 0, 0, 20, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 18, 0, 0, 0, 0, 1, 17, 1, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 8, 7, 0, 0, 0, 0, 3, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 10, 0, 4, 14, 2, 0, 
    
    -- channel=23
    52, 50, 52, 52, 53, 43, 59, 67, 53, 32, 22, 27, 31, 43, 43, 
    52, 55, 56, 55, 51, 5, 43, 33, 16, 0, 0, 0, 3, 25, 37, 
    17, 32, 58, 59, 61, 44, 8, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 53, 52, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 38, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 33, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    7, 5, 2, 6, 7, 4, 7, 7, 10, 22, 18, 3, 0, 12, 12, 
    0, 5, 5, 10, 0, 0, 38, 22, 35, 0, 7, 19, 5, 0, 8, 
    45, 0, 3, 5, 7, 26, 19, 19, 0, 0, 23, 0, 37, 7, 0, 
    76, 0, 12, 0, 22, 0, 14, 22, 5, 0, 21, 22, 12, 22, 0, 
    32, 0, 35, 0, 0, 27, 40, 24, 25, 0, 8, 45, 0, 21, 11, 
    42, 0, 27, 38, 0, 0, 10, 25, 45, 0, 51, 33, 0, 9, 10, 
    15, 41, 0, 40, 0, 0, 28, 9, 50, 0, 41, 26, 0, 0, 20, 
    13, 2, 30, 14, 0, 0, 52, 12, 9, 0, 11, 35, 0, 8, 0, 
    16, 0, 58, 0, 27, 4, 6, 8, 0, 42, 11, 36, 0, 0, 0, 
    0, 0, 51, 0, 47, 6, 0, 12, 37, 16, 37, 2, 0, 0, 18, 
    0, 0, 55, 0, 14, 39, 0, 18, 38, 20, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 121, 15, 3, 2, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 49, 53, 0, 4, 0, 0, 0, 0, 0, 1, 0, 0, 
    4, 0, 0, 40, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 32, 
    15, 0, 0, 10, 11, 0, 0, 0, 0, 0, 9, 0, 0, 14, 23, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 3, 3, 0, 0, 5, 3, 1, 0, 0, 0, 0, 1, 0, 0, 
    3, 10, 7, 0, 8, 29, 0, 0, 0, 4, 0, 0, 0, 8, 0, 
    0, 17, 3, 0, 3, 15, 0, 0, 0, 46, 0, 0, 0, 4, 20, 
    0, 63, 3, 8, 0, 7, 0, 0, 0, 53, 0, 0, 0, 0, 51, 
    0, 59, 0, 46, 27, 0, 0, 0, 0, 56, 0, 0, 3, 0, 8, 
    0, 19, 0, 0, 45, 0, 0, 0, 0, 125, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 61, 24, 0, 0, 0, 107, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 36, 62, 0, 0, 0, 67, 0, 0, 16, 0, 0, 
    0, 2, 0, 33, 0, 0, 0, 0, 27, 0, 9, 0, 5, 27, 16, 
    0, 0, 0, 49, 0, 0, 19, 6, 0, 0, 0, 0, 45, 38, 0, 
    50, 0, 0, 118, 0, 0, 22, 0, 0, 0, 5, 9, 3, 0, 0, 
    37, 8, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 27, 32, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 6, 
    0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 30, 0, 0, 
    
    -- channel=28
    9, 21, 14, 16, 12, 13, 14, 19, 11, 5, 8, 12, 18, 10, 14, 
    15, 17, 13, 16, 15, 43, 0, 5, 10, 12, 0, 0, 0, 17, 15, 
    0, 36, 14, 19, 8, 7, 18, 0, 0, 7, 0, 16, 0, 0, 30, 
    7, 0, 8, 14, 6, 10, 9, 0, 1, 0, 26, 0, 17, 0, 8, 
    31, 0, 0, 0, 53, 0, 4, 0, 0, 0, 5, 0, 6, 14, 0, 
    0, 28, 13, 0, 40, 7, 46, 6, 12, 0, 0, 9, 1, 9, 0, 
    0, 17, 9, 31, 6, 6, 29, 17, 21, 0, 17, 0, 0, 3, 0, 
    0, 46, 0, 30, 0, 4, 16, 7, 30, 0, 29, 0, 0, 0, 24, 
    0, 9, 0, 36, 0, 0, 12, 1, 10, 0, 0, 15, 0, 26, 2, 
    30, 1, 29, 0, 0, 0, 9, 31, 0, 13, 25, 2, 11, 7, 11, 
    36, 0, 23, 0, 61, 0, 0, 29, 27, 0, 0, 0, 0, 0, 0, 
    0, 30, 27, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 83, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    13, 16, 12, 17, 16, 15, 17, 18, 16, 15, 13, 6, 13, 20, 19, 
    13, 19, 11, 20, 9, 11, 40, 20, 21, 0, 23, 19, 0, 1, 18, 
    22, 0, 16, 19, 10, 0, 31, 16, 0, 0, 22, 13, 36, 0, 0, 
    83, 0, 24, 10, 27, 0, 28, 20, 10, 0, 42, 7, 23, 19, 0, 
    68, 0, 48, 0, 39, 31, 48, 32, 19, 0, 25, 50, 5, 35, 0, 
    35, 0, 55, 4, 0, 6, 49, 37, 57, 0, 50, 44, 0, 21, 24, 
    32, 39, 13, 56, 0, 0, 25, 36, 58, 0, 58, 35, 0, 0, 27, 
    27, 37, 27, 45, 0, 0, 54, 6, 30, 0, 30, 40, 0, 1, 14, 
    34, 1, 66, 0, 23, 0, 21, 15, 0, 38, 0, 35, 0, 0, 7, 
    2, 0, 79, 0, 43, 0, 0, 41, 13, 1, 36, 2, 0, 0, 20, 
    0, 5, 73, 0, 91, 39, 0, 13, 48, 30, 0, 0, 0, 0, 7, 
    0, 0, 27, 0, 80, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 23, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 53, 9, 0, 5, 0, 0, 0, 0, 0, 0, 0, 2, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 29, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 13, 6, 3, 28, 25, 25, 0, 0, 
    45, 0, 0, 0, 0, 0, 12, 17, 15, 0, 32, 12, 27, 13, 0, 
    60, 3, 0, 0, 19, 14, 36, 27, 21, 0, 28, 32, 16, 27, 0, 
    46, 19, 0, 0, 0, 21, 38, 32, 37, 0, 38, 39, 12, 26, 21, 
    48, 39, 0, 0, 0, 0, 29, 30, 43, 0, 51, 33, 16, 15, 20, 
    42, 56, 22, 14, 0, 0, 44, 20, 28, 0, 32, 36, 10, 8, 0, 
    52, 42, 53, 11, 5, 16, 26, 18, 7, 17, 2, 31, 4, 0, 0, 
    35, 34, 67, 17, 39, 6, 11, 39, 14, 7, 31, 21, 0, 0, 0, 
    21, 34, 67, 0, 72, 39, 8, 44, 53, 43, 36, 33, 32, 31, 37, 
    31, 33, 49, 0, 77, 68, 51, 53, 55, 49, 51, 54, 59, 57, 62, 
    67, 26, 14, 39, 92, 54, 55, 53, 53, 53, 57, 59, 59, 62, 65, 
    78, 59, 1, 78, 57, 53, 60, 54, 53, 56, 60, 62, 68, 58, 68, 
    78, 64, 52, 64, 52, 45, 50, 53, 52, 61, 64, 59, 53, 77, 84, 
    
    -- channel=32
    4, 2, 5, 0, 0, 4, 2, 0, 0, 0, 0, 6, 2, 0, 0, 
    3, 4, 7, 0, 10, 3, 0, 0, 0, 12, 0, 0, 6, 17, 0, 
    0, 46, 3, 0, 6, 16, 0, 0, 7, 50, 0, 0, 0, 19, 23, 
    0, 68, 0, 9, 0, 19, 0, 0, 0, 82, 0, 0, 0, 0, 71, 
    0, 27, 0, 80, 0, 0, 0, 0, 0, 104, 0, 0, 0, 0, 27, 
    0, 13, 0, 0, 80, 4, 0, 0, 0, 166, 0, 0, 14, 0, 0, 
    0, 0, 4, 0, 73, 47, 0, 0, 0, 133, 0, 0, 4, 14, 0, 
    0, 0, 0, 0, 54, 65, 0, 0, 0, 84, 0, 0, 27, 4, 0, 
    0, 1, 0, 36, 0, 23, 0, 0, 35, 0, 15, 0, 25, 33, 13, 
    0, 4, 0, 63, 0, 0, 42, 0, 0, 0, 0, 2, 40, 31, 0, 
    59, 0, 0, 143, 0, 0, 39, 0, 0, 0, 0, 5, 9, 8, 0, 
    69, 46, 0, 91, 0, 0, 3, 1, 0, 0, 0, 3, 1, 0, 0, 
    0, 66, 95, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 3, 7, 
    0, 2, 125, 0, 0, 4, 0, 0, 3, 1, 0, 1, 0, 17, 0, 
    0, 1, 8, 0, 0, 15, 8, 0, 5, 0, 0, 6, 36, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 10, 12, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 4, 8, 0, 23, 5, 16, 6, 0, 
    29, 0, 0, 0, 0, 0, 18, 15, 16, 0, 5, 16, 3, 13, 0, 
    31, 11, 0, 0, 0, 0, 19, 10, 27, 0, 29, 24, 0, 10, 3, 
    25, 36, 0, 0, 0, 0, 12, 16, 26, 0, 34, 19, 4, 0, 13, 
    21, 30, 0, 0, 0, 0, 42, 13, 18, 0, 23, 25, 0, 9, 1, 
    32, 18, 45, 0, 0, 5, 10, 7, 0, 6, 0, 26, 0, 0, 0, 
    27, 23, 52, 0, 17, 0, 0, 16, 12, 1, 22, 0, 0, 0, 0, 
    2, 16, 52, 0, 41, 8, 0, 25, 31, 15, 6, 5, 7, 0, 2, 
    20, 14, 22, 0, 76, 55, 35, 34, 36, 30, 35, 39, 44, 47, 50, 
    61, 20, 0, 39, 72, 38, 40, 38, 41, 40, 42, 43, 48, 45, 45, 
    67, 44, 0, 73, 45, 38, 45, 39, 38, 42, 51, 53, 55, 45, 72, 
    71, 52, 45, 47, 46, 39, 42, 41, 37, 46, 54, 48, 35, 68, 72, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 28, 13, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 24, 16, 6, 0, 5, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 28, 0, 0, 0, 0, 0, 36, 11, 0, 0, 
    5, 0, 0, 0, 0, 2, 0, 0, 0, 22, 32, 9, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 22, 17, 0, 0, 0, 0, 5, 10, 
    32, 30, 0, 0, 34, 76, 39, 39, 29, 17, 15, 16, 14, 10, 16, 
    14, 28, 15, 0, 71, 13, 13, 14, 12, 9, 7, 2, 13, 22, 4, 
    24, 16, 18, 49, 31, 10, 8, 9, 15, 12, 19, 26, 26, 6, 38, 
    22, 20, 22, 40, 28, 29, 32, 20, 3, 0, 10, 17, 0, 0, 23, 
    
    -- channel=37
    10, 16, 13, 13, 10, 16, 14, 13, 14, 16, 16, 15, 13, 7, 5, 
    9, 16, 15, 14, 14, 23, 12, 23, 20, 9, 0, 0, 4, 8, 6, 
    21, 16, 13, 13, 13, 30, 14, 0, 0, 11, 7, 0, 0, 0, 7, 
    0, 0, 8, 16, 19, 12, 11, 0, 0, 15, 11, 6, 0, 0, 1, 
    5, 6, 5, 24, 38, 22, 20, 3, 0, 3, 12, 0, 0, 0, 0, 
    16, 24, 9, 26, 57, 41, 27, 3, 0, 22, 26, 4, 1, 0, 0, 
    13, 22, 12, 15, 24, 34, 42, 15, 0, 27, 17, 0, 0, 0, 0, 
    28, 24, 0, 9, 9, 52, 28, 18, 3, 20, 19, 0, 1, 6, 0, 
    35, 37, 7, 17, 12, 17, 6, 6, 0, 1, 20, 1, 0, 0, 3, 
    41, 32, 12, 12, 14, 9, 13, 15, 1, 23, 1, 0, 0, 10, 15, 
    42, 35, 13, 33, 18, 8, 39, 44, 15, 0, 0, 0, 0, 4, 3, 
    21, 40, 20, 52, 52, 11, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 31, 60, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    18, 5, 0, 0, 5, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 
    2, 18, 0, 0, 0, 0, 16, 0, 7, 0, 9, 0, 0, 0, 0, 
    5, 11, 0, 0, 0, 17, 28, 6, 0, 0, 0, 0, 0, 4, 0, 
    17, 19, 14, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    14, 14, 21, 0, 16, 0, 0, 0, 0, 15, 18, 1, 0, 0, 0, 
    16, 8, 20, 0, 0, 10, 35, 49, 37, 7, 7, 19, 27, 32, 32, 
    67, 34, 14, 0, 67, 46, 37, 37, 42, 47, 50, 51, 51, 49, 53, 
    63, 50, 3, 41, 56, 44, 47, 43, 42, 44, 48, 51, 61, 61, 52, 
    69, 55, 43, 73, 46, 43, 42, 44, 48, 52, 59, 65, 60, 62, 88, 
    70, 61, 50, 55, 49, 52, 58, 48, 44, 44, 54, 49, 41, 66, 67, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    23, 21, 23, 26, 26, 20, 22, 26, 27, 22, 17, 15, 20, 23, 27, 
    25, 23, 24, 26, 27, 13, 27, 15, 17, 11, 13, 7, 3, 15, 24, 
    8, 15, 23, 26, 23, 8, 16, 16, 13, 2, 12, 21, 18, 7, 13, 
    31, 0, 22, 24, 16, 22, 15, 19, 14, 0, 17, 6, 17, 11, 5, 
    41, 0, 30, 30, 23, 18, 12, 13, 9, 0, 14, 22, 13, 24, 1, 
    17, 0, 29, 0, 0, 7, 10, 24, 20, 0, 13, 22, 10, 23, 20, 
    24, 0, 10, 31, 0, 0, 5, 18, 26, 0, 19, 15, 8, 10, 18, 
    7, 12, 18, 26, 16, 0, 21, 3, 20, 0, 12, 14, 5, 5, 24, 
    7, 0, 13, 0, 7, 2, 11, 5, 13, 11, 0, 19, 2, 12, 17, 
    0, 0, 21, 0, 13, 11, 11, 14, 2, 9, 22, 17, 6, 10, 24, 
    0, 0, 18, 0, 34, 20, 0, 2, 21, 21, 12, 10, 0, 0, 4, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 5, 3, 1, 0, 0, 2, 
    2, 0, 0, 0, 26, 3, 4, 3, 6, 5, 4, 2, 0, 3, 3, 
    6, 0, 0, 0, 13, 4, 6, 2, 3, 1, 0, 0, 3, 0, 0, 
    6, 0, 0, 0, 5, 0, 2, 8, 5, 3, 4, 5, 2, 3, 15, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 0, 1, 41, 10, 0, 0, 0, 16, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 7, 9, 0, 0, 
    24, 19, 3, 0, 3, 0, 31, 9, 1, 0, 0, 0, 0, 0, 0, 
    26, 55, 9, 3, 94, 45, 3, 1, 0, 0, 19, 16, 8, 16, 0, 
    0, 1, 6, 0, 0, 0, 22, 14, 20, 22, 0, 0, 0, 8, 19, 
    0, 0, 0, 4, 0, 5, 4, 7, 10, 5, 0, 0, 0, 8, 14, 
    0, 15, 5, 24, 2, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 1, 0, 0, 6, 6, 0, 0, 0, 0, 0, 15, 
    0, 0, 5, 0, 8, 0, 0, 48, 0, 0, 0, 0, 20, 19, 0, 
    0, 0, 0, 32, 92, 71, 22, 0, 0, 0, 16, 35, 8, 0, 0, 
    0, 0, 14, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 20, 17, 0, 
    
    -- channel=42
    95, 97, 100, 100, 99, 93, 103, 107, 99, 82, 67, 70, 77, 87, 83, 
    98, 102, 105, 103, 100, 105, 95, 87, 57, 35, 31, 33, 43, 64, 81, 
    68, 68, 102, 103, 107, 86, 47, 23, 26, 43, 34, 24, 31, 36, 67, 
    25, 63, 95, 102, 89, 55, 53, 33, 26, 45, 34, 34, 12, 20, 55, 
    14, 72, 86, 85, 81, 77, 41, 27, 19, 36, 43, 33, 27, 18, 40, 
    17, 47, 78, 90, 42, 46, 51, 35, 23, 68, 45, 13, 28, 20, 22, 
    16, 47, 50, 70, 66, 64, 54, 37, 20, 67, 23, 21, 24, 27, 35, 
    31, 25, 41, 48, 66, 76, 33, 33, 20, 74, 33, 17, 24, 37, 49, 
    32, 35, 17, 38, 51, 26, 26, 36, 34, 52, 34, 6, 19, 49, 92, 
    34, 40, 12, 32, 25, 38, 33, 44, 43, 32, 8, 0, 36, 86, 81, 
    30, 40, 10, 60, 49, 43, 53, 21, 5, 0, 0, 0, 4, 0, 0, 
    0, 10, 23, 95, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 4, 4, 0, 0, 1, 5, 4, 0, 0, 0, 8, 10, 
    0, 0, 0, 5, 0, 0, 34, 6, 4, 0, 24, 23, 0, 0, 6, 
    18, 0, 0, 3, 0, 0, 25, 15, 0, 0, 28, 14, 43, 0, 0, 
    94, 0, 8, 0, 20, 0, 26, 28, 12, 0, 42, 9, 24, 27, 0, 
    70, 0, 43, 0, 19, 37, 49, 40, 25, 0, 25, 60, 7, 40, 0, 
    54, 0, 47, 14, 0, 0, 43, 40, 69, 0, 59, 50, 0, 24, 31, 
    49, 40, 0, 46, 0, 0, 12, 37, 61, 0, 61, 46, 3, 0, 34, 
    40, 29, 40, 31, 0, 0, 61, 1, 27, 0, 28, 50, 0, 0, 7, 
    44, 0, 91, 0, 39, 0, 17, 20, 0, 43, 0, 38, 0, 0, 0, 
    0, 0, 89, 0, 45, 6, 0, 36, 34, 0, 33, 0, 0, 0, 9, 
    0, 4, 81, 0, 98, 56, 0, 0, 47, 38, 10, 4, 0, 0, 14, 
    0, 0, 20, 0, 91, 27, 0, 0, 9, 5, 3, 2, 3, 6, 13, 
    32, 0, 0, 27, 80, 7, 13, 8, 10, 6, 2, 6, 7, 0, 0, 
    29, 7, 0, 44, 23, 3, 23, 12, 0, 3, 7, 1, 10, 0, 23, 
    41, 5, 4, 0, 18, 0, 0, 3, 2, 13, 24, 2, 0, 38, 51, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 32, 12, 7, 2, 16, 0, 
    0, 36, 0, 0, 0, 0, 0, 7, 19, 45, 0, 14, 4, 13, 21, 
    0, 29, 0, 0, 0, 0, 0, 0, 13, 45, 0, 0, 14, 0, 27, 
    6, 29, 0, 0, 35, 0, 0, 0, 0, 82, 0, 0, 21, 5, 6, 
    0, 14, 0, 0, 26, 22, 0, 0, 0, 74, 0, 0, 21, 22, 8, 
    8, 0, 0, 0, 13, 42, 0, 13, 0, 50, 0, 0, 28, 26, 0, 
    5, 25, 0, 25, 9, 13, 0, 8, 19, 0, 22, 0, 31, 12, 0, 
    18, 28, 0, 41, 0, 18, 14, 0, 22, 12, 0, 14, 31, 4, 0, 
    53, 20, 0, 72, 0, 7, 57, 22, 1, 5, 30, 43, 50, 42, 30, 
    95, 54, 3, 65, 0, 29, 51, 50, 48, 56, 64, 66, 68, 69, 63, 
    75, 92, 62, 31, 0, 56, 56, 58, 58, 65, 68, 71, 71, 70, 73, 
    69, 73, 115, 14, 41, 61, 53, 58, 63, 67, 74, 77, 71, 89, 84, 
    67, 76, 80, 46, 59, 74, 69, 60, 63, 62, 64, 70, 79, 67, 53, 
    
    -- channel=45
    0, 0, 0, 2, 3, 0, 0, 1, 5, 5, 4, 0, 0, 5, 7, 
    0, 0, 0, 3, 0, 0, 30, 7, 11, 0, 8, 12, 0, 0, 2, 
    20, 0, 0, 1, 0, 0, 35, 13, 1, 0, 18, 8, 29, 0, 0, 
    63, 0, 3, 0, 15, 0, 3, 28, 8, 0, 37, 9, 24, 27, 0, 
    61, 0, 41, 0, 0, 25, 37, 39, 19, 0, 5, 52, 0, 27, 0, 
    77, 0, 54, 34, 0, 22, 24, 26, 42, 0, 59, 58, 0, 16, 24, 
    78, 11, 10, 35, 0, 0, 0, 35, 42, 0, 61, 42, 0, 0, 26, 
    65, 2, 47, 10, 0, 0, 68, 9, 25, 0, 33, 44, 0, 0, 12, 
    51, 0, 104, 0, 47, 0, 17, 5, 0, 21, 0, 49, 0, 0, 0, 
    2, 0, 79, 0, 41, 27, 0, 0, 36, 10, 37, 0, 0, 0, 11, 
    0, 4, 68, 0, 68, 37, 0, 5, 55, 29, 0, 0, 0, 0, 9, 
    0, 0, 19, 0, 92, 57, 0, 2, 13, 0, 0, 0, 0, 0, 9, 
    23, 0, 0, 3, 104, 3, 6, 3, 3, 0, 0, 0, 0, 0, 0, 
    23, 1, 0, 27, 31, 0, 14, 5, 0, 0, 1, 0, 6, 0, 18, 
    33, 0, 4, 0, 16, 0, 0, 1, 0, 0, 14, 0, 0, 14, 41, 
    
    -- channel=46
    12, 9, 10, 12, 14, 10, 9, 15, 16, 13, 10, 7, 8, 9, 13, 
    14, 10, 10, 13, 12, 1, 9, 8, 15, 9, 4, 1, 1, 10, 13, 
    4, 14, 14, 14, 13, 4, 13, 13, 1, 0, 0, 0, 0, 2, 6, 
    10, 0, 12, 14, 10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    28, 29, 26, 30, 30, 23, 31, 33, 30, 35, 40, 32, 30, 30, 29, 
    29, 23, 23, 33, 21, 10, 45, 37, 48, 11, 23, 22, 20, 28, 31, 
    49, 34, 28, 32, 21, 18, 62, 32, 1, 0, 23, 28, 40, 12, 21, 
    74, 0, 34, 23, 38, 12, 18, 22, 21, 0, 61, 14, 39, 30, 0, 
    78, 0, 60, 0, 26, 8, 51, 38, 31, 0, 19, 46, 10, 40, 0, 
    51, 25, 74, 0, 0, 36, 54, 34, 51, 0, 67, 69, 4, 30, 23, 
    45, 50, 53, 59, 0, 0, 46, 52, 63, 0, 80, 39, 5, 0, 31, 
    36, 50, 39, 54, 0, 0, 98, 36, 51, 0, 55, 46, 0, 14, 37, 
    48, 15, 77, 8, 17, 21, 36, 12, 6, 31, 0, 73, 0, 4, 7, 
    34, 13, 94, 0, 51, 17, 0, 24, 12, 41, 76, 16, 0, 0, 44, 
    0, 17, 90, 0, 85, 13, 0, 61, 92, 43, 0, 0, 0, 23, 39, 
    0, 18, 49, 0, 113, 76, 10, 11, 25, 6, 5, 0, 0, 0, 7, 
    20, 0, 0, 32, 121, 7, 9, 6, 4, 0, 0, 0, 7, 6, 0, 
    26, 4, 0, 121, 40, 0, 13, 1, 0, 0, 0, 4, 11, 0, 28, 
    29, 0, 0, 30, 17, 0, 10, 12, 0, 0, 7, 0, 0, 8, 49, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 44, 2, 0, 0, 1, 21, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 
    9, 36, 0, 0, 1, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 37, 0, 0, 50, 21, 0, 0, 0, 8, 13, 6, 3, 8, 0, 
    0, 0, 0, 0, 0, 0, 14, 4, 13, 29, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 3, 0, 10, 4, 
    2, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 11, 1, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 4, 0, 0, 2, 26, 0, 0, 0, 0, 7, 8, 0, 
    0, 0, 0, 42, 74, 45, 0, 0, 0, 0, 26, 31, 7, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 0, 22, 5, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 3, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 0, 2, 0, 0, 0, 
    0, 33, 0, 0, 0, 0, 8, 0, 0, 15, 0, 0, 0, 0, 0, 
    1, 40, 0, 28, 37, 19, 0, 0, 0, 48, 13, 0, 6, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 90, 0, 0, 3, 0, 10, 
    6, 0, 0, 0, 11, 33, 0, 0, 0, 55, 0, 0, 7, 22, 0, 
    9, 0, 0, 0, 26, 18, 0, 0, 0, 22, 0, 0, 10, 0, 0, 
    2, 9, 0, 15, 0, 0, 0, 4, 18, 0, 0, 0, 0, 8, 0, 
    0, 7, 0, 40, 0, 0, 22, 18, 0, 0, 0, 0, 25, 0, 0, 
    20, 4, 0, 103, 32, 39, 20, 0, 0, 0, 31, 42, 23, 0, 0, 
    0, 0, 7, 59, 0, 0, 0, 0, 4, 12, 17, 18, 27, 24, 19, 
    14, 2, 37, 0, 0, 19, 14, 15, 18, 26, 33, 34, 16, 19, 42, 
    13, 22, 29, 0, 0, 22, 19, 19, 21, 24, 19, 14, 17, 45, 0, 
    8, 26, 15, 0, 0, 10, 4, 15, 32, 32, 19, 27, 63, 28, 4, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 2, 6, 4, 10, 5, 1, 0, 0, 
    7, 0, 0, 0, 0, 9, 10, 8, 0, 3, 19, 15, 10, 0, 0, 
    24, 0, 0, 0, 0, 1, 12, 7, 4, 3, 24, 9, 9, 0, 0, 
    40, 11, 0, 0, 38, 21, 33, 14, 7, 0, 23, 16, 5, 7, 0, 
    35, 32, 7, 0, 34, 34, 34, 20, 12, 0, 37, 24, 7, 10, 2, 
    34, 37, 11, 1, 7, 12, 44, 24, 26, 0, 39, 15, 3, 5, 6, 
    38, 46, 20, 11, 0, 26, 43, 21, 16, 0, 27, 18, 6, 7, 0, 
    49, 43, 31, 19, 2, 19, 17, 9, 10, 6, 10, 19, 0, 0, 0, 
    41, 37, 44, 15, 34, 8, 14, 27, 11, 17, 20, 3, 0, 0, 0, 
    31, 37, 45, 8, 51, 27, 25, 51, 43, 15, 7, 8, 16, 21, 21, 
    31, 39, 42, 24, 69, 40, 25, 24, 24, 16, 17, 19, 20, 20, 23, 
    23, 20, 25, 50, 58, 21, 21, 17, 15, 14, 18, 21, 26, 27, 27, 
    29, 22, 15, 65, 25, 20, 20, 18, 18, 20, 21, 24, 24, 21, 32, 
    29, 23, 16, 33, 15, 14, 20, 20, 18, 21, 22, 18, 17, 33, 32, 
    
    -- channel=51
    7, 7, 9, 11, 11, 7, 6, 4, 11, 11, 2, 0, 3, 5, 7, 
    8, 5, 9, 11, 11, 44, 17, 12, 0, 7, 27, 13, 0, 0, 8, 
    16, 0, 7, 7, 10, 1, 1, 0, 5, 31, 35, 25, 29, 0, 0, 
    30, 20, 6, 9, 22, 6, 38, 28, 24, 10, 29, 14, 8, 9, 0, 
    36, 56, 18, 13, 76, 61, 31, 24, 15, 4, 32, 31, 22, 21, 2, 
    31, 38, 13, 25, 0, 8, 44, 25, 32, 39, 46, 11, 15, 24, 19, 
    29, 53, 0, 12, 14, 37, 42, 35, 23, 43, 25, 22, 16, 23, 25, 
    43, 39, 30, 14, 24, 52, 37, 13, 7, 36, 27, 15, 12, 18, 2, 
    56, 45, 41, 20, 38, 0, 0, 33, 14, 22, 0, 0, 0, 6, 25, 
    41, 45, 41, 28, 23, 24, 14, 53, 34, 10, 6, 0, 12, 22, 10, 
    33, 41, 30, 53, 101, 73, 70, 37, 30, 21, 21, 43, 44, 30, 27, 
    20, 26, 34, 90, 46, 0, 1, 0, 15, 29, 35, 35, 37, 41, 37, 
    52, 20, 20, 79, 3, 33, 33, 29, 31, 36, 41, 48, 46, 39, 50, 
    44, 38, 26, 40, 29, 36, 38, 32, 33, 39, 42, 36, 37, 54, 46, 
    49, 40, 35, 0, 25, 23, 27, 34, 44, 47, 42, 34, 53, 71, 40, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 4, 0, 0, 
    0, 4, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 10, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    2, 1, 0, 0, 0, 0, 0, 0, 0, 4, 13, 14, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 15, 0, 0, 20, 18, 0, 
    6, 51, 0, 0, 1, 52, 16, 23, 1, 5, 0, 0, 0, 18, 14, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 42, 0, 5, 2, 0, 39, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 9, 
    0, 3, 0, 13, 109, 21, 0, 0, 0, 35, 0, 0, 8, 0, 0, 
    0, 0, 21, 0, 46, 7, 0, 0, 0, 39, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 18, 0, 27, 0, 32, 0, 0, 16, 4, 0, 
    0, 0, 0, 15, 0, 58, 11, 0, 4, 0, 44, 19, 29, 10, 0, 
    17, 3, 0, 17, 0, 0, 14, 0, 0, 31, 12, 13, 0, 0, 0, 
    45, 0, 0, 20, 0, 0, 0, 17, 0, 0, 0, 0, 0, 19, 13, 
    78, 50, 0, 0, 9, 64, 54, 52, 23, 9, 4, 7, 1, 0, 0, 
    0, 62, 51, 0, 27, 0, 0, 2, 1, 0, 0, 0, 0, 10, 0, 
    0, 0, 76, 31, 8, 1, 0, 0, 4, 0, 5, 17, 8, 1, 12, 
    0, 3, 11, 59, 15, 31, 25, 2, 0, 0, 0, 5, 0, 0, 0, 
    
    -- channel=54
    20, 20, 20, 23, 21, 19, 24, 21, 18, 19, 15, 12, 15, 17, 13, 
    19, 20, 21, 25, 20, 30, 35, 22, 12, 0, 14, 9, 1, 6, 17, 
    22, 3, 22, 21, 21, 21, 9, 0, 0, 11, 33, 18, 21, 0, 8, 
    32, 2, 27, 18, 25, 5, 32, 20, 14, 9, 34, 15, 4, 0, 0, 
    41, 47, 42, 7, 71, 64, 44, 20, 9, 0, 34, 32, 10, 11, 0, 
    43, 43, 46, 20, 3, 27, 46, 27, 24, 0, 61, 20, 9, 14, 7, 
    37, 57, 16, 24, 7, 22, 59, 40, 29, 16, 44, 19, 5, 9, 24, 
    48, 47, 33, 32, 14, 51, 60, 20, 17, 20, 31, 18, 3, 25, 12, 
    57, 50, 46, 14, 37, 6, 10, 18, 10, 31, 4, 9, 0, 1, 23, 
    45, 49, 50, 11, 41, 18, 6, 49, 34, 17, 13, 0, 4, 24, 23, 
    28, 49, 48, 15, 86, 60, 54, 52, 39, 10, 0, 8, 10, 13, 10, 
    19, 29, 48, 69, 82, 0, 0, 0, 0, 5, 9, 9, 11, 16, 15, 
    25, 13, 13, 88, 21, 10, 13, 8, 7, 8, 10, 17, 23, 15, 18, 
    19, 12, 13, 59, 13, 12, 14, 10, 8, 12, 14, 13, 10, 14, 36, 
    28, 10, 11, 4, 7, 1, 8, 11, 15, 18, 19, 8, 15, 43, 22, 
    
    -- channel=55
    26, 25, 25, 25, 25, 23, 31, 34, 27, 22, 21, 23, 21, 24, 23, 
    25, 31, 26, 27, 21, 0, 25, 28, 22, 0, 0, 2, 17, 20, 22, 
    26, 25, 31, 29, 30, 24, 13, 12, 0, 0, 0, 0, 0, 10, 15, 
    0, 0, 30, 26, 24, 1, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 13, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    54, 55, 55, 60, 61, 52, 59, 65, 65, 57, 47, 40, 46, 55, 57, 
    57, 58, 56, 63, 53, 44, 76, 61, 57, 17, 31, 29, 20, 31, 53, 
    58, 18, 60, 63, 60, 29, 63, 31, 14, 0, 22, 11, 40, 11, 24, 
    77, 0, 59, 56, 70, 26, 38, 32, 18, 0, 45, 19, 28, 28, 0, 
    57, 0, 76, 2, 35, 44, 46, 39, 24, 0, 24, 53, 9, 34, 6, 
    43, 0, 77, 68, 0, 24, 48, 35, 50, 0, 56, 47, 0, 22, 26, 
    38, 34, 30, 82, 0, 0, 26, 43, 47, 0, 56, 38, 6, 0, 29, 
    38, 16, 38, 50, 4, 0, 56, 15, 30, 0, 40, 40, 0, 8, 27, 
    36, 0, 72, 0, 52, 1, 27, 25, 0, 51, 2, 39, 0, 0, 38, 
    9, 0, 66, 0, 35, 19, 0, 30, 25, 19, 38, 4, 0, 19, 57, 
    0, 8, 59, 0, 77, 35, 0, 6, 40, 27, 0, 0, 0, 0, 14, 
    0, 0, 15, 0, 78, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 5, 1, 0, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 1, 40, 44, 30, 15, 5, 0, 
    4, 12, 0, 0, 0, 0, 18, 17, 23, 50, 30, 28, 19, 6, 7, 
    27, 51, 0, 0, 34, 28, 36, 20, 22, 26, 37, 16, 24, 9, 4, 
    46, 71, 0, 0, 78, 37, 40, 24, 16, 56, 47, 20, 32, 20, 5, 
    40, 70, 8, 0, 41, 41, 65, 32, 25, 74, 41, 23, 26, 31, 22, 
    50, 68, 17, 3, 20, 81, 50, 42, 25, 61, 39, 27, 33, 40, 12, 
    66, 82, 34, 46, 17, 41, 28, 30, 29, 17, 40, 17, 24, 18, 0, 
    78, 83, 45, 60, 39, 18, 31, 50, 36, 30, 15, 8, 20, 9, 0, 
    89, 73, 50, 86, 50, 41, 73, 76, 37, 16, 26, 33, 46, 44, 32, 
    109, 88, 60, 109, 93, 61, 68, 66, 58, 58, 66, 72, 78, 82, 79, 
    83, 95, 76, 110, 56, 66, 66, 65, 65, 69, 76, 81, 85, 83, 90, 
    88, 76, 103, 99, 58, 72, 66, 66, 69, 76, 84, 90, 82, 96, 103, 
    89, 85, 77, 86, 64, 74, 76, 69, 72, 78, 80, 79, 91, 103, 77, 
    
    -- channel=58
    8, 12, 4, 6, 7, 6, 9, 11, 9, 16, 22, 18, 9, 6, 6, 
    3, 7, 4, 9, 1, 0, 6, 19, 38, 1, 0, 4, 16, 10, 5, 
    34, 25, 7, 9, 6, 61, 37, 26, 0, 0, 0, 0, 4, 4, 8, 
    12, 0, 8, 6, 17, 0, 0, 0, 0, 0, 23, 11, 15, 0, 1, 
    0, 0, 10, 0, 0, 0, 22, 4, 18, 0, 0, 0, 0, 0, 0, 
    5, 12, 12, 18, 56, 19, 12, 0, 9, 0, 27, 25, 0, 0, 0, 
    0, 41, 21, 28, 15, 0, 33, 8, 18, 0, 32, 3, 0, 0, 0, 
    0, 24, 0, 11, 0, 0, 58, 36, 13, 0, 24, 18, 0, 9, 4, 
    7, 12, 11, 0, 0, 46, 20, 2, 0, 34, 19, 48, 6, 0, 0, 
    27, 12, 28, 0, 6, 0, 0, 0, 0, 31, 46, 1, 0, 0, 17, 
    17, 12, 41, 0, 0, 0, 0, 47, 23, 11, 0, 0, 0, 14, 13, 
    36, 26, 0, 0, 105, 62, 39, 34, 8, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 56, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 105, 6, 0, 0, 0, 0, 0, 0, 2, 0, 0, 27, 
    0, 0, 0, 55, 10, 3, 6, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 10, 6, 0, 0, 0, 12, 20, 7, 0, 0, 0, 14, 7, 6, 
    49, 23, 3, 0, 49, 43, 35, 36, 31, 28, 30, 35, 37, 40, 40, 
    49, 45, 16, 26, 43, 30, 31, 29, 29, 31, 35, 39, 44, 45, 41, 
    54, 42, 51, 31, 28, 32, 30, 31, 33, 37, 46, 50, 47, 51, 64, 
    54, 48, 45, 34, 33, 38, 39, 31, 30, 34, 42, 40, 36, 51, 47, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 
    9, 0, 0, 0, 0, 18, 6, 10, 0, 5, 21, 12, 3, 3, 0, 
    1, 0, 0, 0, 0, 0, 0, 9, 8, 18, 17, 19, 14, 6, 0, 
    6, 0, 0, 0, 0, 4, 23, 17, 19, 1, 8, 8, 7, 0, 7, 
    43, 24, 0, 19, 55, 34, 12, 9, 5, 0, 34, 24, 13, 7, 0, 
    35, 29, 1, 0, 17, 10, 27, 13, 13, 13, 28, 16, 11, 5, 6, 
    37, 24, 7, 0, 0, 28, 50, 33, 15, 21, 25, 22, 15, 20, 0, 
    42, 37, 35, 5, 13, 35, 16, 11, 0, 6, 29, 32, 20, 0, 0, 
    44, 41, 28, 16, 23, 23, 9, 0, 28, 29, 22, 7, 0, 0, 0, 
    28, 35, 34, 13, 0, 3, 28, 47, 27, 10, 5, 3, 18, 19, 17, 
    64, 43, 19, 23, 79, 65, 54, 53, 40, 33, 33, 38, 38, 39, 41, 
    41, 58, 32, 58, 72, 35, 36, 34, 32, 31, 33, 36, 42, 43, 37, 
    46, 38, 63, 63, 38, 36, 32, 35, 36, 39, 46, 49, 43, 45, 63, 
    48, 44, 43, 53, 40, 45, 44, 34, 31, 35, 41, 39, 29, 47, 39, 
    
    -- channel=61
    99, 105, 103, 105, 103, 99, 108, 116, 105, 85, 72, 76, 85, 92, 92, 
    101, 111, 109, 109, 106, 94, 95, 88, 72, 40, 26, 27, 41, 72, 88, 
    63, 79, 107, 111, 109, 96, 59, 38, 25, 27, 25, 23, 25, 32, 74, 
    39, 35, 102, 107, 89, 65, 50, 25, 18, 31, 34, 28, 20, 14, 54, 
    29, 39, 89, 85, 74, 50, 42, 23, 16, 18, 41, 30, 23, 21, 21, 
    4, 28, 85, 64, 43, 45, 48, 40, 24, 19, 32, 22, 24, 20, 16, 
    6, 26, 59, 92, 53, 38, 53, 33, 34, 24, 31, 19, 15, 20, 28, 
    7, 32, 20, 65, 55, 48, 29, 28, 33, 42, 34, 22, 17, 29, 57, 
    11, 17, 1, 31, 27, 34, 38, 27, 29, 48, 35, 20, 16, 50, 81, 
    24, 20, 17, 13, 27, 14, 27, 43, 13, 33, 19, 10, 24, 70, 83, 
    14, 22, 20, 15, 31, 14, 5, 13, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 34, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    1, 0, 0, 0, 2, 0, 5, 0, 0, 5, 0, 0, 1, 3, 0, 
    0, 4, 0, 0, 0, 0, 4, 2, 26, 0, 0, 3, 0, 10, 0, 
    0, 11, 0, 0, 0, 19, 0, 15, 0, 0, 0, 0, 0, 4, 0, 
    12, 0, 11, 53, 0, 22, 0, 3, 0, 52, 0, 0, 0, 0, 20, 
    65, 0, 26, 19, 0, 45, 0, 0, 0, 21, 0, 16, 0, 0, 15, 
    98, 0, 25, 0, 0, 21, 0, 10, 0, 0, 0, 4, 2, 0, 0, 
    73, 0, 49, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    24, 0, 41, 0, 37, 0, 0, 0, 15, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 56, 36, 0, 20, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 24, 0, 10, 0, 0, 6, 0, 9, 10, 2, 0, 5, 
    0, 3, 17, 0, 0, 28, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 76, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 36, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 4, 7, 0, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 13, 15, 15, 2, 0, 
    0, 7, 0, 0, 0, 6, 22, 41, 7, 1, 0, 0, 0, 2, 0, 
    2, 13, 0, 2, 0, 29, 0, 0, 0, 0, 0, 0, 8, 0, 5, 
    6, 0, 0, 13, 0, 0, 0, 0, 0, 25, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 2, 0, 0, 0, 8, 0, 0, 0, 
    10, 0, 10, 0, 0, 0, 0, 1, 0, 0, 7, 5, 11, 0, 0, 
    0, 9, 5, 12, 0, 0, 0, 0, 0, 0, 3, 10, 0, 0, 3, 
    0, 0, 0, 0, 0, 25, 22, 0, 4, 33, 0, 10, 6, 1, 0, 
    0, 0, 0, 24, 0, 0, 30, 0, 0, 0, 5, 10, 0, 0, 0, 
    4, 0, 11, 0, 0, 0, 0, 0, 0, 28, 15, 0, 0, 26, 28, 
    0, 5, 0, 0, 0, 43, 35, 34, 13, 4, 0, 4, 3, 1, 0, 
    0, 0, 21, 0, 38, 1, 0, 2, 4, 0, 4, 0, 0, 0, 7, 
    1, 3, 0, 0, 3, 3, 4, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 2, 30, 7, 0, 0, 0, 0, 3, 0, 7, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
