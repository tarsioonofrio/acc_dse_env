library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 8, 11, 8, 7, 6, 3, 9, 0, 0, 0, 0, 8, 5, 
    10, 14, 12, 9, 11, 60, 33, 0, 0, 0, 26, 6, 0, 0, 6, 
    0, 0, 6, 6, 7, 0, 0, 0, 5, 18, 21, 9, 15, 0, 0, 
    37, 31, 10, 8, 14, 0, 48, 25, 3, 0, 0, 0, 0, 0, 0, 
    37, 79, 26, 19, 118, 100, 16, 12, 0, 0, 37, 37, 11, 16, 0, 
    6, 0, 19, 0, 0, 0, 30, 29, 29, 40, 14, 0, 0, 10, 32, 
    27, 0, 0, 4, 0, 22, 0, 17, 10, 11, 0, 12, 0, 14, 28, 
    35, 7, 39, 19, 20, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 7, 21, 0, 40, 0, 0, 17, 2, 0, 0, 0, 0, 0, 33, 
    0, 1, 10, 1, 17, 5, 0, 61, 31, 0, 0, 0, 16, 29, 2, 
    0, 8, 0, 59, 130, 125, 37, 0, 0, 0, 24, 48, 13, 0, 0, 
    0, 0, 17, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 2, 0, 0, 0, 0, 0, 1, 5, 16, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 16, 3, 0, 31, 35, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 5, 0, 0, 10, 6, 0, 0, 0, 0, 11, 11, 0, 0, 0, 
    34, 7, 0, 0, 0, 0, 3, 0, 1, 0, 15, 0, 0, 0, 0, 
    29, 7, 0, 0, 0, 0, 28, 6, 2, 0, 9, 1, 0, 0, 0, 
    33, 20, 29, 0, 0, 6, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    27, 25, 26, 0, 12, 0, 0, 0, 2, 7, 13, 0, 0, 0, 0, 
    8, 13, 27, 0, 3, 3, 20, 41, 41, 0, 6, 15, 24, 8, 9, 
    66, 39, 25, 0, 71, 75, 50, 49, 57, 50, 56, 60, 64, 65, 69, 
    82, 57, 26, 22, 86, 56, 58, 54, 56, 58, 64, 65, 74, 78, 71, 
    92, 68, 54, 61, 64, 57, 56, 55, 60, 64, 76, 82, 79, 79, 100, 
    89, 80, 66, 58, 62, 66, 72, 62, 56, 59, 71, 70, 60, 81, 89, 
    
    -- channel=2
    82, 81, 83, 77, 78, 79, 87, 89, 78, 71, 69, 76, 71, 67, 62, 
    79, 85, 90, 80, 87, 50, 55, 72, 69, 38, 0, 14, 54, 74, 63, 
    51, 114, 87, 82, 92, 99, 28, 27, 25, 44, 0, 0, 0, 53, 71, 
    0, 75, 74, 89, 53, 64, 2, 0, 2, 86, 0, 21, 0, 0, 98, 
    0, 26, 41, 120, 0, 23, 0, 0, 0, 87, 0, 0, 1, 0, 58, 
    0, 16, 27, 84, 94, 45, 0, 0, 0, 124, 0, 0, 21, 0, 0, 
    0, 0, 57, 21, 98, 56, 9, 0, 0, 113, 0, 0, 9, 8, 0, 
    0, 0, 2, 10, 78, 78, 0, 23, 0, 90, 0, 0, 27, 27, 25, 
    0, 3, 0, 30, 15, 59, 1, 0, 33, 23, 38, 0, 36, 39, 60, 
    0, 7, 0, 45, 0, 35, 44, 0, 8, 29, 0, 6, 38, 73, 61, 
    43, 9, 0, 84, 0, 0, 44, 1, 0, 0, 0, 0, 0, 8, 0, 
    45, 33, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    19, 21, 29, 27, 26, 20, 28, 28, 21, 6, 4, 11, 24, 21, 17, 
    28, 27, 28, 27, 29, 60, 24, 13, 0, 0, 6, 0, 0, 7, 21, 
    0, 18, 27, 27, 21, 0, 0, 0, 0, 11, 0, 10, 1, 0, 19, 
    0, 21, 21, 26, 17, 16, 12, 3, 1, 0, 12, 0, 0, 0, 0, 
    22, 31, 32, 28, 82, 57, 0, 0, 0, 7, 0, 4, 0, 5, 0, 
    0, 3, 37, 0, 0, 0, 25, 0, 0, 17, 6, 0, 0, 4, 11, 
    1, 0, 0, 15, 0, 20, 0, 27, 0, 3, 0, 0, 0, 0, 4, 
    6, 4, 6, 20, 4, 0, 11, 0, 0, 0, 0, 0, 0, 0, 15, 
    7, 0, 0, 5, 4, 0, 0, 0, 6, 0, 0, 0, 0, 6, 25, 
    0, 0, 0, 0, 0, 14, 17, 18, 0, 0, 0, 0, 10, 32, 17, 
    0, 0, 0, 18, 100, 20, 23, 0, 10, 2, 0, 7, 0, 0, 0, 
    0, 0, 17, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    90, 93, 99, 96, 95, 93, 102, 105, 96, 69, 57, 68, 81, 85, 81, 
    98, 105, 102, 98, 99, 116, 89, 79, 52, 50, 37, 34, 42, 64, 78, 
    44, 68, 101, 103, 103, 62, 55, 33, 32, 43, 16, 17, 15, 25, 70, 
    16, 67, 94, 101, 85, 71, 52, 20, 16, 26, 30, 22, 13, 9, 52, 
    15, 53, 78, 86, 81, 69, 38, 26, 7, 54, 44, 25, 23, 11, 25, 
    5, 33, 78, 86, 43, 52, 58, 30, 15, 67, 25, 10, 16, 12, 21, 
    20, 23, 54, 75, 49, 75, 28, 40, 7, 53, 20, 20, 23, 28, 22, 
    33, 26, 26, 59, 52, 36, 7, 19, 20, 53, 31, 14, 16, 21, 47, 
    26, 25, 10, 38, 50, 25, 36, 34, 29, 54, 21, 0, 19, 50, 80, 
    31, 26, 6, 39, 7, 25, 47, 43, 20, 6, 0, 1, 28, 77, 74, 
    32, 34, 7, 66, 52, 18, 13, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 4, 18, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 2, 6, 0, 2, 3, 4, 0, 0, 0, 0, 8, 9, 
    2, 0, 0, 4, 0, 0, 38, 2, 5, 0, 21, 20, 0, 0, 5, 
    11, 0, 0, 3, 0, 0, 36, 12, 0, 0, 18, 14, 42, 0, 0, 
    83, 0, 7, 0, 22, 0, 12, 27, 12, 0, 50, 1, 26, 25, 0, 
    71, 0, 53, 0, 0, 46, 48, 45, 22, 0, 13, 60, 0, 37, 0, 
    66, 0, 63, 26, 0, 4, 42, 34, 65, 0, 66, 58, 0, 22, 33, 
    67, 31, 0, 44, 0, 0, 0, 48, 49, 0, 67, 46, 2, 0, 30, 
    56, 21, 51, 26, 0, 0, 80, 2, 22, 0, 33, 48, 0, 0, 16, 
    52, 0, 111, 0, 48, 0, 14, 11, 0, 52, 0, 48, 0, 0, 0, 
    0, 0, 93, 0, 25, 24, 0, 18, 35, 0, 42, 0, 0, 0, 10, 
    0, 1, 84, 0, 112, 38, 0, 0, 53, 48, 0, 0, 0, 0, 11, 
    0, 0, 17, 0, 88, 38, 0, 0, 1, 0, 0, 0, 0, 0, 4, 
    28, 0, 0, 9, 93, 1, 4, 2, 2, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 39, 22, 0, 18, 1, 0, 0, 0, 0, 5, 0, 14, 
    38, 0, 4, 0, 11, 0, 0, 0, 0, 5, 14, 0, 0, 24, 46, 
    
    -- channel=6
    56, 66, 58, 60, 57, 63, 58, 56, 58, 64, 63, 59, 56, 47, 44, 
    53, 57, 59, 62, 61, 106, 58, 68, 68, 69, 67, 47, 47, 52, 48, 
    72, 65, 57, 59, 58, 113, 85, 46, 36, 98, 106, 88, 65, 30, 58, 
    66, 36, 55, 63, 73, 67, 92, 64, 68, 95, 119, 80, 72, 31, 43, 
    122, 111, 66, 77, 163, 108, 124, 79, 65, 64, 116, 75, 69, 49, 13, 
    128, 170, 80, 75, 197, 149, 158, 89, 65, 100, 153, 91, 76, 70, 32, 
    121, 179, 78, 67, 110, 142, 190, 125, 91, 136, 145, 80, 67, 81, 63, 
    151, 180, 73, 79, 75, 184, 163, 125, 87, 121, 146, 84, 75, 88, 63, 
    191, 194, 116, 131, 78, 113, 98, 97, 81, 85, 98, 78, 49, 65, 59, 
    208, 192, 150, 126, 110, 69, 104, 142, 75, 107, 81, 34, 51, 71, 73, 
    200, 181, 151, 159, 200, 105, 164, 199, 128, 67, 47, 65, 87, 107, 99, 
    160, 201, 160, 232, 251, 142, 116, 112, 103, 94, 101, 107, 115, 118, 117, 
    116, 135, 168, 259, 156, 105, 101, 96, 94, 96, 107, 115, 127, 130, 134, 
    126, 108, 139, 253, 120, 108, 104, 95, 102, 109, 118, 127, 122, 130, 150, 
    128, 118, 113, 134, 94, 102, 115, 108, 111, 118, 111, 107, 130, 155, 115, 
    
    -- channel=7
    62, 71, 67, 69, 69, 63, 69, 78, 73, 56, 48, 48, 56, 60, 65, 
    66, 71, 67, 73, 64, 70, 60, 63, 58, 24, 14, 11, 17, 37, 57, 
    55, 41, 70, 77, 68, 59, 71, 28, 1, 0, 7, 9, 17, 0, 41, 
    48, 0, 56, 68, 72, 36, 29, 10, 8, 0, 47, 9, 28, 8, 0, 
    29, 0, 56, 6, 34, 12, 40, 30, 19, 0, 14, 26, 7, 20, 0, 
    2, 0, 63, 65, 16, 30, 58, 23, 38, 0, 38, 37, 0, 13, 4, 
    0, 28, 23, 94, 3, 10, 26, 36, 34, 0, 42, 21, 0, 0, 10, 
    5, 24, 0, 44, 0, 0, 56, 22, 32, 0, 45, 28, 0, 5, 37, 
    18, 0, 32, 0, 22, 15, 28, 21, 0, 43, 1, 45, 1, 16, 35, 
    26, 0, 49, 0, 1, 5, 0, 22, 0, 22, 41, 0, 0, 18, 52, 
    0, 0, 46, 0, 47, 0, 0, 8, 18, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 53, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 3, 6, 7, 3, 1, 2, 7, 0, 0, 0, 0, 8, 12, 
    6, 9, 5, 6, 4, 44, 16, 0, 0, 4, 35, 18, 0, 0, 10, 
    0, 0, 4, 5, 4, 0, 0, 0, 9, 23, 23, 17, 37, 0, 0, 
    62, 21, 6, 4, 15, 1, 44, 23, 19, 0, 16, 2, 10, 16, 0, 
    39, 55, 11, 0, 69, 44, 19, 20, 14, 0, 33, 36, 26, 38, 0, 
    0, 0, 0, 0, 0, 0, 36, 33, 57, 1, 6, 0, 8, 26, 37, 
    0, 32, 0, 23, 0, 0, 4, 16, 34, 4, 4, 23, 17, 22, 28, 
    0, 27, 11, 27, 15, 0, 0, 0, 4, 2, 0, 17, 1, 0, 0, 
    4, 0, 14, 0, 13, 0, 0, 33, 1, 31, 0, 0, 0, 6, 20, 
    0, 0, 28, 15, 5, 0, 0, 65, 11, 0, 0, 5, 21, 21, 5, 
    0, 0, 20, 8, 96, 66, 3, 0, 0, 29, 37, 46, 27, 0, 0, 
    0, 0, 6, 27, 0, 0, 0, 0, 0, 12, 16, 17, 22, 23, 20, 
    29, 0, 0, 10, 0, 17, 20, 18, 23, 26, 29, 31, 18, 10, 28, 
    22, 18, 0, 0, 2, 19, 30, 22, 17, 21, 19, 8, 16, 23, 3, 
    28, 20, 10, 0, 9, 0, 0, 12, 30, 36, 30, 19, 36, 51, 31, 
    
    -- channel=9
    74, 72, 73, 75, 74, 66, 75, 81, 76, 64, 57, 60, 63, 65, 71, 
    73, 71, 72, 75, 74, 63, 59, 61, 54, 44, 25, 30, 44, 60, 69, 
    56, 72, 77, 78, 78, 70, 59, 46, 32, 24, 20, 26, 21, 35, 61, 
    31, 35, 71, 74, 65, 58, 34, 24, 27, 20, 35, 24, 35, 25, 44, 
    17, 8, 59, 49, 24, 7, 26, 29, 30, 21, 23, 21, 29, 27, 24, 
    7, 20, 58, 50, 38, 24, 32, 27, 30, 9, 24, 33, 26, 27, 19, 
    6, 13, 47, 75, 31, 28, 24, 31, 28, 10, 27, 26, 24, 24, 26, 
    1, 20, 6, 54, 26, 15, 39, 33, 40, 30, 33, 30, 21, 29, 52, 
    5, 6, 13, 21, 31, 31, 36, 31, 25, 39, 34, 44, 32, 44, 52, 
    27, 10, 21, 5, 14, 24, 27, 20, 12, 39, 38, 24, 16, 43, 59, 
    18, 11, 24, 5, 2, 0, 0, 15, 13, 21, 8, 0, 0, 11, 17, 
    0, 13, 11, 0, 12, 21, 6, 7, 3, 1, 0, 0, 0, 0, 0, 
    0, 0, 8, 12, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    29, 42, 38, 40, 34, 40, 38, 39, 32, 16, 6, 15, 29, 25, 21, 
    37, 45, 41, 40, 44, 115, 23, 19, 0, 25, 25, 0, 0, 13, 24, 
    0, 15, 37, 41, 36, 47, 10, 0, 0, 75, 57, 49, 14, 0, 34, 
    15, 35, 33, 42, 31, 34, 65, 16, 22, 50, 62, 20, 16, 0, 15, 
    71, 111, 28, 56, 166, 77, 65, 27, 5, 44, 83, 26, 35, 14, 0, 
    29, 120, 41, 1, 115, 69, 119, 51, 26, 106, 68, 15, 33, 28, 4, 
    45, 105, 18, 30, 71, 107, 117, 71, 39, 114, 63, 25, 23, 51, 29, 
    71, 130, 12, 46, 47, 132, 55, 42, 39, 92, 75, 22, 30, 38, 40, 
    107, 123, 25, 91, 16, 26, 43, 52, 52, 24, 29, 0, 2, 52, 46, 
    131, 121, 74, 88, 42, 1, 67, 121, 13, 21, 0, 0, 37, 60, 31, 
    139, 109, 68, 168, 181, 71, 93, 89, 36, 0, 6, 27, 15, 2, 0, 
    39, 107, 106, 202, 73, 0, 8, 4, 12, 12, 25, 29, 45, 47, 41, 
    30, 29, 104, 147, 8, 36, 29, 27, 27, 32, 44, 50, 47, 44, 73, 
    39, 28, 36, 114, 31, 41, 38, 27, 32, 39, 36, 39, 38, 58, 33, 
    42, 43, 22, 29, 5, 17, 29, 39, 52, 59, 38, 40, 89, 84, 32, 
    
    -- channel=11
    0, 2, 0, 0, 0, 0, 0, 0, 0, 9, 23, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 45, 0, 0, 0, 11, 4, 0, 
    44, 30, 0, 0, 0, 65, 26, 12, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 17, 14, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 6, 
    3, 0, 0, 44, 73, 11, 0, 0, 0, 0, 14, 18, 0, 0, 0, 
    0, 20, 6, 9, 23, 0, 15, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 61, 41, 10, 4, 15, 6, 0, 21, 0, 
    0, 0, 1, 0, 0, 54, 1, 0, 0, 8, 34, 62, 24, 0, 0, 
    15, 0, 0, 0, 0, 4, 0, 0, 0, 53, 57, 3, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 47, 18, 0, 0, 0, 0, 0, 2, 
    63, 23, 0, 0, 113, 76, 46, 39, 14, 4, 0, 2, 0, 0, 0, 
    0, 45, 0, 45, 73, 0, 1, 0, 0, 0, 0, 0, 4, 5, 0, 
    2, 0, 26, 101, 16, 0, 0, 0, 0, 0, 7, 16, 4, 0, 59, 
    6, 0, 12, 57, 27, 26, 28, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 32, 24, 22, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 11, 20, 15, 14, 15, 19, 19, 0, 
    32, 28, 0, 0, 0, 0, 15, 16, 25, 6, 18, 16, 19, 21, 1, 
    39, 40, 0, 0, 22, 1, 16, 14, 26, 13, 23, 19, 21, 21, 20, 
    34, 52, 0, 0, 0, 0, 22, 12, 26, 26, 28, 25, 24, 24, 19, 
    37, 45, 19, 0, 0, 19, 23, 21, 15, 8, 19, 26, 24, 19, 0, 
    49, 56, 41, 24, 0, 13, 11, 18, 15, 0, 14, 15, 17, 0, 0, 
    37, 49, 48, 43, 35, 5, 8, 30, 27, 4, 18, 23, 23, 0, 0, 
    52, 40, 48, 36, 46, 46, 47, 51, 46, 35, 54, 62, 70, 61, 54, 
    106, 64, 42, 41, 69, 79, 86, 86, 90, 88, 98, 102, 108, 108, 107, 
    125, 97, 46, 60, 72, 94, 96, 93, 93, 99, 108, 112, 113, 111, 119, 
    130, 117, 86, 81, 79, 97, 98, 97, 97, 105, 114, 120, 119, 127, 133, 
    126, 123, 111, 99, 92, 99, 98, 95, 97, 106, 112, 109, 111, 131, 126, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 19, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 36, 34, 27, 15, 0, 0, 
    12, 23, 0, 0, 0, 0, 23, 24, 19, 15, 14, 7, 5, 3, 0, 
    35, 56, 0, 0, 56, 54, 19, 20, 8, 23, 33, 23, 24, 17, 0, 
    38, 32, 0, 0, 0, 0, 26, 24, 24, 60, 27, 4, 18, 23, 23, 
    48, 30, 0, 0, 0, 33, 18, 26, 14, 50, 14, 23, 23, 30, 24, 
    53, 41, 30, 0, 13, 36, 11, 0, 3, 30, 10, 13, 19, 14, 0, 
    55, 50, 37, 17, 28, 0, 0, 26, 20, 2, 0, 0, 3, 0, 0, 
    36, 49, 31, 44, 20, 22, 26, 49, 37, 0, 0, 1, 18, 2, 0, 
    38, 46, 23, 92, 91, 82, 62, 23, 20, 26, 48, 65, 57, 27, 20, 
    41, 34, 43, 88, 10, 2, 25, 26, 38, 54, 63, 67, 76, 78, 76, 
    87, 47, 50, 51, 12, 64, 62, 61, 64, 73, 81, 90, 78, 75, 99, 
    85, 74, 61, 12, 48, 71, 70, 65, 66, 76, 79, 73, 76, 103, 70, 
    88, 80, 64, 24, 51, 55, 54, 64, 78, 85, 79, 78, 105, 110, 74, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 24, 22, 10, 0, 0, 15, 0, 10, 0, 0, 
    58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 4, 14, 0, 0, 
    22, 0, 0, 0, 0, 0, 44, 19, 21, 0, 2, 17, 0, 0, 0, 
    32, 8, 0, 13, 22, 0, 39, 6, 38, 0, 58, 35, 0, 0, 0, 
    0, 77, 0, 21, 0, 0, 47, 17, 41, 0, 58, 20, 0, 0, 0, 
    14, 43, 0, 2, 0, 0, 82, 25, 15, 0, 34, 37, 0, 0, 0, 
    46, 25, 62, 0, 6, 12, 14, 15, 0, 33, 16, 46, 0, 0, 0, 
    40, 22, 79, 0, 30, 0, 0, 21, 8, 15, 40, 0, 0, 0, 0, 
    4, 22, 87, 0, 27, 0, 0, 54, 42, 16, 0, 0, 0, 16, 30, 
    24, 7, 0, 0, 183, 84, 50, 45, 27, 13, 9, 14, 12, 13, 21, 
    30, 7, 0, 114, 117, 10, 16, 10, 9, 2, 1, 5, 20, 16, 0, 
    36, 12, 0, 154, 31, 5, 16, 11, 5, 9, 23, 27, 23, 4, 71, 
    45, 17, 20, 62, 31, 13, 14, 4, 0, 11, 26, 3, 0, 46, 44, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 26, 27, 12, 0, 0, 
    12, 0, 0, 0, 0, 0, 7, 16, 14, 0, 21, 3, 13, 0, 0, 
    55, 23, 0, 0, 38, 33, 22, 19, 5, 12, 26, 20, 14, 15, 0, 
    49, 29, 0, 0, 0, 19, 34, 20, 18, 18, 30, 18, 10, 21, 17, 
    60, 31, 0, 0, 0, 20, 20, 29, 20, 17, 32, 22, 15, 22, 13, 
    61, 52, 21, 0, 0, 13, 25, 7, 10, 0, 27, 16, 12, 5, 0, 
    68, 55, 45, 19, 5, 0, 7, 15, 12, 0, 0, 0, 0, 0, 0, 
    48, 51, 51, 38, 22, 11, 25, 41, 15, 0, 4, 6, 7, 0, 0, 
    38, 45, 45, 55, 101, 58, 45, 40, 41, 31, 39, 55, 46, 25, 24, 
    36, 49, 56, 52, 43, 45, 41, 43, 55, 59, 66, 71, 81, 80, 81, 
    89, 39, 54, 41, 59, 70, 68, 66, 67, 73, 83, 86, 81, 85, 99, 
    96, 79, 39, 47, 64, 72, 76, 67, 72, 78, 83, 80, 88, 97, 80, 
    97, 89, 72, 40, 57, 58, 63, 71, 79, 86, 82, 83, 100, 107, 93, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 22, 0, 0, 0, 0, 0, 
    0, 72, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 12, 0, 65, 13, 0, 0, 0, 0, 95, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 27, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 28, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 20, 0, 0, 42, 0, 0, 0, 0, 0, 31, 0, 0, 
    0, 0, 0, 129, 3, 0, 0, 0, 0, 0, 35, 39, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 0, 
    
    -- channel=17
    1, 0, 0, 0, 5, 3, 0, 3, 11, 10, 8, 4, 3, 2, 5, 
    5, 3, 0, 0, 0, 0, 18, 9, 23, 30, 31, 36, 29, 6, 1, 
    5, 1, 6, 3, 8, 18, 31, 55, 21, 4, 0, 0, 8, 13, 0, 
    25, 14, 9, 10, 19, 34, 8, 0, 0, 0, 0, 5, 7, 0, 0, 
    6, 0, 5, 9, 0, 6, 7, 1, 2, 18, 14, 5, 0, 0, 16, 
    21, 0, 0, 39, 0, 2, 0, 7, 6, 0, 0, 8, 0, 0, 2, 
    16, 6, 10, 9, 5, 7, 0, 5, 0, 0, 15, 15, 18, 4, 0, 
    15, 1, 22, 24, 9, 0, 0, 2, 0, 0, 3, 19, 0, 0, 0, 
    9, 5, 18, 0, 25, 31, 25, 15, 0, 68, 5, 1, 5, 0, 0, 
    0, 0, 0, 33, 0, 1, 18, 3, 8, 0, 1, 11, 0, 0, 15, 
    12, 14, 20, 0, 0, 0, 0, 0, 0, 40, 27, 5, 17, 48, 58, 
    7, 0, 0, 0, 37, 46, 53, 48, 17, 13, 3, 11, 7, 7, 7, 
    7, 10, 4, 10, 27, 2, 1, 6, 8, 5, 6, 1, 0, 4, 2, 
    1, 9, 2, 0, 4, 5, 10, 4, 0, 0, 8, 1, 12, 0, 0, 
    0, 0, 23, 26, 18, 1, 0, 0, 0, 7, 5, 4, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 14, 0, 11, 41, 21, 0, 0, 0, 7, 10, 0, 0, 0, 0, 
    15, 1, 0, 0, 6, 9, 9, 0, 0, 18, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 26, 20, 0, 0, 21, 0, 0, 0, 0, 0, 
    25, 22, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 32, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    17, 26, 0, 30, 0, 0, 11, 10, 0, 0, 0, 0, 0, 0, 0, 
    22, 25, 4, 51, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 32, 46, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 42, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    11, 7, 9, 10, 10, 6, 12, 11, 7, 7, 6, 6, 7, 7, 7, 
    13, 8, 8, 11, 10, 11, 7, 4, 3, 1, 5, 2, 2, 11, 10, 
    1, 16, 13, 10, 12, 0, 2, 0, 0, 4, 0, 0, 6, 7, 13, 
    0, 17, 18, 9, 4, 2, 4, 0, 7, 4, 2, 0, 0, 5, 12, 
    0, 18, 14, 0, 6, 0, 0, 0, 1, 3, 0, 0, 1, 4, 1, 
    0, 11, 13, 0, 0, 0, 2, 0, 3, 7, 0, 0, 1, 1, 2, 
    0, 12, 12, 4, 0, 2, 3, 3, 0, 10, 0, 0, 2, 5, 6, 
    0, 0, 2, 13, 5, 4, 0, 1, 2, 5, 4, 0, 0, 6, 6, 
    0, 0, 0, 10, 4, 0, 0, 2, 7, 8, 0, 0, 0, 10, 13, 
    0, 0, 2, 3, 0, 0, 0, 8, 0, 0, 1, 0, 11, 17, 10, 
    11, 0, 0, 0, 14, 2, 6, 0, 0, 0, 0, 5, 2, 11, 10, 
    5, 6, 3, 14, 0, 0, 0, 0, 0, 2, 6, 3, 3, 5, 3, 
    11, 4, 3, 8, 0, 1, 1, 2, 3, 4, 4, 4, 5, 2, 4, 
    6, 7, 0, 8, 2, 1, 3, 1, 1, 1, 3, 4, 5, 3, 10, 
    5, 3, 9, 0, 5, 3, 4, 4, 3, 3, 3, 3, 6, 5, 7, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 1, 4, 
    0, 0, 0, 0, 0, 0, 32, 6, 17, 0, 18, 17, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 43, 19, 0, 0, 32, 15, 54, 0, 0, 
    123, 0, 0, 0, 18, 0, 17, 30, 12, 0, 60, 11, 40, 38, 0, 
    98, 0, 45, 0, 0, 11, 62, 52, 35, 0, 18, 74, 1, 53, 0, 
    71, 0, 58, 0, 0, 2, 54, 46, 85, 0, 78, 77, 0, 28, 31, 
    59, 54, 5, 58, 0, 0, 25, 42, 89, 0, 91, 57, 0, 0, 38, 
    46, 39, 41, 34, 0, 0, 92, 13, 44, 0, 47, 68, 0, 0, 8, 
    54, 0, 120, 0, 27, 0, 27, 17, 0, 32, 0, 70, 0, 0, 0, 
    1, 0, 130, 0, 70, 0, 0, 32, 27, 15, 65, 6, 0, 0, 11, 
    0, 0, 117, 0, 114, 52, 0, 25, 89, 45, 1, 0, 0, 0, 19, 
    0, 0, 30, 0, 156, 71, 2, 6, 25, 6, 4, 0, 0, 4, 18, 
    38, 0, 0, 32, 144, 9, 18, 10, 12, 3, 0, 0, 10, 2, 0, 
    45, 7, 0, 101, 42, 0, 27, 14, 1, 1, 6, 6, 15, 0, 41, 
    56, 7, 2, 14, 26, 0, 0, 7, 0, 7, 29, 0, 0, 39, 79, 
    
    -- channel=21
    3, 0, 6, 0, 0, 5, 0, 0, 0, 0, 0, 6, 2, 0, 0, 
    3, 3, 9, 0, 12, 14, 0, 0, 0, 19, 0, 0, 9, 11, 0, 
    0, 28, 4, 0, 10, 0, 0, 0, 23, 59, 0, 0, 0, 21, 12, 
    0, 85, 0, 11, 0, 27, 0, 0, 0, 83, 0, 0, 0, 0, 59, 
    0, 40, 0, 95, 0, 19, 0, 0, 0, 115, 0, 0, 0, 0, 42, 
    0, 1, 0, 35, 44, 1, 0, 0, 0, 198, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 66, 67, 0, 0, 0, 148, 0, 0, 10, 21, 0, 
    0, 0, 0, 0, 70, 75, 0, 0, 0, 89, 0, 0, 29, 2, 0, 
    0, 2, 0, 25, 7, 3, 0, 0, 31, 0, 14, 0, 22, 15, 17, 
    0, 5, 0, 66, 0, 25, 46, 0, 3, 0, 0, 0, 42, 39, 0, 
    51, 5, 0, 172, 0, 0, 71, 0, 0, 0, 15, 34, 32, 17, 0, 
    61, 32, 0, 118, 0, 0, 0, 0, 0, 6, 7, 10, 8, 8, 0, 
    0, 67, 102, 0, 0, 0, 0, 0, 0, 10, 14, 15, 3, 9, 18, 
    0, 8, 152, 0, 0, 10, 0, 1, 10, 10, 7, 2, 0, 37, 0, 
    0, 4, 18, 0, 0, 17, 4, 0, 17, 3, 0, 9, 52, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    50, 57, 55, 57, 57, 51, 59, 65, 64, 55, 50, 48, 53, 54, 56, 
    59, 60, 55, 61, 53, 51, 63, 61, 58, 25, 24, 19, 19, 42, 53, 
    50, 42, 58, 63, 53, 22, 63, 26, 11, 0, 5, 15, 29, 7, 40, 
    55, 0, 56, 58, 64, 32, 29, 18, 13, 0, 41, 8, 28, 22, 5, 
    50, 0, 64, 14, 42, 13, 31, 28, 17, 0, 15, 35, 9, 35, 0, 
    5, 0, 70, 21, 0, 22, 47, 27, 39, 0, 30, 40, 0, 21, 22, 
    9, 17, 40, 81, 0, 0, 22, 35, 42, 0, 42, 24, 0, 0, 19, 
    8, 22, 15, 57, 0, 0, 36, 12, 32, 0, 34, 24, 0, 0, 33, 
    11, 0, 34, 7, 16, 0, 24, 14, 0, 25, 0, 39, 0, 11, 31, 
    3, 0, 52, 0, 22, 5, 0, 24, 0, 26, 44, 14, 0, 26, 59, 
    0, 0, 41, 0, 68, 4, 0, 13, 44, 25, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 32, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 5, 9, 0, 
    0, 47, 0, 0, 0, 45, 0, 0, 0, 14, 0, 0, 0, 19, 3, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 84, 0, 6, 0, 0, 51, 
    0, 0, 0, 48, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 18, 
    0, 21, 0, 0, 115, 34, 0, 0, 0, 94, 0, 0, 14, 0, 0, 
    0, 0, 21, 0, 61, 17, 11, 0, 0, 92, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 81, 0, 28, 0, 66, 0, 0, 24, 14, 0, 
    0, 22, 0, 25, 0, 59, 0, 0, 19, 0, 42, 0, 19, 5, 0, 
    21, 29, 0, 33, 0, 8, 22, 0, 0, 41, 0, 0, 9, 4, 0, 
    63, 18, 0, 79, 0, 0, 49, 46, 0, 0, 0, 0, 6, 24, 2, 
    135, 81, 0, 64, 4, 33, 42, 41, 16, 14, 16, 18, 11, 17, 11, 
    0, 110, 97, 16, 0, 7, 7, 9, 7, 8, 10, 9, 23, 31, 11, 
    5, 16, 160, 9, 2, 15, 0, 7, 18, 16, 20, 35, 17, 27, 37, 
    0, 19, 25, 58, 15, 44, 45, 16, 8, 0, 1, 19, 22, 0, 0, 
    
    -- channel=25
    15, 12, 21, 17, 19, 19, 13, 17, 21, 5, 0, 11, 19, 12, 15, 
    24, 19, 20, 12, 29, 48, 0, 2, 0, 46, 21, 10, 14, 22, 15, 
    0, 28, 20, 18, 19, 0, 0, 16, 38, 48, 0, 11, 0, 12, 24, 
    0, 75, 10, 29, 6, 57, 8, 0, 3, 29, 0, 0, 0, 0, 41, 
    0, 18, 0, 92, 23, 6, 0, 0, 0, 98, 8, 0, 15, 0, 15, 
    0, 0, 0, 0, 6, 2, 0, 0, 0, 120, 0, 0, 12, 5, 15, 
    14, 0, 6, 0, 19, 57, 0, 0, 0, 66, 0, 0, 20, 31, 0, 
    3, 0, 4, 5, 39, 0, 0, 0, 0, 28, 0, 0, 21, 0, 13, 
    0, 0, 0, 27, 4, 0, 3, 4, 41, 0, 0, 0, 18, 32, 17, 
    0, 0, 0, 48, 0, 14, 64, 0, 0, 0, 0, 17, 30, 23, 5, 
    27, 0, 0, 126, 0, 0, 0, 0, 0, 5, 39, 35, 14, 15, 10, 
    0, 14, 0, 32, 0, 0, 0, 0, 0, 7, 4, 5, 11, 1, 0, 
    0, 0, 82, 0, 0, 5, 0, 1, 5, 11, 16, 11, 0, 0, 27, 
    0, 0, 34, 0, 0, 9, 0, 0, 5, 5, 0, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 11, 10, 0, 12, 47, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 14, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 53, 20, 0, 0, 0, 8, 12, 0, 0, 0, 0, 
    0, 33, 0, 0, 25, 0, 45, 0, 0, 38, 2, 0, 0, 0, 0, 
    0, 26, 0, 0, 2, 61, 22, 10, 0, 25, 0, 0, 0, 1, 0, 
    19, 41, 0, 9, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 39, 0, 19, 1, 0, 0, 5, 0, 1, 0, 0, 0, 0, 0, 
    41, 30, 2, 22, 0, 0, 46, 54, 4, 0, 0, 0, 0, 0, 0, 
    61, 47, 24, 73, 61, 0, 2, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 39, 25, 67, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 1, 
    0, 1, 50, 51, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 32, 
    3, 4, 3, 22, 0, 0, 7, 0, 0, 0, 0, 0, 4, 16, 0, 
    
    -- channel=28
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 4, 9, 0, 
    0, 40, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 14, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 5, 0, 0, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 11, 
    0, 0, 0, 16, 102, 13, 0, 0, 0, 29, 0, 0, 1, 0, 0, 
    0, 0, 12, 0, 42, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 40, 0, 20, 0, 43, 0, 0, 9, 15, 1, 
    0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 46, 8, 25, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    14, 0, 0, 1, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    75, 26, 0, 0, 0, 20, 21, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 60, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 83, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 35, 0, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 2, 0, 0, 
    8, 0, 0, 0, 0, 20, 23, 19, 0, 0, 9, 1, 8, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 3, 2, 0, 16, 18, 26, 15, 0, 
    7, 0, 0, 0, 0, 0, 18, 17, 22, 0, 0, 12, 0, 11, 0, 
    16, 0, 1, 20, 31, 23, 7, 9, 16, 0, 12, 30, 2, 6, 0, 
    6, 11, 5, 24, 0, 0, 9, 1, 27, 0, 27, 15, 1, 0, 3, 
    1, 9, 0, 0, 0, 0, 26, 24, 22, 0, 21, 28, 4, 9, 11, 
    2, 0, 22, 0, 0, 34, 25, 4, 0, 6, 31, 45, 15, 0, 0, 
    9, 0, 30, 0, 20, 0, 0, 0, 0, 28, 34, 20, 0, 0, 0, 
    0, 0, 34, 0, 0, 0, 0, 17, 16, 4, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 67, 60, 35, 35, 21, 5, 1, 3, 1, 2, 7, 
    0, 2, 0, 6, 67, 7, 11, 9, 8, 1, 0, 0, 1, 3, 0, 
    10, 0, 0, 48, 18, 0, 5, 9, 7, 3, 4, 11, 9, 0, 21, 
    12, 8, 6, 38, 17, 15, 14, 5, 0, 0, 9, 4, 0, 0, 19, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 49, 0, 1, 49, 22, 0, 0, 0, 32, 18, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 21, 0, 0, 84, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 46, 0, 0, 0, 58, 0, 0, 0, 9, 0, 
    21, 24, 0, 0, 0, 14, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    27, 31, 0, 12, 0, 0, 0, 2, 4, 0, 0, 0, 0, 4, 0, 
    24, 33, 0, 42, 0, 0, 23, 28, 0, 0, 0, 0, 0, 0, 0, 
    33, 25, 0, 131, 75, 27, 10, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 10, 12, 102, 0, 0, 0, 0, 0, 0, 0, 4, 18, 22, 11, 
    10, 0, 53, 10, 0, 8, 0, 2, 4, 13, 23, 29, 8, 5, 48, 
    9, 10, 17, 0, 0, 15, 12, 4, 4, 14, 11, 5, 10, 43, 0, 
    9, 19, 4, 0, 0, 0, 0, 5, 23, 33, 11, 21, 67, 42, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 1, 7, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 3, 7, 3, 0, 6, 1, 6, 0, 
    6, 10, 0, 0, 0, 0, 2, 4, 11, 0, 0, 5, 1, 5, 0, 
    21, 20, 0, 0, 5, 0, 0, 0, 9, 0, 16, 1, 4, 3, 0, 
    6, 39, 0, 0, 0, 0, 20, 0, 12, 7, 9, 6, 0, 3, 6, 
    16, 17, 0, 0, 0, 28, 13, 6, 0, 0, 2, 6, 7, 11, 0, 
    26, 30, 27, 3, 0, 0, 0, 4, 0, 0, 13, 1, 0, 0, 0, 
    18, 26, 29, 4, 29, 0, 0, 13, 15, 10, 5, 2, 3, 0, 0, 
    29, 20, 24, 3, 20, 36, 49, 45, 35, 6, 24, 38, 44, 31, 30, 
    81, 36, 17, 27, 68, 44, 47, 47, 56, 58, 67, 67, 71, 73, 74, 
    90, 70, 9, 61, 39, 61, 65, 60, 61, 66, 70, 77, 83, 77, 75, 
    92, 79, 65, 67, 53, 61, 63, 65, 66, 72, 80, 86, 78, 91, 109, 
    92, 85, 77, 59, 63, 70, 72, 63, 64, 67, 78, 69, 68, 96, 87, 
    
    -- channel=32
    12, 11, 11, 11, 11, 10, 10, 11, 11, 11, 8, 10, 11, 11, 11, 
    9, 9, 9, 9, 8, 9, 8, 8, 8, 0, 0, 0, 10, 9, 10, 
    1, 4, 8, 9, 11, 10, 2, 0, 0, 0, 0, 0, 8, 8, 9, 
    10, 13, 9, 9, 9, 0, 0, 9, 42, 62, 74, 54, 7, 9, 9, 
    0, 0, 0, 0, 4, 7, 35, 16, 33, 20, 0, 0, 0, 0, 0, 
    116, 120, 40, 0, 0, 0, 0, 0, 0, 0, 54, 96, 95, 78, 4, 
    0, 0, 0, 0, 27, 0, 0, 34, 71, 0, 0, 0, 0, 0, 0, 
    0, 90, 0, 0, 0, 108, 153, 40, 0, 0, 0, 16, 41, 62, 63, 
    91, 48, 96, 83, 24, 0, 0, 0, 29, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 9, 
    0, 0, 18, 26, 0, 0, 45, 130, 72, 71, 85, 99, 26, 0, 22, 
    31, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 15, 25, 27, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 57, 7, 10, 7, 
    0, 25, 17, 10, 11, 12, 3, 0, 46, 68, 25, 0, 11, 19, 18, 
    
    -- channel=33
    27, 26, 26, 26, 27, 27, 27, 26, 26, 28, 30, 26, 26, 26, 26, 
    28, 27, 27, 27, 26, 26, 27, 26, 26, 42, 34, 24, 26, 26, 26, 
    30, 28, 26, 26, 26, 27, 30, 36, 52, 52, 41, 33, 27, 27, 27, 
    29, 30, 27, 26, 26, 30, 27, 30, 29, 25, 14, 14, 31, 30, 28, 
    61, 58, 30, 26, 28, 26, 15, 27, 29, 44, 66, 68, 63, 47, 30, 
    22, 13, 18, 38, 39, 78, 79, 73, 59, 38, 25, 14, 11, 4, 31, 
    71, 62, 51, 28, 27, 41, 11, 0, 1, 42, 64, 71, 66, 61, 54, 
    28, 0, 22, 11, 28, 15, 6, 38, 45, 34, 21, 9, 3, 5, 23, 
    0, 23, 15, 14, 37, 47, 56, 66, 48, 67, 65, 71, 73, 67, 52, 
    45, 79, 78, 79, 73, 66, 60, 49, 51, 53, 55, 53, 44, 39, 30, 
    28, 30, 43, 55, 60, 69, 84, 81, 75, 68, 60, 45, 31, 18, 16, 
    5, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 11, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 7, 15, 
    
    -- channel=34
    5, 8, 8, 8, 9, 8, 9, 8, 10, 6, 7, 8, 8, 8, 9, 
    6, 8, 8, 8, 9, 8, 9, 8, 4, 0, 33, 20, 7, 8, 8, 
    12, 12, 9, 7, 9, 4, 13, 0, 5, 0, 40, 48, 8, 9, 9, 
    7, 2, 10, 10, 10, 0, 32, 0, 0, 0, 0, 24, 3, 6, 8, 
    29, 51, 41, 17, 10, 0, 18, 0, 2, 0, 0, 15, 25, 67, 10, 
    0, 0, 12, 26, 22, 28, 59, 54, 50, 0, 0, 0, 0, 32, 13, 
    31, 70, 31, 13, 0, 0, 0, 0, 24, 7, 18, 26, 33, 32, 58, 
    45, 0, 0, 65, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 1, 
    96, 0, 0, 10, 20, 2, 13, 0, 0, 0, 0, 0, 18, 22, 1, 
    74, 21, 22, 14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    2, 18, 2, 19, 35, 42, 22, 21, 5, 0, 0, 0, 0, 0, 13, 
    0, 46, 0, 0, 0, 12, 2, 0, 0, 0, 0, 0, 14, 10, 22, 
    0, 25, 33, 2, 0, 6, 170, 51, 48, 43, 59, 44, 15, 25, 27, 
    0, 2, 12, 4, 4, 4, 111, 130, 112, 74, 27, 32, 16, 25, 28, 
    0, 0, 0, 0, 0, 0, 37, 64, 28, 43, 23, 12, 17, 19, 22, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 4, 1, 8, 0, 0, 0, 0, 0, 0, 
    71, 75, 8, 0, 0, 0, 0, 0, 0, 0, 9, 35, 41, 10, 0, 
    0, 0, 0, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 0, 0, 50, 72, 3, 0, 0, 0, 0, 0, 1, 0, 
    21, 24, 64, 47, 16, 0, 0, 0, 29, 5, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 6, 0, 0, 46, 5, 0, 0, 7, 10, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 37, 20, 0, 0, 0, 6, 2, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 8, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 30, 6, 0, 0, 2, 0, 
    
    -- channel=36
    42, 42, 42, 42, 42, 42, 42, 43, 44, 40, 39, 42, 42, 42, 42, 
    42, 43, 43, 42, 43, 42, 43, 43, 40, 19, 30, 43, 43, 43, 43, 
    39, 42, 44, 43, 44, 41, 38, 26, 4, 0, 5, 33, 42, 42, 43, 
    35, 37, 39, 44, 45, 36, 41, 29, 31, 28, 40, 43, 34, 37, 39, 
    0, 0, 33, 42, 42, 34, 47, 38, 40, 21, 0, 0, 0, 13, 36, 
    24, 41, 35, 21, 21, 0, 0, 0, 5, 23, 29, 36, 38, 54, 33, 
    0, 0, 0, 30, 17, 0, 17, 52, 54, 17, 0, 0, 0, 0, 7, 
    0, 41, 12, 41, 29, 42, 49, 13, 6, 16, 22, 29, 34, 36, 24, 
    65, 11, 34, 35, 23, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 19, 
    0, 0, 1, 0, 0, 0, 44, 29, 19, 23, 37, 30, 19, 24, 36, 
    0, 3, 5, 1, 0, 2, 31, 74, 86, 68, 44, 42, 42, 32, 33, 
    0, 1, 3, 1, 0, 1, 57, 147, 113, 74, 61, 44, 27, 27, 25, 
    0, 10, 6, 4, 8, 7, 27, 59, 60, 58, 37, 20, 24, 26, 28, 
    
    -- channel=37
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 0, 30, 9, 28, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 8, 5, 0, 0, 0, 0, 
    14, 5, 0, 0, 0, 0, 0, 0, 0, 14, 19, 21, 58, 0, 0, 
    0, 0, 0, 0, 33, 116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 0, 0, 29, 0, 42, 0, 8, 29, 9, 2, 0, 0, 
    0, 0, 5, 0, 0, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 4, 0, 19, 0, 4, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 19, 39, 16, 0, 0, 73, 30, 19, 5, 0, 0, 0, 0, 
    58, 0, 0, 9, 6, 0, 0, 0, 4, 10, 5, 0, 0, 0, 0, 
    98, 3, 0, 4, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    77, 19, 9, 8, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    256, 255, 255, 255, 255, 257, 257, 256, 255, 256, 258, 256, 256, 255, 256, 
    257, 256, 256, 256, 256, 256, 256, 256, 255, 250, 244, 251, 256, 256, 257, 
    257, 256, 257, 257, 256, 258, 256, 256, 239, 218, 210, 254, 257, 258, 259, 
    252, 256, 257, 258, 259, 258, 245, 243, 214, 203, 189, 217, 261, 260, 261, 
    194, 204, 258, 256, 258, 254, 240, 253, 249, 255, 253, 239, 223, 235, 263, 
    186, 197, 233, 229, 252, 235, 249, 254, 261, 258, 211, 193, 181, 196, 258, 
    179, 187, 212, 218, 231, 115, 95, 117, 177, 251, 252, 240, 237, 235, 233, 
    76, 134, 131, 181, 221, 186, 189, 215, 210, 187, 149, 133, 137, 159, 179, 
    70, 222, 192, 213, 246, 257, 259, 236, 205, 208, 222, 212, 206, 201, 187, 
    171, 201, 204, 205, 205, 202, 193, 163, 169, 146, 147, 132, 120, 125, 141, 
    34, 59, 60, 67, 79, 100, 124, 126, 126, 110, 98, 93, 98, 104, 126, 
    5, 14, 42, 4, 0, 0, 55, 27, 32, 36, 48, 77, 114, 122, 130, 
    0, 0, 6, 0, 0, 0, 44, 126, 107, 105, 105, 95, 88, 120, 159, 
    20, 0, 0, 0, 0, 0, 0, 43, 41, 40, 43, 83, 116, 134, 180, 
    31, 0, 0, 0, 0, 0, 0, 17, 14, 57, 105, 115, 126, 149, 186, 
    
    -- channel=39
    5, 4, 4, 4, 4, 4, 4, 6, 6, 4, 2, 4, 5, 4, 4, 
    5, 4, 4, 5, 4, 4, 4, 5, 6, 22, 0, 0, 5, 4, 4, 
    6, 5, 5, 6, 4, 7, 0, 13, 3, 5, 0, 0, 4, 4, 4, 
    0, 0, 0, 5, 6, 27, 0, 20, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 6, 4, 15, 0, 5, 0, 0, 0, 3, 1, 0, 0, 
    0, 0, 0, 2, 9, 0, 0, 0, 0, 13, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 13, 24, 0, 0, 0, 0, 3, 10, 1, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    10, 0, 5, 16, 3, 0, 0, 73, 68, 60, 52, 33, 0, 0, 0, 
    41, 0, 0, 3, 0, 0, 0, 97, 102, 56, 6, 0, 1, 0, 0, 
    33, 3, 0, 0, 0, 0, 0, 31, 12, 0, 5, 1, 0, 0, 0, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 20, 40, 47, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 2, 0, 0, 0, 0, 0, 0, 
    55, 56, 18, 0, 0, 0, 0, 0, 0, 0, 30, 52, 68, 29, 0, 
    0, 0, 0, 0, 30, 15, 20, 39, 22, 0, 0, 0, 0, 0, 0, 
    0, 63, 0, 0, 0, 58, 75, 23, 0, 0, 5, 25, 35, 42, 25, 
    22, 33, 39, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 21, 8, 
    11, 1, 32, 45, 30, 17, 67, 114, 78, 71, 71, 58, 13, 0, 15, 
    53, 12, 0, 3, 19, 25, 0, 0, 0, 0, 0, 0, 11, 21, 13, 
    52, 29, 21, 22, 26, 27, 0, 0, 0, 0, 33, 40, 14, 7, 2, 
    29, 50, 46, 41, 41, 43, 17, 0, 35, 45, 25, 7, 11, 12, 7, 
    
    -- channel=41
    9, 9, 9, 9, 9, 9, 9, 10, 10, 9, 8, 10, 10, 9, 9, 
    10, 9, 9, 10, 10, 10, 9, 10, 10, 12, 16, 9, 9, 10, 9, 
    10, 9, 10, 10, 9, 10, 9, 11, 15, 17, 5, 12, 10, 10, 9, 
    5, 7, 10, 10, 8, 14, 14, 17, 5, 0, 0, 0, 10, 10, 10, 
    23, 23, 21, 11, 10, 16, 5, 11, 3, 5, 7, 18, 22, 21, 13, 
    0, 0, 0, 12, 21, 14, 23, 21, 17, 17, 9, 0, 0, 0, 8, 
    18, 15, 16, 15, 8, 15, 6, 5, 0, 5, 11, 17, 21, 16, 15, 
    6, 1, 15, 12, 21, 4, 0, 0, 16, 17, 12, 7, 3, 1, 0, 
    0, 0, 0, 0, 0, 8, 12, 14, 3, 0, 2, 1, 7, 16, 18, 
    0, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 5, 
    21, 19, 10, 13, 18, 14, 2, 0, 3, 1, 1, 0, 0, 1, 6, 
    29, 21, 20, 17, 20, 18, 4, 0, 0, 0, 0, 0, 0, 16, 12, 
    24, 24, 27, 30, 28, 26, 3, 8, 0, 0, 10, 28, 19, 16, 14, 
    34, 26, 25, 27, 27, 27, 2, 0, 2, 26, 22, 14, 26, 21, 17, 
    45, 32, 31, 30, 28, 27, 17, 21, 27, 18, 24, 31, 26, 21, 16, 
    
    -- channel=42
    170, 171, 171, 171, 171, 171, 172, 172, 172, 170, 171, 171, 172, 171, 172, 
    170, 171, 171, 171, 170, 170, 170, 171, 164, 131, 148, 169, 170, 171, 172, 
    167, 169, 172, 172, 173, 170, 167, 146, 111, 109, 110, 164, 171, 172, 173, 
    166, 166, 171, 173, 173, 160, 163, 159, 159, 155, 150, 158, 170, 171, 174, 
    43, 67, 173, 167, 169, 175, 170, 174, 174, 162, 125, 95, 74, 128, 176, 
    164, 177, 161, 114, 141, 69, 87, 105, 141, 170, 162, 164, 148, 160, 171, 
    20, 41, 96, 150, 148, 16, 45, 99, 146, 153, 121, 94, 109, 97, 112, 
    36, 123, 56, 109, 155, 175, 188, 121, 83, 78, 70, 83, 95, 128, 119, 
    99, 169, 158, 159, 157, 144, 137, 126, 127, 104, 123, 94, 77, 64, 74, 
    71, 48, 51, 53, 61, 71, 74, 65, 69, 50, 46, 41, 45, 51, 73, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 13, 48, 65, 77, 
    0, 0, 18, 0, 0, 0, 94, 45, 34, 42, 70, 83, 66, 66, 92, 
    0, 0, 0, 0, 0, 0, 18, 100, 97, 68, 22, 27, 53, 78, 111, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 32, 58, 64, 82, 119, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 58, 63, 58, 77, 97, 127, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 49, 31, 30, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    104, 83, 14, 0, 0, 0, 0, 0, 0, 0, 56, 90, 100, 40, 0, 
    0, 0, 0, 38, 43, 114, 129, 107, 57, 0, 0, 0, 0, 0, 0, 
    128, 105, 53, 0, 0, 0, 0, 0, 0, 21, 73, 102, 85, 96, 57, 
    0, 0, 11, 16, 0, 0, 0, 12, 64, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 49, 29, 0, 31, 29, 57, 82, 92, 55, 
    67, 108, 103, 95, 80, 56, 42, 16, 22, 16, 40, 29, 5, 10, 6, 
    67, 58, 79, 106, 125, 131, 126, 116, 102, 86, 59, 31, 0, 0, 0, 
    19, 6, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 1, 1, 0, 
    0, 20, 40, 30, 7, 5, 41, 49, 23, 43, 81, 35, 0, 0, 0, 
    0, 0, 2, 4, 0, 0, 0, 16, 51, 2, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    49, 49, 49, 49, 49, 49, 49, 49, 47, 50, 52, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 50, 60, 55, 52, 49, 49, 50, 
    48, 48, 48, 49, 49, 50, 50, 56, 62, 67, 60, 52, 50, 49, 50, 
    60, 57, 53, 48, 49, 54, 47, 53, 59, 67, 66, 64, 57, 54, 53, 
    72, 64, 55, 46, 49, 52, 49, 51, 55, 63, 69, 67, 64, 52, 55, 
    57, 55, 59, 46, 50, 55, 56, 54, 54, 64, 63, 60, 62, 56, 57, 
    74, 66, 63, 46, 67, 62, 67, 64, 60, 58, 56, 55, 52, 58, 56, 
    48, 58, 50, 44, 55, 53, 55, 65, 62, 64, 65, 62, 59, 61, 63, 
    37, 63, 49, 50, 59, 62, 64, 61, 61, 69, 72, 74, 70, 70, 68, 
    71, 80, 87, 91, 91, 90, 93, 87, 88, 82, 85, 80, 75, 67, 61, 
    54, 58, 68, 67, 64, 67, 86, 85, 83, 81, 78, 74, 70, 61, 49, 
    22, 25, 27, 27, 25, 26, 45, 69, 71, 68, 56, 51, 41, 35, 35, 
    20, 19, 17, 13, 16, 17, 16, 0, 0, 0, 0, 11, 20, 29, 39, 
    23, 16, 15, 16, 15, 15, 0, 0, 0, 0, 2, 15, 24, 32, 43, 
    21, 11, 14, 17, 15, 16, 13, 0, 0, 1, 11, 24, 27, 34, 45, 
    
    -- channel=45
    60, 60, 60, 60, 60, 59, 60, 58, 59, 61, 60, 60, 59, 60, 60, 
    59, 59, 59, 59, 59, 59, 59, 58, 59, 39, 37, 55, 60, 59, 60, 
    55, 56, 59, 60, 60, 59, 58, 51, 33, 37, 47, 47, 59, 59, 60, 
    65, 65, 61, 59, 58, 48, 52, 59, 80, 90, 95, 92, 63, 63, 62, 
    0, 6, 43, 53, 57, 56, 72, 62, 76, 71, 47, 23, 9, 27, 62, 
    108, 111, 75, 31, 37, 7, 0, 9, 30, 60, 87, 101, 92, 100, 65, 
    0, 0, 17, 58, 64, 41, 47, 78, 95, 58, 33, 14, 14, 18, 25, 
    22, 95, 38, 37, 52, 100, 126, 69, 17, 20, 41, 58, 72, 83, 89, 
    106, 77, 92, 87, 70, 51, 47, 45, 76, 60, 59, 48, 29, 18, 22, 
    46, 5, 14, 13, 20, 28, 37, 45, 43, 44, 39, 32, 47, 44, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 12, 24, 44, 56, 47, 
    0, 18, 22, 21, 6, 10, 65, 97, 73, 72, 79, 81, 39, 27, 49, 
    15, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 26, 45, 61, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 42, 33, 45, 57, 
    2, 14, 13, 10, 9, 12, 0, 0, 11, 40, 32, 28, 40, 53, 64, 
    
    -- channel=46
    45, 43, 43, 43, 43, 44, 43, 44, 41, 46, 44, 43, 44, 43, 43, 
    46, 44, 44, 45, 44, 45, 44, 44, 53, 98, 37, 32, 45, 44, 44, 
    46, 44, 44, 45, 42, 51, 41, 79, 78, 71, 25, 15, 46, 44, 44, 
    38, 46, 43, 44, 45, 86, 22, 65, 15, 22, 4, 0, 46, 46, 44, 
    86, 49, 20, 42, 46, 54, 24, 43, 32, 58, 80, 86, 87, 6, 41, 
    0, 0, 42, 57, 63, 93, 70, 60, 33, 60, 18, 0, 23, 0, 36, 
    88, 48, 44, 0, 77, 75, 0, 0, 0, 57, 75, 81, 54, 79, 27, 
    0, 0, 26, 3, 27, 0, 0, 69, 75, 66, 47, 10, 0, 0, 4, 
    0, 27, 0, 0, 32, 70, 68, 54, 18, 34, 30, 59, 53, 67, 55, 
    16, 77, 81, 81, 77, 69, 78, 53, 52, 48, 51, 41, 14, 8, 4, 
    34, 15, 48, 46, 45, 45, 60, 55, 56, 51, 32, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 9, 33, 9, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    64, 64, 64, 64, 63, 64, 64, 63, 63, 64, 65, 63, 63, 64, 64, 
    64, 64, 64, 63, 63, 63, 63, 63, 61, 53, 51, 60, 64, 64, 64, 
    62, 62, 64, 63, 64, 63, 63, 57, 50, 55, 44, 56, 63, 63, 64, 
    67, 68, 62, 62, 64, 58, 55, 68, 81, 87, 87, 68, 65, 65, 64, 
    23, 26, 49, 59, 63, 66, 63, 67, 73, 72, 58, 42, 30, 43, 63, 
    93, 93, 62, 40, 45, 26, 25, 33, 52, 74, 84, 88, 88, 70, 65, 
    21, 22, 35, 66, 66, 62, 51, 65, 64, 58, 47, 37, 36, 37, 43, 
    40, 65, 37, 32, 63, 94, 94, 61, 38, 46, 55, 59, 62, 72, 66, 
    57, 70, 83, 72, 69, 61, 52, 65, 73, 65, 68, 59, 47, 39, 43, 
    38, 43, 46, 50, 55, 60, 67, 65, 60, 64, 55, 54, 56, 49, 49, 
    2, 14, 13, 9, 2, 9, 26, 31, 36, 38, 40, 44, 55, 52, 43, 
    3, 2, 25, 18, 4, 4, 68, 80, 66, 67, 67, 62, 40, 37, 41, 
    1, 0, 0, 0, 0, 0, 0, 12, 24, 16, 2, 6, 23, 33, 43, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 24, 31, 44, 
    7, 0, 0, 0, 0, 0, 0, 0, 4, 9, 18, 20, 26, 37, 49, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 27, 90, 37, 0, 0, 0, 0, 0, 0, 
    52, 33, 0, 0, 0, 47, 43, 0, 0, 0, 0, 18, 27, 35, 0, 
    215, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 13, 0, 0, 0, 10, 163, 79, 70, 82, 96, 35, 0, 0, 14, 
    0, 0, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    0, 8, 4, 3, 9, 9, 42, 0, 0, 5, 72, 9, 0, 0, 0, 
    0, 24, 25, 24, 29, 32, 35, 16, 83, 41, 0, 0, 0, 0, 0, 
    
    -- channel=49
    7, 6, 6, 6, 6, 6, 6, 5, 6, 6, 6, 6, 6, 6, 6, 
    8, 8, 8, 8, 9, 9, 9, 11, 14, 17, 18, 11, 10, 10, 10, 
    5, 6, 8, 9, 8, 7, 9, 15, 22, 5, 0, 0, 9, 8, 8, 
    19, 17, 11, 7, 8, 13, 7, 9, 4, 12, 28, 26, 11, 12, 10, 
    57, 34, 0, 7, 10, 7, 14, 5, 5, 0, 0, 5, 18, 8, 6, 
    0, 0, 6, 9, 0, 0, 0, 0, 0, 14, 10, 0, 10, 10, 7, 
    30, 44, 4, 0, 9, 58, 69, 83, 22, 0, 0, 0, 0, 0, 4, 
    0, 0, 28, 31, 13, 0, 0, 1, 44, 70, 75, 58, 52, 28, 7, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 7, 23, 
    0, 0, 13, 17, 26, 28, 39, 41, 30, 22, 19, 10, 1, 0, 1, 
    43, 39, 36, 19, 7, 2, 0, 0, 0, 5, 7, 10, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 45, 40, 29, 8, 0, 0, 1, 8, 
    9, 8, 10, 4, 0, 0, 0, 0, 0, 0, 0, 33, 13, 6, 6, 
    0, 0, 1, 3, 0, 0, 0, 2, 38, 60, 27, 3, 8, 7, 4, 
    0, 2, 3, 2, 4, 7, 17, 53, 23, 0, 0, 5, 1, 2, 5, 
    
    -- channel=50
    58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 57, 58, 58, 58, 
    59, 59, 59, 58, 58, 58, 59, 58, 56, 50, 54, 57, 58, 58, 59, 
    60, 59, 59, 59, 59, 58, 59, 54, 51, 30, 45, 59, 59, 59, 59, 
    53, 55, 59, 60, 60, 51, 59, 43, 32, 24, 21, 53, 57, 58, 60, 
    51, 57, 57, 60, 60, 44, 53, 50, 54, 53, 54, 55, 55, 63, 60, 
    7, 17, 49, 54, 55, 55, 58, 59, 61, 45, 27, 18, 5, 40, 59, 
    37, 49, 43, 33, 25, 0, 0, 8, 39, 56, 58, 56, 47, 52, 59, 
    0, 0, 18, 45, 38, 4, 16, 39, 44, 28, 10, 0, 4, 5, 29, 
    0, 19, 5, 23, 47, 50, 55, 25, 22, 25, 24, 25, 30, 39, 30, 
    25, 36, 41, 40, 39, 32, 23, 16, 15, 4, 9, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 6, 7, 4, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 22, 17, 10, 5, 4, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 30, 
    
    -- channel=51
    2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 3, 2, 2, 2, 
    1, 2, 2, 2, 2, 2, 2, 2, 1, 2, 4, 2, 1, 2, 2, 
    1, 1, 2, 2, 1, 1, 2, 2, 0, 0, 4, 5, 3, 2, 2, 
    4, 4, 5, 2, 1, 3, 3, 0, 4, 5, 7, 6, 6, 5, 5, 
    0, 0, 10, 2, 0, 3, 5, 3, 3, 1, 4, 5, 0, 2, 8, 
    8, 9, 8, 0, 0, 0, 1, 2, 5, 7, 6, 7, 6, 9, 7, 
    0, 0, 0, 2, 10, 0, 4, 1, 1, 2, 0, 0, 0, 0, 0, 
    0, 10, 1, 0, 1, 6, 10, 8, 0, 0, 0, 0, 2, 3, 4, 
    0, 4, 8, 4, 2, 5, 3, 3, 2, 3, 4, 3, 4, 2, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 8, 11, 
    8, 6, 4, 4, 2, 1, 4, 0, 0, 2, 4, 9, 10, 10, 12, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 29, 18, 36, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 0, 38, 0, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 0, 3, 0, 17, 28, 15, 6, 0, 0, 
    1, 0, 0, 5, 0, 39, 0, 0, 0, 16, 14, 7, 47, 0, 0, 
    0, 0, 0, 0, 48, 124, 0, 0, 0, 2, 16, 18, 0, 3, 0, 
    0, 0, 12, 0, 0, 23, 0, 46, 6, 14, 27, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 44, 0, 11, 0, 27, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 10, 1, 31, 7, 23, 0, 0, 0, 
    23, 0, 17, 2, 0, 0, 0, 0, 4, 15, 5, 0, 0, 0, 0, 
    38, 0, 30, 47, 25, 0, 0, 47, 10, 0, 0, 0, 0, 0, 0, 
    71, 0, 0, 28, 17, 4, 0, 0, 1, 20, 16, 0, 0, 0, 0, 
    132, 10, 1, 12, 8, 6, 0, 0, 24, 0, 0, 0, 0, 0, 0, 
    110, 21, 11, 10, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 20, 17, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 4, 0, 0, 0, 38, 41, 0, 0, 0, 
    12, 1, 2, 0, 0, 0, 31, 0, 2, 0, 10, 68, 0, 1, 0, 
    0, 25, 40, 2, 0, 0, 27, 0, 13, 0, 0, 0, 0, 58, 6, 
    14, 39, 11, 0, 0, 0, 2, 6, 22, 0, 0, 2, 0, 97, 12, 
    0, 34, 11, 30, 0, 0, 25, 57, 96, 0, 0, 0, 0, 0, 40, 
    69, 55, 0, 72, 0, 0, 52, 0, 0, 0, 0, 2, 26, 22, 47, 
    237, 0, 20, 36, 25, 0, 0, 0, 7, 1, 3, 0, 0, 0, 0, 
    78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 23, 
    0, 14, 0, 0, 1, 11, 0, 0, 0, 0, 0, 7, 25, 13, 30, 
    0, 63, 0, 0, 0, 26, 78, 0, 5, 16, 35, 34, 17, 0, 44, 
    0, 26, 4, 0, 0, 7, 165, 0, 0, 0, 0, 0, 25, 37, 54, 
    0, 2, 9, 0, 3, 5, 95, 12, 0, 9, 38, 48, 12, 39, 44, 
    0, 0, 3, 1, 5, 8, 44, 18, 35, 63, 17, 6, 24, 33, 42, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 35, 35, 55, 40, 28, 29, 25, 0, 0, 0, 0, 
    27, 30, 8, 13, 35, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 44, 45, 43, 45, 46, 77, 89, 50, 37, 25, 0, 0, 0, 0, 
    0, 41, 40, 43, 49, 48, 52, 55, 51, 5, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 1, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 29, 24, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 7, 24, 18, 12, 0, 37, 34, 35, 29, 14, 2, 0, 0, 
    61, 15, 13, 18, 15, 15, 0, 81, 86, 45, 13, 0, 0, 0, 0, 
    53, 20, 14, 14, 14, 11, 6, 32, 16, 0, 3, 0, 0, 0, 0, 
    
    -- channel=56
    28, 31, 31, 31, 32, 32, 32, 29, 31, 30, 33, 31, 31, 31, 31, 
    30, 31, 31, 31, 32, 31, 33, 30, 27, 21, 74, 48, 30, 31, 31, 
    37, 36, 32, 30, 31, 29, 40, 25, 59, 32, 85, 85, 31, 33, 33, 
    36, 28, 34, 33, 32, 6, 63, 0, 0, 0, 0, 39, 35, 33, 34, 
    106, 131, 89, 41, 36, 9, 29, 21, 24, 24, 59, 85, 97, 134, 44, 
    0, 0, 23, 62, 65, 108, 147, 135, 113, 14, 0, 0, 0, 30, 48, 
    111, 145, 99, 43, 0, 0, 1, 0, 31, 52, 81, 96, 108, 89, 123, 
    77, 0, 12, 84, 32, 0, 0, 0, 63, 30, 0, 0, 0, 0, 13, 
    70, 9, 0, 8, 45, 46, 77, 39, 27, 55, 61, 56, 88, 91, 63, 
    103, 107, 108, 103, 91, 76, 39, 28, 40, 13, 41, 26, 24, 32, 37, 
    29, 49, 43, 75, 100, 119, 113, 108, 84, 66, 52, 39, 21, 0, 24, 
    0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 14, 18, 
    0, 0, 20, 0, 0, 0, 148, 30, 5, 14, 40, 34, 0, 10, 29, 
    0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 5, 27, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 22, 37, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 13, 7, 28, 27, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 
    14, 22, 0, 0, 0, 0, 0, 0, 0, 0, 20, 22, 0, 43, 0, 
    0, 0, 0, 31, 0, 0, 47, 91, 56, 0, 0, 0, 0, 0, 0, 
    61, 37, 0, 22, 17, 34, 35, 0, 0, 0, 14, 37, 44, 44, 9, 
    173, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 14, 11, 
    0, 36, 0, 0, 5, 24, 113, 40, 48, 54, 63, 25, 0, 6, 36, 
    0, 15, 4, 0, 14, 17, 50, 0, 0, 0, 0, 11, 38, 25, 33, 
    0, 17, 18, 16, 18, 19, 48, 0, 0, 36, 64, 27, 11, 26, 21, 
    0, 25, 27, 27, 29, 32, 37, 39, 68, 44, 4, 12, 20, 23, 21, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    61, 61, 61, 61, 61, 62, 62, 62, 61, 60, 62, 61, 62, 61, 62, 
    61, 61, 61, 61, 61, 61, 61, 60, 57, 58, 60, 60, 61, 61, 61, 
    64, 64, 61, 61, 62, 61, 63, 58, 56, 41, 62, 73, 61, 62, 62, 
    56, 57, 62, 63, 64, 57, 57, 44, 33, 28, 17, 45, 60, 60, 62, 
    39, 48, 62, 65, 61, 55, 57, 57, 57, 56, 71, 66, 57, 65, 62, 
    32, 40, 71, 61, 60, 80, 87, 87, 83, 52, 21, 22, 15, 37, 66, 
    43, 55, 51, 37, 50, 0, 0, 0, 23, 74, 80, 75, 73, 77, 68, 
    9, 0, 12, 42, 36, 2, 26, 58, 47, 19, 0, 0, 0, 2, 26, 
    0, 70, 27, 57, 75, 68, 69, 52, 47, 65, 63, 64, 65, 56, 33, 
    87, 63, 66, 63, 59, 51, 44, 23, 33, 13, 30, 14, 10, 18, 23, 
    0, 0, 0, 0, 11, 24, 36, 38, 31, 21, 8, 5, 2, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 10, 5, 
    0, 0, 0, 0, 0, 0, 55, 70, 63, 51, 38, 0, 0, 4, 15, 
    0, 0, 0, 0, 0, 0, 0, 36, 13, 0, 0, 0, 0, 4, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 30, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 89, 31, 0, 0, 0, 0, 0, 0, 0, 15, 46, 66, 66, 0, 
    0, 0, 0, 19, 22, 72, 102, 86, 48, 0, 0, 0, 0, 0, 0, 
    96, 106, 62, 0, 0, 0, 0, 0, 0, 4, 40, 63, 69, 54, 64, 
    39, 0, 0, 42, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 0, 0, 6, 9, 17, 50, 56, 33, 
    61, 81, 78, 73, 59, 38, 9, 0, 9, 0, 18, 9, 0, 5, 5, 
    50, 58, 65, 97, 118, 127, 114, 103, 80, 62, 45, 26, 1, 0, 0, 
    1, 37, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 16, 43, 15, 1, 0, 143, 85, 53, 51, 62, 34, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 41, 57, 44, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 17, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 35, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 40, 1, 0, 
    0, 0, 0, 13, 6, 41, 31, 23, 1, 0, 0, 0, 0, 0, 0, 
    63, 50, 26, 0, 0, 29, 1, 0, 0, 0, 20, 35, 28, 27, 10, 
    9, 0, 9, 3, 0, 0, 0, 0, 30, 31, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 8, 19, 30, 31, 
    0, 53, 49, 52, 46, 37, 34, 28, 25, 29, 31, 36, 13, 9, 4, 
    65, 55, 76, 83, 85, 84, 83, 74, 67, 67, 52, 36, 15, 5, 0, 
    33, 2, 16, 20, 26, 25, 0, 0, 3, 1, 0, 0, 13, 12, 0, 
    19, 22, 46, 48, 29, 24, 10, 98, 81, 78, 74, 50, 2, 0, 0, 
    30, 20, 22, 26, 22, 21, 10, 102, 106, 46, 0, 0, 0, 0, 0, 
    27, 3, 5, 8, 10, 8, 0, 30, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    51, 52, 52, 52, 52, 51, 51, 51, 52, 51, 51, 50, 51, 52, 52, 
    50, 52, 52, 51, 52, 52, 52, 52, 47, 5, 34, 56, 52, 53, 53, 
    44, 48, 53, 53, 54, 50, 48, 24, 0, 0, 11, 42, 51, 52, 53, 
    55, 52, 51, 52, 52, 29, 54, 43, 70, 76, 91, 90, 50, 52, 53, 
    0, 0, 52, 45, 50, 46, 64, 51, 64, 45, 0, 0, 0, 21, 55, 
    78, 92, 51, 0, 16, 0, 0, 0, 0, 46, 80, 89, 74, 101, 53, 
    0, 0, 0, 53, 27, 0, 37, 105, 108, 26, 0, 0, 0, 0, 3, 
    4, 90, 9, 39, 56, 98, 116, 17, 0, 7, 29, 52, 65, 80, 60, 
    137, 40, 68, 53, 35, 12, 6, 0, 24, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 6, 0, 0, 0, 2, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 34, 24, 
    0, 0, 0, 0, 0, 0, 85, 80, 62, 65, 81, 67, 0, 9, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 22, 47, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 5, 24, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 27, 2, 0, 15, 30, 47, 
    
    -- channel=63
    28, 28, 28, 28, 28, 28, 28, 28, 26, 30, 31, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 26, 30, 46, 28, 27, 28, 27, 28, 
    28, 28, 27, 27, 27, 30, 28, 41, 42, 43, 47, 27, 29, 27, 28, 
    34, 33, 30, 27, 28, 37, 24, 28, 30, 33, 27, 35, 34, 32, 30, 
    41, 35, 31, 25, 28, 25, 28, 29, 34, 49, 63, 53, 47, 24, 33, 
    40, 36, 42, 34, 38, 64, 58, 54, 37, 34, 28, 30, 30, 35, 35, 
    53, 33, 42, 21, 48, 23, 14, 1, 32, 51, 57, 54, 49, 49, 35, 
    8, 39, 17, 18, 19, 25, 36, 55, 31, 20, 17, 17, 16, 23, 45, 
    1, 43, 34, 40, 48, 50, 57, 55, 54, 71, 67, 74, 67, 52, 37, 
    71, 62, 65, 66, 61, 57, 56, 50, 55, 50, 58, 48, 49, 47, 35, 
    24, 20, 38, 41, 43, 47, 64, 64, 62, 55, 51, 42, 30, 33, 25, 
    9, 11, 14, 11, 7, 7, 0, 20, 19, 18, 11, 32, 36, 7, 8, 
    3, 4, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 8, 17, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 12, 22, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 10, 14, 24, 
    
    -- channel=64
    14, 17, 15, 12, 12, 10, 9, 9, 10, 9, 0, 8, 15, 13, 14, 
    6, 9, 3, 8, 2, 3, 0, 0, 6, 0, 0, 2, 9, 1, 7, 
    0, 1, 0, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 26, 0, 0, 
    5, 27, 11, 0, 38, 33, 12, 0, 0, 9, 49, 92, 72, 0, 19, 
    3, 0, 0, 0, 0, 14, 31, 47, 72, 60, 50, 0, 0, 0, 0, 
    35, 53, 78, 83, 46, 33, 26, 14, 0, 0, 0, 0, 0, 17, 91, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 32, 62, 20, 0, 4, 0, 
    6, 52, 23, 0, 0, 26, 21, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    60, 52, 51, 54, 48, 45, 37, 35, 32, 36, 41, 30, 35, 30, 30, 
    51, 45, 40, 44, 34, 35, 32, 31, 31, 43, 33, 25, 34, 30, 29, 
    42, 41, 29, 29, 21, 27, 24, 34, 37, 48, 31, 42, 35, 24, 27, 
    38, 32, 25, 22, 15, 19, 21, 24, 47, 41, 26, 35, 37, 28, 28, 
    41, 34, 28, 26, 27, 31, 37, 46, 45, 39, 39, 12, 6, 0, 16, 
    14, 20, 25, 12, 7, 18, 37, 49, 37, 31, 14, 0, 0, 0, 24, 
    33, 32, 32, 26, 33, 38, 36, 32, 19, 19, 10, 14, 15, 13, 37, 
    37, 22, 25, 33, 44, 51, 56, 58, 57, 49, 24, 9, 14, 10, 0, 
    62, 61, 49, 59, 70, 72, 63, 43, 31, 22, 1, 11, 21, 24, 18, 
    41, 36, 50, 57, 53, 44, 45, 54, 52, 32, 26, 34, 42, 36, 22, 
    58, 56, 58, 64, 63, 55, 48, 38, 23, 41, 49, 41, 34, 25, 17, 
    42, 56, 53, 40, 30, 33, 59, 44, 29, 29, 38, 29, 18, 18, 9, 
    47, 64, 64, 53, 45, 37, 30, 30, 36, 29, 23, 20, 21, 12, 7, 
    27, 29, 26, 25, 26, 26, 23, 20, 13, 19, 16, 13, 12, 8, 7, 
    6, 4, 6, 6, 10, 12, 18, 15, 14, 26, 9, 9, 10, 8, 7, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 3, 0, 13, 5, 11, 11, 0, 0, 14, 
    0, 11, 10, 0, 2, 4, 7, 6, 15, 0, 52, 26, 2, 6, 23, 
    0, 24, 27, 1, 11, 7, 0, 33, 39, 0, 76, 53, 5, 18, 33, 
    0, 34, 40, 44, 28, 28, 2, 0, 4, 0, 19, 49, 88, 42, 69, 
    27, 36, 28, 60, 51, 57, 38, 0, 0, 0, 0, 0, 44, 0, 44, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 26, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 20, 29, 0, 33, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 33, 9, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 8, 6, 1, 0, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 5, 0, 17, 
    0, 0, 0, 0, 8, 8, 0, 0, 22, 12, 5, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 13, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 
    
    -- channel=67
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 53, 24, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 6, 0, 0, 0, 0, 
    0, 14, 27, 29, 10, 1, 0, 0, 0, 0, 0, 0, 0, 15, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 21, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=68
    0, 5, 12, 13, 22, 26, 32, 31, 37, 36, 32, 42, 37, 40, 43, 
    1, 15, 23, 24, 32, 33, 35, 35, 38, 18, 31, 47, 40, 40, 47, 
    10, 18, 33, 36, 39, 37, 32, 22, 26, 0, 23, 24, 34, 40, 45, 
    13, 28, 34, 44, 44, 45, 31, 25, 0, 0, 6, 0, 11, 25, 36, 
    0, 3, 0, 6, 9, 10, 4, 0, 0, 0, 0, 11, 26, 37, 21, 
    1, 0, 0, 9, 19, 2, 0, 0, 0, 0, 18, 47, 40, 38, 2, 
    0, 0, 0, 5, 2, 3, 1, 4, 12, 11, 34, 36, 25, 10, 0, 
    0, 7, 10, 8, 2, 0, 0, 0, 0, 0, 16, 36, 31, 29, 59, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 34, 28, 22, 17, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 17, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=69
    20, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 
    22, 0, 0, 4, 0, 2, 0, 0, 0, 40, 0, 0, 11, 0, 0, 
    21, 0, 0, 7, 0, 1, 7, 0, 0, 88, 0, 0, 12, 0, 0, 
    14, 0, 0, 0, 0, 0, 3, 18, 35, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 0, 0, 28, 0, 
    0, 0, 21, 0, 0, 3, 0, 13, 0, 3, 0, 0, 93, 0, 60, 
    0, 13, 7, 0, 0, 13, 6, 21, 21, 9, 0, 0, 22, 7, 77, 
    2, 11, 0, 0, 0, 0, 0, 13, 0, 36, 0, 0, 1, 93, 20, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 28, 0, 3, 3, 10, 0, 
    26, 0, 0, 4, 0, 0, 0, 2, 0, 0, 0, 7, 6, 15, 0, 
    0, 0, 0, 2, 0, 0, 34, 31, 0, 0, 0, 10, 6, 5, 4, 
    0, 0, 32, 10, 0, 0, 5, 10, 0, 0, 2, 7, 8, 7, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 32, 1, 4, 4, 0, 2, 
    1, 0, 0, 0, 0, 0, 0, 7, 0, 42, 0, 2, 0, 0, 26, 
    
    -- channel=70
    223, 189, 244, 247, 259, 250, 262, 265, 257, 270, 260, 267, 258, 270, 257, 
    223, 189, 241, 241, 257, 242, 256, 265, 253, 258, 215, 263, 258, 271, 257, 
    221, 176, 229, 233, 247, 235, 243, 228, 236, 228, 183, 256, 255, 256, 253, 
    211, 163, 216, 226, 230, 224, 224, 209, 180, 143, 115, 119, 200, 231, 215, 
    146, 128, 141, 151, 166, 173, 179, 180, 135, 123, 112, 95, 122, 166, 131, 
    89, 87, 117, 94, 125, 115, 146, 137, 121, 119, 105, 163, 140, 169, 98, 
    112, 102, 102, 113, 148, 155, 151, 138, 130, 135, 150, 193, 186, 126, 100, 
    127, 128, 139, 160, 186, 198, 202, 195, 197, 175, 154, 170, 173, 116, 79, 
    150, 157, 159, 199, 205, 204, 193, 175, 161, 162, 141, 164, 169, 154, 161, 
    121, 133, 172, 177, 174, 172, 181, 180, 171, 183, 176, 176, 159, 129, 100, 
    166, 166, 169, 165, 166, 183, 172, 110, 96, 165, 161, 134, 101, 75, 66, 
    137, 160, 155, 104, 104, 135, 157, 116, 104, 108, 97, 83, 59, 48, 30, 
    118, 140, 134, 110, 104, 98, 88, 84, 86, 81, 60, 53, 52, 31, 25, 
    52, 51, 51, 52, 62, 64, 63, 56, 55, 58, 45, 36, 30, 26, 26, 
    24, 22, 27, 31, 37, 41, 48, 42, 54, 52, 31, 26, 24, 28, 17, 
    
    -- channel=71
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 1, 0, 1, 4, 0, 
    0, 0, 0, 0, 0, 0, 5, 7, 0, 29, 0, 0, 6, 9, 0, 
    5, 0, 0, 6, 7, 8, 20, 0, 0, 60, 0, 0, 18, 14, 0, 
    19, 0, 6, 17, 25, 16, 20, 19, 18, 13, 0, 0, 0, 17, 7, 
    5, 0, 4, 0, 13, 8, 4, 10, 0, 0, 0, 0, 0, 39, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 6, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 9, 40, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 2, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 15, 1, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 4, 
    
    -- channel=72
    15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 2, 10, 8, 8, 0, 
    23, 16, 27, 11, 42, 26, 16, 3, 8, 23, 21, 53, 56, 7, 21, 
    19, 3, 1, 7, 2, 23, 35, 44, 61, 51, 18, 0, 0, 0, 0, 
    29, 42, 50, 49, 26, 19, 15, 7, 0, 0, 0, 0, 0, 31, 81, 
    0, 0, 0, 0, 0, 0, 0, 1, 8, 31, 33, 9, 0, 0, 0, 
    24, 32, 19, 0, 0, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 2, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 6, 
    2, 0, 14, 2, 21, 4, 0, 0, 2, 0, 0, 0, 13, 10, 11, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 9, 8, 10, 16, 22, 
    0, 0, 2, 6, 5, 1, 3, 10, 16, 35, 9, 16, 16, 24, 24, 
    20, 24, 26, 26, 26, 28, 21, 12, 0, 14, 18, 17, 21, 20, 22, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 4, 9, 5, 5, 8, 9, 6, 7, 4, 
    3, 0, 2, 3, 9, 7, 10, 13, 7, 12, 14, 9, 8, 11, 7, 
    10, 1, 9, 13, 17, 14, 17, 16, 16, 27, 5, 13, 18, 20, 10, 
    16, 4, 11, 18, 23, 18, 23, 14, 15, 31, 10, 21, 27, 25, 24, 
    25, 17, 25, 22, 29, 25, 23, 23, 14, 6, 4, 10, 5, 31, 20, 
    8, 3, 9, 10, 1, 1, 0, 4, 7, 11, 2, 0, 12, 28, 11, 
    0, 6, 11, 0, 1, 0, 0, 0, 0, 0, 0, 14, 25, 13, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 20, 18, 16, 19, 17, 
    0, 2, 0, 0, 0, 0, 9, 12, 3, 11, 0, 9, 13, 13, 23, 
    0, 0, 0, 0, 5, 0, 0, 5, 12, 13, 6, 11, 16, 26, 26, 
    0, 0, 0, 0, 2, 11, 10, 17, 9, 11, 19, 27, 24, 26, 19, 
    0, 0, 5, 7, 3, 0, 13, 11, 12, 20, 20, 25, 19, 19, 24, 
    2, 8, 15, 9, 17, 21, 17, 14, 16, 24, 22, 17, 21, 19, 18, 
    18, 22, 22, 18, 18, 21, 22, 22, 18, 12, 21, 17, 20, 18, 20, 
    22, 21, 21, 20, 19, 17, 19, 22, 18, 22, 15, 18, 18, 18, 22, 
    
    -- channel=74
    141, 114, 170, 162, 176, 163, 176, 180, 175, 182, 164, 184, 170, 186, 174, 
    139, 111, 165, 155, 177, 154, 165, 179, 168, 137, 119, 179, 165, 183, 170, 
    137, 95, 153, 153, 169, 150, 154, 125, 136, 108, 100, 150, 154, 169, 166, 
    117, 82, 124, 137, 144, 145, 141, 121, 40, 26, 17, 0, 93, 127, 114, 
    27, 14, 25, 30, 40, 45, 53, 63, 51, 49, 44, 63, 67, 89, 19, 
    46, 39, 54, 45, 84, 56, 72, 53, 52, 64, 86, 155, 85, 135, 23, 
    52, 29, 28, 51, 79, 92, 98, 96, 100, 102, 111, 115, 118, 31, 0, 
    76, 90, 114, 120, 126, 127, 128, 107, 108, 72, 70, 97, 97, 57, 94, 
    59, 51, 74, 115, 103, 93, 93, 101, 101, 113, 106, 96, 92, 81, 76, 
    60, 92, 102, 84, 99, 112, 110, 80, 70, 107, 101, 87, 52, 21, 8, 
    91, 89, 84, 68, 59, 91, 77, 20, 31, 73, 48, 29, 14, 4, 0, 
    74, 77, 65, 30, 50, 69, 58, 37, 31, 32, 12, 9, 0, 0, 0, 
    39, 36, 33, 21, 15, 14, 21, 20, 5, 5, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 3, 0, 43, 8, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 13, 37, 21, 60, 9, 32, 17, 13, 0, 
    32, 1, 34, 29, 25, 11, 13, 12, 83, 60, 37, 90, 72, 57, 49, 
    83, 63, 67, 78, 84, 83, 66, 64, 17, 10, 9, 0, 0, 23, 48, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 2, 
    0, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 36, 58, 
    0, 0, 0, 0, 0, 0, 0, 1, 19, 50, 35, 4, 0, 0, 0, 
    19, 52, 11, 0, 18, 40, 30, 0, 0, 0, 0, 0, 0, 0, 38, 
    0, 0, 0, 19, 0, 0, 0, 38, 39, 3, 0, 22, 58, 66, 46, 
    3, 0, 6, 34, 60, 32, 30, 26, 0, 41, 68, 57, 39, 26, 35, 
    6, 10, 23, 3, 0, 0, 54, 26, 17, 22, 38, 31, 11, 20, 12, 
    31, 64, 69, 49, 54, 44, 13, 12, 40, 36, 12, 15, 24, 6, 0, 
    43, 39, 25, 16, 24, 32, 25, 17, 0, 6, 15, 10, 6, 0, 2, 
    6, 0, 0, 0, 0, 0, 8, 22, 12, 17, 8, 5, 3, 0, 27, 
    
    -- channel=76
    94, 79, 87, 82, 78, 67, 62, 61, 58, 60, 53, 51, 55, 58, 52, 
    82, 65, 69, 64, 61, 54, 55, 55, 53, 64, 45, 49, 50, 53, 47, 
    66, 52, 52, 47, 46, 45, 51, 48, 46, 62, 49, 48, 47, 43, 43, 
    49, 37, 36, 27, 26, 29, 36, 43, 57, 64, 64, 55, 41, 34, 21, 
    49, 44, 48, 42, 36, 35, 42, 59, 62, 69, 66, 45, 33, 37, 31, 
    60, 52, 58, 49, 60, 61, 74, 79, 67, 63, 50, 42, 37, 28, 35, 
    73, 60, 62, 65, 76, 79, 87, 82, 78, 73, 53, 39, 33, 27, 24, 
    80, 71, 73, 82, 86, 87, 90, 86, 78, 68, 43, 32, 34, 36, 33, 
    90, 81, 82, 91, 96, 92, 87, 76, 65, 57, 44, 43, 48, 42, 35, 
    87, 84, 88, 89, 85, 82, 75, 68, 57, 60, 56, 55, 50, 46, 39, 
    89, 94, 90, 82, 78, 74, 79, 65, 55, 61, 58, 56, 49, 44, 42, 
    82, 85, 90, 76, 74, 74, 67, 56, 55, 57, 54, 52, 49, 44, 38, 
    71, 73, 71, 65, 63, 61, 57, 55, 54, 53, 48, 44, 45, 42, 40, 
    53, 51, 51, 50, 48, 47, 50, 50, 43, 52, 43, 41, 41, 41, 39, 
    35, 35, 40, 41, 44, 45, 47, 43, 37, 49, 41, 39, 40, 40, 36, 
    
    -- channel=77
    79, 83, 87, 81, 78, 72, 68, 65, 68, 66, 56, 64, 66, 67, 65, 
    70, 70, 72, 67, 64, 58, 55, 54, 62, 41, 37, 59, 60, 57, 61, 
    58, 57, 59, 56, 55, 50, 46, 32, 43, 24, 44, 39, 46, 43, 52, 
    33, 43, 31, 24, 27, 37, 35, 45, 9, 0, 23, 0, 0, 15, 14, 
    0, 0, 0, 0, 0, 0, 1, 12, 36, 46, 39, 56, 48, 22, 1, 
    50, 56, 46, 46, 61, 63, 62, 49, 49, 55, 77, 84, 57, 18, 32, 
    54, 42, 34, 53, 59, 69, 81, 85, 94, 85, 75, 40, 21, 24, 0, 
    75, 80, 91, 103, 91, 88, 86, 75, 56, 33, 15, 24, 34, 31, 69, 
    56, 33, 56, 68, 67, 55, 53, 57, 65, 60, 71, 51, 40, 38, 18, 
    68, 87, 78, 61, 66, 80, 73, 48, 31, 48, 50, 36, 14, 0, 3, 
    65, 74, 68, 46, 38, 44, 43, 23, 47, 31, 14, 10, 14, 15, 9, 
    61, 59, 49, 41, 55, 61, 26, 33, 36, 28, 22, 18, 23, 17, 9, 
    44, 30, 19, 27, 21, 15, 25, 36, 22, 17, 25, 27, 12, 18, 19, 
    11, 8, 17, 25, 24, 18, 21, 21, 39, 37, 17, 18, 18, 23, 23, 
    15, 21, 25, 28, 32, 35, 31, 15, 26, 17, 17, 16, 21, 22, 1, 
    
    -- channel=78
    58, 0, 27, 40, 44, 37, 42, 60, 35, 48, 46, 38, 45, 52, 30, 
    61, 0, 24, 42, 44, 43, 54, 50, 36, 112, 4, 33, 51, 57, 32, 
    59, 0, 16, 37, 44, 40, 70, 48, 28, 138, 0, 26, 61, 51, 31, 
    59, 0, 36, 29, 48, 32, 50, 57, 94, 81, 38, 61, 6, 52, 22, 
    53, 31, 54, 44, 56, 53, 48, 79, 29, 23, 1, 0, 0, 67, 35, 
    0, 0, 23, 0, 0, 1, 19, 35, 7, 4, 0, 0, 54, 0, 36, 
    3, 9, 22, 0, 12, 19, 16, 0, 0, 0, 0, 26, 46, 37, 55, 
    0, 0, 0, 0, 7, 22, 28, 43, 34, 75, 9, 9, 27, 36, 0, 
    34, 41, 14, 26, 52, 55, 49, 30, 5, 20, 0, 19, 28, 24, 32, 
    21, 0, 13, 47, 24, 11, 21, 48, 16, 24, 24, 50, 52, 58, 23, 
    5, 26, 34, 44, 41, 19, 74, 45, 0, 32, 55, 55, 29, 9, 16, 
    0, 26, 66, 21, 0, 0, 53, 14, 6, 23, 25, 14, 9, 0, 0, 
    0, 37, 44, 18, 26, 26, 8, 2, 15, 16, 0, 0, 11, 0, 0, 
    12, 4, 0, 0, 0, 0, 2, 3, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 9, 
    
    -- channel=79
    89, 82, 89, 86, 84, 77, 73, 72, 69, 70, 65, 68, 72, 71, 70, 
    77, 70, 72, 72, 67, 63, 60, 63, 65, 55, 45, 63, 66, 63, 65, 
    67, 59, 58, 60, 52, 57, 50, 40, 47, 52, 35, 49, 55, 49, 57, 
    49, 45, 36, 38, 36, 43, 44, 46, 31, 27, 29, 0, 8, 26, 23, 
    14, 16, 10, 2, 2, 6, 23, 33, 50, 51, 48, 47, 33, 23, 8, 
    45, 44, 46, 45, 58, 53, 61, 59, 52, 54, 59, 67, 48, 22, 36, 
    51, 45, 42, 53, 59, 78, 81, 86, 82, 71, 55, 38, 41, 10, 25, 
    75, 76, 86, 93, 90, 89, 87, 77, 66, 45, 24, 29, 39, 54, 49, 
    63, 55, 61, 79, 78, 71, 66, 64, 59, 65, 53, 46, 45, 41, 21, 
    77, 78, 79, 69, 76, 76, 68, 51, 46, 52, 52, 44, 29, 17, 13, 
    75, 79, 71, 60, 47, 58, 55, 40, 36, 34, 31, 26, 22, 21, 11, 
    56, 67, 64, 52, 58, 46, 43, 44, 37, 31, 25, 26, 22, 19, 12, 
    41, 42, 38, 39, 31, 25, 32, 32, 24, 24, 24, 22, 20, 18, 18, 
    16, 16, 20, 22, 21, 19, 22, 20, 33, 29, 19, 18, 18, 19, 16, 
    13, 15, 18, 20, 23, 25, 23, 13, 19, 25, 16, 17, 17, 19, 3, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 
    16, 8, 0, 16, 9, 0, 0, 0, 0, 0, 68, 31, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 20, 29, 6, 6, 0, 0, 0, 0, 
    0, 15, 37, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 5, 0, 0, 0, 0, 0, 0, 6, 0, 2, 3, 8, 5, 7, 
    1, 6, 0, 0, 0, 6, 2, 0, 7, 21, 23, 9, 10, 2, 10, 
    0, 6, 0, 1, 0, 6, 4, 8, 1, 18, 0, 0, 4, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 50, 58, 78, 80, 0, 0, 0, 
    17, 30, 39, 32, 27, 25, 28, 15, 0, 0, 0, 0, 0, 27, 42, 
    13, 0, 0, 21, 22, 18, 4, 0, 0, 0, 0, 0, 15, 0, 13, 
    2, 12, 15, 26, 28, 24, 23, 21, 22, 10, 0, 7, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 12, 11, 38, 29, 
    0, 6, 22, 0, 0, 0, 15, 19, 5, 0, 0, 11, 13, 0, 0, 
    33, 0, 0, 14, 16, 0, 0, 0, 0, 0, 6, 0, 0, 10, 19, 
    0, 5, 0, 0, 0, 0, 18, 42, 27, 0, 2, 15, 1, 0, 0, 
    2, 6, 19, 33, 26, 0, 0, 0, 11, 12, 0, 13, 6, 3, 3, 
    0, 0, 0, 0, 8, 23, 6, 0, 0, 11, 0, 0, 0, 0, 1, 
    15, 9, 2, 0, 0, 0, 13, 8, 0, 0, 0, 2, 0, 0, 0, 
    0, 4, 7, 9, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 
    
    -- channel=82
    26, 38, 48, 54, 56, 59, 60, 53, 60, 64, 64, 64, 61, 60, 63, 
    32, 40, 54, 54, 56, 56, 57, 55, 60, 49, 60, 64, 63, 61, 67, 
    33, 43, 54, 51, 53, 51, 44, 55, 61, 24, 46, 65, 59, 58, 65, 
    31, 38, 47, 51, 49, 49, 39, 25, 29, 5, 11, 36, 44, 48, 61, 
    12, 10, 12, 23, 26, 31, 28, 13, 0, 0, 0, 0, 13, 12, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 19, 39, 7, 21, 0, 
    0, 0, 0, 0, 13, 20, 22, 24, 26, 15, 23, 22, 20, 0, 0, 
    5, 9, 23, 25, 29, 30, 28, 16, 16, 0, 4, 16, 18, 10, 16, 
    0, 0, 8, 21, 16, 12, 16, 21, 22, 19, 21, 16, 13, 0, 0, 
    6, 9, 12, 7, 19, 22, 7, 0, 5, 14, 14, 0, 0, 0, 0, 
    7, 11, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    5, 0, 4, 2, 2, 0, 3, 4, 3, 2, 2, 3, 1, 4, 0, 
    5, 1, 4, 2, 4, 1, 1, 4, 2, 6, 0, 2, 0, 3, 0, 
    4, 0, 4, 3, 7, 2, 4, 0, 0, 4, 1, 3, 3, 4, 0, 
    0, 0, 0, 0, 1, 0, 1, 5, 2, 0, 1, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 3, 2, 0, 
    1, 1, 5, 0, 5, 0, 1, 0, 4, 6, 3, 11, 9, 8, 0, 
    3, 2, 0, 1, 0, 2, 0, 2, 7, 8, 9, 2, 0, 0, 0, 
    0, 2, 0, 2, 2, 3, 4, 4, 3, 5, 2, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 2, 6, 6, 3, 4, 6, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 5, 6, 5, 4, 5, 0, 0, 2, 0, 0, 
    2, 1, 0, 1, 0, 4, 8, 0, 0, 6, 2, 0, 3, 2, 5, 
    4, 1, 5, 0, 0, 2, 0, 3, 5, 2, 5, 7, 1, 4, 0, 
    1, 0, 0, 2, 4, 0, 0, 4, 4, 4, 3, 4, 0, 0, 1, 
    0, 0, 1, 2, 4, 6, 4, 5, 3, 6, 2, 0, 0, 1, 2, 
    1, 2, 5, 5, 4, 6, 6, 5, 1, 2, 1, 0, 1, 2, 3, 
    
    -- channel=84
    36, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 3, 0, 0, 
    35, 0, 0, 3, 0, 0, 0, 0, 0, 64, 0, 0, 8, 0, 0, 
    35, 0, 0, 3, 0, 0, 19, 0, 0, 129, 0, 0, 14, 0, 0, 
    32, 0, 0, 0, 0, 0, 18, 31, 48, 44, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 37, 24, 22, 0, 0, 0, 29, 0, 
    0, 0, 32, 0, 0, 2, 0, 32, 5, 10, 0, 0, 88, 0, 77, 
    0, 12, 20, 0, 0, 10, 5, 13, 6, 2, 0, 0, 54, 18, 93, 
    0, 1, 0, 0, 0, 0, 4, 20, 0, 60, 0, 0, 4, 95, 1, 
    12, 4, 0, 0, 11, 9, 5, 8, 0, 40, 0, 0, 3, 22, 0, 
    26, 0, 0, 7, 0, 0, 3, 21, 0, 0, 0, 27, 29, 42, 1, 
    0, 1, 7, 26, 0, 0, 55, 44, 0, 0, 20, 35, 31, 21, 25, 
    0, 0, 53, 16, 0, 0, 46, 23, 0, 11, 28, 15, 26, 17, 27, 
    0, 8, 27, 9, 4, 3, 9, 8, 13, 9, 21, 0, 36, 10, 12, 
    7, 3, 5, 0, 4, 3, 1, 15, 0, 46, 10, 14, 14, 4, 10, 
    10, 0, 1, 0, 0, 4, 7, 22, 0, 66, 6, 12, 6, 0, 50, 
    
    -- channel=85
    0, 44, 23, 6, 4, 6, 5, 0, 17, 3, 0, 8, 0, 0, 15, 
    0, 42, 27, 0, 1, 0, 0, 0, 13, 0, 50, 22, 0, 0, 20, 
    0, 39, 31, 0, 0, 0, 0, 4, 27, 0, 104, 32, 0, 0, 23, 
    0, 40, 14, 10, 0, 5, 0, 0, 0, 0, 19, 19, 61, 0, 24, 
    0, 10, 0, 19, 0, 7, 1, 0, 0, 0, 8, 26, 50, 0, 20, 
    28, 35, 0, 27, 13, 14, 15, 0, 0, 0, 66, 39, 0, 6, 0, 
    19, 2, 0, 53, 25, 0, 1, 0, 8, 6, 64, 13, 0, 0, 0, 
    12, 8, 29, 39, 21, 11, 1, 0, 0, 0, 25, 21, 0, 0, 3, 
    2, 0, 41, 21, 0, 0, 0, 0, 17, 0, 42, 9, 0, 0, 0, 
    0, 48, 22, 0, 1, 10, 3, 0, 11, 1, 5, 0, 0, 0, 0, 
    26, 3, 0, 0, 9, 19, 0, 0, 61, 8, 0, 0, 0, 0, 0, 
    58, 3, 0, 0, 9, 51, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 11, 3, 1, 1, 0, 31, 0, 0, 0, 0, 4, 0, 
    0, 10, 7, 9, 8, 8, 3, 0, 57, 0, 2, 0, 4, 9, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 2, 0, 6, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 2, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 5, 
    0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 3, 0, 18, 0, 2, 0, 0, 18, 
    
    -- channel=88
    3, 47, 43, 39, 36, 39, 40, 19, 44, 41, 46, 41, 28, 27, 41, 
    6, 49, 54, 33, 38, 34, 39, 41, 44, 10, 93, 51, 29, 35, 46, 
    9, 53, 57, 25, 34, 29, 17, 70, 80, 0, 116, 97, 34, 44, 54, 
    26, 51, 62, 65, 42, 42, 27, 3, 37, 33, 38, 93, 156, 72, 94, 
    74, 64, 60, 89, 84, 91, 80, 40, 16, 7, 24, 3, 32, 0, 54, 
    3, 13, 0, 11, 0, 0, 10, 9, 15, 0, 17, 0, 0, 33, 0, 
    17, 8, 8, 31, 31, 0, 0, 0, 0, 0, 24, 39, 0, 36, 0, 
    0, 0, 0, 0, 9, 14, 16, 17, 46, 13, 70, 46, 16, 0, 0, 
    34, 55, 63, 48, 42, 54, 44, 18, 22, 0, 0, 7, 15, 7, 48, 
    0, 10, 24, 31, 27, 13, 20, 41, 71, 32, 22, 19, 41, 31, 37, 
    48, 20, 26, 36, 73, 72, 0, 5, 48, 58, 52, 32, 19, 12, 6, 
    63, 35, 0, 9, 0, 50, 36, 18, 22, 20, 22, 13, 0, 0, 0, 
    65, 60, 54, 42, 42, 38, 16, 13, 27, 21, 1, 15, 0, 0, 0, 
    22, 28, 16, 19, 19, 22, 16, 4, 11, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 
    0, 12, 2, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 5, 0, 0, 
    35, 25, 0, 39, 24, 15, 0, 0, 0, 6, 64, 30, 0, 9, 0, 
    0, 1, 0, 32, 19, 14, 14, 25, 30, 19, 28, 0, 0, 0, 0, 
    13, 23, 30, 14, 3, 0, 0, 0, 0, 0, 5, 8, 0, 0, 60, 
    0, 0, 22, 0, 0, 0, 0, 3, 10, 0, 22, 0, 0, 0, 0, 
    17, 29, 0, 0, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 3, 0, 0, 42, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 8, 24, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 3, 0, 9, 12, 
    0, 1, 4, 8, 0, 0, 6, 1, 43, 0, 5, 2, 9, 14, 7, 
    9, 19, 18, 20, 20, 13, 3, 0, 32, 0, 5, 9, 11, 17, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    45, 39, 61, 64, 66, 63, 67, 63, 66, 69, 70, 66, 61, 67, 65, 
    43, 36, 62, 56, 63, 57, 63, 67, 64, 59, 47, 68, 61, 70, 63, 
    45, 35, 57, 49, 60, 49, 54, 64, 58, 37, 43, 79, 57, 64, 65, 
    49, 29, 63, 62, 62, 53, 52, 34, 33, 0, 0, 8, 58, 68, 65, 
    23, 12, 15, 31, 33, 39, 32, 32, 5, 8, 10, 0, 28, 10, 4, 
    0, 0, 4, 0, 0, 0, 16, 13, 5, 0, 0, 24, 0, 36, 0, 
    12, 0, 0, 4, 15, 6, 10, 0, 0, 2, 22, 45, 27, 30, 0, 
    9, 1, 13, 29, 39, 38, 38, 38, 47, 32, 28, 27, 25, 0, 0, 
    27, 37, 23, 43, 50, 49, 33, 16, 19, 10, 17, 24, 24, 15, 41, 
    0, 10, 42, 37, 17, 20, 33, 41, 38, 31, 31, 30, 31, 9, 0, 
    26, 26, 27, 33, 44, 36, 20, 0, 0, 35, 30, 6, 0, 0, 0, 
    26, 21, 12, 0, 0, 24, 33, 6, 0, 0, 0, 0, 0, 0, 0, 
    22, 30, 25, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 26, 24, 0, 56, 33, 0, 0, 0, 
    0, 10, 28, 26, 9, 4, 0, 0, 17, 24, 15, 81, 115, 40, 52, 
    61, 43, 45, 68, 65, 66, 46, 20, 0, 0, 0, 0, 0, 0, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 38, 11, 0, 0, 0, 
    7, 24, 19, 0, 0, 12, 4, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 9, 27, 0, 0, 0, 22, 26, 28, 
    1, 0, 0, 8, 42, 26, 0, 0, 12, 30, 32, 21, 11, 4, 10, 
    22, 0, 0, 0, 0, 15, 20, 0, 0, 5, 11, 3, 0, 0, 0, 
    36, 41, 42, 27, 30, 28, 5, 0, 16, 13, 0, 5, 0, 0, 0, 
    29, 32, 15, 13, 11, 14, 8, 2, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 25, 0, 0, 0, 0, 0, 0, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 4, 9, 0, 42, 0, 0, 0, 0, 0, 
    19, 0, 9, 9, 10, 2, 8, 1, 38, 58, 21, 52, 29, 13, 13, 
    47, 35, 39, 35, 42, 38, 31, 36, 19, 10, 7, 0, 0, 16, 25, 
    0, 0, 2, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 4, 20, 
    0, 10, 22, 0, 1, 0, 0, 0, 0, 0, 0, 0, 20, 13, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 28, 14, 6, 4, 14, 0, 
    17, 26, 7, 2, 8, 14, 11, 3, 0, 0, 0, 0, 2, 7, 15, 
    8, 0, 0, 10, 3, 0, 0, 9, 8, 0, 0, 15, 27, 40, 28, 
    0, 0, 4, 20, 21, 6, 22, 35, 0, 13, 30, 35, 27, 20, 27, 
    0, 9, 23, 21, 3, 0, 33, 13, 6, 18, 21, 18, 23, 21, 27, 
    7, 27, 39, 24, 29, 33, 24, 9, 19, 23, 19, 12, 28, 18, 14, 
    38, 38, 25, 16, 13, 16, 18, 20, 0, 10, 20, 21, 19, 12, 15, 
    17, 11, 8, 7, 5, 2, 7, 21, 3, 30, 20, 22, 14, 11, 35, 
    
    -- channel=94
    44, 55, 72, 60, 66, 58, 58, 52, 61, 57, 39, 61, 55, 60, 61, 
    39, 47, 62, 49, 57, 45, 44, 48, 53, 6, 35, 57, 48, 51, 59, 
    30, 31, 52, 45, 47, 40, 29, 11, 28, 0, 34, 21, 30, 38, 49, 
    0, 20, 9, 15, 13, 28, 17, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 13, 9, 0, 
    20, 11, 0, 19, 37, 22, 14, 0, 1, 11, 60, 76, 22, 19, 0, 
    7, 0, 0, 22, 33, 41, 53, 57, 69, 59, 62, 24, 3, 0, 0, 
    34, 49, 60, 64, 55, 51, 47, 28, 16, 0, 0, 15, 11, 2, 77, 
    0, 0, 30, 39, 19, 4, 16, 33, 41, 32, 49, 23, 15, 5, 0, 
    36, 52, 30, 16, 41, 49, 30, 0, 0, 22, 24, 0, 0, 0, 0, 
    29, 31, 21, 0, 0, 12, 0, 0, 22, 0, 0, 0, 0, 0, 0, 
    28, 19, 0, 4, 25, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    66, 48, 57, 55, 51, 41, 40, 39, 35, 40, 32, 30, 32, 36, 28, 
    55, 38, 43, 42, 38, 32, 36, 34, 31, 50, 15, 27, 29, 34, 24, 
    45, 27, 30, 25, 29, 23, 35, 29, 27, 43, 33, 32, 29, 25, 23, 
    36, 19, 31, 14, 17, 15, 20, 37, 38, 23, 26, 26, 25, 29, 12, 
    28, 24, 22, 24, 18, 22, 22, 41, 39, 49, 39, 19, 17, 14, 13, 
    26, 31, 39, 13, 28, 35, 51, 54, 43, 36, 17, 22, 24, 8, 19, 
    48, 37, 32, 33, 40, 41, 48, 40, 39, 40, 32, 20, 11, 24, 11, 
    48, 39, 46, 57, 59, 60, 63, 65, 57, 53, 17, 11, 15, 0, 0, 
    71, 54, 44, 60, 72, 67, 55, 39, 37, 28, 24, 23, 24, 30, 21, 
    40, 58, 64, 60, 46, 53, 56, 60, 38, 35, 33, 42, 39, 28, 16, 
    56, 62, 65, 65, 63, 45, 55, 27, 24, 50, 42, 32, 33, 23, 30, 
    53, 54, 58, 36, 35, 55, 56, 41, 32, 32, 40, 24, 28, 25, 15, 
    55, 61, 56, 50, 41, 30, 29, 39, 38, 28, 27, 27, 24, 19, 17, 
    28, 25, 27, 29, 32, 29, 25, 26, 17, 36, 20, 22, 19, 19, 21, 
    15, 13, 16, 17, 21, 25, 29, 25, 17, 25, 21, 17, 20, 18, 21, 
    
    -- channel=96
    3, 7, 16, 6, 0, 5, 9, 9, 17, 11, 11, 7, 16, 25, 16, 
    1, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 14, 39, 22, 28, 36, 43, 40, 42, 0, 6, 6, 
    9, 0, 0, 37, 14, 12, 28, 21, 10, 0, 0, 7, 19, 0, 0, 
    17, 5, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 22, 6, 4, 
    10, 8, 0, 0, 50, 48, 46, 42, 44, 42, 41, 28, 2, 7, 12, 
    7, 18, 31, 0, 0, 0, 7, 11, 14, 14, 7, 5, 1, 0, 0, 
    6, 11, 36, 112, 39, 0, 0, 0, 2, 0, 7, 7, 9, 8, 7, 
    5, 7, 9, 11, 42, 0, 0, 0, 0, 0, 0, 10, 6, 2, 3, 
    1, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 3, 1, 115, 168, 92, 110, 145, 125, 140, 115, 95, 58, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 
    0, 0, 0, 0, 0, 9, 18, 15, 17, 20, 12, 2, 9, 62, 0, 
    
    -- channel=97
    29, 35, 33, 17, 22, 20, 18, 18, 16, 16, 17, 18, 15, 21, 29, 
    41, 51, 47, 0, 2, 21, 17, 11, 16, 21, 21, 16, 37, 36, 33, 
    42, 51, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 39, 37, 
    41, 50, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 42, 
    41, 47, 44, 35, 31, 32, 31, 26, 36, 30, 22, 28, 32, 41, 45, 
    39, 53, 62, 40, 31, 31, 29, 31, 32, 33, 29, 35, 43, 38, 40, 
    33, 34, 10, 37, 64, 48, 39, 41, 40, 41, 41, 44, 43, 43, 44, 
    34, 43, 29, 0, 9, 41, 53, 40, 38, 39, 37, 40, 40, 41, 43, 
    33, 38, 36, 30, 29, 0, 11, 46, 63, 54, 41, 36, 40, 43, 44, 
    29, 33, 36, 41, 45, 1, 0, 0, 0, 17, 46, 67, 66, 51, 42, 
    29, 32, 36, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 28, 
    62, 70, 73, 72, 74, 75, 59, 51, 63, 61, 54, 56, 51, 58, 59, 
    19, 18, 20, 19, 17, 21, 24, 31, 42, 44, 46, 48, 53, 54, 50, 
    15, 10, 13, 5, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    
    -- channel=98
    21, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 3, 3, 1, 
    14, 0, 0, 0, 53, 57, 42, 54, 47, 49, 44, 50, 16, 4, 4, 
    13, 0, 0, 24, 21, 42, 39, 53, 33, 26, 32, 40, 37, 0, 4, 
    3, 0, 0, 29, 30, 23, 18, 40, 30, 17, 37, 26, 45, 0, 1, 
    0, 0, 0, 0, 1, 2, 0, 2, 1, 0, 7, 20, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 46, 68, 17, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    13, 0, 0, 0, 0, 85, 65, 7, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 24, 66, 81, 69, 33, 18, 0, 0, 0, 0, 
    20, 5, 0, 0, 0, 22, 28, 20, 28, 33, 86, 78, 69, 33, 3, 
    25, 1, 1, 0, 0, 0, 0, 12, 0, 0, 0, 0, 24, 7, 7, 
    63, 43, 46, 49, 56, 14, 33, 59, 24, 8, 23, 7, 21, 17, 18, 
    8, 0, 0, 0, 1, 0, 5, 23, 7, 18, 19, 25, 26, 22, 27, 
    15, 21, 13, 17, 11, 13, 13, 15, 7, 6, 10, 9, 9, 7, 0, 
    0, 6, 5, 10, 5, 5, 0, 6, 0, 0, 0, 3, 11, 0, 0, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 32, 30, 32, 30, 40, 35, 34, 32, 1, 0, 0, 
    0, 0, 0, 12, 0, 0, 10, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 6, 13, 16, 16, 15, 16, 14, 14, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 44, 75, 3, 12, 73, 36, 60, 19, 3, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=100
    20, 18, 20, 30, 35, 35, 36, 36, 38, 39, 38, 35, 38, 38, 32, 
    16, 6, 15, 63, 74, 58, 59, 62, 60, 57, 55, 49, 40, 30, 33, 
    13, 6, 9, 56, 61, 71, 71, 77, 65, 62, 62, 65, 37, 29, 28, 
    16, 7, 33, 107, 78, 72, 74, 87, 86, 85, 87, 78, 74, 26, 24, 
    18, 10, 8, 15, 20, 19, 19, 25, 19, 18, 26, 25, 32, 21, 21, 
    20, 2, 0, 16, 22, 23, 27, 27, 26, 21, 25, 28, 21, 25, 26, 
    27, 27, 36, 0, 0, 19, 28, 27, 26, 23, 23, 20, 20, 20, 22, 
    29, 23, 20, 46, 18, 0, 10, 28, 27, 26, 26, 23, 23, 22, 20, 
    31, 28, 29, 26, 5, 22, 20, 0, 0, 7, 24, 30, 25, 21, 20, 
    34, 33, 31, 19, 0, 5, 16, 26, 27, 7, 0, 0, 0, 11, 25, 
    32, 33, 31, 32, 58, 63, 61, 69, 64, 47, 66, 59, 62, 50, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 13, 8, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 11, 7, 10, 10, 10, 11, 11, 8, 9, 9, 9, 11, 14, 15, 
    14, 13, 12, 14, 14, 23, 22, 24, 22, 22, 14, 13, 19, 0, 0, 
    
    -- channel=101
    0, 0, 38, 6, 0, 2, 9, 0, 10, 4, 3, 5, 0, 0, 0, 
    0, 0, 5, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 20, 12, 0, 14, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 24, 24, 0, 0, 14, 0, 3, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 4, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 9, 4, 0, 3, 9, 5, 0, 0, 0, 0, 0, 
    0, 48, 73, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 10, 103, 48, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 159, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 18, 142, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 44, 48, 134, 32, 0, 47, 76, 36, 61, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 3, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    19, 4, 1, 0, 4, 0, 11, 1, 13, 10, 9, 3, 0, 0, 24, 
    
    -- channel=102
    197, 220, 194, 178, 193, 200, 197, 190, 191, 193, 198, 195, 198, 218, 228, 
    198, 227, 222, 158, 161, 182, 179, 177, 184, 190, 190, 186, 232, 232, 233, 
    197, 223, 217, 161, 165, 154, 141, 153, 167, 168, 171, 175, 224, 234, 238, 
    194, 219, 206, 142, 159, 161, 159, 159, 166, 167, 163, 178, 174, 230, 234, 
    207, 217, 216, 205, 187, 186, 184, 189, 196, 191, 187, 202, 221, 228, 232, 
    222, 219, 211, 223, 206, 204, 209, 215, 211, 208, 209, 217, 229, 227, 229, 
    227, 206, 143, 138, 209, 234, 229, 233, 231, 229, 228, 231, 230, 232, 235, 
    233, 240, 220, 157, 82, 155, 229, 241, 233, 228, 225, 227, 228, 226, 228, 
    236, 244, 241, 231, 122, 72, 100, 160, 212, 230, 228, 228, 227, 227, 230, 
    237, 239, 242, 237, 133, 43, 59, 69, 77, 92, 122, 186, 220, 231, 231, 
    233, 235, 238, 223, 130, 76, 44, 75, 127, 70, 81, 60, 113, 175, 208, 
    212, 221, 218, 215, 213, 200, 178, 194, 206, 193, 194, 195, 197, 200, 203, 
    114, 118, 112, 107, 103, 102, 101, 113, 122, 119, 121, 121, 128, 128, 122, 
    69, 72, 71, 62, 58, 53, 51, 53, 54, 44, 41, 43, 42, 42, 57, 
    44, 43, 43, 41, 40, 41, 40, 40, 42, 37, 36, 39, 48, 74, 94, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 31, 37, 44, 34, 43, 41, 35, 16, 2, 0, 0, 
    0, 0, 0, 33, 41, 29, 41, 31, 29, 30, 32, 22, 2, 0, 0, 
    0, 0, 9, 38, 20, 14, 26, 23, 21, 35, 24, 30, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 63, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 82, 0, 0, 6, 7, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 4, 29, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 4, 8, 8, 6, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 2, 0, 0, 9, 3, 
    16, 9, 11, 6, 10, 8, 4, 4, 5, 6, 1, 1, 1, 0, 0, 
    14, 3, 1, 0, 4, 1, 2, 0, 4, 0, 0, 1, 0, 0, 0, 
    
    -- channel=104
    0, 0, 9, 1, 0, 3, 6, 1, 8, 5, 5, 1, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 9, 0, 0, 0, 
    14, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 22, 18, 15, 13, 16, 16, 13, 7, 0, 0, 0, 
    3, 24, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 84, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 41, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 70, 137, 89, 62, 103, 87, 108, 96, 54, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 2, 8, 7, 8, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 6, 12, 12, 14, 13, 19, 44, 
    14, 16, 16, 17, 16, 27, 32, 29, 35, 34, 28, 22, 33, 51, 12, 
    
    -- channel=105
    0, 0, 0, 2, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 8, 3, 4, 4, 6, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 4, 3, 0, 0, 0, 0, 
    2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 1, 8, 10, 12, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 5, 7, 0, 12, 10, 2, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 1, 7, 14, 20, 20, 24, 21, 9, 0, 0, 0, 0, 0, 
    6, 2, 1, 6, 33, 19, 24, 21, 21, 27, 23, 28, 22, 8, 0, 
    5, 0, 1, 9, 1, 0, 0, 0, 0, 3, 0, 1, 0, 0, 0, 
    15, 12, 18, 20, 20, 25, 9, 1, 5, 0, 0, 0, 0, 0, 0, 
    10, 4, 4, 9, 12, 13, 7, 6, 13, 13, 14, 15, 16, 16, 16, 
    29, 27, 27, 29, 33, 30, 28, 29, 31, 32, 30, 29, 29, 29, 34, 
    29, 26, 25, 27, 30, 27, 23, 27, 28, 27, 26, 33, 30, 27, 38, 
    
    -- channel=106
    125, 139, 111, 110, 117, 125, 123, 120, 121, 122, 126, 119, 130, 146, 146, 
    126, 138, 144, 93, 112, 113, 102, 110, 112, 116, 114, 113, 153, 146, 147, 
    124, 135, 136, 86, 107, 101, 88, 99, 106, 113, 109, 108, 144, 149, 152, 
    123, 137, 133, 86, 104, 103, 97, 104, 104, 106, 111, 123, 109, 146, 143, 
    137, 136, 134, 114, 100, 96, 101, 107, 106, 102, 103, 128, 137, 146, 144, 
    153, 130, 101, 153, 143, 143, 147, 149, 145, 144, 144, 141, 144, 145, 149, 
    155, 135, 81, 24, 93, 146, 150, 153, 153, 148, 146, 145, 143, 142, 141, 
    161, 158, 162, 136, 9, 49, 125, 153, 145, 142, 143, 144, 146, 143, 142, 
    165, 163, 158, 157, 38, 23, 11, 33, 87, 123, 141, 147, 143, 142, 143, 
    165, 155, 156, 135, 18, 0, 10, 26, 13, 0, 0, 41, 95, 132, 146, 
    158, 150, 153, 152, 136, 86, 55, 104, 139, 72, 109, 65, 119, 128, 132, 
    85, 75, 66, 60, 55, 60, 65, 74, 67, 73, 76, 85, 79, 72, 77, 
    53, 58, 52, 48, 45, 44, 43, 39, 38, 33, 30, 28, 31, 31, 19, 
    0, 1, 2, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 1, 37, 
    0, 0, 0, 0, 0, 15, 12, 15, 15, 12, 3, 2, 19, 47, 15, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 24, 55, 54, 45, 51, 50, 51, 24, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 10, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 76, 84, 17, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 1, 80, 57, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 61, 114, 105, 58, 6, 0, 0, 0, 0, 
    0, 0, 0, 25, 62, 22, 11, 0, 20, 80, 121, 141, 104, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    102, 115, 127, 133, 137, 111, 78, 77, 87, 55, 59, 40, 52, 60, 59, 
    3, 0, 0, 2, 6, 9, 12, 34, 54, 61, 69, 75, 81, 85, 84, 
    42, 43, 40, 28, 27, 24, 19, 17, 12, 10, 5, 5, 5, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    
    -- channel=108
    60, 77, 72, 54, 56, 62, 59, 57, 57, 58, 58, 57, 55, 57, 58, 
    69, 83, 78, 30, 14, 15, 14, 13, 14, 15, 18, 18, 55, 62, 60, 
    69, 82, 78, 16, 23, 16, 8, 5, 21, 24, 21, 23, 46, 66, 63, 
    70, 81, 74, 13, 26, 32, 29, 29, 31, 31, 24, 35, 31, 66, 68, 
    72, 81, 78, 73, 64, 64, 64, 63, 64, 63, 59, 61, 64, 70, 71, 
    67, 76, 70, 69, 71, 69, 68, 68, 68, 68, 66, 68, 72, 68, 69, 
    62, 74, 63, 55, 54, 65, 71, 72, 70, 69, 68, 69, 69, 69, 69, 
    63, 73, 62, 44, 42, 49, 53, 63, 67, 65, 65, 67, 69, 70, 73, 
    61, 63, 62, 58, 46, 27, 32, 43, 45, 53, 61, 68, 70, 70, 71, 
    56, 58, 60, 62, 43, 26, 21, 18, 25, 41, 49, 47, 45, 54, 65, 
    56, 62, 63, 62, 39, 40, 40, 31, 37, 35, 36, 37, 41, 52, 62, 
    49, 56, 53, 53, 53, 53, 49, 54, 67, 64, 66, 65, 71, 76, 73, 
    37, 47, 48, 44, 40, 40, 42, 48, 52, 51, 51, 53, 54, 55, 51, 
    23, 31, 31, 26, 21, 23, 24, 22, 22, 20, 20, 20, 20, 22, 28, 
    13, 22, 22, 19, 18, 19, 20, 16, 17, 17, 17, 15, 20, 38, 38, 
    
    -- channel=109
    60, 66, 64, 49, 51, 54, 53, 54, 58, 56, 56, 54, 60, 63, 62, 
    66, 71, 64, 13, 12, 0, 0, 3, 1, 4, 3, 17, 56, 57, 61, 
    64, 72, 59, 0, 11, 18, 7, 13, 21, 26, 30, 35, 45, 64, 63, 
    68, 72, 37, 15, 22, 29, 21, 22, 25, 11, 15, 20, 48, 61, 62, 
    71, 72, 67, 50, 44, 41, 47, 47, 45, 41, 44, 54, 64, 66, 67, 
    67, 66, 44, 61, 82, 79, 79, 76, 76, 77, 76, 74, 63, 65, 71, 
    66, 66, 57, 8, 4, 50, 66, 67, 68, 66, 64, 63, 63, 60, 60, 
    67, 69, 71, 79, 42, 5, 19, 55, 60, 58, 62, 63, 66, 66, 68, 
    65, 64, 64, 58, 32, 14, 3, 0, 0, 26, 51, 65, 64, 63, 66, 
    60, 59, 61, 51, 0, 0, 4, 12, 11, 0, 0, 0, 0, 34, 60, 
    58, 58, 61, 47, 84, 94, 66, 84, 95, 85, 90, 80, 85, 77, 61, 
    7, 0, 0, 0, 0, 0, 13, 18, 9, 19, 27, 29, 34, 23, 23, 
    32, 33, 35, 30, 30, 28, 30, 25, 12, 9, 5, 4, 1, 0, 0, 
    0, 0, 0, 0, 0, 1, 3, 5, 6, 7, 8, 9, 9, 12, 57, 
    8, 11, 10, 12, 9, 21, 22, 22, 24, 25, 19, 14, 29, 68, 23, 
    
    -- channel=110
    11, 34, 50, 31, 22, 35, 40, 26, 32, 32, 35, 35, 18, 28, 33, 
    19, 33, 40, 50, 31, 34, 47, 28, 39, 40, 39, 9, 34, 41, 39, 
    16, 38, 54, 13, 20, 7, 11, 0, 6, 17, 12, 9, 23, 39, 38, 
    22, 34, 53, 10, 22, 17, 18, 18, 26, 41, 24, 34, 7, 42, 42, 
    36, 34, 33, 63, 38, 38, 33, 34, 43, 44, 35, 9, 38, 39, 40, 
    34, 52, 48, 20, 23, 17, 17, 25, 26, 23, 19, 30, 40, 40, 36, 
    31, 56, 61, 57, 18, 28, 37, 42, 39, 44, 38, 42, 43, 45, 43, 
    29, 44, 26, 25, 36, 14, 11, 39, 49, 46, 38, 41, 39, 41, 40, 
    29, 40, 42, 44, 101, 0, 19, 42, 34, 40, 27, 43, 45, 42, 40, 
    29, 42, 44, 82, 124, 0, 0, 0, 7, 59, 41, 51, 31, 27, 36, 
    30, 42, 44, 65, 0, 9, 0, 0, 0, 0, 0, 0, 0, 6, 33, 
    51, 71, 77, 77, 75, 70, 30, 33, 75, 46, 50, 39, 56, 67, 59, 
    5, 6, 8, 3, 0, 0, 0, 8, 30, 22, 28, 28, 31, 39, 33, 
    22, 15, 17, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    
    -- channel=111
    63, 76, 75, 55, 62, 64, 62, 61, 63, 62, 62, 61, 64, 68, 69, 
    69, 79, 78, 32, 27, 32, 30, 29, 31, 35, 36, 37, 76, 69, 71, 
    67, 78, 67, 39, 40, 39, 25, 38, 45, 42, 46, 49, 60, 72, 73, 
    71, 79, 59, 39, 42, 44, 44, 37, 47, 36, 35, 45, 51, 70, 74, 
    76, 78, 77, 67, 58, 57, 60, 59, 60, 57, 54, 63, 75, 74, 78, 
    73, 70, 59, 79, 84, 82, 82, 83, 83, 81, 78, 78, 75, 75, 77, 
    69, 85, 57, 6, 33, 72, 78, 79, 79, 77, 74, 75, 73, 71, 73, 
    69, 78, 78, 83, 27, 10, 46, 71, 73, 72, 71, 74, 76, 76, 78, 
    66, 71, 72, 69, 54, 11, 0, 0, 21, 51, 70, 77, 75, 74, 77, 
    62, 65, 71, 57, 35, 0, 5, 13, 11, 0, 0, 0, 26, 57, 75, 
    60, 69, 70, 73, 83, 81, 48, 53, 78, 66, 70, 57, 54, 67, 65, 
    24, 28, 22, 19, 18, 25, 33, 38, 41, 51, 48, 56, 56, 53, 54, 
    36, 42, 42, 36, 31, 33, 34, 32, 29, 25, 24, 21, 22, 22, 18, 
    6, 3, 4, 3, 0, 2, 4, 3, 3, 2, 1, 2, 4, 8, 27, 
    8, 6, 8, 5, 5, 12, 14, 11, 12, 12, 8, 3, 18, 27, 7, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 92, 46, 93, 151, 60, 66, 110, 75, 94, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 73, 
    0, 0, 0, 0, 0, 16, 3, 14, 3, 9, 0, 0, 43, 25, 0, 
    
    -- channel=113
    6, 8, 23, 11, 19, 29, 31, 29, 31, 34, 29, 30, 20, 5, 5, 
    8, 5, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 
    6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 
    9, 7, 13, 63, 44, 43, 41, 56, 60, 57, 55, 49, 51, 12, 13, 
    7, 9, 0, 9, 18, 19, 19, 14, 10, 15, 23, 5, 13, 2, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 13, 12, 
    8, 40, 62, 32, 0, 0, 8, 6, 2, 0, 0, 0, 3, 5, 11, 
    6, 5, 0, 0, 37, 0, 0, 0, 11, 9, 8, 6, 5, 9, 12, 
    1, 1, 3, 0, 4, 9, 39, 0, 0, 0, 0, 9, 8, 6, 7, 
    3, 8, 7, 0, 7, 12, 0, 0, 35, 64, 34, 0, 0, 0, 0, 
    8, 10, 8, 27, 12, 47, 75, 28, 12, 40, 30, 69, 26, 32, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 28, 21, 18, 19, 21, 15, 12, 7, 10, 7, 3, 6, 19, 17, 
    9, 7, 6, 7, 7, 10, 8, 8, 12, 8, 0, 0, 22, 0, 0, 
    
    -- channel=114
    29, 32, 25, 26, 29, 28, 27, 28, 29, 30, 30, 30, 33, 38, 42, 
    35, 41, 33, 21, 37, 51, 46, 49, 48, 47, 48, 46, 44, 45, 47, 
    33, 40, 43, 16, 2, 2, 5, 6, 3, 5, 7, 20, 45, 45, 48, 
    31, 37, 22, 0, 15, 17, 3, 13, 20, 15, 18, 14, 36, 46, 48, 
    31, 37, 32, 22, 22, 24, 26, 27, 28, 23, 24, 34, 35, 44, 45, 
    35, 39, 41, 28, 23, 22, 27, 27, 25, 25, 26, 39, 41, 42, 45, 
    40, 25, 5, 40, 46, 44, 44, 45, 43, 41, 43, 42, 43, 45, 47, 
    46, 47, 21, 0, 0, 40, 49, 48, 45, 41, 41, 41, 40, 40, 42, 
    49, 51, 48, 36, 0, 0, 17, 45, 48, 45, 45, 42, 43, 43, 44, 
    47, 50, 49, 45, 0, 0, 0, 0, 0, 9, 37, 44, 47, 45, 44, 
    48, 46, 50, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 40, 
    48, 46, 48, 47, 48, 24, 15, 33, 38, 20, 28, 18, 31, 36, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 7, 10, 8, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 7, 0, 9, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 2, 6, 9, 
    0, 0, 1, 2, 3, 0, 1, 3, 4, 4, 4, 6, 9, 17, 28, 
    
    -- channel=116
    0, 0, 36, 1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 59, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 25, 12, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 12, 0, 0, 13, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 34, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 11, 4, 0, 3, 0, 0, 0, 6, 1, 0, 0, 0, 0, 0, 
    0, 44, 69, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 24, 100, 46, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 197, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 41, 107, 0, 0, 22, 50, 2, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 0, 0, 1, 6, 0, 0, 0, 0, 0, 
    0, 3, 12, 9, 6, 8, 0, 0, 12, 0, 3, 0, 0, 7, 0, 
    18, 1, 8, 0, 12, 4, 2, 0, 8, 11, 1, 4, 2, 0, 0, 
    27, 5, 5, 0, 7, 0, 9, 0, 9, 7, 12, 7, 0, 0, 29, 
    
    -- channel=117
    46, 11, 0, 0, 21, 0, 0, 6, 1, 4, 1, 0, 19, 14, 9, 
    42, 18, 0, 0, 16, 2, 0, 7, 0, 0, 0, 21, 20, 3, 8, 
    39, 15, 0, 0, 0, 20, 0, 29, 11, 1, 13, 31, 29, 5, 9, 
    30, 15, 0, 7, 11, 7, 0, 18, 11, 0, 8, 0, 60, 4, 10, 
    9, 15, 0, 0, 2, 3, 3, 7, 0, 0, 6, 35, 9, 4, 8, 
    6, 0, 0, 3, 2, 8, 13, 4, 0, 2, 8, 18, 1, 1, 10, 
    17, 0, 0, 18, 44, 16, 7, 1, 0, 0, 4, 0, 1, 1, 7, 
    28, 0, 0, 0, 0, 69, 46, 5, 0, 0, 3, 0, 1, 0, 8, 
    27, 5, 0, 0, 0, 18, 44, 37, 24, 6, 18, 0, 0, 0, 6, 
    25, 5, 0, 0, 0, 5, 18, 11, 13, 0, 46, 19, 24, 16, 10, 
    32, 1, 1, 0, 0, 0, 16, 93, 0, 0, 18, 0, 99, 35, 20, 
    23, 0, 0, 0, 0, 0, 1, 35, 0, 0, 4, 0, 7, 0, 2, 
    11, 0, 0, 0, 0, 0, 6, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 2, 8, 49, 
    0, 0, 0, 6, 0, 12, 0, 12, 0, 1, 0, 1, 29, 39, 0, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 38, 15, 0, 0, 19, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 33, 31, 19, 29, 16, 23, 19, 10, 1, 0, 0, 0, 
    0, 0, 12, 38, 13, 6, 28, 12, 9, 27, 15, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 81, 0, 1, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 28, 44, 0, 0, 18, 12, 11, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 1, 1, 8, 4, 4, 4, 10, 11, 8, 9, 7, 8, 0, 
    17, 8, 9, 6, 12, 4, 9, 5, 9, 7, 9, 12, 2, 0, 0, 
    
    -- channel=120
    43, 28, 0, 7, 29, 9, 0, 11, 0, 5, 5, 8, 18, 18, 25, 
    44, 46, 17, 0, 33, 61, 48, 57, 51, 53, 56, 71, 36, 32, 32, 
    47, 40, 22, 19, 0, 0, 0, 0, 0, 0, 0, 0, 57, 32, 34, 
    32, 38, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 32, 36, 39, 
    13, 33, 24, 0, 21, 26, 24, 22, 28, 19, 22, 47, 14, 30, 34, 
    23, 31, 63, 31, 0, 0, 5, 2, 0, 3, 7, 19, 29, 23, 27, 
    30, 0, 0, 88, 145, 62, 28, 24, 22, 19, 31, 30, 33, 36, 41, 
    40, 23, 0, 0, 0, 136, 124, 42, 26, 25, 27, 25, 25, 23, 30, 
    42, 34, 28, 10, 0, 10, 65, 142, 142, 84, 56, 20, 24, 30, 33, 
    42, 33, 31, 17, 0, 19, 18, 1, 8, 44, 142, 163, 141, 81, 38, 
    47, 30, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    121, 116, 120, 126, 133, 99, 86, 99, 89, 68, 75, 62, 62, 74, 81, 
    8, 7, 0, 6, 9, 11, 17, 40, 39, 55, 56, 67, 72, 64, 73, 
    10, 27, 20, 19, 7, 7, 8, 8, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    
    -- channel=121
    18, 0, 0, 0, 8, 0, 0, 8, 5, 6, 2, 2, 16, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 1, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 16, 6, 5, 2, 10, 5, 0, 5, 0, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 11, 1, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 57, 12, 65, 111, 34, 46, 63, 53, 80, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 6, 6, 7, 6, 7, 12, 10, 11, 25, 75, 
    7, 12, 11, 13, 14, 32, 17, 28, 21, 23, 11, 11, 51, 37, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    43, 56, 32, 37, 40, 39, 34, 33, 31, 33, 35, 36, 39, 54, 53, 
    44, 56, 53, 48, 56, 77, 67, 70, 76, 75, 71, 67, 60, 60, 58, 
    43, 49, 65, 54, 52, 39, 47, 46, 47, 51, 45, 44, 74, 56, 60, 
    41, 51, 56, 10, 31, 32, 22, 33, 30, 33, 33, 42, 29, 57, 57, 
    40, 49, 48, 48, 38, 39, 34, 41, 46, 38, 38, 50, 54, 57, 55, 
    49, 55, 64, 51, 42, 43, 49, 52, 48, 47, 47, 53, 54, 51, 52, 
    50, 25, 0, 35, 73, 65, 57, 58, 56, 56, 58, 58, 58, 60, 59, 
    55, 57, 42, 0, 0, 53, 80, 63, 57, 54, 53, 54, 55, 53, 54, 
    58, 61, 59, 53, 0, 0, 10, 49, 76, 74, 65, 56, 55, 55, 55, 
    59, 59, 58, 56, 0, 0, 0, 0, 0, 0, 28, 63, 77, 72, 59, 
    59, 59, 59, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 45, 
    79, 82, 78, 76, 77, 61, 63, 73, 67, 54, 66, 58, 67, 64, 62, 
    8, 13, 12, 13, 10, 9, 14, 25, 24, 25, 26, 27, 30, 31, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 47, 69, 57, 64, 62, 60, 57, 47, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 79, 108, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 112, 76, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 58, 131, 115, 47, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 17, 0, 3, 54, 137, 150, 107, 36, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    90, 91, 98, 105, 112, 84, 60, 63, 63, 40, 41, 27, 26, 44, 47, 
    0, 0, 0, 0, 0, 2, 7, 29, 40, 54, 57, 69, 74, 72, 74, 
    16, 33, 29, 22, 12, 12, 12, 10, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    
    -- channel=125
    0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 55, 63, 65, 61, 66, 59, 62, 47, 1, 0, 0, 
    0, 0, 8, 57, 23, 11, 29, 20, 10, 11, 6, 7, 12, 0, 0, 
    0, 0, 16, 23, 20, 17, 13, 17, 22, 35, 27, 18, 8, 0, 0, 
    0, 0, 0, 9, 9, 12, 8, 8, 12, 10, 5, 0, 0, 0, 0, 
    0, 3, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 13, 51, 40, 5, 0, 1, 0, 1, 0, 0, 0, 2, 2, 
    0, 0, 0, 0, 17, 35, 18, 2, 5, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 40, 15, 29, 58, 45, 22, 5, 1, 2, 1, 1, 
    0, 0, 0, 13, 76, 30, 18, 14, 18, 56, 68, 67, 36, 10, 2, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    30, 48, 50, 53, 55, 55, 24, 20, 46, 34, 26, 25, 24, 42, 38, 
    8, 16, 12, 10, 6, 11, 13, 20, 40, 41, 44, 48, 51, 57, 58, 
    38, 45, 43, 32, 30, 30, 28, 24, 19, 16, 13, 11, 12, 2, 0, 
    17, 12, 13, 10, 11, 3, 6, 0, 2, 1, 6, 5, 0, 0, 4, 
    
    -- channel=126
    43, 45, 38, 33, 45, 42, 43, 46, 48, 49, 47, 43, 54, 50, 47, 
    45, 48, 45, 4, 11, 2, 0, 6, 1, 1, 2, 15, 50, 43, 45, 
    43, 47, 33, 0, 12, 15, 0, 18, 16, 16, 19, 24, 35, 47, 46, 
    46, 48, 35, 25, 26, 31, 24, 29, 33, 23, 31, 28, 50, 42, 46, 
    51, 50, 46, 21, 21, 18, 29, 33, 20, 21, 24, 48, 40, 49, 47, 
    51, 28, 0, 52, 60, 57, 59, 56, 52, 52, 55, 51, 48, 50, 56, 
    54, 55, 40, 0, 0, 37, 55, 54, 53, 47, 46, 42, 41, 40, 41, 
    57, 55, 54, 54, 0, 0, 4, 45, 45, 40, 45, 44, 48, 47, 48, 
    58, 53, 50, 44, 0, 0, 0, 0, 0, 0, 39, 51, 47, 44, 47, 
    54, 45, 47, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 45, 
    51, 47, 48, 39, 92, 69, 71, 105, 84, 67, 89, 73, 96, 68, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    
    -- channel=127
    34, 47, 39, 29, 26, 30, 27, 24, 24, 24, 27, 25, 24, 35, 35, 
    44, 52, 49, 2, 9, 6, 6, 5, 8, 12, 11, 4, 35, 36, 35, 
    42, 53, 55, 1, 2, 0, 0, 0, 2, 10, 9, 14, 26, 41, 37, 
    43, 51, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 42, 
    44, 50, 48, 46, 35, 36, 33, 34, 39, 33, 30, 31, 39, 45, 44, 
    41, 59, 54, 38, 45, 43, 43, 42, 43, 44, 40, 46, 43, 39, 41, 
    36, 29, 27, 38, 40, 39, 41, 43, 42, 44, 43, 45, 45, 44, 43, 
    37, 43, 35, 21, 28, 37, 36, 36, 40, 40, 39, 41, 43, 43, 45, 
    37, 38, 38, 30, 33, 10, 13, 34, 41, 39, 33, 41, 43, 44, 44, 
    33, 35, 36, 53, 22, 7, 4, 2, 4, 14, 29, 46, 40, 37, 39, 
    31, 37, 38, 22, 0, 4, 0, 0, 9, 0, 0, 0, 10, 22, 35, 
    49, 57, 55, 54, 53, 52, 53, 48, 51, 55, 53, 54, 53, 53, 54, 
    21, 26, 30, 29, 30, 29, 32, 36, 40, 39, 38, 40, 40, 40, 33, 
    2, 7, 7, 2, 1, 1, 4, 2, 3, 1, 0, 2, 1, 0, 0, 
    0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 27, 30, 
    
    -- channel=128
    19, 23, 39, 5, 0, 9, 14, 0, 0, 0, 0, 2, 7, 0, 10, 
    16, 43, 9, 6, 0, 0, 0, 14, 5, 19, 0, 12, 22, 71, 28, 
    0, 0, 0, 0, 0, 30, 65, 20, 0, 0, 0, 29, 24, 24, 22, 
    0, 37, 35, 0, 19, 50, 0, 0, 17, 5, 48, 34, 0, 18, 0, 
    13, 4, 29, 12, 21, 20, 0, 53, 39, 51, 15, 0, 2, 4, 0, 
    0, 0, 0, 65, 58, 2, 23, 46, 32, 1, 0, 45, 0, 0, 0, 
    30, 15, 0, 11, 5, 1, 28, 22, 0, 0, 16, 30, 0, 16, 3, 
    0, 0, 20, 0, 26, 23, 0, 18, 26, 60, 40, 0, 43, 0, 0, 
    25, 42, 0, 0, 0, 30, 26, 5, 24, 0, 0, 19, 0, 0, 1, 
    20, 0, 0, 0, 0, 0, 11, 30, 13, 13, 4, 5, 0, 7, 12, 
    0, 0, 17, 3, 36, 9, 2, 15, 8, 0, 0, 0, 12, 14, 41, 
    56, 128, 83, 41, 0, 8, 6, 0, 0, 7, 20, 8, 0, 1, 0, 
    0, 0, 12, 65, 30, 1, 0, 0, 0, 3, 6, 3, 0, 0, 0, 
    0, 0, 0, 0, 60, 38, 2, 18, 56, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 65, 50, 19, 0, 0, 0, 0, 56, 44, 61, 
    
    -- channel=129
    0, 0, 0, 4, 7, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 
    0, 0, 1, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 10, 4, 10, 5, 0, 0, 3, 6, 8, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 1, 8, 0, 0, 0, 0, 7, 2, 13, 
    6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 10, 17, 
    14, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 7, 
    1, 0, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 
    7, 0, 1, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 
    0, 0, 19, 14, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 5, 
    11, 16, 12, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 
    21, 18, 0, 0, 0, 7, 0, 0, 4, 0, 0, 0, 0, 8, 17, 
    0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    7, 0, 0, 1, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    
    -- channel=130
    0, 0, 0, 0, 0, 39, 0, 22, 13, 24, 0, 66, 0, 44, 0, 
    0, 0, 0, 0, 0, 41, 5, 25, 0, 12, 0, 83, 0, 17, 0, 
    4, 17, 0, 0, 0, 16, 0, 0, 23, 0, 9, 80, 0, 0, 0, 
    0, 26, 0, 0, 0, 22, 0, 0, 36, 0, 22, 49, 0, 0, 0, 
    0, 58, 0, 0, 40, 5, 0, 16, 0, 8, 0, 58, 0, 0, 0, 
    0, 72, 0, 0, 17, 20, 0, 29, 0, 11, 0, 51, 0, 5, 0, 
    0, 37, 37, 0, 8, 43, 20, 30, 24, 39, 33, 33, 0, 7, 0, 
    0, 27, 12, 0, 11, 23, 56, 32, 29, 20, 24, 58, 0, 7, 0, 
    0, 4, 9, 10, 61, 0, 54, 38, 34, 41, 26, 46, 11, 24, 0, 
    0, 5, 0, 21, 16, 79, 31, 32, 35, 21, 31, 20, 0, 0, 13, 
    0, 26, 0, 16, 3, 0, 76, 27, 19, 23, 38, 23, 0, 2, 0, 
    0, 0, 0, 11, 0, 24, 53, 41, 32, 4, 32, 29, 16, 33, 0, 
    48, 91, 0, 0, 0, 31, 41, 36, 90, 24, 43, 11, 1, 48, 0, 
    0, 80, 102, 11, 0, 0, 12, 0, 44, 51, 36, 14, 0, 33, 1, 
    0, 0, 99, 100, 15, 0, 0, 0, 14, 52, 64, 20, 0, 0, 66, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 11, 14, 5, 
    0, 0, 0, 0, 0, 9, 12, 0, 0, 0, 0, 5, 3, 0, 0, 
    0, 7, 0, 0, 0, 7, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 27, 7, 0, 4, 17, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 0, 0, 1, 49, 15, 0, 0, 14, 0, 0, 0, 
    6, 0, 0, 1, 3, 20, 22, 0, 0, 5, 24, 11, 0, 0, 0, 
    0, 0, 0, 0, 52, 0, 4, 1, 46, 29, 0, 4, 20, 0, 0, 
    4, 1, 0, 0, 0, 62, 3, 16, 13, 0, 0, 10, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 42, 23, 0, 17, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 0, 15, 11, 0, 7, 0, 0, 0, 3, 
    27, 64, 27, 0, 0, 0, 16, 0, 0, 3, 21, 0, 0, 0, 0, 
    0, 0, 31, 18, 3, 0, 6, 0, 0, 17, 0, 8, 0, 0, 0, 
    0, 0, 0, 15, 23, 9, 0, 10, 1, 0, 11, 0, 0, 0, 21, 
    0, 18, 0, 0, 15, 38, 10, 0, 0, 0, 0, 0, 9, 5, 0, 
    
    -- channel=132
    6, 1, 4, 0, 0, 7, 0, 0, 0, 0, 0, 18, 0, 6, 10, 
    4, 6, 0, 0, 0, 0, 0, 10, 0, 0, 0, 27, 8, 21, 0, 
    0, 0, 0, 0, 0, 22, 8, 0, 0, 0, 6, 27, 12, 3, 0, 
    0, 26, 0, 5, 10, 9, 0, 0, 18, 5, 26, 21, 0, 7, 0, 
    0, 14, 1, 0, 24, 1, 0, 26, 1, 14, 0, 0, 9, 1, 0, 
    0, 5, 0, 11, 17, 30, 23, 28, 14, 18, 14, 33, 0, 0, 0, 
    1, 11, 0, 3, 27, 54, 63, 56, 43, 47, 54, 59, 15, 2, 0, 
    0, 8, 14, 1, 59, 38, 64, 57, 66, 78, 63, 51, 54, 10, 0, 
    9, 8, 0, 0, 17, 62, 55, 58, 72, 68, 53, 58, 18, 0, 0, 
    0, 0, 0, 1, 11, 7, 60, 70, 57, 60, 58, 51, 37, 16, 6, 
    0, 19, 0, 2, 1, 24, 51, 57, 61, 47, 58, 57, 41, 10, 4, 
    31, 58, 23, 3, 0, 12, 52, 62, 53, 46, 69, 58, 36, 21, 0, 
    0, 4, 26, 17, 5, 0, 24, 23, 34, 59, 54, 57, 41, 5, 0, 
    0, 0, 9, 23, 17, 11, 7, 16, 39, 54, 61, 42, 6, 5, 6, 
    0, 7, 0, 11, 19, 25, 10, 15, 10, 26, 21, 31, 27, 21, 40, 
    
    -- channel=133
    2, 29, 0, 0, 53, 0, 5, 0, 0, 0, 30, 0, 96, 0, 0, 
    9, 29, 11, 0, 63, 0, 0, 0, 0, 0, 28, 0, 81, 0, 23, 
    6, 0, 0, 9, 55, 0, 0, 12, 0, 44, 0, 0, 41, 6, 3, 
    30, 0, 26, 32, 7, 0, 21, 40, 0, 36, 0, 0, 0, 0, 57, 
    39, 0, 61, 20, 0, 0, 81, 0, 0, 0, 4, 0, 3, 0, 102, 
    59, 0, 0, 94, 0, 0, 11, 0, 23, 6, 14, 0, 29, 0, 111, 
    53, 0, 0, 9, 20, 0, 11, 8, 0, 0, 0, 12, 10, 0, 86, 
    32, 0, 0, 0, 1, 44, 0, 0, 11, 18, 19, 0, 61, 0, 94, 
    0, 0, 0, 0, 0, 43, 0, 0, 14, 0, 0, 5, 4, 10, 62, 
    0, 14, 25, 0, 0, 0, 10, 0, 0, 16, 8, 11, 45, 11, 0, 
    57, 0, 37, 0, 4, 30, 0, 8, 10, 7, 3, 5, 24, 0, 0, 
    0, 3, 72, 0, 8, 0, 0, 0, 0, 28, 0, 6, 25, 0, 1, 
    0, 0, 20, 43, 36, 0, 0, 16, 0, 0, 0, 36, 29, 0, 0, 
    35, 0, 0, 0, 55, 22, 0, 19, 0, 0, 0, 29, 64, 0, 0, 
    40, 25, 0, 0, 0, 48, 35, 10, 1, 0, 0, 7, 51, 8, 0, 
    
    -- channel=134
    64, 16, 44, 55, 30, 11, 53, 41, 77, 81, 80, 61, 97, 37, 46, 
    75, 43, 68, 65, 20, 16, 44, 34, 79, 64, 78, 68, 112, 47, 87, 
    84, 77, 69, 57, 14, 11, 45, 65, 76, 51, 74, 78, 152, 98, 110, 
    49, 60, 66, 55, 3, 69, 90, 33, 42, 55, 72, 100, 174, 124, 126, 
    53, 111, 120, 41, 62, 99, 64, 20, 85, 84, 117, 100, 149, 138, 98, 
    53, 107, 149, 76, 73, 92, 77, 111, 107, 103, 95, 89, 145, 140, 85, 
    55, 85, 122, 143, 103, 98, 89, 94, 98, 105, 105, 105, 125, 125, 90, 
    75, 94, 111, 143, 137, 59, 109, 115, 117, 99, 97, 143, 127, 131, 68, 
    86, 99, 112, 120, 127, 139, 105, 129, 128, 134, 125, 126, 137, 111, 75, 
    113, 109, 84, 103, 120, 115, 139, 145, 140, 155, 122, 129, 112, 69, 72, 
    103, 87, 77, 91, 82, 105, 131, 166, 162, 139, 132, 123, 103, 88, 124, 
    94, 130, 102, 90, 120, 98, 144, 162, 157, 132, 136, 124, 107, 110, 126, 
    130, 181, 177, 125, 108, 124, 142, 137, 132, 146, 144, 122, 99, 67, 117, 
    82, 53, 157, 176, 134, 111, 115, 105, 75, 145, 145, 119, 86, 64, 101, 
    82, 32, 40, 161, 191, 150, 128, 122, 99, 129, 135, 113, 55, 60, 106, 
    
    -- channel=135
    1, 0, 0, 0, 13, 0, 0, 0, 0, 0, 16, 0, 63, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 17, 0, 58, 0, 2, 
    1, 5, 0, 0, 12, 0, 0, 0, 0, 3, 0, 0, 31, 0, 0, 
    4, 0, 0, 16, 0, 0, 4, 17, 0, 17, 0, 0, 20, 0, 39, 
    0, 0, 26, 0, 0, 0, 36, 0, 0, 0, 0, 0, 9, 0, 59, 
    13, 0, 0, 21, 0, 6, 14, 0, 2, 3, 13, 0, 19, 0, 62, 
    7, 0, 0, 0, 17, 29, 33, 18, 22, 20, 20, 10, 13, 0, 42, 
    3, 0, 0, 0, 34, 10, 21, 22, 38, 27, 22, 8, 43, 0, 34, 
    0, 0, 0, 0, 0, 60, 2, 27, 31, 32, 26, 24, 31, 14, 32, 
    0, 0, 3, 0, 8, 0, 37, 23, 20, 41, 25, 34, 53, 1, 0, 
    25, 0, 5, 0, 0, 21, 0, 31, 35, 30, 36, 36, 32, 0, 0, 
    0, 0, 21, 0, 0, 0, 9, 33, 29, 33, 32, 32, 43, 0, 0, 
    0, 0, 23, 7, 10, 0, 6, 44, 10, 34, 19, 47, 40, 0, 0, 
    19, 0, 0, 8, 15, 0, 0, 22, 0, 25, 32, 38, 59, 0, 0, 
    23, 20, 0, 0, 8, 9, 0, 4, 4, 21, 24, 37, 14, 0, 0, 
    
    -- channel=136
    46, 40, 57, 36, 39, 25, 37, 13, 22, 0, 29, 1, 59, 9, 28, 
    35, 38, 40, 34, 30, 20, 11, 22, 35, 31, 33, 6, 66, 59, 51, 
    0, 0, 22, 16, 20, 48, 69, 38, 3, 18, 18, 13, 52, 37, 37, 
    37, 54, 46, 30, 24, 63, 31, 2, 26, 31, 67, 24, 18, 28, 37, 
    34, 23, 58, 25, 22, 38, 46, 40, 61, 46, 37, 0, 24, 18, 40, 
    14, 3, 13, 73, 65, 7, 11, 42, 34, 21, 19, 14, 23, 11, 54, 
    42, 34, 0, 16, 8, 0, 24, 28, 0, 0, 7, 25, 11, 23, 37, 
    16, 21, 19, 4, 29, 6, 0, 1, 18, 40, 21, 0, 38, 14, 13, 
    30, 40, 0, 0, 0, 21, 6, 0, 16, 0, 0, 5, 0, 0, 32, 
    20, 0, 7, 1, 5, 0, 0, 14, 0, 10, 0, 3, 24, 33, 20, 
    18, 15, 37, 32, 28, 21, 0, 5, 4, 0, 0, 4, 21, 22, 50, 
    41, 99, 83, 44, 21, 9, 5, 0, 0, 1, 15, 1, 2, 10, 18, 
    0, 0, 27, 57, 45, 9, 0, 0, 0, 0, 1, 5, 17, 0, 16, 
    35, 0, 0, 13, 60, 47, 20, 40, 25, 0, 0, 0, 0, 9, 23, 
    29, 50, 0, 0, 8, 61, 57, 41, 0, 0, 0, 0, 59, 78, 44, 
    
    -- channel=137
    40, 40, 40, 46, 45, 41, 46, 44, 54, 59, 57, 40, 63, 46, 45, 
    41, 39, 49, 43, 43, 38, 49, 42, 51, 45, 60, 34, 67, 30, 45, 
    46, 57, 47, 39, 43, 47, 47, 47, 52, 42, 64, 31, 57, 48, 52, 
    50, 43, 38, 43, 40, 53, 72, 64, 44, 48, 44, 51, 60, 45, 47, 
    44, 43, 47, 37, 45, 54, 61, 42, 57, 53, 66, 66, 60, 42, 55, 
    42, 42, 55, 46, 45, 47, 36, 36, 53, 55, 58, 45, 66, 48, 53, 
    40, 37, 44, 46, 44, 39, 40, 33, 39, 33, 28, 33, 55, 47, 57, 
    50, 43, 40, 47, 32, 23, 38, 35, 35, 29, 28, 23, 35, 48, 49, 
    41, 42, 43, 52, 34, 36, 17, 27, 27, 33, 37, 28, 40, 49, 54, 
    37, 52, 49, 50, 47, 26, 33, 20, 26, 27, 30, 35, 38, 35, 51, 
    49, 47, 53, 46, 46, 44, 28, 29, 21, 31, 30, 36, 42, 41, 39, 
    43, 33, 65, 48, 49, 43, 31, 34, 27, 28, 29, 30, 51, 44, 65, 
    48, 66, 73, 74, 65, 40, 39, 38, 40, 29, 21, 33, 36, 53, 65, 
    49, 51, 82, 73, 79, 73, 67, 58, 26, 29, 30, 35, 47, 53, 75, 
    57, 59, 49, 79, 71, 72, 75, 75, 47, 40, 35, 51, 48, 48, 44, 
    
    -- channel=138
    33, 0, 21, 13, 0, 0, 14, 1, 20, 17, 21, 34, 33, 0, 11, 
    40, 6, 19, 23, 0, 0, 0, 2, 36, 20, 26, 44, 74, 42, 42, 
    0, 10, 22, 0, 0, 12, 36, 8, 24, 0, 47, 53, 100, 52, 69, 
    3, 60, 22, 11, 0, 52, 24, 0, 18, 26, 67, 58, 103, 75, 44, 
    2, 85, 74, 0, 38, 61, 13, 22, 60, 58, 58, 37, 88, 74, 16, 
    0, 64, 93, 49, 57, 59, 40, 91, 67, 62, 52, 62, 68, 79, 20, 
    12, 53, 60, 88, 56, 58, 66, 60, 50, 59, 69, 68, 66, 71, 30, 
    14, 51, 55, 79, 114, 0, 68, 77, 89, 86, 58, 95, 80, 69, 0, 
    54, 60, 33, 51, 49, 105, 65, 84, 82, 80, 74, 71, 55, 24, 26, 
    49, 24, 7, 43, 58, 40, 90, 104, 89, 99, 68, 74, 52, 22, 44, 
    23, 55, 27, 60, 30, 55, 99, 110, 103, 71, 76, 76, 56, 50, 75, 
    94, 145, 79, 47, 58, 55, 99, 107, 93, 76, 102, 71, 49, 50, 56, 
    27, 87, 125, 87, 58, 72, 75, 29, 55, 100, 91, 67, 43, 0, 42, 
    23, 0, 73, 128, 96, 66, 59, 65, 44, 85, 93, 49, 0, 12, 75, 
    19, 7, 0, 84, 131, 114, 85, 78, 32, 52, 38, 43, 32, 56, 93, 
    
    -- channel=139
    0, 0, 0, 0, 19, 0, 0, 0, 24, 26, 21, 0, 28, 13, 0, 
    0, 0, 2, 0, 12, 17, 21, 0, 0, 0, 18, 0, 0, 0, 0, 
    52, 37, 0, 16, 9, 0, 0, 13, 19, 38, 0, 0, 0, 0, 0, 
    4, 0, 0, 2, 0, 0, 34, 43, 0, 0, 0, 0, 22, 0, 52, 
    0, 0, 0, 4, 0, 0, 14, 0, 0, 0, 11, 20, 8, 0, 52, 
    23, 13, 0, 0, 0, 0, 0, 0, 0, 6, 8, 0, 20, 11, 25, 
    0, 0, 8, 0, 8, 0, 0, 0, 3, 0, 0, 0, 10, 0, 7, 
    7, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 45, 
    0, 0, 28, 22, 21, 0, 0, 0, 0, 0, 0, 0, 38, 55, 0, 
    2, 41, 25, 21, 20, 31, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 5, 0, 0, 0, 0, 13, 8, 11, 
    76, 64, 0, 0, 0, 0, 15, 75, 47, 0, 0, 0, 11, 21, 29, 
    23, 87, 71, 0, 0, 0, 0, 0, 0, 13, 0, 16, 60, 6, 0, 
    29, 0, 41, 56, 0, 0, 0, 0, 21, 41, 71, 16, 0, 0, 0, 
    
    -- channel=140
    23, 16, 20, 30, 33, 11, 17, 14, 14, 10, 23, 9, 19, 10, 13, 
    24, 15, 23, 31, 26, 12, 19, 13, 19, 17, 21, 10, 16, 18, 27, 
    25, 10, 22, 29, 19, 10, 19, 24, 18, 25, 14, 11, 23, 24, 26, 
    28, 19, 27, 20, 10, 13, 14, 10, 16, 17, 17, 9, 27, 25, 40, 
    26, 24, 34, 24, 1, 10, 13, 5, 16, 12, 13, 0, 17, 32, 42, 
    19, 24, 31, 26, 16, 5, 0, 5, 4, 0, 0, 0, 13, 36, 33, 
    21, 25, 26, 28, 0, 0, 0, 0, 0, 0, 0, 0, 3, 25, 28, 
    22, 24, 27, 29, 4, 0, 0, 0, 0, 0, 0, 3, 6, 16, 30, 
    20, 24, 27, 26, 18, 2, 0, 0, 0, 0, 0, 0, 11, 8, 19, 
    30, 22, 24, 23, 22, 21, 0, 7, 1, 3, 0, 0, 7, 22, 17, 
    31, 14, 18, 26, 22, 18, 12, 8, 10, 9, 0, 0, 1, 16, 35, 
    17, 11, 7, 21, 30, 21, 9, 0, 6, 7, 1, 0, 0, 3, 31, 
    24, 8, 0, 1, 14, 24, 15, 3, 1, 2, 7, 0, 0, 0, 29, 
    26, 6, 0, 0, 0, 7, 14, 13, 15, 5, 0, 0, 4, 11, 13, 
    24, 6, 4, 0, 2, 0, 5, 10, 7, 5, 5, 0, 11, 20, 10, 
    
    -- channel=141
    30, 26, 45, 41, 11, 32, 29, 26, 28, 16, 20, 40, 13, 10, 31, 
    40, 43, 36, 41, 9, 14, 4, 37, 29, 40, 19, 47, 25, 59, 42, 
    11, 4, 32, 26, 5, 40, 58, 37, 21, 11, 19, 55, 39, 50, 48, 
    16, 53, 42, 21, 26, 58, 33, 0, 43, 19, 53, 58, 26, 48, 16, 
    32, 55, 42, 20, 41, 46, 16, 51, 49, 55, 44, 27, 38, 46, 3, 
    14, 40, 47, 56, 61, 21, 20, 53, 47, 32, 19, 55, 37, 38, 8, 
    32, 48, 42, 45, 18, 2, 15, 23, 7, 5, 16, 38, 21, 56, 18, 
    25, 40, 53, 35, 19, 10, 4, 13, 14, 31, 28, 9, 36, 37, 0, 
    46, 62, 31, 28, 18, 25, 19, 9, 19, 5, 4, 24, 0, 12, 21, 
    49, 17, 20, 28, 9, 0, 22, 27, 18, 16, 12, 10, 0, 26, 50, 
    14, 29, 37, 41, 59, 30, 26, 27, 16, 6, 5, 5, 15, 40, 61, 
    62, 88, 60, 61, 28, 44, 26, 7, 16, 14, 21, 6, 1, 31, 47, 
    11, 0, 41, 61, 47, 35, 18, 0, 0, 14, 11, 6, 0, 18, 44, 
    14, 0, 0, 38, 62, 50, 28, 28, 50, 5, 9, 2, 0, 36, 43, 
    13, 20, 18, 9, 36, 72, 59, 44, 12, 0, 0, 0, 42, 54, 67, 
    
    -- channel=142
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 23, 0, 83, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 18, 0, 53, 0, 1, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 47, 0, 4, 
    4, 0, 5, 0, 0, 0, 16, 4, 0, 0, 0, 0, 37, 0, 90, 
    0, 0, 27, 1, 0, 0, 42, 0, 0, 0, 3, 0, 19, 6, 107, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 36, 0, 88, 
    0, 0, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 11, 0, 53, 
    0, 0, 0, 9, 0, 5, 0, 0, 0, 0, 1, 0, 32, 1, 61, 
    0, 0, 2, 0, 0, 0, 0, 0, 4, 10, 0, 0, 44, 20, 5, 
    0, 11, 12, 0, 0, 0, 0, 0, 2, 23, 0, 17, 38, 0, 0, 
    51, 0, 1, 0, 0, 0, 0, 18, 18, 32, 5, 9, 15, 0, 0, 
    0, 0, 5, 0, 4, 0, 0, 14, 17, 20, 0, 11, 13, 0, 0, 
    22, 0, 0, 0, 3, 0, 0, 63, 0, 0, 9, 19, 29, 0, 6, 
    31, 0, 0, 0, 8, 0, 0, 0, 0, 9, 0, 34, 61, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 7, 10, 25, 3, 0, 0, 0, 
    
    -- channel=143
    10, 9, 7, 10, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 7, 
    16, 13, 6, 12, 0, 0, 0, 0, 5, 3, 0, 4, 16, 13, 15, 
    0, 0, 11, 6, 1, 5, 8, 0, 4, 0, 0, 8, 21, 16, 11, 
    3, 11, 7, 10, 10, 0, 0, 0, 0, 18, 6, 0, 11, 19, 7, 
    8, 12, 30, 0, 7, 5, 3, 9, 4, 4, 0, 0, 9, 22, 5, 
    8, 1, 25, 36, 3, 0, 13, 20, 14, 0, 3, 9, 4, 20, 9, 
    18, 8, 12, 20, 0, 0, 6, 1, 0, 1, 13, 11, 11, 17, 14, 
    9, 9, 19, 12, 19, 0, 0, 0, 13, 15, 6, 14, 23, 18, 1, 
    21, 17, 8, 8, 0, 36, 4, 12, 10, 3, 4, 8, 0, 6, 18, 
    15, 4, 2, 0, 8, 0, 21, 23, 13, 16, 10, 6, 11, 11, 13, 
    8, 6, 9, 12, 7, 19, 2, 20, 24, 6, 9, 5, 8, 22, 21, 
    34, 36, 20, 6, 13, 7, 7, 7, 20, 16, 14, 3, 0, 11, 12, 
    0, 0, 15, 11, 5, 5, 0, 0, 0, 20, 8, 10, 0, 0, 0, 
    0, 0, 0, 8, 12, 0, 0, 12, 4, 2, 15, 0, 0, 0, 16, 
    0, 0, 0, 0, 8, 22, 6, 0, 0, 0, 0, 5, 19, 15, 0, 
    
    -- channel=144
    0, 16, 14, 0, 0, 62, 0, 13, 0, 0, 0, 68, 0, 4, 24, 
    0, 17, 0, 0, 0, 0, 0, 40, 0, 0, 0, 73, 0, 57, 0, 
    0, 0, 0, 0, 0, 90, 47, 0, 0, 0, 19, 64, 0, 0, 0, 
    0, 85, 0, 0, 66, 24, 0, 0, 35, 23, 21, 22, 0, 0, 0, 
    0, 28, 0, 0, 64, 0, 0, 111, 0, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 9, 0, 0, 0, 0, 0, 0, 54, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 7, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 
    0, 28, 0, 8, 0, 0, 5, 0, 0, 0, 0, 0, 0, 9, 0, 
    90, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 19, 0, 0, 0, 0, 13, 45, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 37, 36, 
    
    -- channel=145
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 9, 
    7, 5, 3, 0, 0, 0, 7, 8, 0, 0, 0, 3, 2, 0, 0, 
    0, 0, 2, 0, 0, 9, 0, 0, 0, 14, 0, 8, 0, 8, 0, 
    10, 12, 7, 2, 9, 0, 0, 21, 7, 0, 7, 9, 0, 0, 0, 
    0, 0, 1, 2, 0, 0, 19, 0, 0, 0, 0, 1, 1, 2, 0, 
    0, 0, 0, 16, 10, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    3, 6, 6, 0, 0, 0, 5, 21, 4, 0, 0, 19, 3, 0, 0, 
    8, 9, 15, 0, 0, 36, 16, 0, 0, 22, 23, 0, 10, 0, 24, 
    0, 2, 1, 0, 0, 0, 1, 0, 23, 30, 2, 10, 0, 0, 0, 
    0, 9, 12, 0, 8, 0, 0, 7, 4, 4, 15, 3, 20, 24, 6, 
    11, 0, 0, 1, 9, 6, 1, 3, 7, 11, 8, 10, 5, 2, 0, 
    0, 0, 10, 13, 0, 4, 0, 0, 10, 0, 3, 1, 0, 1, 4, 
    0, 0, 0, 0, 10, 0, 0, 1, 0, 0, 1, 15, 0, 30, 0, 
    2, 20, 0, 0, 0, 14, 11, 15, 17, 3, 0, 2, 19, 0, 12, 
    0, 0, 12, 0, 0, 3, 7, 25, 0, 0, 0, 21, 28, 37, 8, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 4, 1, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 2, 4, 0, 
    0, 0, 13, 1, 0, 0, 0, 1, 0, 0, 0, 9, 0, 3, 0, 
    0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 5, 5, 0, 1, 0, 
    0, 0, 5, 3, 21, 0, 4, 2, 6, 13, 3, 15, 8, 3, 0, 
    0, 0, 0, 0, 0, 17, 4, 6, 15, 8, 7, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 21, 10, 11, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 14, 19, 19, 2, 3, 2, 0, 0, 0, 
    23, 37, 8, 0, 0, 0, 12, 8, 21, 5, 12, 0, 0, 0, 0, 
    0, 7, 27, 13, 0, 0, 0, 0, 0, 13, 7, 4, 0, 0, 0, 
    0, 0, 1, 32, 18, 6, 0, 2, 1, 3, 8, 0, 0, 0, 6, 
    
    -- channel=147
    20, 15, 26, 29, 24, 19, 27, 21, 32, 31, 30, 24, 30, 22, 17, 
    23, 20, 28, 29, 18, 19, 22, 20, 33, 29, 31, 25, 29, 25, 30, 
    22, 25, 23, 18, 15, 21, 35, 31, 30, 24, 30, 27, 31, 33, 31, 
    27, 32, 22, 17, 11, 45, 48, 24, 22, 21, 34, 44, 33, 31, 28, 
    25, 35, 36, 14, 23, 41, 30, 20, 43, 41, 39, 43, 33, 27, 22, 
    15, 28, 33, 30, 39, 23, 0, 28, 35, 33, 27, 34, 33, 33, 24, 
    20, 27, 28, 35, 16, 9, 2, 8, 1, 3, 0, 9, 23, 34, 22, 
    24, 28, 28, 30, 20, 0, 6, 0, 4, 1, 0, 1, 8, 23, 22, 
    23, 31, 23, 29, 9, 7, 0, 0, 1, 0, 0, 1, 0, 8, 28, 
    24, 23, 26, 29, 36, 1, 0, 2, 0, 0, 0, 2, 4, 14, 20, 
    27, 29, 26, 30, 22, 31, 6, 0, 1, 0, 0, 0, 1, 10, 40, 
    22, 39, 42, 33, 37, 19, 18, 1, 0, 0, 0, 0, 6, 18, 43, 
    27, 27, 47, 50, 41, 31, 18, 0, 0, 0, 0, 0, 6, 9, 49, 
    30, 20, 40, 47, 51, 52, 43, 23, 15, 1, 2, 0, 0, 23, 43, 
    29, 30, 25, 45, 43, 54, 58, 53, 24, 1, 3, 3, 14, 31, 49, 
    
    -- channel=148
    9, 32, 0, 0, 89, 0, 13, 0, 0, 0, 55, 0, 146, 0, 0, 
    2, 25, 20, 0, 94, 0, 0, 0, 14, 0, 52, 0, 120, 0, 27, 
    25, 0, 2, 19, 75, 0, 0, 27, 0, 67, 0, 0, 71, 0, 19, 
    54, 0, 39, 34, 0, 0, 38, 54, 0, 41, 0, 0, 32, 0, 104, 
    52, 0, 82, 45, 0, 0, 102, 0, 0, 0, 8, 0, 13, 2, 164, 
    78, 0, 0, 93, 0, 0, 29, 0, 14, 0, 24, 0, 41, 0, 178, 
    64, 0, 0, 17, 27, 0, 0, 0, 2, 0, 0, 0, 25, 0, 136, 
    39, 0, 0, 0, 0, 39, 0, 0, 0, 0, 3, 0, 56, 0, 133, 
    0, 0, 7, 0, 0, 35, 0, 0, 0, 0, 8, 0, 36, 16, 77, 
    3, 19, 38, 0, 0, 0, 0, 0, 0, 13, 0, 15, 63, 16, 0, 
    81, 0, 50, 0, 0, 12, 0, 0, 11, 19, 0, 8, 33, 0, 0, 
    0, 0, 76, 0, 30, 0, 0, 0, 0, 35, 0, 13, 32, 0, 6, 
    0, 0, 23, 44, 36, 0, 0, 46, 0, 0, 0, 34, 53, 0, 11, 
    61, 0, 0, 0, 56, 16, 0, 28, 0, 0, 0, 44, 99, 0, 0, 
    82, 21, 0, 0, 0, 32, 35, 2, 23, 0, 0, 12, 49, 0, 0, 
    
    -- channel=149
    0, 0, 27, 8, 0, 76, 0, 34, 4, 16, 0, 102, 0, 44, 13, 
    0, 3, 0, 7, 0, 48, 0, 56, 0, 26, 0, 127, 0, 64, 0, 
    0, 2, 0, 0, 0, 57, 32, 0, 22, 0, 15, 122, 0, 7, 0, 
    0, 73, 0, 0, 20, 55, 0, 0, 80, 0, 47, 86, 0, 1, 0, 
    0, 96, 0, 0, 77, 3, 0, 77, 1, 38, 0, 48, 0, 0, 0, 
    0, 96, 0, 0, 47, 9, 0, 41, 0, 0, 0, 95, 0, 5, 0, 
    0, 61, 47, 0, 0, 6, 0, 7, 0, 12, 13, 26, 0, 27, 0, 
    0, 47, 37, 0, 0, 0, 29, 7, 0, 7, 10, 36, 0, 8, 0, 
    17, 27, 0, 0, 38, 0, 32, 1, 7, 4, 0, 24, 0, 0, 0, 
    11, 0, 0, 28, 0, 41, 9, 18, 2, 0, 2, 0, 0, 0, 44, 
    0, 46, 0, 28, 25, 0, 77, 0, 0, 0, 0, 0, 0, 11, 22, 
    20, 27, 0, 40, 0, 34, 35, 0, 0, 0, 7, 0, 0, 42, 0, 
    21, 52, 0, 0, 0, 40, 6, 0, 44, 0, 0, 0, 0, 45, 0, 
    0, 57, 74, 0, 0, 0, 0, 0, 66, 11, 5, 0, 0, 67, 11, 
    0, 0, 99, 80, 0, 0, 0, 0, 0, 7, 0, 0, 0, 1, 115, 
    
    -- channel=150
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=151
    11, 17, 0, 0, 33, 0, 11, 0, 0, 0, 22, 0, 66, 0, 2, 
    0, 5, 3, 0, 38, 0, 5, 0, 15, 0, 27, 0, 70, 0, 8, 
    2, 11, 0, 0, 36, 0, 0, 0, 0, 12, 0, 0, 36, 0, 5, 
    23, 0, 1, 20, 4, 0, 8, 30, 0, 36, 0, 0, 20, 0, 35, 
    15, 0, 42, 6, 0, 0, 43, 0, 1, 0, 0, 0, 3, 0, 62, 
    28, 0, 0, 44, 0, 1, 25, 0, 6, 1, 14, 0, 15, 0, 78, 
    30, 0, 0, 4, 21, 26, 30, 4, 10, 17, 21, 0, 16, 0, 62, 
    15, 0, 0, 0, 43, 9, 10, 18, 37, 21, 3, 7, 31, 0, 47, 
    0, 0, 0, 0, 0, 59, 0, 23, 16, 13, 24, 4, 22, 5, 49, 
    0, 3, 9, 0, 17, 0, 27, 13, 11, 27, 16, 23, 49, 5, 0, 
    25, 0, 17, 0, 0, 23, 0, 13, 24, 15, 22, 25, 25, 0, 0, 
    0, 0, 33, 0, 12, 0, 0, 15, 11, 29, 16, 25, 35, 0, 0, 
    0, 0, 31, 15, 12, 0, 2, 31, 0, 27, 9, 34, 41, 0, 0, 
    25, 0, 0, 12, 22, 5, 2, 32, 0, 10, 22, 28, 58, 0, 0, 
    36, 31, 0, 0, 14, 16, 10, 0, 8, 10, 15, 37, 28, 0, 0, 
    
    -- channel=152
    0, 0, 0, 0, 0, 27, 0, 25, 17, 41, 0, 63, 0, 36, 0, 
    0, 0, 0, 1, 0, 30, 12, 18, 0, 7, 0, 69, 0, 0, 0, 
    20, 34, 0, 8, 0, 0, 0, 0, 40, 0, 20, 65, 0, 0, 0, 
    0, 3, 0, 0, 0, 7, 0, 0, 26, 0, 2, 40, 6, 4, 0, 
    0, 67, 0, 0, 26, 3, 0, 0, 0, 0, 2, 77, 5, 11, 0, 
    0, 89, 25, 0, 0, 6, 0, 7, 0, 7, 0, 38, 0, 33, 0, 
    0, 32, 67, 1, 0, 4, 0, 0, 4, 13, 0, 0, 8, 26, 0, 
    0, 34, 16, 23, 0, 0, 14, 0, 0, 0, 0, 39, 0, 24, 0, 
    0, 2, 40, 41, 65, 0, 16, 2, 0, 2, 4, 3, 22, 32, 0, 
    10, 32, 0, 40, 20, 96, 0, 0, 6, 0, 0, 0, 0, 0, 26, 
    0, 29, 0, 24, 5, 0, 61, 0, 0, 4, 4, 0, 0, 4, 5, 
    0, 0, 0, 8, 3, 30, 25, 19, 11, 0, 0, 0, 0, 34, 28, 
    76, 138, 0, 0, 0, 51, 36, 27, 88, 0, 14, 0, 0, 56, 27, 
    0, 96, 147, 23, 0, 0, 13, 0, 4, 22, 6, 0, 0, 34, 16, 
    0, 0, 101, 133, 32, 0, 0, 0, 18, 47, 61, 9, 0, 0, 53, 
    
    -- channel=153
    14, 24, 29, 25, 0, 65, 8, 35, 0, 21, 0, 82, 0, 40, 43, 
    24, 27, 7, 19, 0, 24, 17, 56, 11, 24, 0, 88, 0, 55, 0, 
    0, 18, 25, 0, 0, 79, 49, 0, 34, 0, 45, 84, 0, 23, 2, 
    0, 82, 0, 8, 60, 39, 0, 3, 61, 29, 38, 56, 0, 13, 0, 
    0, 61, 0, 0, 70, 17, 0, 92, 18, 44, 0, 44, 0, 6, 0, 
    0, 45, 19, 17, 32, 24, 7, 23, 5, 11, 0, 68, 0, 12, 0, 
    8, 38, 29, 0, 0, 7, 28, 7, 6, 6, 23, 20, 0, 21, 0, 
    6, 42, 34, 0, 21, 0, 30, 10, 13, 31, 12, 21, 0, 7, 0, 
    40, 24, 0, 7, 7, 18, 6, 7, 5, 10, 3, 4, 0, 0, 3, 
    0, 0, 0, 17, 6, 0, 23, 13, 4, 0, 11, 0, 0, 16, 68, 
    0, 46, 0, 39, 24, 23, 47, 0, 0, 0, 2, 0, 0, 38, 1, 
    81, 35, 1, 37, 0, 35, 11, 0, 0, 0, 11, 0, 0, 21, 14, 
    0, 25, 10, 6, 11, 18, 0, 0, 22, 9, 0, 0, 0, 39, 0, 
    0, 0, 44, 33, 0, 19, 15, 34, 47, 0, 8, 0, 0, 46, 74, 
    0, 24, 30, 39, 22, 18, 10, 20, 0, 0, 0, 15, 38, 48, 58, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 25, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 17, 15, 3, 5, 0, 5, 13, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 12, 17, 18, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 25, 19, 15, 8, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 25, 20, 6, 9, 7, 0, 0, 0, 
    1, 26, 0, 0, 0, 0, 20, 21, 24, 11, 34, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 24, 11, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 12, 31, 0, 0, 0, 0, 
    
    -- channel=156
    0, 0, 0, 0, 0, 4, 0, 0, 0, 11, 0, 11, 0, 16, 0, 
    0, 0, 0, 0, 0, 20, 5, 0, 0, 0, 0, 12, 0, 0, 0, 
    17, 19, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 4, 2, 31, 0, 0, 0, 0, 0, 0, 0, 20, 16, 0, 
    0, 5, 0, 14, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    50, 80, 0, 0, 0, 9, 5, 30, 65, 0, 0, 0, 0, 18, 0, 
    0, 80, 92, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 17, 0, 
    0, 0, 66, 69, 0, 0, 0, 0, 2, 35, 52, 0, 0, 0, 0, 
    
    -- channel=157
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 15, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 39, 
    10, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 9, 0, 29, 2, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 2, 2, 7, 24, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 4, 18, 7, 12, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 6, 12, 0, 10, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 36, 13, 3, 5, 13, 18, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 21, 45, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 9, 0, 0, 0, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 26, 0, 
    0, 0, 0, 0, 0, 18, 19, 0, 0, 0, 0, 35, 0, 7, 2, 
    0, 39, 0, 0, 0, 13, 0, 0, 20, 0, 29, 28, 0, 8, 0, 
    0, 33, 0, 0, 10, 0, 0, 34, 0, 23, 0, 0, 0, 4, 0, 
    0, 10, 12, 14, 23, 8, 0, 14, 2, 0, 0, 35, 0, 0, 0, 
    0, 14, 1, 5, 0, 0, 5, 9, 0, 0, 2, 16, 0, 16, 0, 
    0, 8, 18, 1, 17, 0, 2, 2, 5, 34, 18, 4, 7, 0, 0, 
    12, 19, 0, 0, 0, 20, 2, 0, 13, 5, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 26, 8, 5, 0, 0, 0, 0, 23, 
    0, 7, 0, 7, 11, 4, 32, 17, 9, 0, 0, 0, 0, 11, 7, 
    60, 74, 18, 20, 0, 19, 15, 7, 6, 0, 23, 0, 0, 0, 0, 
    0, 0, 9, 18, 6, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 19, 9, 0, 4, 30, 0, 5, 0, 0, 0, 28, 
    0, 0, 0, 0, 7, 34, 13, 14, 0, 0, 0, 0, 10, 30, 50, 
    
    -- channel=159
    7, 0, 10, 14, 18, 0, 8, 1, 12, 0, 15, 0, 19, 0, 0, 
    1, 1, 9, 17, 11, 4, 2, 0, 8, 8, 11, 0, 0, 4, 15, 
    26, 1, 7, 16, 1, 0, 1, 23, 0, 19, 0, 0, 14, 8, 21, 
    8, 0, 17, 2, 0, 9, 20, 0, 5, 0, 1, 3, 14, 13, 37, 
    12, 12, 16, 12, 0, 2, 0, 0, 2, 2, 12, 0, 9, 17, 32, 
    9, 16, 15, 0, 9, 0, 0, 6, 4, 0, 0, 0, 9, 19, 22, 
    4, 9, 11, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 11, 
    6, 7, 12, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 11, 
    0, 11, 15, 11, 4, 0, 0, 0, 0, 0, 0, 0, 1, 6, 3, 
    25, 8, 15, 17, 5, 6, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    18, 2, 7, 2, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 
    0, 0, 0, 4, 17, 1, 0, 0, 0, 0, 0, 0, 0, 3, 13, 
    26, 0, 0, 1, 0, 18, 3, 6, 0, 0, 0, 0, 0, 0, 29, 
    17, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    19, 0, 1, 0, 0, 0, 2, 0, 4, 0, 7, 0, 0, 0, 10, 
    
    -- channel=160
    33, 86, 13, 19, 13, 15, 6, 13, 0, 0, 0, 9, 10, 16, 2, 
    15, 3, 16, 18, 18, 28, 28, 20, 18, 12, 0, 0, 5, 8, 3, 
    7, 0, 21, 9, 17, 12, 20, 14, 23, 65, 63, 35, 1, 0, 12, 
    0, 6, 5, 12, 11, 6, 5, 7, 0, 5, 24, 19, 0, 7, 0, 
    0, 10, 14, 11, 12, 14, 6, 37, 19, 0, 1, 0, 0, 0, 0, 
    0, 18, 28, 19, 0, 27, 43, 0, 0, 5, 0, 0, 0, 0, 0, 
    41, 0, 8, 4, 26, 24, 0, 51, 86, 61, 6, 0, 0, 2, 0, 
    15, 0, 1, 0, 26, 27, 47, 17, 11, 12, 36, 0, 0, 34, 28, 
    23, 22, 21, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 19, 
    4, 9, 5, 0, 0, 0, 0, 38, 36, 0, 9, 28, 0, 13, 35, 
    16, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    0, 21, 0, 69, 55, 67, 68, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 14, 0, 42, 0, 10, 47, 50, 45, 37, 28, 14, 0, 0, 
    0, 0, 0, 0, 0, 17, 12, 7, 28, 45, 47, 69, 63, 55, 0, 
    1, 43, 7, 33, 37, 29, 5, 0, 0, 2, 18, 17, 24, 16, 28, 
    
    -- channel=161
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=162
    11, 53, 67, 74, 62, 72, 59, 67, 13, 46, 45, 31, 34, 56, 18, 
    60, 53, 71, 68, 74, 68, 66, 77, 24, 27, 59, 55, 58, 40, 43, 
    35, 65, 71, 80, 77, 76, 62, 89, 65, 0, 46, 37, 61, 59, 49, 
    32, 71, 72, 83, 77, 85, 77, 75, 91, 72, 60, 25, 51, 60, 56, 
    68, 65, 70, 78, 76, 77, 61, 51, 48, 100, 76, 3, 62, 58, 57, 
    130, 51, 65, 71, 74, 74, 11, 60, 39, 77, 49, 4, 60, 53, 62, 
    112, 100, 53, 47, 62, 65, 35, 0, 22, 32, 1, 2, 42, 46, 54, 
    32, 127, 45, 65, 74, 35, 54, 59, 40, 29, 0, 1, 56, 46, 12, 
    43, 109, 42, 39, 74, 82, 29, 86, 75, 73, 17, 12, 75, 78, 0, 
    45, 115, 41, 0, 137, 91, 17, 70, 10, 27, 10, 11, 76, 103, 0, 
    47, 106, 45, 0, 46, 71, 65, 110, 33, 30, 39, 44, 58, 138, 0, 
    65, 69, 59, 0, 17, 22, 38, 19, 8, 14, 8, 45, 72, 100, 49, 
    75, 69, 56, 85, 22, 56, 63, 10, 0, 0, 0, 4, 51, 45, 73, 
    56, 101, 44, 74, 32, 49, 83, 36, 37, 24, 20, 31, 16, 43, 35, 
    57, 70, 53, 64, 44, 59, 70, 70, 63, 56, 69, 70, 52, 40, 59, 
    
    -- channel=163
    36, 48, 24, 30, 29, 21, 18, 16, 0, 1, 6, 6, 0, 4, 8, 
    23, 27, 29, 26, 27, 32, 35, 36, 16, 0, 0, 0, 22, 14, 2, 
    6, 15, 29, 25, 28, 27, 31, 18, 38, 51, 31, 25, 8, 7, 18, 
    12, 18, 21, 26, 24, 33, 21, 29, 20, 29, 24, 4, 4, 1, 5, 
    10, 15, 29, 24, 23, 27, 25, 33, 10, 10, 19, 7, 8, 7, 10, 
    0, 20, 8, 24, 14, 26, 27, 0, 28, 20, 0, 0, 0, 5, 5, 
    0, 19, 18, 23, 23, 5, 4, 47, 29, 25, 3, 0, 0, 4, 0, 
    12, 6, 16, 4, 33, 28, 41, 20, 14, 24, 12, 0, 7, 32, 0, 
    19, 35, 17, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 
    16, 0, 12, 0, 0, 25, 2, 57, 12, 0, 0, 12, 6, 19, 18, 
    19, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 6, 
    14, 17, 1, 43, 31, 45, 42, 5, 0, 0, 0, 0, 0, 0, 0, 
    28, 15, 0, 0, 36, 41, 23, 25, 28, 17, 0, 2, 0, 0, 0, 
    3, 4, 9, 13, 0, 16, 13, 22, 20, 30, 38, 44, 42, 28, 11, 
    11, 28, 21, 28, 40, 24, 12, 12, 16, 10, 26, 26, 24, 21, 21, 
    
    -- channel=164
    81, 97, 92, 103, 101, 102, 95, 89, 57, 48, 60, 64, 64, 68, 53, 
    88, 86, 100, 103, 109, 110, 109, 114, 91, 48, 57, 59, 74, 72, 63, 
    73, 88, 102, 106, 109, 111, 114, 108, 105, 87, 87, 76, 75, 71, 75, 
    64, 82, 98, 107, 104, 117, 109, 103, 101, 106, 103, 77, 71, 79, 75, 
    66, 91, 101, 107, 110, 105, 94, 106, 87, 102, 95, 53, 61, 64, 72, 
    79, 98, 107, 100, 93, 92, 63, 37, 56, 86, 75, 34, 50, 60, 69, 
    74, 86, 82, 88, 93, 81, 65, 83, 86, 77, 52, 37, 45, 62, 62, 
    72, 94, 81, 72, 91, 83, 98, 84, 64, 70, 54, 26, 41, 78, 50, 
    92, 102, 83, 60, 73, 83, 75, 63, 59, 39, 9, 24, 50, 79, 39, 
    99, 99, 70, 38, 28, 72, 57, 104, 74, 38, 44, 46, 54, 85, 36, 
    95, 91, 60, 27, 59, 25, 48, 76, 35, 31, 18, 38, 62, 75, 34, 
    89, 102, 71, 85, 68, 81, 81, 55, 25, 13, 8, 15, 47, 59, 58, 
    109, 100, 88, 64, 67, 75, 99, 81, 56, 43, 32, 34, 42, 53, 59, 
    90, 94, 80, 87, 63, 91, 99, 96, 83, 74, 76, 83, 77, 78, 56, 
    100, 111, 100, 102, 96, 102, 96, 86, 90, 90, 98, 100, 94, 86, 86, 
    
    -- channel=165
    52, 5, 6, 0, 11, 7, 10, 2, 34, 0, 0, 17, 2, 0, 25, 
    4, 16, 9, 5, 0, 6, 21, 5, 42, 24, 0, 0, 0, 16, 0, 
    34, 0, 8, 0, 0, 10, 21, 0, 7, 58, 0, 27, 0, 0, 4, 
    33, 0, 1, 0, 4, 7, 8, 14, 0, 2, 25, 41, 3, 0, 0, 
    0, 0, 3, 7, 0, 7, 8, 7, 34, 0, 0, 58, 0, 0, 0, 
    0, 28, 0, 4, 14, 0, 45, 0, 22, 0, 19, 47, 0, 0, 0, 
    0, 0, 10, 16, 0, 0, 16, 42, 0, 11, 57, 39, 0, 0, 0, 
    33, 0, 14, 0, 0, 12, 26, 0, 2, 9, 69, 39, 0, 0, 46, 
    13, 0, 4, 42, 0, 0, 38, 0, 0, 0, 35, 16, 0, 0, 96, 
    32, 0, 0, 125, 0, 0, 45, 0, 76, 23, 12, 18, 0, 0, 119, 
    25, 0, 0, 96, 9, 0, 0, 0, 16, 23, 0, 0, 0, 0, 68, 
    8, 0, 0, 45, 44, 11, 11, 46, 30, 0, 4, 0, 0, 0, 0, 
    0, 0, 18, 0, 41, 23, 0, 43, 43, 32, 31, 2, 0, 5, 0, 
    12, 0, 21, 11, 11, 0, 0, 34, 8, 23, 20, 4, 28, 5, 2, 
    0, 0, 13, 0, 21, 4, 3, 0, 10, 6, 0, 0, 15, 24, 0, 
    
    -- channel=166
    60, 48, 66, 68, 66, 55, 50, 43, 47, 26, 34, 27, 21, 38, 40, 
    99, 97, 63, 72, 74, 65, 54, 53, 43, 8, 29, 37, 50, 48, 35, 
    101, 94, 77, 81, 85, 77, 69, 52, 65, 40, 33, 34, 42, 48, 46, 
    89, 92, 87, 88, 91, 84, 80, 67, 72, 75, 55, 45, 37, 33, 48, 
    84, 92, 91, 87, 89, 94, 89, 84, 61, 73, 78, 72, 39, 48, 52, 
    46, 89, 94, 100, 89, 111, 121, 112, 94, 74, 75, 41, 30, 36, 45, 
    36, 112, 129, 118, 89, 130, 119, 97, 78, 90, 75, 28, 17, 30, 40, 
    49, 86, 130, 109, 134, 138, 105, 143, 144, 142, 96, 37, 22, 56, 31, 
    63, 95, 129, 93, 158, 120, 121, 117, 128, 116, 85, 14, 8, 84, 62, 
    69, 90, 153, 98, 96, 124, 103, 99, 61, 28, 6, 9, 16, 97, 100, 
    83, 89, 142, 72, 1, 40, 54, 70, 64, 13, 17, 24, 16, 90, 135, 
    77, 83, 106, 68, 31, 18, 23, 38, 0, 0, 0, 0, 18, 43, 116, 
    69, 87, 77, 109, 74, 73, 58, 39, 13, 0, 0, 0, 6, 13, 51, 
    79, 75, 89, 64, 82, 53, 71, 69, 45, 38, 25, 31, 26, 28, 57, 
    68, 74, 75, 67, 67, 74, 71, 73, 62, 49, 55, 66, 63, 57, 42, 
    
    -- channel=167
    71, 32, 63, 64, 74, 69, 72, 53, 61, 30, 37, 41, 31, 25, 48, 
    54, 71, 64, 66, 70, 71, 80, 75, 83, 33, 26, 34, 43, 53, 37, 
    63, 53, 62, 66, 69, 75, 85, 62, 78, 73, 30, 51, 46, 48, 45, 
    57, 44, 65, 61, 71, 81, 81, 75, 62, 74, 66, 69, 51, 37, 44, 
    41, 46, 63, 68, 68, 73, 63, 59, 61, 56, 60, 82, 35, 42, 46, 
    0, 60, 47, 62, 64, 36, 48, 31, 73, 39, 55, 61, 17, 39, 39, 
    0, 39, 58, 66, 36, 40, 60, 65, 13, 26, 60, 42, 12, 33, 38, 
    56, 0, 62, 40, 31, 52, 57, 45, 38, 47, 67, 41, 7, 28, 41, 
    66, 17, 48, 48, 52, 38, 72, 61, 58, 51, 79, 40, 0, 16, 76, 
    81, 6, 42, 103, 0, 37, 86, 46, 75, 44, 23, 31, 0, 1, 91, 
    76, 27, 51, 98, 12, 13, 47, 37, 72, 37, 18, 26, 16, 0, 87, 
    70, 54, 41, 58, 52, 37, 34, 63, 29, 9, 9, 0, 9, 12, 52, 
    61, 65, 48, 30, 59, 71, 55, 63, 41, 23, 16, 4, 0, 30, 17, 
    68, 41, 72, 49, 63, 49, 44, 81, 49, 45, 43, 34, 43, 31, 49, 
    64, 52, 71, 52, 59, 60, 64, 66, 64, 58, 55, 55, 60, 65, 39, 
    
    -- channel=168
    24, 47, 0, 2, 6, 5, 3, 6, 14, 0, 6, 20, 15, 8, 8, 
    0, 0, 0, 6, 6, 6, 9, 8, 29, 16, 0, 0, 3, 10, 4, 
    8, 0, 0, 0, 0, 0, 7, 0, 9, 52, 37, 18, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 3, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 6, 0, 0, 9, 0, 0, 0, 
    0, 14, 8, 0, 0, 4, 27, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 7, 0, 49, 58, 33, 12, 13, 9, 10, 0, 
    17, 0, 0, 0, 0, 3, 8, 2, 0, 7, 30, 8, 0, 30, 23, 
    6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 31, 
    6, 0, 0, 20, 0, 0, 0, 21, 30, 0, 17, 40, 0, 0, 60, 
    3, 0, 0, 10, 28, 0, 0, 0, 0, 0, 0, 0, 15, 0, 26, 
    0, 3, 0, 40, 43, 43, 35, 23, 9, 8, 16, 0, 0, 0, 0, 
    0, 0, 1, 0, 1, 0, 1, 35, 48, 52, 53, 46, 19, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 5, 17, 31, 35, 48, 44, 31, 14, 
    0, 13, 0, 6, 13, 12, 0, 0, 0, 0, 3, 2, 8, 13, 8, 
    
    -- channel=169
    50, 27, 36, 35, 43, 40, 41, 37, 40, 27, 27, 27, 28, 19, 28, 
    39, 48, 43, 40, 40, 42, 41, 37, 44, 28, 28, 24, 24, 25, 27, 
    37, 49, 40, 42, 41, 44, 44, 40, 47, 37, 21, 21, 22, 28, 24, 
    50, 39, 43, 41, 43, 44, 40, 40, 37, 42, 36, 35, 28, 24, 25, 
    34, 37, 43, 45, 46, 40, 34, 32, 30, 33, 36, 44, 32, 27, 26, 
    37, 35, 37, 40, 45, 46, 24, 29, 46, 26, 27, 43, 26, 31, 26, 
    7, 42, 37, 40, 37, 35, 45, 29, 18, 24, 30, 28, 24, 32, 25, 
    25, 21, 35, 36, 32, 35, 29, 32, 30, 32, 30, 29, 27, 26, 21, 
    25, 17, 29, 32, 43, 39, 31, 47, 41, 36, 50, 40, 22, 29, 32, 
    26, 19, 27, 38, 33, 28, 39, 22, 25, 33, 26, 21, 18, 27, 36, 
    22, 22, 33, 49, 19, 34, 35, 27, 42, 32, 30, 30, 17, 20, 46, 
    26, 19, 32, 36, 22, 16, 13, 27, 33, 31, 27, 27, 31, 19, 46, 
    19, 23, 25, 31, 34, 27, 23, 25, 23, 23, 24, 26, 18, 29, 29, 
    19, 22, 27, 25, 32, 28, 16, 26, 24, 18, 25, 20, 23, 20, 26, 
    27, 10, 23, 19, 22, 19, 24, 27, 26, 23, 22, 24, 23, 27, 22, 
    
    -- channel=170
    46, 62, 40, 48, 48, 36, 32, 27, 13, 0, 8, 5, 8, 17, 8, 
    61, 61, 41, 56, 58, 54, 38, 45, 27, 0, 2, 8, 32, 21, 11, 
    47, 69, 51, 56, 61, 54, 51, 31, 53, 49, 48, 15, 13, 17, 24, 
    39, 62, 57, 62, 62, 56, 49, 35, 40, 58, 34, 11, 8, 12, 20, 
    34, 66, 65, 57, 67, 51, 50, 66, 21, 38, 38, 13, 10, 12, 22, 
    26, 59, 77, 65, 40, 90, 71, 30, 34, 45, 21, 0, 0, 3, 17, 
    23, 67, 81, 74, 64, 82, 69, 90, 88, 70, 21, 0, 0, 8, 7, 
    22, 66, 81, 58, 103, 105, 76, 108, 96, 102, 50, 0, 0, 59, 0, 
    43, 80, 90, 21, 100, 64, 49, 37, 52, 12, 0, 0, 0, 66, 6, 
    37, 67, 100, 5, 36, 60, 40, 113, 17, 0, 0, 0, 1, 88, 51, 
    48, 49, 74, 7, 0, 0, 0, 1, 0, 0, 0, 0, 0, 55, 80, 
    38, 53, 65, 74, 29, 43, 35, 0, 0, 0, 0, 0, 0, 0, 78, 
    47, 60, 36, 58, 31, 30, 46, 31, 13, 0, 0, 0, 0, 0, 2, 
    33, 36, 44, 20, 35, 43, 53, 41, 37, 35, 37, 53, 38, 29, 32, 
    56, 63, 51, 54, 55, 62, 37, 33, 31, 24, 41, 51, 43, 34, 30, 
    
    -- channel=171
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 49, 29, 0, 5, 26, 0, 0, 0, 
    0, 1, 0, 0, 0, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 15, 38, 0, 22, 70, 62, 90, 104, 25, 0, 0, 1, 
    0, 0, 0, 47, 54, 23, 29, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 31, 30, 0, 68, 47, 52, 60, 22, 33, 4, 0, 1, 18, 
    0, 0, 0, 0, 0, 0, 0, 11, 9, 7, 9, 18, 0, 28, 18, 
    0, 0, 0, 13, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    2, 0, 8, 3, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=172
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=173
    0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 7, 0, 13, 35, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 1, 0, 7, 10, 7, 3, 0, 0, 2, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 14, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 9, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=174
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 26, 9, 0, 12, 30, 0, 0, 0, 
    0, 0, 11, 7, 0, 12, 4, 0, 0, 0, 28, 2, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 6, 5, 43, 9, 0, 0, 6, 
    0, 0, 2, 18, 20, 0, 52, 28, 20, 44, 72, 0, 0, 0, 53, 
    8, 0, 12, 108, 0, 0, 40, 0, 41, 0, 0, 0, 0, 0, 87, 
    11, 0, 33, 74, 0, 16, 1, 8, 35, 0, 0, 0, 0, 0, 76, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 15, 0, 11, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23, 13, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 4, 8, 12, 7, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 10, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    93, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 20, 0, 0, 15, 41, 0, 0, 0, 5, 0, 0, 
    0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 33, 0, 
    0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 12, 0, 
    0, 19, 0, 0, 0, 0, 0, 25, 0, 0, 24, 0, 23, 41, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 23, 0, 46, 8, 0, 0, 0, 0, 0, 23, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 11, 30, 23, 47, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 23, 30, 22, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    
    -- channel=177
    9, 0, 0, 0, 0, 3, 0, 2, 0, 0, 4, 14, 11, 0, 0, 
    0, 0, 5, 2, 2, 0, 0, 0, 12, 16, 2, 0, 0, 0, 0, 
    14, 0, 5, 4, 6, 6, 7, 5, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 3, 0, 0, 0, 0, 0, 1, 0, 19, 15, 12, 12, 4, 
    4, 0, 0, 14, 0, 13, 21, 22, 19, 5, 3, 0, 0, 0, 2, 
    9, 34, 18, 9, 20, 10, 2, 0, 0, 11, 21, 22, 0, 1, 1, 
    0, 0, 0, 9, 16, 7, 0, 10, 10, 11, 14, 15, 5, 3, 3, 
    5, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 4, 9, 0, 27, 0, 0, 0, 0, 3, 11, 2, 1, 7, 
    23, 16, 0, 14, 0, 0, 0, 0, 13, 19, 4, 0, 0, 0, 4, 
    1, 6, 2, 12, 44, 40, 16, 30, 6, 15, 3, 0, 0, 1, 0, 
    1, 8, 8, 0, 0, 0, 0, 17, 35, 12, 4, 16, 7, 9, 0, 
    0, 11, 19, 0, 0, 0, 8, 0, 0, 2, 7, 0, 0, 21, 24, 
    10, 7, 0, 14, 0, 5, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 3, 0, 
    
    -- channel=178
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 7, 0, 0, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 4, 5, 12, 6, 2, 13, 14, 4, 0, 0, 0, 0, 0, 
    0, 2, 3, 0, 11, 22, 0, 13, 8, 9, 0, 0, 0, 0, 0, 
    0, 7, 12, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=179
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=180
    49, 0, 2, 0, 3, 0, 9, 0, 47, 0, 0, 8, 0, 0, 30, 
    0, 16, 0, 0, 0, 0, 12, 0, 45, 25, 0, 0, 0, 12, 0, 
    45, 0, 0, 0, 0, 0, 14, 0, 0, 45, 0, 20, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 7, 4, 0, 0, 7, 49, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 31, 0, 0, 85, 0, 0, 0, 
    0, 8, 0, 0, 8, 0, 48, 9, 28, 0, 23, 69, 0, 0, 0, 
    0, 0, 7, 11, 0, 0, 22, 37, 0, 0, 70, 51, 0, 0, 0, 
    24, 0, 16, 0, 0, 15, 10, 0, 0, 5, 94, 56, 0, 0, 56, 
    14, 0, 4, 43, 0, 0, 64, 0, 0, 16, 84, 28, 0, 0, 124, 
    27, 0, 0, 166, 0, 0, 73, 0, 80, 29, 11, 21, 0, 0, 159, 
    27, 0, 6, 148, 0, 0, 0, 0, 62, 26, 2, 0, 0, 0, 114, 
    8, 0, 0, 42, 42, 0, 0, 49, 35, 8, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 51, 16, 0, 43, 39, 22, 26, 0, 0, 0, 0, 
    15, 0, 32, 0, 34, 0, 0, 36, 0, 17, 7, 0, 13, 0, 14, 
    0, 0, 9, 0, 3, 0, 0, 1, 2, 1, 0, 0, 7, 23, 0, 
    
    -- channel=181
    0, 35, 0, 9, 0, 0, 0, 16, 0, 9, 6, 0, 9, 30, 0, 
    5, 0, 5, 0, 1, 0, 0, 5, 0, 0, 23, 9, 14, 0, 4, 
    0, 6, 7, 5, 5, 0, 0, 15, 0, 0, 27, 0, 8, 4, 8, 
    0, 5, 0, 15, 0, 0, 0, 0, 15, 0, 0, 0, 0, 22, 9, 
    4, 15, 1, 7, 0, 1, 0, 5, 0, 28, 13, 0, 20, 5, 7, 
    116, 0, 17, 2, 0, 49, 0, 0, 0, 32, 0, 0, 25, 7, 17, 
    120, 47, 0, 0, 28, 17, 0, 0, 27, 16, 0, 0, 20, 12, 7, 
    0, 107, 0, 4, 44, 0, 0, 17, 0, 0, 0, 0, 33, 27, 0, 
    0, 88, 0, 0, 15, 27, 0, 0, 0, 0, 0, 0, 74, 60, 0, 
    0, 98, 0, 0, 81, 36, 0, 34, 0, 0, 0, 0, 62, 98, 0, 
    0, 64, 0, 0, 46, 14, 0, 38, 0, 0, 1, 4, 42, 116, 0, 
    0, 22, 6, 0, 0, 10, 20, 0, 0, 0, 0, 28, 47, 58, 0, 
    20, 0, 11, 18, 0, 0, 14, 0, 0, 0, 0, 14, 41, 13, 39, 
    0, 43, 0, 28, 0, 8, 31, 0, 1, 0, 0, 18, 0, 25, 0, 
    0, 28, 0, 17, 0, 0, 2, 0, 0, 0, 14, 14, 0, 0, 28, 
    
    -- channel=182
    0, 15, 0, 1, 0, 4, 2, 9, 0, 10, 19, 25, 29, 16, 3, 
    0, 0, 0, 0, 0, 0, 10, 18, 9, 20, 19, 9, 14, 9, 14, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 22, 34, 24, 19, 7, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 18, 29, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 2, 6, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 12, 
    25, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 22, 20, 11, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 17, 4, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 36, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 41, 33, 0, 0, 
    0, 0, 0, 0, 51, 0, 0, 0, 0, 14, 1, 18, 40, 0, 0, 
    0, 0, 0, 0, 18, 54, 48, 13, 23, 25, 26, 28, 26, 0, 0, 
    10, 0, 0, 0, 0, 0, 29, 24, 39, 50, 52, 53, 31, 30, 0, 
    0, 0, 0, 0, 0, 20, 7, 2, 22, 23, 38, 43, 38, 34, 0, 
    8, 16, 1, 11, 9, 6, 0, 0, 2, 17, 21, 11, 7, 7, 24, 
    
    -- channel=183
    67, 29, 54, 51, 59, 51, 59, 35, 50, 30, 34, 35, 26, 19, 46, 
    44, 60, 51, 49, 54, 58, 65, 58, 69, 31, 22, 31, 36, 44, 33, 
    52, 39, 48, 52, 52, 58, 68, 47, 64, 62, 28, 46, 36, 40, 38, 
    45, 33, 49, 47, 49, 64, 62, 62, 48, 57, 50, 59, 44, 28, 34, 
    35, 36, 48, 46, 54, 60, 56, 49, 50, 42, 46, 76, 31, 36, 37, 
    0, 43, 34, 49, 54, 25, 40, 21, 69, 32, 44, 56, 20, 36, 30, 
    0, 25, 40, 50, 29, 11, 46, 60, 15, 16, 55, 44, 16, 30, 32, 
    42, 0, 46, 29, 16, 44, 47, 20, 22, 34, 64, 44, 14, 30, 42, 
    53, 1, 37, 38, 20, 16, 56, 26, 34, 32, 67, 38, 0, 5, 75, 
    60, 0, 25, 90, 0, 21, 76, 42, 56, 38, 31, 35, 3, 0, 87, 
    57, 5, 25, 96, 0, 0, 38, 8, 73, 37, 21, 34, 16, 0, 78, 
    54, 31, 27, 57, 48, 39, 32, 53, 28, 17, 24, 3, 10, 0, 39, 
    47, 45, 23, 27, 63, 60, 43, 56, 44, 30, 21, 13, 3, 28, 0, 
    49, 22, 56, 27, 57, 35, 26, 67, 40, 41, 42, 31, 43, 27, 46, 
    44, 34, 56, 39, 47, 43, 47, 53, 47, 46, 44, 42, 49, 56, 32, 
    
    -- channel=184
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 1, 0, 35, 0, 0, 0, 0, 6, 0, 0, 
    37, 45, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 59, 0, 12, 7, 0, 0, 2, 1, 0, 0, 0, 9, 0, 0, 
    0, 28, 0, 0, 28, 37, 0, 44, 44, 54, 10, 0, 20, 19, 0, 
    0, 44, 0, 0, 142, 35, 0, 0, 0, 0, 0, 0, 18, 45, 0, 
    0, 37, 10, 0, 0, 55, 26, 49, 2, 0, 7, 1, 0, 86, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 7, 24, 40, 23, 
    0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=185
    18, 22, 2, 10, 6, 4, 4, 18, 0, 11, 15, 14, 30, 16, 0, 
    6, 0, 20, 9, 9, 13, 3, 12, 0, 8, 21, 7, 11, 0, 17, 
    0, 18, 13, 10, 13, 5, 4, 16, 16, 16, 27, 2, 0, 9, 12, 
    11, 0, 6, 15, 0, 5, 0, 2, 8, 9, 16, 0, 8, 24, 11, 
    0, 16, 8, 15, 10, 2, 13, 26, 0, 15, 12, 0, 19, 2, 9, 
    103, 8, 26, 4, 0, 62, 0, 0, 0, 25, 0, 0, 14, 10, 14, 
    37, 39, 0, 0, 46, 0, 0, 22, 40, 20, 0, 0, 23, 20, 4, 
    0, 55, 0, 3, 33, 0, 0, 7, 0, 0, 0, 0, 35, 38, 0, 
    0, 46, 1, 0, 0, 36, 0, 0, 0, 0, 0, 6, 55, 43, 0, 
    0, 52, 0, 0, 20, 0, 0, 31, 0, 3, 30, 0, 36, 66, 0, 
    0, 26, 0, 0, 29, 0, 0, 0, 0, 0, 0, 19, 26, 48, 0, 
    0, 4, 11, 23, 0, 32, 15, 0, 11, 18, 7, 16, 45, 4, 10, 
    12, 7, 0, 5, 0, 0, 32, 0, 12, 25, 22, 40, 16, 35, 9, 
    0, 26, 0, 12, 0, 24, 11, 0, 22, 5, 23, 27, 21, 17, 0, 
    21, 8, 5, 13, 17, 0, 0, 0, 0, 11, 13, 15, 4, 0, 31, 
    
    -- channel=186
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=187
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 3, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 26, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 16, 2, 0, 18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 14, 10, 11, 17, 5, 22, 24, 18, 0, 0, 0, 0, 0, 
    0, 17, 11, 0, 27, 8, 10, 23, 23, 26, 1, 0, 0, 0, 0, 
    0, 11, 21, 0, 48, 26, 8, 20, 0, 0, 0, 0, 0, 11, 0, 
    5, 15, 23, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 29, 0, 
    12, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 
    0, 12, 0, 26, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 13, 10, 0, 1, 0, 14, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 7, 2, 2, 0, 11, 3, 8, 0, 0, 0, 2, 0, 0, 0, 
    
    -- channel=188
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 15, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 1, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 23, 1, 0, 12, 9, 3, 
    57, 0, 0, 0, 0, 0, 0, 43, 2, 0, 0, 0, 17, 5, 8, 
    27, 31, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 40, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 8, 0, 0, 29, 21, 0, 60, 56, 67, 48, 9, 20, 9, 0, 
    0, 27, 0, 0, 118, 22, 0, 0, 0, 5, 0, 0, 21, 17, 0, 
    0, 34, 14, 0, 0, 74, 52, 69, 34, 1, 27, 18, 0, 63, 0, 
    7, 0, 8, 0, 0, 0, 0, 0, 0, 6, 0, 19, 32, 50, 29, 
    0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 31, 
    0, 34, 2, 7, 7, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 14, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=189
    15, 0, 22, 16, 22, 24, 33, 22, 39, 24, 27, 26, 23, 20, 35, 
    7, 13, 15, 15, 18, 16, 23, 24, 39, 27, 25, 34, 27, 32, 29, 
    20, 6, 9, 16, 11, 21, 24, 18, 21, 13, 6, 27, 34, 35, 25, 
    17, 4, 16, 11, 16, 25, 31, 25, 22, 28, 21, 35, 35, 26, 30, 
    20, 8, 9, 11, 14, 15, 13, 3, 25, 28, 21, 41, 22, 30, 29, 
    0, 12, 2, 8, 17, 0, 3, 34, 32, 8, 32, 51, 20, 27, 27, 
    0, 8, 10, 13, 0, 0, 31, 4, 0, 0, 35, 38, 15, 21, 30, 
    33, 0, 19, 14, 0, 3, 4, 4, 6, 6, 29, 36, 10, 0, 30, 
    39, 0, 7, 24, 9, 17, 42, 44, 45, 57, 85, 47, 1, 0, 42, 
    46, 0, 4, 64, 22, 4, 58, 2, 42, 47, 23, 25, 8, 0, 37, 
    42, 19, 27, 76, 11, 58, 60, 51, 76, 35, 37, 32, 10, 0, 45, 
    48, 27, 22, 4, 24, 15, 13, 44, 38, 32, 29, 19, 21, 27, 34, 
    31, 37, 25, 26, 13, 29, 28, 35, 22, 13, 18, 8, 12, 27, 22, 
    44, 33, 48, 26, 50, 23, 28, 49, 26, 25, 19, 5, 11, 10, 37, 
    40, 22, 41, 26, 19, 30, 39, 43, 39, 40, 28, 25, 30, 34, 18, 
    
    -- channel=190
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 11, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 10, 0, 0, 21, 45, 24, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 22, 3, 0, 11, 2, 5, 0, 0, 0, 7, 0, 
    0, 22, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 19, 4, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=191
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=192
    60, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 0, 17, 10, 
    0, 0, 0, 0, 0, 0, 1, 5, 10, 13, 18, 0, 29, 33, 10, 
    0, 0, 4, 6, 10, 11, 20, 30, 30, 25, 0, 0, 0, 0, 0, 
    7, 6, 4, 4, 6, 18, 6, 10, 57, 107, 58, 43, 10, 0, 0, 
    8, 7, 6, 2, 3, 43, 101, 60, 0, 0, 72, 87, 0, 8, 0, 
    8, 7, 1, 0, 31, 0, 0, 0, 0, 0, 35, 65, 46, 0, 0, 
    4, 3, 19, 54, 0, 5, 0, 93, 218, 219, 34, 0, 0, 3, 76, 
    2, 5, 8, 0, 0, 0, 0, 85, 5, 0, 0, 0, 38, 142, 62, 
    3, 124, 58, 0, 0, 0, 1, 0, 0, 0, 0, 82, 122, 29, 0, 
    13, 0, 0, 0, 0, 30, 73, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 23, 12, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 79, 107, 72, 0, 0, 8, 47, 7, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 12, 58, 26, 28, 24, 11, 3, 0, 0, 0, 0, 0, 3, 
    
    -- channel=193
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 53, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 26, 2, 0, 7, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 69, 9, 0, 0, 
    0, 0, 0, 5, 19, 1, 0, 1, 44, 46, 38, 17, 0, 0, 0, 
    0, 0, 20, 5, 14, 0, 11, 32, 47, 78, 73, 11, 0, 23, 34, 
    0, 51, 50, 8, 1, 0, 0, 39, 59, 52, 18, 50, 62, 53, 46, 
    0, 13, 14, 12, 0, 0, 17, 44, 50, 0, 0, 9, 37, 39, 0, 
    0, 6, 15, 9, 0, 0, 4, 41, 44, 0, 0, 0, 24, 39, 0, 
    0, 3, 37, 48, 51, 73, 81, 84, 65, 1, 17, 4, 2, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 4, 0, 0, 0, 
    
    -- channel=194
    160, 169, 187, 188, 172, 163, 164, 140, 144, 109, 97, 80, 39, 66, 67, 
    179, 153, 157, 158, 148, 135, 135, 119, 114, 99, 95, 45, 0, 63, 77, 
    144, 132, 129, 124, 120, 111, 111, 105, 100, 103, 67, 11, 26, 71, 76, 
    104, 108, 108, 104, 111, 109, 107, 98, 97, 91, 1, 48, 66, 88, 86, 
    102, 110, 111, 108, 116, 105, 105, 99, 74, 0, 0, 33, 71, 88, 89, 
    108, 109, 107, 106, 114, 81, 46, 53, 81, 44, 0, 0, 69, 40, 81, 
    112, 109, 98, 106, 87, 85, 14, 3, 16, 88, 45, 0, 0, 45, 62, 
    112, 104, 96, 52, 10, 34, 0, 0, 0, 17, 0, 0, 0, 21, 8, 
    107, 102, 41, 29, 0, 34, 66, 51, 22, 4, 0, 0, 16, 5, 20, 
    116, 71, 0, 16, 0, 38, 114, 18, 0, 4, 59, 0, 0, 0, 0, 
    142, 94, 0, 0, 0, 15, 82, 0, 0, 0, 53, 123, 0, 0, 0, 
    99, 3, 0, 0, 3, 36, 69, 0, 0, 0, 0, 109, 3, 0, 0, 
    73, 14, 0, 0, 10, 0, 30, 0, 0, 24, 0, 13, 65, 0, 32, 
    52, 33, 19, 5, 68, 68, 69, 62, 0, 46, 0, 0, 35, 0, 17, 
    43, 4, 0, 0, 0, 0, 0, 0, 0, 51, 2, 0, 0, 2, 11, 
    
    -- channel=195
    87, 68, 60, 52, 47, 40, 38, 36, 25, 0, 12, 11, 0, 0, 20, 
    48, 48, 44, 36, 31, 29, 30, 27, 26, 28, 29, 0, 0, 22, 26, 
    23, 12, 20, 26, 25, 29, 30, 30, 32, 35, 2, 8, 20, 32, 28, 
    18, 26, 31, 31, 35, 36, 43, 43, 38, 30, 0, 0, 20, 17, 17, 
    31, 32, 31, 31, 35, 36, 38, 37, 49, 18, 0, 22, 25, 20, 20, 
    33, 33, 31, 29, 32, 33, 43, 61, 20, 0, 92, 5, 0, 38, 16, 
    33, 31, 28, 30, 10, 0, 0, 0, 0, 0, 0, 52, 0, 0, 8, 
    31, 31, 31, 26, 0, 0, 0, 54, 57, 64, 1, 0, 31, 0, 39, 
    30, 34, 0, 0, 0, 0, 0, 41, 5, 0, 0, 0, 9, 41, 27, 
    39, 57, 14, 0, 0, 0, 11, 0, 0, 0, 0, 98, 45, 0, 0, 
    7, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 28, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=196
    222, 213, 219, 216, 207, 193, 187, 173, 163, 117, 125, 108, 40, 42, 99, 
    212, 196, 189, 187, 175, 161, 158, 149, 141, 131, 129, 78, 23, 72, 116, 
    144, 146, 153, 151, 145, 143, 146, 141, 138, 136, 74, 18, 56, 98, 111, 
    131, 139, 141, 141, 146, 150, 157, 153, 141, 123, 17, 27, 100, 117, 118, 
    134, 145, 145, 144, 147, 140, 121, 141, 157, 126, 30, 40, 97, 113, 114, 
    144, 146, 143, 140, 142, 129, 74, 27, 0, 0, 42, 9, 12, 80, 104, 
    147, 145, 139, 133, 96, 34, 7, 0, 11, 46, 32, 17, 10, 9, 64, 
    145, 144, 123, 88, 30, 35, 17, 70, 93, 79, 23, 0, 8, 23, 65, 
    143, 137, 56, 5, 0, 1, 19, 45, 18, 21, 29, 13, 73, 70, 35, 
    147, 127, 0, 4, 0, 0, 29, 15, 10, 0, 0, 36, 40, 17, 1, 
    118, 0, 0, 0, 0, 28, 40, 11, 0, 0, 0, 0, 0, 0, 0, 
    95, 17, 0, 0, 11, 10, 29, 10, 0, 14, 0, 8, 3, 0, 13, 
    69, 12, 0, 0, 36, 39, 41, 15, 0, 14, 11, 8, 0, 0, 17, 
    66, 17, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 6, 
    58, 31, 9, 7, 0, 2, 2, 3, 3, 0, 0, 0, 1, 2, 6, 
    
    -- channel=197
    5, 12, 0, 4, 9, 6, 0, 13, 0, 0, 7, 0, 22, 0, 13, 
    0, 9, 15, 5, 1, 5, 0, 6, 3, 9, 0, 30, 27, 0, 12, 
    0, 5, 0, 6, 0, 4, 5, 4, 4, 0, 0, 28, 20, 0, 15, 
    0, 1, 4, 8, 2, 2, 1, 9, 6, 5, 43, 0, 1, 7, 8, 
    0, 3, 4, 6, 0, 0, 0, 0, 6, 56, 54, 3, 8, 7, 2, 
    1, 5, 6, 5, 0, 0, 0, 0, 0, 0, 0, 185, 0, 29, 6, 
    3, 6, 11, 0, 0, 0, 5, 23, 0, 0, 0, 194, 56, 0, 0, 
    3, 9, 0, 13, 25, 0, 23, 20, 0, 0, 0, 98, 80, 0, 0, 
    6, 0, 25, 0, 35, 0, 0, 0, 0, 0, 59, 145, 0, 0, 0, 
    0, 0, 156, 0, 55, 0, 0, 0, 0, 8, 0, 68, 10, 10, 27, 
    0, 0, 68, 29, 26, 0, 0, 0, 60, 68, 0, 0, 24, 20, 74, 
    0, 7, 0, 72, 0, 0, 0, 0, 157, 0, 17, 0, 0, 103, 6, 
    0, 0, 0, 77, 0, 3, 0, 0, 161, 0, 58, 16, 0, 91, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 23, 0, 17, 41, 0, 9, 0, 
    0, 22, 12, 31, 10, 9, 14, 14, 14, 0, 1, 35, 1, 1, 0, 
    
    -- channel=198
    6, 11, 15, 12, 12, 5, 7, 2, 2, 19, 4, 7, 22, 0, 0, 
    13, 12, 4, 0, 0, 0, 0, 0, 0, 0, 4, 4, 1, 0, 0, 
    21, 12, 0, 0, 0, 0, 0, 0, 0, 0, 57, 40, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 1, 3, 4, 17, 44, 0, 2, 1, 0, 
    0, 0, 0, 0, 0, 15, 36, 37, 40, 51, 33, 0, 11, 0, 0, 
    0, 0, 0, 0, 6, 40, 100, 138, 175, 190, 184, 25, 19, 23, 0, 
    0, 0, 0, 1, 42, 89, 111, 52, 45, 46, 217, 152, 0, 36, 0, 
    0, 0, 17, 39, 58, 44, 62, 34, 42, 144, 239, 195, 51, 0, 40, 
    0, 12, 33, 68, 63, 33, 42, 216, 257, 264, 249, 72, 33, 44, 141, 
    0, 103, 80, 38, 13, 8, 82, 228, 229, 223, 238, 179, 143, 168, 157, 
    24, 166, 140, 36, 0, 10, 74, 217, 215, 84, 52, 183, 209, 167, 87, 
    24, 45, 119, 24, 0, 66, 146, 221, 156, 29, 14, 40, 168, 96, 0, 
    6, 56, 115, 30, 44, 103, 162, 212, 131, 45, 42, 5, 118, 47, 0, 
    2, 46, 91, 62, 89, 135, 151, 154, 108, 61, 64, 1, 13, 0, 0, 
    16, 24, 14, 5, 0, 1, 0, 0, 0, 14, 53, 0, 0, 0, 0, 
    
    -- channel=199
    150, 163, 163, 168, 168, 153, 142, 143, 123, 102, 103, 76, 48, 26, 74, 
    157, 149, 148, 147, 137, 125, 118, 117, 105, 100, 80, 63, 40, 16, 83, 
    120, 124, 117, 118, 109, 106, 105, 103, 98, 89, 46, 35, 34, 47, 90, 
    95, 97, 100, 101, 100, 103, 102, 99, 94, 80, 60, 0, 61, 87, 93, 
    91, 100, 102, 103, 97, 92, 84, 83, 67, 61, 22, 0, 64, 82, 85, 
    99, 102, 102, 102, 86, 48, 0, 7, 13, 22, 14, 38, 0, 67, 74, 
    102, 103, 104, 85, 43, 33, 35, 22, 23, 0, 0, 100, 0, 5, 44, 
    101, 103, 64, 42, 35, 0, 19, 0, 0, 0, 0, 54, 60, 0, 0, 
    102, 79, 33, 0, 17, 0, 0, 0, 0, 0, 40, 72, 2, 0, 0, 
    78, 4, 54, 0, 16, 0, 0, 0, 0, 0, 0, 34, 0, 0, 13, 
    30, 0, 57, 2, 8, 0, 0, 0, 35, 46, 0, 0, 9, 10, 55, 
    55, 0, 0, 14, 0, 0, 0, 0, 79, 0, 0, 0, 0, 43, 9, 
    38, 0, 0, 4, 0, 0, 0, 0, 69, 0, 11, 0, 0, 44, 0, 
    37, 0, 0, 0, 0, 0, 0, 6, 50, 0, 12, 8, 0, 9, 0, 
    32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 0, 0, 0, 
    
    -- channel=200
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 17, 8, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 30, 14, 2, 
    0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 36, 82, 67, 25, 2, 0, 0, 
    0, 0, 0, 0, 0, 21, 37, 0, 0, 0, 63, 70, 0, 8, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 25, 78, 46, 0, 0, 
    0, 0, 0, 25, 12, 5, 34, 97, 149, 116, 10, 0, 10, 24, 60, 
    0, 0, 16, 0, 10, 0, 0, 39, 0, 0, 10, 0, 47, 79, 40, 
    0, 58, 66, 8, 7, 0, 0, 0, 0, 0, 0, 43, 70, 19, 0, 
    0, 0, 0, 26, 6, 47, 22, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 34, 32, 34, 33, 0, 5, 32, 25, 28, 0, 0, 15, 1, 
    0, 10, 26, 40, 67, 89, 45, 0, 38, 22, 58, 15, 0, 0, 6, 
    13, 6, 0, 0, 0, 0, 0, 0, 0, 1, 3, 22, 0, 0, 20, 
    12, 31, 44, 70, 47, 50, 48, 40, 36, 0, 0, 6, 32, 31, 29, 
    
    -- channel=201
    40, 47, 53, 56, 57, 49, 48, 48, 39, 44, 44, 31, 20, 30, 28, 
    45, 44, 39, 36, 34, 32, 32, 35, 33, 31, 27, 25, 36, 14, 22, 
    34, 34, 28, 26, 28, 24, 24, 31, 28, 27, 16, 30, 25, 16, 27, 
    25, 20, 20, 21, 22, 21, 19, 24, 28, 26, 37, 24, 22, 27, 29, 
    16, 17, 17, 19, 17, 21, 26, 21, 17, 14, 17, 3, 18, 26, 25, 
    15, 16, 18, 20, 15, 16, 0, 2, 15, 31, 20, 5, 26, 22, 22, 
    17, 16, 18, 18, 10, 20, 32, 35, 36, 10, 0, 22, 3, 20, 22, 
    16, 17, 14, 5, 31, 17, 21, 17, 0, 0, 0, 16, 30, 15, 7, 
    14, 14, 11, 27, 23, 26, 15, 0, 0, 10, 6, 27, 1, 0, 0, 
    10, 0, 13, 11, 24, 18, 0, 3, 4, 2, 25, 4, 0, 1, 12, 
    8, 13, 36, 15, 28, 18, 0, 3, 12, 44, 18, 17, 8, 19, 39, 
    16, 15, 19, 19, 20, 3, 0, 0, 30, 17, 22, 5, 19, 20, 28, 
    19, 14, 13, 14, 3, 0, 0, 4, 25, 11, 13, 11, 22, 33, 22, 
    17, 12, 19, 26, 22, 31, 34, 36, 47, 16, 21, 21, 29, 33, 22, 
    15, 17, 19, 12, 15, 16, 18, 19, 23, 18, 19, 34, 26, 26, 25, 
    
    -- channel=202
    56, 25, 21, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 11, 13, 11, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 8, 21, 27, 55, 49, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 45, 87, 65, 47, 62, 186, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 31, 173, 97, 0, 0, 0, 
    0, 0, 8, 2, 0, 10, 21, 83, 135, 169, 165, 63, 4, 0, 67, 
    0, 2, 0, 0, 0, 0, 17, 194, 152, 164, 146, 0, 49, 71, 116, 
    0, 125, 2, 0, 0, 0, 44, 146, 137, 67, 113, 142, 113, 101, 57, 
    0, 26, 51, 0, 0, 14, 60, 139, 80, 0, 0, 87, 93, 51, 0, 
    0, 0, 82, 0, 0, 34, 109, 141, 45, 0, 0, 0, 96, 0, 0, 
    0, 9, 73, 0, 60, 112, 127, 128, 36, 25, 14, 0, 43, 0, 0, 
    0, 2, 6, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=203
    0, 0, 0, 2, 7, 4, 3, 2, 4, 36, 9, 0, 30, 12, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    26, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 83, 97, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 71, 92, 92, 57, 0, 0, 0, 0, 29, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 89, 15, 0, 0, 
    0, 0, 0, 21, 49, 25, 0, 0, 19, 13, 31, 10, 0, 0, 0, 
    0, 0, 0, 1, 26, 9, 0, 7, 0, 107, 88, 0, 0, 0, 48, 
    0, 129, 44, 16, 7, 0, 0, 0, 97, 94, 79, 76, 51, 75, 120, 
    12, 0, 0, 8, 0, 0, 0, 0, 63, 0, 0, 30, 20, 63, 0, 
    1, 1, 1, 0, 0, 0, 0, 0, 22, 0, 0, 5, 69, 59, 7, 
    0, 18, 79, 81, 126, 179, 194, 199, 129, 16, 26, 12, 60, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 53, 19, 0, 0, 0, 
    
    -- channel=204
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 15, 30, 45, 32, 6, 0, 0, 
    0, 0, 0, 0, 0, 4, 37, 39, 26, 22, 70, 55, 24, 21, 0, 
    0, 0, 0, 0, 14, 11, 24, 29, 31, 49, 72, 72, 20, 9, 20, 
    0, 0, 0, 28, 39, 25, 21, 54, 61, 65, 72, 32, 10, 22, 44, 
    0, 0, 44, 39, 31, 21, 31, 74, 72, 72, 50, 44, 54, 63, 54, 
    0, 40, 58, 43, 20, 25, 48, 73, 83, 43, 43, 55, 72, 64, 39, 
    0, 27, 62, 41, 22, 49, 53, 72, 72, 32, 31, 30, 60, 61, 12, 
    0, 30, 62, 43, 42, 62, 69, 73, 66, 34, 41, 28, 49, 40, 10, 
    0, 17, 49, 40, 50, 57, 56, 57, 47, 36, 44, 31, 31, 21, 16, 
    0, 12, 38, 40, 35, 36, 34, 31, 25, 28, 34, 19, 18, 16, 16, 
    
    -- channel=205
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 33, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 24, 0, 0, 81, 38, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 83, 41, 24, 0, 0, 
    0, 0, 0, 0, 0, 7, 14, 72, 132, 150, 84, 3, 0, 12, 40, 
    0, 0, 0, 0, 0, 0, 41, 97, 64, 55, 43, 0, 21, 90, 63, 
    0, 56, 39, 20, 0, 12, 55, 64, 65, 23, 0, 69, 92, 61, 26, 
    0, 0, 7, 16, 0, 44, 95, 67, 27, 0, 0, 0, 36, 20, 0, 
    0, 23, 36, 11, 25, 52, 78, 76, 6, 16, 15, 27, 31, 0, 0, 
    0, 19, 38, 32, 79, 100, 98, 66, 20, 33, 40, 20, 7, 0, 0, 
    0, 7, 6, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    0, 7, 31, 44, 31, 33, 28, 19, 11, 10, 0, 0, 5, 6, 11, 
    
    -- channel=206
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 41, 0, 74, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 79, 62, 19, 0, 0, 115, 0, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 40, 162, 17, 0, 0, 
    0, 0, 21, 0, 42, 0, 0, 0, 50, 54, 115, 91, 0, 0, 0, 
    0, 0, 94, 0, 15, 0, 0, 39, 40, 111, 17, 1, 0, 27, 74, 
    0, 61, 84, 13, 0, 0, 0, 33, 157, 74, 26, 0, 76, 86, 98, 
    0, 0, 19, 28, 0, 0, 0, 33, 172, 0, 0, 0, 14, 110, 0, 
    0, 0, 4, 0, 0, 0, 0, 39, 139, 0, 10, 0, 2, 62, 0, 
    0, 0, 28, 15, 23, 69, 81, 91, 84, 0, 26, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    
    -- channel=207
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 17, 2, 20, 81, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 57, 81, 8, 0, 0, 
    0, 0, 0, 0, 3, 5, 25, 62, 77, 85, 79, 36, 25, 13, 25, 
    0, 0, 0, 5, 7, 0, 25, 65, 64, 70, 64, 27, 27, 58, 48, 
    0, 35, 48, 16, 7, 0, 40, 60, 71, 33, 36, 91, 72, 57, 29, 
    0, 3, 47, 15, 2, 30, 49, 68, 38, 15, 0, 15, 59, 30, 0, 
    0, 28, 38, 18, 16, 27, 59, 75, 43, 17, 12, 2, 49, 24, 0, 
    0, 24, 37, 42, 51, 76, 66, 71, 51, 26, 34, 8, 5, 13, 0, 
    0, 12, 8, 8, 0, 0, 0, 0, 3, 15, 18, 4, 0, 0, 0, 
    0, 17, 26, 27, 20, 21, 15, 12, 4, 0, 7, 1, 0, 0, 0, 
    
    -- channel=208
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 37, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 20, 13, 0, 
    0, 0, 0, 0, 0, 0, 10, 7, 4, 0, 0, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 97, 40, 22, 28, 0, 0, 0, 
    0, 0, 0, 0, 16, 82, 36, 0, 0, 0, 58, 0, 4, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 160, 0, 0, 0, 0, 0, 
    0, 0, 45, 0, 0, 16, 0, 195, 244, 99, 0, 0, 0, 45, 117, 
    0, 37, 0, 0, 0, 0, 117, 3, 0, 0, 0, 0, 89, 141, 0, 
    51, 135, 0, 0, 0, 7, 109, 0, 0, 0, 0, 23, 8, 0, 0, 
    32, 0, 0, 0, 0, 116, 118, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 66, 11, 79, 0, 0, 19, 0, 0, 0, 0, 27, 
    0, 0, 0, 17, 141, 86, 12, 0, 0, 50, 0, 0, 0, 0, 1, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 52, 37, 36, 39, 24, 16, 12, 0, 0, 0, 15, 18, 30, 
    
    -- channel=209
    0, 0, 1, 10, 15, 17, 15, 17, 22, 16, 14, 7, 30, 0, 0, 
    33, 20, 18, 23, 22, 18, 14, 15, 11, 4, 26, 34, 0, 0, 0, 
    14, 25, 18, 18, 12, 7, 6, 4, 0, 6, 5, 5, 1, 0, 0, 
    9, 2, 1, 2, 1, 1, 10, 11, 6, 12, 33, 0, 0, 0, 4, 
    0, 0, 1, 1, 2, 0, 2, 37, 80, 88, 31, 0, 21, 14, 3, 
    0, 2, 2, 5, 23, 47, 0, 0, 0, 0, 0, 35, 0, 3, 7, 
    4, 2, 4, 17, 4, 29, 47, 49, 32, 48, 8, 1, 32, 0, 10, 
    2, 8, 21, 32, 35, 0, 19, 58, 52, 4, 5, 0, 0, 15, 6, 
    2, 35, 67, 16, 2, 25, 16, 0, 0, 8, 33, 45, 38, 12, 0, 
    33, 20, 27, 9, 2, 0, 0, 13, 4, 0, 0, 0, 8, 7, 0, 
    10, 1, 0, 2, 3, 25, 29, 8, 0, 35, 54, 0, 0, 0, 10, 
    35, 19, 0, 6, 9, 5, 0, 0, 1, 11, 3, 18, 0, 8, 0, 
    27, 6, 1, 30, 31, 30, 34, 24, 2, 2, 8, 14, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 8, 19, 0, 0, 
    2, 35, 42, 17, 12, 13, 12, 11, 9, 2, 0, 0, 0, 0, 0, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 51, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 24, 57, 59, 40, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 8, 43, 44, 50, 42, 0, 0, 11, 13, 
    0, 32, 0, 0, 0, 0, 13, 35, 25, 0, 2, 41, 26, 16, 0, 
    0, 0, 0, 0, 0, 0, 25, 38, 0, 0, 0, 8, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 38, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 27, 34, 36, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=211
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 1, 17, 3, 0, 0, 0, 2, 
    0, 0, 0, 0, 1, 0, 0, 16, 6, 0, 9, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 2, 0, 1, 0, 5, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 6, 2, 4, 3, 2, 0, 0, 0, 1, 0, 
    0, 0, 7, 0, 5, 8, 9, 1, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 3, 4, 3, 0, 0, 0, 0, 0, 0, 1, 1, 
    
    -- channel=212
    0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 1, 0, 41, 0, 6, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 37, 36, 0, 3, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 10, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 68, 0, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 202, 0, 24, 0, 
    0, 0, 5, 0, 0, 0, 29, 52, 5, 0, 0, 246, 56, 0, 2, 
    0, 0, 0, 4, 27, 0, 28, 0, 0, 0, 0, 200, 92, 0, 0, 
    0, 0, 20, 0, 67, 0, 0, 0, 0, 0, 74, 192, 0, 0, 0, 
    0, 0, 183, 0, 82, 0, 0, 0, 0, 62, 0, 66, 0, 8, 53, 
    0, 0, 119, 43, 40, 0, 0, 0, 116, 98, 0, 0, 50, 58, 124, 
    0, 0, 0, 100, 0, 0, 0, 0, 244, 0, 35, 0, 0, 162, 14, 
    0, 0, 0, 84, 0, 0, 0, 0, 237, 0, 66, 6, 0, 143, 0, 
    0, 0, 0, 29, 0, 0, 0, 0, 101, 0, 46, 69, 0, 33, 0, 
    0, 15, 7, 38, 8, 7, 13, 17, 19, 0, 30, 51, 6, 3, 0, 
    
    -- channel=213
    15, 1, 6, 2, 0, 0, 5, 0, 14, 0, 0, 6, 0, 12, 0, 
    9, 0, 0, 0, 0, 0, 5, 0, 4, 0, 22, 0, 0, 39, 0, 
    3, 0, 0, 0, 6, 4, 4, 4, 5, 16, 36, 0, 0, 24, 0, 
    4, 10, 8, 4, 11, 9, 12, 7, 9, 22, 0, 31, 5, 0, 0, 
    10, 10, 9, 5, 17, 18, 15, 16, 34, 0, 0, 28, 0, 0, 3, 
    11, 8, 6, 4, 32, 55, 60, 28, 23, 0, 0, 0, 43, 0, 1, 
    11, 7, 0, 22, 54, 18, 0, 0, 0, 156, 82, 0, 0, 3, 0, 
    10, 4, 40, 23, 0, 34, 0, 28, 84, 144, 8, 0, 0, 34, 48, 
    7, 36, 12, 13, 0, 28, 119, 112, 15, 0, 0, 0, 34, 92, 37, 
    45, 129, 0, 31, 0, 57, 189, 28, 5, 0, 10, 0, 40, 0, 0, 
    124, 18, 0, 0, 0, 71, 190, 11, 0, 0, 47, 127, 0, 0, 0, 
    52, 26, 0, 0, 35, 83, 147, 5, 0, 13, 0, 140, 11, 0, 0, 
    39, 26, 10, 0, 96, 35, 99, 0, 0, 54, 0, 28, 58, 0, 19, 
    24, 31, 0, 0, 41, 2, 0, 0, 0, 63, 0, 0, 12, 0, 16, 
    13, 0, 0, 0, 10, 8, 2, 0, 0, 56, 0, 0, 5, 8, 23, 
    
    -- channel=214
    114, 101, 98, 95, 91, 95, 93, 90, 90, 42, 68, 65, 18, 37, 81, 
    106, 97, 102, 111, 108, 103, 103, 96, 96, 93, 97, 46, 25, 82, 98, 
    67, 77, 100, 108, 105, 107, 108, 100, 98, 99, 16, 0, 56, 78, 75, 
    102, 112, 111, 110, 113, 111, 117, 104, 92, 70, 0, 25, 61, 74, 87, 
    113, 117, 114, 110, 111, 88, 60, 75, 96, 66, 15, 43, 75, 87, 91, 
    116, 116, 111, 107, 105, 82, 0, 0, 0, 0, 0, 0, 0, 64, 86, 
    115, 112, 104, 103, 45, 0, 0, 0, 0, 13, 0, 0, 26, 0, 62, 
    111, 108, 91, 54, 0, 0, 0, 73, 83, 0, 0, 0, 0, 40, 61, 
    110, 102, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 52, 0, 
    116, 56, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74, 0, 0, 0, 12, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 0, 0, 0, 39, 0, 0, 0, 0, 8, 2, 0, 0, 0, 21, 
    62, 0, 0, 0, 33, 0, 0, 0, 0, 2, 1, 10, 0, 0, 38, 
    65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 41, 
    49, 27, 23, 33, 32, 33, 30, 31, 34, 0, 0, 7, 42, 42, 38, 
    
    -- channel=215
    116, 126, 126, 129, 131, 119, 112, 115, 91, 69, 77, 75, 48, 28, 66, 
    124, 120, 120, 117, 109, 100, 95, 94, 85, 81, 70, 54, 35, 21, 72, 
    93, 97, 97, 94, 86, 83, 83, 80, 79, 77, 35, 49, 37, 45, 77, 
    76, 77, 78, 81, 80, 82, 82, 82, 76, 69, 37, 0, 53, 70, 78, 
    73, 79, 79, 82, 79, 78, 69, 73, 62, 55, 33, 21, 70, 75, 71, 
    79, 81, 82, 81, 72, 41, 22, 28, 9, 23, 23, 58, 3, 68, 66, 
    80, 81, 85, 76, 35, 5, 2, 5, 12, 0, 0, 121, 5, 19, 52, 
    79, 85, 62, 46, 24, 10, 24, 11, 0, 0, 0, 55, 66, 3, 12, 
    81, 69, 16, 0, 23, 0, 0, 0, 0, 0, 10, 77, 12, 0, 0, 
    75, 0, 60, 0, 33, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 
    13, 0, 59, 10, 28, 0, 0, 0, 8, 35, 0, 0, 0, 0, 48, 
    30, 0, 0, 33, 2, 0, 0, 0, 83, 6, 13, 0, 0, 46, 27, 
    24, 0, 0, 32, 0, 0, 0, 0, 83, 0, 23, 0, 0, 60, 13, 
    27, 0, 0, 5, 0, 0, 0, 0, 53, 0, 17, 25, 0, 27, 10, 
    34, 21, 3, 14, 5, 5, 5, 9, 13, 0, 21, 35, 13, 12, 5, 
    
    -- channel=216
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 79, 94, 0, 0, 51, 0, 0, 
    0, 0, 0, 0, 0, 40, 33, 29, 23, 78, 64, 0, 0, 28, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 30, 72, 50, 55, 54, 0, 0, 0, 0, 1, 
    0, 0, 0, 14, 0, 35, 112, 56, 42, 78, 154, 0, 0, 0, 8, 
    34, 128, 0, 0, 0, 0, 66, 37, 0, 15, 64, 211, 30, 30, 7, 
    0, 0, 0, 0, 0, 27, 91, 27, 0, 0, 0, 109, 48, 0, 0, 
    0, 7, 18, 0, 0, 0, 26, 25, 0, 13, 0, 0, 99, 0, 0, 
    0, 18, 56, 48, 118, 157, 166, 162, 43, 38, 0, 0, 34, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 10, 0, 0, 0, 0, 
    
    -- channel=217
    5, 0, 0, 1, 0, 0, 4, 0, 7, 0, 5, 16, 0, 25, 6, 
    15, 8, 0, 0, 1, 3, 4, 6, 8, 7, 39, 0, 6, 31, 8, 
    0, 0, 5, 2, 10, 10, 8, 13, 12, 23, 4, 0, 22, 16, 0, 
    12, 12, 11, 9, 13, 11, 22, 19, 19, 17, 0, 36, 4, 0, 5, 
    10, 9, 9, 6, 15, 10, 10, 29, 82, 38, 20, 17, 6, 5, 10, 
    10, 9, 7, 6, 30, 78, 37, 0, 0, 0, 45, 0, 36, 0, 7, 
    11, 7, 0, 26, 20, 0, 0, 0, 0, 148, 18, 0, 0, 0, 7, 
    9, 5, 50, 14, 0, 29, 4, 127, 152, 68, 0, 0, 0, 44, 80, 
    3, 45, 0, 21, 0, 24, 116, 28, 0, 0, 0, 0, 71, 94, 6, 
    50, 111, 0, 19, 0, 32, 112, 0, 0, 0, 0, 15, 15, 0, 0, 
    63, 0, 0, 0, 13, 95, 112, 0, 0, 0, 0, 48, 0, 0, 0, 
    18, 35, 0, 0, 58, 34, 95, 0, 0, 26, 7, 46, 14, 0, 28, 
    29, 21, 5, 13, 107, 63, 39, 0, 0, 53, 0, 6, 0, 0, 17, 
    21, 3, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 13, 22, 
    14, 18, 48, 24, 31, 33, 24, 20, 17, 19, 0, 2, 22, 24, 34, 
    
    -- channel=218
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=219
    1, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 42, 73, 73, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 2, 0, 0, 0, 74, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 58, 53, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 66, 80, 68, 57, 0, 0, 0, 41, 
    0, 0, 0, 0, 0, 0, 4, 64, 48, 79, 91, 0, 17, 29, 25, 
    0, 89, 0, 0, 0, 0, 0, 50, 45, 0, 0, 68, 47, 27, 4, 
    0, 0, 5, 0, 0, 0, 18, 51, 7, 0, 0, 4, 19, 0, 0, 
    0, 0, 13, 0, 0, 0, 30, 34, 0, 0, 0, 0, 29, 0, 0, 
    0, 0, 18, 0, 26, 47, 51, 50, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=220
    8, 13, 31, 32, 28, 26, 30, 17, 28, 40, 23, 5, 0, 33, 9, 
    16, 6, 18, 25, 25, 20, 23, 15, 15, 11, 0, 0, 0, 9, 1, 
    36, 38, 27, 20, 20, 13, 14, 10, 7, 3, 0, 0, 0, 0, 2, 
    20, 17, 13, 9, 12, 9, 0, 0, 0, 0, 0, 38, 25, 17, 14, 
    14, 15, 15, 13, 14, 4, 0, 0, 0, 0, 0, 0, 0, 5, 10, 
    14, 12, 10, 13, 3, 0, 0, 0, 55, 68, 0, 0, 44, 0, 6, 
    11, 13, 11, 4, 0, 49, 52, 58, 47, 16, 0, 0, 0, 37, 8, 
    15, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 30, 2, 24, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 31, 37, 2, 0, 59, 97, 0, 0, 0, 6, 
    44, 108, 0, 0, 0, 0, 0, 0, 7, 35, 71, 155, 4, 28, 40, 
    33, 0, 0, 0, 0, 2, 16, 0, 0, 0, 0, 75, 21, 0, 2, 
    21, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86, 0, 15, 
    5, 28, 61, 59, 117, 161, 169, 169, 75, 29, 1, 0, 50, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 26, 0, 0, 0, 0, 
    
    -- channel=221
    58, 65, 67, 72, 78, 75, 70, 73, 70, 77, 68, 55, 42, 35, 58, 
    67, 67, 76, 84, 82, 76, 72, 70, 66, 64, 39, 48, 48, 20, 58, 
    72, 87, 81, 79, 73, 71, 71, 63, 61, 55, 24, 27, 21, 31, 61, 
    72, 71, 69, 70, 67, 69, 56, 51, 48, 45, 57, 26, 58, 64, 68, 
    68, 73, 73, 74, 68, 55, 38, 39, 3, 3, 7, 0, 33, 58, 59, 
    72, 74, 72, 71, 58, 8, 0, 0, 8, 36, 0, 27, 20, 32, 58, 
    72, 75, 77, 61, 26, 42, 71, 79, 63, 0, 0, 33, 16, 37, 40, 
    74, 76, 35, 15, 23, 8, 16, 0, 0, 0, 0, 77, 43, 13, 0, 
    78, 53, 32, 31, 41, 20, 0, 0, 0, 0, 25, 90, 8, 0, 0, 
    62, 0, 25, 15, 46, 13, 0, 0, 0, 43, 26, 0, 0, 0, 29, 
    38, 49, 50, 26, 36, 0, 0, 0, 52, 85, 43, 25, 27, 40, 88, 
    62, 20, 8, 35, 0, 0, 0, 0, 74, 14, 24, 0, 14, 66, 32, 
    49, 19, 1, 15, 0, 0, 0, 0, 62, 0, 9, 17, 22, 71, 25, 
    42, 33, 38, 49, 44, 81, 86, 94, 100, 6, 47, 42, 38, 44, 17, 
    35, 25, 3, 0, 0, 0, 5, 14, 18, 15, 41, 37, 16, 14, 6, 
    
    -- channel=222
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 31, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 22, 0, 0, 0, 82, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 77, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 104, 172, 142, 67, 0, 0, 0, 58, 
    0, 0, 0, 0, 0, 0, 31, 88, 25, 40, 18, 0, 41, 84, 43, 
    0, 91, 0, 0, 0, 0, 43, 44, 43, 0, 0, 52, 57, 28, 0, 
    0, 0, 0, 0, 0, 30, 89, 44, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 14, 82, 45, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 8, 0, 73, 94, 89, 48, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=223
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 24, 41, 29, 18, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 10, 0, 0, 45, 28, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 45, 76, 5, 0, 0, 
    0, 0, 0, 4, 27, 1, 0, 49, 51, 37, 49, 0, 0, 0, 24, 
    0, 0, 28, 17, 12, 9, 4, 48, 45, 85, 37, 15, 34, 38, 49, 
    0, 38, 37, 27, 0, 0, 16, 46, 87, 3, 26, 31, 56, 58, 18, 
    0, 5, 38, 19, 0, 31, 21, 50, 53, 7, 10, 13, 32, 44, 0, 
    0, 11, 34, 6, 0, 18, 40, 40, 47, 4, 16, 16, 37, 18, 0, 
    0, 11, 47, 35, 48, 51, 53, 52, 30, 14, 15, 14, 11, 1, 0, 
    0, 0, 0, 16, 10, 9, 9, 6, 2, 11, 28, 0, 0, 0, 0, 
    
    -- channel=224
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 18, 34, 45, 46, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 42, 29, 21, 8, 0, 0, 
    0, 2, 22, 16, 0, 5, 13, 8, 0, 0, 0, 0, 0, 3, 7, 
    69, 90, 69, 6, 3, 0, 32, 20, 4, 2, 0, 0, 13, 25, 30, 
    30, 8, 0, 21, 16, 29, 1, 0, 7, 9, 4, 0, 1, 4, 5, 
    0, 0, 0, 53, 0, 0, 0, 0, 10, 14, 2, 1, 0, 0, 0, 
    4, 20, 18, 4, 76, 66, 29, 11, 10, 10, 5, 4, 0, 0, 10, 
    25, 40, 89, 117, 39, 55, 5, 25, 0, 0, 12, 10, 0, 3, 0, 
    119, 91, 0, 0, 0, 0, 0, 2, 3, 1, 10, 9, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 23, 
    0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 14, 13, 4, 0, 14, 
    0, 0, 0, 0, 10, 33, 0, 0, 10, 12, 23, 2, 11, 3, 0, 
    0, 3, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=225
    4, 4, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 39, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 36, 40, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 50, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=226
    0, 0, 15, 8, 17, 12, 0, 1, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 11, 14, 14, 41, 15, 12, 6, 3, 0, 0, 0, 0, 0, 
    2, 0, 2, 28, 16, 29, 39, 36, 27, 4, 8, 10, 14, 14, 13, 
    2, 3, 0, 17, 23, 22, 29, 46, 49, 44, 26, 13, 15, 6, 12, 
    0, 0, 0, 0, 26, 41, 17, 19, 39, 42, 48, 29, 29, 17, 23, 
    16, 13, 0, 0, 6, 43, 16, 12, 30, 34, 36, 49, 52, 39, 29, 
    18, 13, 0, 0, 29, 62, 14, 27, 29, 17, 25, 53, 39, 48, 21, 
    11, 10, 3, 4, 0, 21, 5, 39, 33, 4, 18, 34, 31, 33, 12, 
    17, 16, 0, 0, 0, 0, 20, 19, 35, 9, 12, 16, 38, 33, 35, 
    0, 13, 27, 0, 40, 0, 49, 7, 28, 17, 15, 8, 34, 15, 32, 
    12, 0, 0, 12, 38, 28, 39, 44, 34, 30, 26, 12, 27, 23, 26, 
    31, 16, 0, 0, 0, 32, 30, 0, 39, 34, 22, 11, 26, 63, 8, 
    7, 18, 10, 13, 0, 4, 48, 1, 27, 44, 5, 14, 17, 54, 45, 
    12, 18, 25, 34, 41, 23, 29, 25, 33, 50, 38, 14, 25, 49, 62, 
    26, 37, 36, 33, 61, 48, 29, 36, 43, 35, 48, 45, 31, 53, 52, 
    
    -- channel=227
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 4, 12, 16, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 19, 15, 8, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 2, 
    21, 35, 25, 9, 0, 13, 24, 13, 5, 4, 0, 3, 8, 11, 17, 
    12, 0, 0, 0, 16, 0, 0, 3, 7, 8, 4, 0, 0, 10, 3, 
    0, 0, 0, 26, 0, 0, 3, 4, 4, 6, 3, 0, 2, 0, 0, 
    0, 0, 0, 14, 60, 0, 10, 6, 7, 8, 5, 1, 0, 0, 0, 
    11, 19, 37, 18, 44, 22, 15, 10, 0, 0, 7, 4, 0, 0, 0, 
    47, 44, 0, 19, 0, 0, 0, 9, 0, 0, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 20, 5, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 3, 11, 0, 2, 19, 
    0, 0, 0, 0, 9, 27, 0, 0, 0, 8, 10, 0, 22, 0, 4, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 
    
    -- channel=228
    4, 3, 12, 7, 11, 19, 12, 5, 5, 6, 2, 0, 2, 10, 12, 
    4, 4, 11, 7, 12, 10, 13, 17, 9, 16, 24, 29, 28, 30, 27, 
    2, 3, 0, 11, 9, 16, 19, 27, 30, 28, 29, 30, 24, 21, 20, 
    7, 13, 26, 17, 8, 22, 30, 35, 39, 20, 21, 23, 30, 27, 33, 
    41, 43, 23, 11, 7, 20, 27, 27, 32, 33, 25, 26, 42, 53, 54, 
    34, 27, 8, 11, 26, 32, 11, 14, 28, 33, 32, 28, 43, 59, 50, 
    19, 22, 22, 36, 14, 10, 11, 21, 26, 24, 26, 25, 33, 38, 25, 
    28, 36, 29, 21, 44, 47, 35, 34, 22, 14, 20, 24, 22, 30, 37, 
    40, 59, 70, 50, 47, 45, 44, 33, 16, 11, 19, 18, 18, 22, 35, 
    69, 60, 21, 13, 15, 18, 30, 26, 17, 11, 18, 14, 15, 30, 52, 
    45, 30, 5, 0, 4, 0, 9, 15, 21, 14, 20, 20, 25, 51, 53, 
    0, 0, 8, 11, 9, 7, 24, 23, 18, 18, 23, 26, 36, 53, 56, 
    2, 8, 18, 25, 15, 23, 24, 17, 14, 19, 17, 12, 39, 57, 53, 
    20, 24, 19, 21, 37, 44, 38, 25, 22, 16, 1, 8, 23, 51, 56, 
    17, 26, 41, 50, 57, 51, 43, 48, 56, 46, 37, 34, 42, 59, 59, 
    
    -- channel=229
    0, 5, 0, 0, 0, 0, 9, 0, 8, 4, 5, 9, 7, 1, 13, 
    1, 7, 0, 5, 1, 0, 0, 6, 3, 4, 10, 9, 8, 8, 14, 
    0, 0, 9, 0, 2, 0, 0, 0, 0, 2, 5, 5, 4, 6, 10, 
    0, 0, 41, 8, 0, 0, 0, 0, 0, 0, 0, 13, 0, 12, 10, 
    0, 0, 50, 55, 0, 0, 1, 25, 0, 0, 0, 0, 0, 11, 9, 
    0, 0, 52, 54, 8, 0, 9, 15, 0, 7, 4, 0, 0, 0, 9, 
    0, 0, 5, 115, 0, 0, 10, 0, 0, 15, 10, 0, 0, 0, 11, 
    0, 0, 7, 0, 96, 0, 26, 0, 0, 18, 16, 1, 0, 0, 5, 
    0, 0, 13, 69, 12, 59, 0, 31, 0, 8, 13, 12, 0, 0, 15, 
    0, 0, 0, 58, 0, 25, 0, 38, 0, 0, 5, 21, 0, 23, 4, 
    0, 15, 119, 0, 0, 0, 0, 0, 0, 0, 7, 16, 1, 0, 22, 
    3, 5, 18, 19, 57, 0, 0, 53, 0, 0, 0, 18, 15, 0, 41, 
    0, 0, 0, 0, 14, 28, 0, 12, 0, 0, 3, 8, 24, 0, 0, 
    0, 0, 1, 7, 0, 0, 14, 0, 4, 0, 0, 9, 7, 2, 0, 
    4, 5, 1, 7, 0, 0, 11, 14, 9, 2, 0, 0, 9, 0, 0, 
    
    -- channel=230
    78, 72, 76, 81, 75, 76, 66, 66, 55, 48, 41, 31, 20, 14, 8, 
    77, 72, 72, 49, 64, 62, 70, 53, 48, 43, 32, 28, 28, 34, 35, 
    70, 70, 57, 47, 41, 33, 35, 37, 51, 70, 68, 70, 64, 64, 51, 
    62, 63, 43, 4, 25, 26, 23, 31, 44, 74, 82, 73, 65, 52, 40, 
    76, 97, 115, 24, 21, 56, 63, 38, 39, 40, 56, 70, 67, 57, 52, 
    146, 159, 151, 19, 33, 49, 69, 58, 49, 35, 39, 50, 64, 77, 71, 
    153, 150, 141, 63, 35, 71, 74, 54, 64, 51, 41, 38, 66, 79, 70, 
    135, 139, 146, 123, 76, 23, 54, 49, 80, 72, 44, 37, 58, 51, 48, 
    146, 160, 168, 117, 162, 115, 96, 54, 76, 76, 54, 42, 47, 50, 51, 
    197, 236, 247, 235, 154, 157, 86, 72, 71, 75, 68, 50, 42, 33, 15, 
    274, 272, 163, 131, 102, 97, 76, 63, 71, 74, 69, 48, 32, 42, 14, 
    249, 203, 135, 106, 49, 28, 55, 36, 41, 52, 67, 59, 30, 46, 38, 
    118, 110, 98, 88, 79, 43, 56, 57, 40, 61, 94, 71, 48, 31, 52, 
    74, 76, 80, 68, 47, 52, 31, 42, 35, 51, 84, 65, 47, 27, 33, 
    66, 51, 33, 18, 17, 49, 43, 27, 14, 19, 22, 35, 27, 12, 20, 
    
    -- channel=231
    0, 0, 0, 0, 0, 12, 8, 5, 1, 0, 3, 2, 2, 0, 2, 
    0, 0, 0, 0, 7, 3, 22, 17, 9, 3, 5, 2, 0, 1, 6, 
    0, 0, 4, 1, 8, 10, 14, 20, 12, 4, 5, 13, 11, 15, 19, 
    0, 0, 21, 0, 5, 9, 9, 13, 28, 14, 11, 26, 19, 15, 19, 
    0, 0, 27, 16, 0, 0, 8, 18, 24, 25, 17, 27, 23, 27, 27, 
    0, 1, 45, 1, 9, 0, 6, 20, 17, 19, 27, 15, 20, 37, 34, 
    3, 7, 12, 49, 0, 0, 24, 15, 10, 15, 24, 6, 29, 27, 30, 
    0, 0, 10, 10, 52, 0, 18, 8, 8, 17, 19, 17, 21, 18, 21, 
    0, 0, 3, 0, 34, 44, 19, 18, 4, 11, 14, 18, 6, 17, 45, 
    0, 0, 0, 65, 4, 56, 0, 33, 5, 5, 12, 20, 13, 39, 38, 
    4, 21, 59, 21, 9, 28, 20, 13, 11, 11, 21, 23, 18, 36, 37, 
    29, 32, 21, 16, 20, 2, 2, 22, 0, 1, 4, 21, 29, 23, 57, 
    8, 8, 9, 6, 19, 12, 6, 27, 0, 0, 7, 10, 45, 33, 36, 
    6, 5, 18, 35, 33, 27, 15, 18, 18, 5, 8, 15, 29, 44, 33, 
    21, 34, 36, 35, 25, 29, 33, 43, 39, 31, 19, 26, 42, 40, 45, 
    
    -- channel=232
    16, 15, 10, 7, 7, 18, 24, 16, 20, 20, 17, 18, 22, 25, 34, 
    16, 20, 15, 0, 20, 3, 16, 30, 20, 25, 36, 44, 47, 46, 41, 
    12, 14, 7, 0, 17, 24, 21, 20, 30, 41, 31, 28, 15, 10, 7, 
    18, 24, 48, 32, 25, 37, 36, 27, 21, 4, 11, 15, 14, 18, 21, 
    56, 62, 67, 21, 27, 24, 44, 35, 28, 26, 15, 18, 21, 25, 26, 
    18, 5, 30, 22, 43, 41, 25, 23, 32, 29, 31, 18, 6, 6, 9, 
    0, 0, 9, 59, 12, 0, 15, 26, 34, 33, 33, 19, 10, 0, 0, 
    9, 14, 13, 0, 84, 52, 42, 25, 30, 34, 32, 31, 22, 16, 20, 
    17, 26, 60, 55, 37, 53, 21, 33, 23, 27, 36, 39, 27, 10, 0, 
    54, 31, 0, 0, 0, 19, 6, 23, 30, 26, 32, 37, 24, 11, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 17, 18, 31, 25, 25, 24, 
    0, 0, 0, 17, 28, 13, 26, 36, 10, 16, 30, 38, 19, 2, 23, 
    0, 0, 0, 8, 23, 34, 8, 25, 33, 24, 41, 22, 26, 11, 5, 
    7, 11, 0, 0, 0, 15, 26, 17, 11, 0, 0, 12, 12, 1, 0, 
    0, 0, 0, 7, 2, 9, 12, 3, 12, 17, 9, 0, 1, 1, 4, 
    
    -- channel=233
    30, 31, 29, 27, 45, 55, 42, 35, 31, 34, 34, 33, 32, 29, 29, 
    31, 32, 31, 38, 54, 69, 73, 61, 39, 35, 34, 31, 27, 22, 23, 
    33, 33, 34, 45, 70, 80, 87, 90, 59, 33, 32, 33, 29, 28, 32, 
    34, 33, 34, 41, 81, 83, 82, 84, 84, 66, 56, 50, 31, 30, 33, 
    23, 18, 27, 50, 73, 74, 73, 81, 93, 93, 86, 72, 39, 32, 32, 
    20, 24, 40, 36, 67, 64, 78, 88, 86, 89, 95, 87, 51, 35, 31, 
    26, 27, 32, 30, 42, 67, 85, 88, 78, 78, 92, 88, 66, 40, 34, 
    30, 25, 27, 35, 34, 34, 63, 79, 80, 80, 90, 91, 79, 51, 35, 
    25, 21, 18, 20, 44, 36, 52, 73, 84, 83, 87, 94, 82, 54, 39, 
    2, 1, 10, 48, 53, 59, 55, 81, 85, 83, 86, 94, 83, 55, 33, 
    11, 16, 43, 69, 70, 89, 75, 74, 84, 81, 82, 92, 76, 47, 29, 
    34, 45, 35, 40, 63, 81, 70, 49, 76, 82, 71, 78, 63, 43, 40, 
    38, 35, 36, 32, 38, 45, 60, 68, 69, 74, 68, 78, 68, 43, 44, 
    36, 33, 41, 44, 45, 41, 45, 59, 67, 67, 77, 82, 72, 49, 41, 
    36, 42, 45, 39, 33, 40, 46, 47, 45, 49, 52, 55, 56, 41, 38, 
    
    -- channel=234
    27, 20, 28, 25, 22, 36, 21, 19, 9, 5, 0, 0, 0, 0, 0, 
    26, 23, 24, 0, 20, 12, 29, 19, 6, 10, 11, 17, 20, 24, 17, 
    17, 21, 0, 0, 0, 0, 0, 12, 35, 48, 39, 38, 23, 15, 2, 
    17, 25, 21, 0, 0, 2, 3, 8, 10, 29, 39, 25, 25, 17, 13, 
    75, 97, 82, 0, 0, 33, 40, 5, 11, 12, 21, 35, 42, 39, 34, 
    98, 94, 87, 0, 17, 35, 18, 14, 20, 7, 7, 17, 34, 42, 29, 
    76, 76, 89, 24, 0, 12, 25, 23, 35, 15, 8, 7, 20, 24, 4, 
    83, 94, 88, 79, 61, 21, 28, 22, 45, 32, 9, 2, 23, 14, 24, 
    103, 129, 163, 80, 131, 73, 70, 15, 32, 33, 21, 9, 17, 10, 0, 
    184, 188, 133, 132, 77, 92, 39, 22, 32, 35, 34, 12, 5, 0, 0, 
    184, 164, 25, 37, 20, 16, 12, 5, 30, 29, 22, 12, 5, 29, 0, 
    84, 59, 52, 49, 0, 0, 35, 0, 0, 15, 33, 28, 0, 20, 11, 
    36, 36, 39, 43, 41, 14, 13, 20, 9, 33, 55, 25, 19, 2, 26, 
    29, 35, 24, 3, 0, 27, 0, 10, 0, 0, 19, 17, 6, 0, 0, 
    8, 0, 0, 0, 0, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=235
    1, 4, 0, 13, 13, 0, 3, 5, 1, 5, 9, 9, 3, 0, 0, 
    1, 1, 6, 5, 13, 28, 17, 3, 3, 0, 0, 0, 0, 0, 0, 
    8, 6, 29, 21, 14, 8, 19, 5, 0, 0, 0, 0, 0, 8, 14, 
    0, 0, 0, 0, 6, 0, 0, 0, 15, 23, 7, 9, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 3, 10, 17, 4, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 10, 6, 0, 0, 9, 8, 0, 0, 0, 
    15, 12, 0, 0, 9, 41, 27, 4, 0, 0, 6, 4, 10, 17, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 7, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 0, 1, 1, 10, 40, 
    0, 0, 37, 46, 33, 31, 4, 5, 4, 2, 0, 5, 10, 14, 0, 
    0, 25, 74, 69, 58, 69, 36, 32, 14, 16, 20, 4, 0, 0, 0, 
    133, 108, 19, 10, 14, 16, 0, 1, 16, 0, 0, 0, 1, 0, 0, 
    41, 37, 12, 0, 0, 0, 24, 3, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 30, 51, 28, 0, 0, 12, 19, 40, 52, 18, 15, 9, 11, 
    36, 46, 19, 0, 0, 3, 4, 7, 1, 2, 17, 30, 19, 1, 7, 
    
    -- channel=236
    28, 27, 24, 27, 13, 3, 15, 20, 22, 20, 20, 20, 19, 17, 17, 
    28, 27, 24, 15, 2, 0, 0, 0, 11, 15, 11, 10, 9, 11, 12, 
    26, 26, 22, 5, 0, 0, 0, 0, 0, 9, 8, 6, 7, 12, 9, 
    21, 22, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 0, 
    20, 22, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 29, 34, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 30, 28, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    27, 26, 25, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 23, 27, 16, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 37, 41, 30, 12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 51, 29, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 44, 25, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 25, 23, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=237
    26, 24, 23, 16, 14, 14, 19, 16, 18, 15, 12, 10, 9, 12, 14, 
    25, 23, 19, 13, 9, 3, 3, 12, 10, 14, 20, 26, 30, 31, 25, 
    21, 19, 8, 0, 0, 1, 0, 0, 17, 34, 25, 20, 13, 6, 0, 
    21, 24, 23, 13, 3, 7, 6, 0, 0, 0, 10, 5, 7, 9, 4, 
    59, 70, 46, 7, 11, 13, 23, 5, 0, 0, 0, 1, 8, 9, 8, 
    48, 40, 18, 15, 18, 30, 16, 3, 5, 0, 0, 0, 0, 0, 0, 
    26, 26, 30, 31, 8, 0, 0, 6, 13, 8, 0, 4, 0, 0, 0, 
    36, 42, 36, 18, 37, 42, 18, 8, 19, 15, 3, 2, 0, 1, 6, 
    46, 56, 77, 79, 38, 33, 10, 13, 16, 14, 12, 6, 8, 1, 0, 
    98, 88, 42, 14, 14, 0, 10, 4, 18, 18, 15, 9, 6, 0, 0, 
    62, 46, 0, 0, 0, 0, 0, 0, 10, 10, 0, 4, 3, 0, 0, 
    0, 0, 7, 16, 12, 0, 15, 9, 0, 6, 18, 12, 0, 0, 0, 
    6, 9, 11, 18, 15, 22, 0, 4, 17, 25, 30, 10, 0, 0, 0, 
    13, 17, 2, 0, 0, 0, 6, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=238
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 19, 13, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 18, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 2, 30, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 5, 61, 91, 13, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 85, 111, 53, 7, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    108, 93, 26, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=239
    15, 13, 12, 12, 0, 0, 1, 6, 9, 4, 4, 3, 1, 3, 6, 
    15, 13, 7, 2, 0, 0, 0, 0, 0, 5, 5, 10, 12, 14, 12, 
    10, 10, 0, 0, 0, 0, 0, 0, 0, 12, 8, 5, 4, 3, 0, 
    9, 12, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 
    34, 41, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 30, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 25, 29, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 30, 24, 20, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 44, 62, 37, 25, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 67, 40, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 53, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 12, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 10, 9, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=240
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 30, 31, 21, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 1, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    60, 49, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=241
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 10, 3, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 6, 20, 15, 4, 14, 10, 0, 9, 0, 0, 1, 2, 0, 0, 
    8, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 5, 8, 8, 0, 3, 3, 5, 6, 0, 0, 2, 
    5, 7, 0, 23, 0, 0, 0, 0, 2, 5, 3, 0, 0, 5, 9, 
    6, 5, 0, 0, 11, 22, 3, 0, 0, 0, 0, 5, 1, 15, 0, 
    7, 26, 26, 17, 0, 0, 0, 6, 5, 0, 1, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, 1, 4, 2, 
    8, 0, 50, 33, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 3, 
    0, 27, 0, 0, 20, 13, 0, 24, 25, 12, 1, 4, 1, 0, 1, 
    0, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    5, 0, 0, 0, 5, 0, 11, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 
    
    -- channel=242
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 16, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 45, 64, 15, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 60, 29, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=243
    11, 11, 8, 7, 15, 23, 13, 8, 9, 10, 6, 6, 5, 3, 2, 
    11, 11, 11, 5, 25, 29, 32, 24, 8, 9, 8, 6, 6, 3, 2, 
    11, 11, 7, 17, 30, 39, 43, 39, 20, 12, 12, 8, 2, 0, 0, 
    11, 12, 7, 14, 41, 44, 42, 43, 35, 21, 22, 12, 0, 0, 1, 
    11, 13, 18, 15, 38, 41, 43, 44, 44, 43, 38, 30, 7, 0, 0, 
    9, 8, 15, 8, 35, 38, 39, 48, 45, 46, 46, 43, 14, 0, 0, 
    7, 5, 7, 9, 13, 32, 44, 47, 42, 42, 45, 44, 26, 0, 0, 
    11, 7, 9, 5, 15, 13, 30, 39, 43, 46, 48, 48, 38, 14, 0, 
    12, 9, 9, 7, 25, 15, 21, 33, 44, 48, 49, 51, 42, 21, 0, 
    9, 9, 3, 22, 22, 23, 19, 35, 46, 49, 48, 52, 45, 15, 0, 
    4, 5, 2, 15, 33, 32, 35, 30, 43, 45, 42, 47, 37, 10, 0, 
    8, 0, 5, 19, 26, 41, 34, 20, 36, 42, 37, 43, 24, 1, 0, 
    6, 10, 4, 7, 8, 21, 27, 24, 36, 44, 41, 43, 30, 0, 0, 
    6, 7, 9, 3, 0, 1, 9, 22, 24, 29, 32, 43, 32, 0, 0, 
    5, 0, 0, 0, 0, 0, 6, 0, 0, 4, 11, 13, 9, 0, 0, 
    
    -- channel=244
    4, 10, 0, 8, 0, 0, 18, 9, 14, 10, 13, 18, 13, 1, 13, 
    5, 14, 0, 4, 10, 0, 9, 8, 12, 4, 5, 4, 1, 0, 11, 
    4, 6, 27, 0, 10, 0, 0, 0, 0, 0, 3, 5, 7, 13, 18, 
    2, 0, 42, 7, 0, 0, 0, 0, 0, 0, 0, 18, 3, 15, 10, 
    0, 0, 71, 55, 0, 0, 0, 23, 0, 0, 0, 0, 0, 6, 4, 
    0, 0, 89, 58, 0, 0, 12, 20, 0, 2, 3, 0, 0, 0, 12, 
    0, 0, 14, 113, 0, 0, 20, 0, 0, 15, 13, 0, 0, 0, 25, 
    0, 0, 13, 13, 90, 0, 21, 0, 0, 24, 18, 0, 0, 0, 7, 
    0, 0, 0, 52, 14, 66, 0, 25, 0, 13, 14, 15, 0, 0, 27, 
    0, 0, 17, 103, 0, 71, 0, 41, 0, 0, 6, 26, 0, 30, 9, 
    0, 35, 139, 23, 1, 20, 0, 0, 0, 0, 10, 17, 0, 1, 25, 
    38, 33, 49, 30, 61, 0, 0, 46, 0, 0, 0, 15, 19, 0, 43, 
    15, 3, 1, 0, 33, 21, 0, 24, 0, 0, 5, 16, 29, 0, 0, 
    0, 0, 10, 18, 0, 0, 0, 5, 0, 0, 0, 10, 16, 3, 0, 
    15, 12, 3, 9, 0, 0, 10, 14, 3, 0, 0, 0, 13, 0, 0, 
    
    -- channel=245
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 7, 3, 0, 13, 0, 0, 0, 0, 0, 4, 9, 11, 0, 
    0, 0, 0, 13, 0, 1, 1, 5, 24, 10, 3, 0, 0, 0, 0, 
    1, 4, 0, 13, 1, 4, 10, 11, 10, 13, 3, 0, 0, 0, 0, 
    29, 31, 0, 0, 13, 32, 5, 0, 0, 4, 12, 0, 6, 0, 1, 
    18, 5, 0, 0, 0, 50, 0, 0, 1, 0, 0, 17, 21, 1, 0, 
    1, 0, 0, 0, 18, 32, 0, 0, 10, 0, 0, 29, 3, 8, 0, 
    8, 12, 0, 0, 0, 46, 0, 17, 16, 0, 0, 5, 0, 6, 0, 
    21, 30, 3, 0, 0, 0, 0, 0, 15, 0, 0, 0, 16, 4, 0, 
    43, 33, 0, 0, 0, 0, 17, 0, 12, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 7, 26, 0, 16, 16, 9, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 0, 18, 0, 16, 43, 0, 0, 0, 13, 1, 
    0, 7, 0, 0, 0, 0, 8, 0, 3, 25, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 27, 11, 0, 0, 0, 0, 14, 0, 0, 6, 2, 
    
    -- channel=246
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 7, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 20, 0, 0, 0, 12, 1, 0, 0, 0, 19, 19, 
    
    -- channel=247
    1, 4, 0, 3, 4, 15, 9, 8, 9, 8, 9, 12, 12, 9, 14, 
    2, 7, 1, 1, 16, 6, 27, 17, 12, 12, 12, 13, 13, 13, 17, 
    1, 5, 10, 12, 18, 20, 19, 22, 15, 11, 15, 17, 17, 18, 21, 
    4, 3, 28, 1, 18, 21, 23, 25, 21, 8, 12, 21, 16, 17, 24, 
    0, 0, 34, 36, 13, 11, 23, 34, 32, 26, 17, 28, 18, 27, 29, 
    0, 0, 46, 24, 23, 0, 11, 34, 28, 32, 33, 17, 16, 32, 31, 
    0, 0, 10, 57, 0, 3, 33, 24, 17, 29, 34, 13, 28, 22, 28, 
    0, 0, 4, 26, 61, 0, 27, 18, 13, 30, 34, 25, 24, 14, 21, 
    0, 0, 5, 3, 35, 40, 27, 27, 7, 23, 29, 31, 13, 20, 40, 
    0, 0, 0, 61, 0, 55, 0, 41, 8, 14, 23, 33, 17, 40, 40, 
    0, 0, 40, 4, 9, 23, 21, 26, 16, 17, 28, 32, 24, 41, 39, 
    2, 3, 30, 25, 28, 16, 9, 25, 3, 10, 17, 30, 35, 20, 56, 
    3, 2, 3, 7, 32, 25, 9, 35, 8, 0, 14, 22, 52, 29, 36, 
    5, 5, 14, 25, 24, 30, 18, 20, 21, 2, 6, 24, 35, 42, 24, 
    18, 25, 31, 37, 24, 23, 31, 42, 36, 29, 15, 22, 41, 39, 39, 
    
    -- channel=248
    1, 0, 10, 9, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 10, 1, 30, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 19, 3, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 27, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 19, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    6, 17, 0, 0, 0, 10, 1, 0, 0, 0, 0, 12, 7, 0, 0, 
    29, 22, 0, 0, 15, 58, 3, 1, 0, 0, 0, 16, 0, 11, 0, 
    11, 4, 0, 8, 0, 0, 0, 4, 8, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 8, 0, 0, 
    0, 0, 58, 0, 52, 0, 27, 0, 8, 5, 0, 0, 2, 0, 0, 
    36, 27, 0, 44, 49, 42, 24, 31, 14, 13, 4, 0, 0, 0, 0, 
    98, 77, 8, 0, 0, 14, 4, 0, 23, 15, 0, 0, 0, 8, 0, 
    34, 29, 13, 2, 0, 0, 24, 0, 4, 23, 0, 0, 0, 0, 0, 
    2, 1, 11, 15, 11, 0, 0, 0, 4, 34, 50, 4, 0, 0, 0, 
    9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 0, 
    
    -- channel=249
    7, 4, 16, 0, 4, 19, 3, 8, 6, 4, 6, 4, 11, 21, 23, 
    8, 4, 6, 17, 0, 11, 9, 14, 12, 18, 28, 33, 32, 26, 16, 
    6, 6, 0, 13, 13, 25, 21, 35, 45, 22, 13, 9, 5, 0, 0, 
    13, 20, 19, 16, 31, 40, 43, 29, 23, 19, 12, 1, 14, 5, 11, 
    55, 45, 0, 4, 25, 44, 30, 15, 28, 25, 25, 21, 21, 15, 14, 
    8, 0, 0, 4, 40, 52, 11, 18, 33, 26, 23, 37, 25, 10, 1, 
    0, 0, 1, 0, 5, 16, 1, 27, 33, 20, 17, 41, 15, 7, 0, 
    15, 18, 0, 7, 0, 58, 12, 31, 30, 9, 18, 27, 24, 24, 19, 
    22, 44, 52, 6, 3, 0, 19, 8, 30, 16, 23, 21, 35, 9, 0, 
    41, 2, 0, 0, 0, 0, 14, 5, 30, 24, 21, 14, 28, 4, 13, 
    0, 0, 0, 0, 0, 0, 9, 15, 21, 16, 9, 23, 28, 24, 3, 
    0, 0, 0, 0, 0, 30, 50, 0, 32, 43, 32, 17, 12, 23, 1, 
    0, 0, 7, 7, 0, 3, 7, 15, 28, 54, 14, 7, 12, 14, 18, 
    15, 6, 0, 0, 9, 16, 23, 4, 15, 11, 6, 16, 4, 12, 12, 
    0, 0, 9, 11, 25, 11, 5, 6, 13, 15, 15, 4, 5, 13, 9, 
    
    -- channel=250
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=251
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 13, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 55, 79, 29, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    69, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    1, 0, 0, 0, 12, 35, 0, 0, 0, 0, 0, 0, 0, 9, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 12, 0, 17, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 33, 35, 9, 15, 0, 0, 0, 0, 0, 0, 0, 
    71, 60, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 12, 0, 
    26, 17, 4, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 15, 31, 26, 0, 0, 4, 4, 25, 35, 0, 0, 5, 16, 
    20, 32, 18, 0, 9, 7, 0, 0, 0, 0, 16, 25, 7, 7, 7, 
    
    -- channel=253
    0, 0, 0, 8, 0, 0, 0, 4, 3, 5, 10, 14, 13, 10, 10, 
    0, 0, 1, 1, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 
    1, 2, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 21, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 14, 
    0, 2, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 11, 0, 9, 0, 0, 0, 0, 0, 0, 0, 11, 32, 
    0, 3, 46, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 
    41, 49, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 
    23, 13, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 
    5, 1, 12, 32, 33, 12, 0, 0, 0, 0, 0, 0, 0, 18, 20, 
    22, 36, 32, 25, 17, 13, 8, 21, 19, 12, 5, 14, 21, 24, 30, 
    
    -- channel=254
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 55, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 12, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 28, 8, 0, 3, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 62, 93, 49, 24, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    103, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=255
    12, 11, 7, 13, 1, 0, 1, 3, 7, 8, 5, 5, 2, 0, 0, 
    11, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 4, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 26, 43, 30, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 42, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 20, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=256
    0, 0, 0, 8, 8, 0, 17, 20, 40, 46, 0, 44, 35, 31, 26, 
    0, 0, 0, 0, 31, 32, 0, 13, 13, 10, 67, 31, 29, 23, 19, 
    0, 0, 0, 32, 7, 20, 0, 0, 0, 0, 54, 0, 14, 29, 38, 
    144, 109, 121, 13, 0, 19, 77, 35, 7, 14, 0, 21, 39, 7, 0, 
    54, 89, 26, 8, 8, 0, 6, 0, 0, 0, 0, 27, 17, 8, 0, 
    14, 15, 0, 22, 21, 0, 0, 0, 34, 25, 0, 0, 10, 22, 15, 
    11, 7, 0, 0, 9, 0, 13, 9, 28, 11, 12, 8, 8, 26, 48, 
    6, 0, 5, 0, 32, 5, 0, 39, 0, 18, 0, 0, 0, 0, 0, 
    10, 0, 21, 42, 10, 58, 57, 12, 1, 0, 5, 21, 0, 0, 0, 
    18, 40, 18, 11, 0, 0, 0, 32, 78, 20, 0, 0, 36, 19, 0, 
    7, 16, 0, 27, 28, 9, 0, 0, 0, 2, 0, 25, 11, 0, 0, 
    2, 3, 7, 6, 5, 0, 27, 14, 5, 0, 19, 0, 0, 12, 2, 
    3, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 15, 76, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 7, 17, 0, 
    
    -- channel=257
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 10, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 8, 0, 0, 0, 0, 7, 0, 6, 16, 5, 
    0, 0, 0, 0, 0, 12, 9, 7, 0, 0, 3, 0, 8, 6, 0, 
    0, 0, 0, 0, 0, 16, 10, 0, 0, 0, 3, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 4, 2, 1, 3, 0, 10, 2, 0, 
    0, 0, 0, 0, 7, 10, 13, 2, 4, 4, 10, 21, 14, 15, 9, 
    0, 0, 0, 0, 9, 0, 3, 1, 0, 0, 0, 0, 0, 14, 2, 
    0, 0, 0, 2, 5, 22, 23, 5, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 6, 2, 14, 8, 0, 0, 0, 0, 0, 0, 
    4, 2, 0, 11, 9, 9, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 12, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=258
    0, 133, 70, 38, 37, 62, 47, 49, 0, 0, 96, 45, 47, 50, 47, 
    3, 82, 99, 58, 4, 17, 50, 47, 26, 0, 103, 28, 33, 42, 44, 
    4, 32, 118, 52, 39, 0, 33, 66, 42, 28, 47, 39, 22, 24, 21, 
    0, 11, 60, 13, 71, 0, 0, 0, 22, 79, 21, 52, 12, 5, 45, 
    0, 37, 15, 0, 67, 19, 0, 0, 26, 62, 44, 54, 11, 0, 55, 
    15, 31, 17, 0, 46, 21, 0, 0, 4, 39, 43, 65, 12, 0, 23, 
    19, 30, 17, 29, 10, 18, 0, 38, 0, 29, 33, 63, 22, 0, 0, 
    11, 41, 0, 88, 0, 15, 0, 3, 36, 34, 21, 103, 73, 11, 24, 
    0, 38, 7, 63, 3, 0, 0, 0, 79, 20, 15, 3, 106, 43, 84, 
    0, 19, 29, 19, 31, 31, 15, 0, 0, 34, 18, 37, 32, 22, 71, 
    12, 0, 41, 15, 13, 0, 51, 33, 0, 9, 35, 39, 34, 13, 31, 
    21, 0, 60, 20, 13, 13, 32, 24, 11, 0, 57, 31, 34, 11, 10, 
    14, 2, 59, 16, 0, 60, 47, 35, 16, 11, 52, 30, 40, 35, 21, 
    11, 4, 64, 25, 0, 24, 32, 35, 21, 32, 43, 29, 12, 54, 29, 
    23, 9, 55, 44, 2, 5, 19, 43, 11, 45, 37, 30, 15, 39, 41, 
    
    -- channel=259
    0, 0, 21, 12, 7, 12, 21, 18, 36, 0, 6, 30, 30, 28, 26, 
    0, 0, 0, 0, 21, 0, 8, 25, 7, 14, 32, 26, 18, 17, 20, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 14, 10, 0, 9, 19, 27, 
    45, 30, 40, 0, 0, 15, 40, 7, 0, 0, 2, 13, 23, 5, 1, 
    35, 55, 12, 4, 0, 0, 0, 0, 0, 0, 0, 19, 6, 0, 0, 
    9, 4, 3, 14, 6, 0, 0, 0, 7, 3, 0, 0, 6, 13, 0, 
    4, 3, 0, 15, 0, 0, 0, 10, 10, 5, 0, 7, 1, 22, 24, 
    0, 4, 14, 2, 6, 10, 0, 7, 3, 0, 0, 0, 11, 0, 11, 
    4, 0, 19, 2, 16, 34, 12, 0, 0, 8, 4, 21, 0, 0, 0, 
    10, 16, 12, 11, 0, 0, 1, 25, 30, 0, 0, 2, 22, 5, 0, 
    5, 0, 1, 8, 13, 0, 0, 0, 5, 0, 0, 9, 9, 0, 0, 
    0, 4, 0, 3, 1, 4, 19, 6, 0, 0, 7, 0, 5, 6, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 11, 46, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    
    -- channel=260
    3, 45, 80, 65, 62, 71, 76, 72, 68, 39, 63, 80, 90, 87, 87, 
    5, 28, 68, 60, 51, 45, 49, 64, 58, 35, 82, 69, 77, 82, 83, 
    7, 14, 69, 74, 51, 32, 36, 37, 32, 48, 61, 49, 57, 62, 65, 
    60, 66, 72, 38, 46, 40, 54, 44, 43, 54, 43, 59, 54, 38, 46, 
    42, 64, 48, 37, 55, 42, 37, 28, 37, 45, 43, 64, 55, 35, 45, 
    47, 47, 41, 48, 49, 34, 34, 34, 45, 49, 46, 57, 47, 41, 42, 
    47, 50, 38, 66, 52, 47, 32, 40, 34, 41, 44, 61, 47, 46, 45, 
    38, 46, 58, 74, 37, 41, 28, 43, 42, 35, 35, 17, 46, 39, 45, 
    37, 46, 66, 68, 44, 56, 49, 35, 47, 49, 49, 65, 44, 25, 45, 
    37, 45, 51, 53, 43, 31, 37, 44, 65, 60, 39, 58, 67, 53, 52, 
    41, 36, 48, 55, 53, 38, 49, 44, 37, 40, 48, 58, 58, 47, 44, 
    40, 33, 49, 46, 46, 41, 61, 54, 46, 37, 61, 46, 53, 48, 47, 
    39, 29, 44, 45, 41, 59, 60, 49, 41, 40, 52, 44, 36, 43, 52, 
    35, 31, 40, 43, 41, 81, 47, 50, 42, 39, 49, 48, 39, 52, 51, 
    27, 36, 31, 40, 42, 42, 32, 47, 38, 50, 44, 48, 47, 50, 45, 
    
    -- channel=261
    2, 0, 0, 6, 8, 0, 5, 0, 33, 87, 0, 0, 4, 4, 8, 
    1, 0, 0, 0, 1, 24, 0, 0, 5, 81, 0, 5, 10, 5, 6, 
    2, 0, 0, 0, 0, 81, 8, 0, 0, 0, 0, 0, 0, 0, 10, 
    105, 0, 0, 34, 0, 27, 58, 41, 0, 0, 0, 0, 6, 23, 0, 
    27, 0, 3, 65, 0, 0, 20, 54, 0, 0, 0, 0, 5, 54, 0, 
    3, 0, 4, 38, 0, 0, 38, 24, 0, 0, 0, 0, 5, 56, 4, 
    9, 0, 34, 0, 21, 0, 33, 0, 19, 0, 0, 0, 0, 18, 42, 
    19, 0, 70, 0, 18, 10, 0, 32, 0, 0, 8, 0, 0, 9, 0, 
    46, 0, 0, 0, 0, 9, 35, 54, 0, 24, 0, 61, 0, 0, 0, 
    23, 6, 0, 4, 0, 0, 0, 31, 72, 0, 23, 0, 1, 7, 0, 
    2, 37, 0, 8, 0, 50, 0, 0, 13, 35, 0, 0, 0, 21, 0, 
    0, 36, 0, 0, 11, 14, 0, 0, 15, 53, 0, 0, 0, 22, 24, 
    9, 16, 0, 0, 47, 0, 0, 0, 17, 25, 0, 0, 0, 0, 10, 
    16, 24, 0, 0, 33, 15, 15, 3, 13, 9, 0, 1, 19, 0, 0, 
    7, 7, 0, 0, 16, 23, 24, 0, 28, 0, 0, 0, 14, 0, 0, 
    
    -- channel=262
    0, 17, 137, 134, 123, 126, 127, 130, 129, 61, 82, 150, 149, 148, 146, 
    0, 4, 126, 130, 159, 127, 149, 158, 165, 110, 114, 185, 175, 167, 164, 
    0, 3, 89, 117, 193, 161, 109, 133, 149, 126, 165, 199, 204, 200, 192, 
    17, 8, 116, 143, 194, 188, 123, 104, 96, 124, 203, 207, 229, 226, 214, 
    160, 148, 183, 133, 158, 195, 183, 134, 111, 126, 185, 227, 240, 200, 183, 
    191, 183, 195, 144, 174, 189, 173, 115, 124, 129, 173, 232, 249, 209, 169, 
    189, 179, 159, 178, 158, 154, 160, 134, 159, 157, 165, 226, 249, 241, 183, 
    188, 181, 146, 178, 187, 185, 170, 141, 170, 143, 180, 187, 252, 250, 219, 
    190, 155, 165, 166, 210, 203, 174, 160, 112, 141, 166, 109, 137, 197, 205, 
    201, 165, 195, 196, 195, 217, 222, 184, 128, 145, 148, 132, 117, 140, 145, 
    213, 185, 199, 196, 202, 182, 181, 197, 195, 154, 124, 133, 152, 136, 124, 
    210, 194, 191, 221, 216, 180, 179, 185, 182, 132, 119, 143, 162, 138, 117, 
    202, 184, 186, 218, 198, 113, 185, 177, 166, 123, 127, 130, 139, 134, 121, 
    195, 170, 165, 219, 189, 138, 161, 148, 129, 97, 115, 116, 106, 106, 131, 
    174, 165, 137, 215, 199, 178, 138, 126, 104, 85, 106, 116, 103, 106, 125, 
    
    -- channel=263
    0, 0, 35, 44, 28, 32, 42, 31, 50, 39, 0, 23, 44, 45, 51, 
    0, 0, 16, 25, 11, 11, 19, 25, 35, 65, 0, 25, 36, 38, 45, 
    0, 0, 0, 19, 0, 46, 15, 11, 39, 15, 0, 9, 21, 19, 25, 
    26, 0, 0, 36, 0, 28, 24, 27, 7, 0, 15, 0, 11, 27, 9, 
    29, 0, 15, 49, 0, 9, 27, 43, 6, 0, 0, 0, 17, 40, 3, 
    22, 9, 26, 35, 0, 10, 41, 22, 7, 0, 0, 0, 15, 41, 13, 
    24, 18, 39, 37, 22, 0, 26, 0, 15, 0, 0, 0, 11, 24, 14, 
    24, 20, 71, 0, 16, 18, 13, 16, 18, 0, 25, 0, 20, 28, 12, 
    41, 11, 36, 0, 17, 11, 10, 42, 0, 32, 28, 48, 0, 31, 0, 
    27, 6, 15, 24, 5, 10, 19, 20, 30, 10, 37, 32, 18, 25, 14, 
    16, 27, 3, 14, 13, 38, 2, 10, 32, 41, 27, 13, 23, 35, 22, 
    12, 39, 0, 12, 26, 31, 14, 19, 28, 52, 3, 23, 22, 32, 36, 
    16, 27, 0, 16, 55, 16, 20, 28, 41, 39, 14, 24, 21, 29, 29, 
    21, 30, 0, 7, 35, 20, 33, 36, 38, 26, 15, 23, 32, 9, 20, 
    23, 28, 0, 1, 22, 32, 40, 33, 44, 12, 19, 22, 28, 11, 22, 
    
    -- channel=264
    24, 0, 0, 0, 0, 0, 3, 4, 35, 40, 0, 19, 8, 5, 2, 
    23, 0, 0, 0, 20, 8, 0, 0, 1, 21, 19, 9, 6, 1, 0, 
    23, 9, 0, 7, 0, 19, 0, 0, 0, 0, 31, 0, 0, 2, 9, 
    125, 75, 69, 0, 0, 11, 46, 36, 12, 0, 0, 0, 3, 0, 0, 
    33, 42, 13, 10, 0, 0, 0, 7, 0, 0, 0, 3, 0, 6, 0, 
    4, 0, 0, 3, 4, 0, 0, 0, 29, 4, 0, 0, 0, 18, 9, 
    2, 0, 0, 0, 13, 0, 13, 0, 23, 7, 0, 0, 0, 11, 23, 
    0, 0, 1, 0, 7, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 7, 9, 0, 33, 27, 25, 0, 0, 10, 19, 0, 0, 0, 
    14, 10, 0, 3, 0, 0, 0, 16, 45, 3, 0, 0, 12, 12, 0, 
    0, 5, 0, 5, 3, 8, 0, 0, 0, 5, 0, 9, 2, 0, 0, 
    0, 10, 0, 0, 0, 0, 6, 0, 0, 0, 5, 0, 0, 1, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 1, 0, 0, 5, 19, 0, 0, 0, 0, 2, 0, 0, 0, 1, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 8, 0, 
    
    -- channel=265
    21, 8, 41, 31, 29, 37, 37, 36, 33, 21, 21, 24, 33, 37, 38, 
    21, 11, 42, 28, 13, 19, 29, 33, 28, 33, 8, 29, 31, 33, 33, 
    21, 16, 34, 23, 8, 17, 20, 29, 37, 29, 15, 33, 28, 27, 28, 
    19, 15, 4, 35, 14, 17, 12, 17, 20, 9, 26, 23, 15, 26, 36, 
    39, 18, 34, 38, 10, 15, 17, 21, 19, 12, 25, 28, 29, 47, 44, 
    39, 33, 40, 37, 13, 13, 24, 23, 15, 9, 17, 33, 35, 51, 53, 
    44, 37, 37, 37, 22, 17, 17, 8, 18, 15, 17, 32, 34, 39, 41, 
    46, 35, 29, 20, 18, 17, 18, 8, 31, 18, 28, 32, 48, 39, 45, 
    51, 34, 19, 7, 22, 10, 6, 20, 16, 29, 29, 32, 30, 54, 44, 
    50, 31, 21, 22, 22, 21, 21, 16, 14, 23, 29, 33, 23, 26, 32, 
    43, 37, 27, 21, 22, 26, 22, 17, 26, 26, 35, 22, 22, 29, 26, 
    42, 48, 22, 17, 19, 21, 21, 21, 23, 36, 24, 25, 24, 26, 31, 
    44, 56, 34, 20, 23, 15, 26, 28, 31, 31, 29, 27, 26, 34, 27, 
    46, 58, 43, 24, 26, 4, 26, 33, 34, 34, 28, 29, 30, 26, 27, 
    50, 58, 42, 25, 24, 27, 33, 33, 34, 31, 30, 29, 30, 23, 30, 
    
    -- channel=266
    0, 0, 103, 77, 64, 76, 81, 85, 96, 2, 65, 122, 112, 109, 105, 
    0, 0, 89, 74, 116, 63, 87, 110, 109, 57, 112, 133, 121, 116, 112, 
    0, 0, 77, 71, 141, 85, 32, 47, 54, 84, 126, 127, 137, 140, 135, 
    41, 56, 126, 65, 130, 134, 93, 60, 56, 79, 136, 158, 161, 137, 138, 
    128, 125, 129, 64, 112, 122, 112, 58, 60, 70, 129, 172, 166, 118, 110, 
    128, 118, 125, 86, 122, 110, 90, 56, 89, 84, 107, 168, 167, 136, 105, 
    122, 116, 76, 130, 93, 96, 91, 86, 104, 103, 106, 169, 171, 176, 122, 
    110, 110, 79, 144, 119, 112, 107, 76, 114, 80, 100, 74, 163, 155, 147, 
    115, 90, 128, 110, 150, 162, 120, 101, 57, 73, 120, 58, 51, 92, 130, 
    138, 109, 132, 129, 118, 119, 143, 133, 86, 104, 75, 85, 84, 89, 66, 
    142, 104, 140, 135, 143, 106, 116, 116, 127, 78, 70, 90, 97, 72, 63, 
    133, 121, 132, 145, 135, 107, 130, 122, 112, 63, 82, 80, 109, 79, 66, 
    126, 110, 121, 143, 110, 36, 125, 101, 86, 55, 76, 67, 63, 70, 71, 
    117, 95, 97, 150, 127, 103, 89, 76, 57, 35, 67, 61, 48, 59, 84, 
    86, 101, 63, 144, 126, 102, 54, 62, 37, 42, 53, 67, 59, 61, 66, 
    
    -- channel=267
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 22, 45, 57, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 11, 0, 0, 0, 0, 0, 6, 0, 0, 18, 2, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 5, 7, 
    0, 0, 6, 0, 0, 9, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 5, 3, 0, 0, 2, 0, 0, 7, 0, 26, 81, 39, 25, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 72, 21, 
    0, 0, 0, 0, 3, 33, 6, 0, 0, 0, 24, 0, 0, 0, 33, 
    0, 2, 0, 0, 0, 7, 4, 9, 0, 26, 0, 0, 0, 0, 5, 
    2, 4, 0, 0, 7, 7, 0, 0, 3, 8, 0, 3, 0, 0, 0, 
    3, 12, 0, 0, 28, 10, 6, 17, 26, 12, 1, 5, 31, 14, 0, 
    9, 15, 0, 0, 0, 0, 19, 21, 24, 8, 0, 0, 6, 0, 0, 
    31, 7, 7, 10, 0, 8, 36, 21, 22, 0, 2, 0, 0, 0, 11, 
    
    -- channel=268
    22, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    21, 9, 0, 0, 26, 13, 1, 0, 4, 7, 6, 6, 0, 0, 0, 
    18, 17, 0, 0, 34, 35, 17, 9, 8, 6, 25, 16, 13, 12, 8, 
    16, 8, 14, 4, 31, 35, 21, 19, 17, 15, 30, 18, 29, 30, 16, 
    7, 6, 16, 5, 27, 36, 31, 23, 21, 20, 24, 19, 27, 16, 7, 
    11, 14, 13, 2, 23, 34, 30, 20, 28, 24, 26, 20, 26, 14, 2, 
    6, 6, 2, 3, 26, 31, 36, 21, 33, 31, 28, 20, 23, 21, 8, 
    8, 6, 1, 6, 29, 32, 35, 31, 18, 17, 22, 9, 8, 25, 13, 
    12, 9, 13, 16, 30, 35, 37, 37, 8, 4, 15, 0, 6, 10, 2, 
    13, 10, 24, 22, 29, 37, 35, 33, 18, 9, 12, 0, 0, 5, 1, 
    16, 18, 23, 23, 21, 27, 25, 27, 26, 15, 0, 6, 11, 8, 5, 
    17, 17, 22, 31, 28, 14, 15, 19, 21, 7, 1, 9, 13, 8, 4, 
    15, 9, 13, 35, 32, 1, 13, 11, 11, 4, 4, 7, 13, 5, 6, 
    12, 3, 2, 33, 26, 7, 10, 3, 3, 0, 5, 5, 7, 2, 6, 
    8, 3, 0, 34, 28, 21, 5, 0, 3, 0, 3, 5, 3, 5, 5, 
    
    -- channel=269
    4, 10, 0, 3, 7, 0, 2, 10, 19, 20, 19, 26, 11, 10, 4, 
    5, 8, 0, 7, 42, 30, 8, 22, 19, 5, 61, 33, 22, 16, 9, 
    4, 4, 0, 24, 45, 30, 0, 0, 0, 15, 61, 31, 35, 39, 37, 
    69, 68, 76, 17, 28, 40, 53, 26, 18, 38, 34, 53, 56, 37, 30, 
    43, 67, 42, 12, 42, 35, 29, 11, 17, 29, 35, 57, 48, 31, 33, 
    34, 38, 28, 27, 42, 33, 16, 18, 41, 44, 36, 48, 50, 40, 35, 
    33, 31, 7, 19, 35, 35, 30, 30, 43, 38, 44, 52, 52, 54, 54, 
    31, 22, 1, 27, 45, 38, 29, 43, 15, 37, 25, 0, 21, 36, 43, 
    31, 22, 19, 50, 44, 65, 61, 24, 22, 16, 21, 17, 2, 0, 24, 
    42, 47, 37, 35, 38, 27, 32, 48, 51, 28, 5, 3, 30, 21, 9, 
    42, 38, 36, 48, 47, 31, 28, 31, 22, 12, 2, 25, 22, 8, 9, 
    40, 31, 44, 41, 36, 12, 43, 35, 27, 0, 25, 15, 19, 18, 11, 
    37, 26, 39, 41, 13, 0, 19, 14, 3, 0, 12, 9, 3, 0, 13, 
    31, 22, 32, 42, 29, 42, 14, 0, 0, 0, 11, 10, 4, 11, 16, 
    13, 19, 30, 36, 35, 23, 0, 0, 0, 9, 7, 12, 13, 18, 6, 
    
    -- channel=270
    0, 0, 0, 8, 7, 0, 0, 0, 7, 43, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 16, 0, 0, 23, 43, 0, 8, 14, 8, 10, 
    0, 0, 0, 0, 0, 68, 22, 19, 42, 0, 0, 9, 21, 13, 13, 
    0, 0, 0, 35, 0, 31, 4, 19, 0, 0, 30, 0, 27, 60, 6, 
    3, 0, 15, 39, 0, 27, 42, 50, 0, 0, 0, 0, 35, 60, 2, 
    18, 9, 29, 12, 0, 30, 60, 12, 0, 0, 0, 0, 38, 54, 10, 
    22, 8, 50, 5, 33, 2, 52, 0, 29, 0, 0, 0, 30, 35, 14, 
    34, 9, 55, 0, 34, 29, 22, 31, 0, 0, 37, 13, 9, 66, 5, 
    52, 2, 7, 0, 14, 11, 25, 59, 0, 10, 19, 13, 2, 50, 0, 
    31, 0, 17, 23, 28, 51, 28, 18, 20, 0, 43, 0, 0, 15, 12, 
    24, 43, 0, 21, 15, 59, 7, 26, 37, 57, 0, 0, 9, 25, 11, 
    26, 49, 0, 30, 49, 26, 4, 17, 37, 42, 0, 13, 7, 19, 11, 
    29, 36, 0, 35, 88, 0, 18, 28, 45, 23, 0, 8, 28, 6, 8, 
    32, 33, 0, 23, 42, 0, 40, 24, 31, 0, 0, 2, 16, 0, 0, 
    29, 19, 0, 13, 34, 49, 38, 9, 31, 0, 0, 0, 0, 0, 3, 
    
    -- channel=271
    3, 0, 0, 4, 3, 0, 0, 1, 20, 13, 9, 11, 4, 1, 0, 
    2, 0, 0, 11, 45, 16, 7, 15, 15, 26, 24, 23, 14, 8, 5, 
    2, 0, 0, 10, 47, 43, 5, 0, 0, 28, 30, 23, 30, 31, 29, 
    38, 33, 24, 9, 34, 54, 47, 25, 16, 22, 34, 37, 52, 36, 27, 
    32, 35, 25, 18, 28, 41, 37, 27, 18, 24, 29, 36, 42, 23, 8, 
    24, 24, 18, 24, 33, 38, 31, 28, 33, 34, 30, 29, 41, 29, 7, 
    17, 19, 2, 24, 31, 36, 34, 36, 40, 36, 33, 31, 39, 44, 32, 
    14, 14, 16, 23, 41, 41, 42, 33, 27, 23, 24, 0, 25, 29, 33, 
    19, 11, 30, 32, 50, 61, 56, 38, 4, 22, 19, 15, 0, 0, 10, 
    26, 26, 32, 39, 30, 30, 48, 57, 38, 21, 8, 6, 22, 13, 0, 
    29, 26, 32, 40, 43, 33, 25, 35, 36, 11, 11, 16, 21, 14, 5, 
    24, 24, 27, 44, 37, 30, 34, 34, 28, 15, 10, 15, 21, 18, 15, 
    22, 11, 20, 43, 26, 11, 21, 17, 13, 9, 6, 12, 4, 9, 13, 
    19, 5, 8, 39, 38, 36, 13, 6, 2, 3, 5, 10, 7, 6, 14, 
    6, 5, 1, 35, 39, 22, 3, 1, 0, 2, 5, 8, 13, 7, 7, 
    
    -- channel=272
    0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 85, 0, 0, 0, 0, 
    1, 31, 0, 0, 0, 0, 0, 0, 0, 0, 87, 0, 0, 0, 0, 
    0, 3, 45, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    53, 176, 39, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=273
    0, 3, 0, 11, 18, 10, 12, 12, 17, 32, 2, 0, 5, 4, 4, 
    0, 6, 0, 11, 4, 15, 0, 0, 0, 0, 0, 10, 19, 14, 9, 
    0, 1, 8, 29, 0, 9, 27, 11, 7, 6, 18, 16, 14, 11, 12, 
    39, 21, 0, 3, 0, 0, 5, 19, 14, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 16, 8, 0, 6, 5, 12, 0, 6, 9, 11, 12, 
    0, 3, 0, 3, 0, 0, 12, 18, 6, 11, 13, 8, 10, 11, 13, 
    9, 8, 5, 0, 43, 33, 10, 0, 0, 8, 9, 3, 3, 0, 15, 
    5, 0, 3, 1, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    12, 21, 0, 21, 0, 3, 18, 11, 11, 8, 0, 28, 37, 2, 0, 
    2, 2, 1, 10, 20, 4, 0, 4, 27, 0, 4, 1, 7, 0, 24, 
    4, 10, 3, 13, 0, 13, 11, 6, 0, 2, 2, 4, 6, 13, 0, 
    6, 2, 7, 0, 0, 0, 0, 2, 0, 7, 2, 3, 0, 0, 8, 
    7, 0, 4, 9, 15, 31, 0, 3, 2, 2, 3, 5, 2, 1, 10, 
    3, 3, 13, 4, 0, 0, 7, 8, 5, 10, 7, 8, 5, 9, 0, 
    6, 3, 13, 0, 5, 3, 0, 0, 9, 4, 7, 0, 5, 0, 6, 
    
    -- channel=274
    0, 0, 2, 2, 0, 2, 2, 3, 0, 0, 2, 12, 14, 15, 13, 
    0, 0, 1, 12, 4, 8, 10, 17, 20, 0, 14, 25, 24, 23, 20, 
    0, 0, 0, 12, 30, 2, 4, 16, 11, 0, 26, 37, 32, 29, 25, 
    0, 0, 0, 10, 37, 10, 0, 0, 0, 21, 31, 43, 47, 44, 46, 
    0, 13, 27, 0, 29, 32, 17, 0, 0, 16, 32, 51, 52, 33, 43, 
    29, 35, 29, 8, 25, 31, 16, 0, 0, 12, 31, 55, 55, 28, 28, 
    32, 33, 28, 13, 21, 22, 6, 6, 7, 14, 30, 56, 60, 41, 27, 
    32, 33, 1, 24, 24, 26, 11, 14, 14, 27, 28, 56, 62, 56, 47, 
    21, 25, 3, 36, 28, 22, 21, 0, 23, 14, 8, 0, 46, 41, 53, 
    26, 24, 31, 27, 43, 50, 37, 16, 0, 9, 12, 1, 3, 6, 32, 
    39, 28, 36, 36, 33, 24, 36, 42, 19, 13, 3, 6, 13, 5, 3, 
    44, 21, 41, 42, 39, 23, 27, 31, 26, 0, 6, 13, 13, 6, 0, 
    39, 27, 41, 43, 23, 28, 28, 31, 19, 0, 7, 7, 14, 5, 0, 
    34, 21, 34, 41, 16, 5, 22, 16, 5, 0, 0, 1, 0, 2, 1, 
    29, 13, 27, 43, 31, 22, 8, 2, 0, 0, 0, 0, 0, 0, 6, 
    
    -- channel=275
    0, 0, 4, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 1, 4, 0, 0, 5, 8, 2, 1, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 12, 11, 7, 6, 6, 
    4, 0, 20, 2, 0, 0, 0, 0, 0, 0, 8, 8, 3, 11, 12, 
    12, 17, 14, 5, 0, 0, 0, 0, 0, 0, 5, 17, 11, 15, 18, 
    14, 11, 17, 3, 0, 0, 0, 0, 0, 0, 4, 16, 18, 26, 27, 
    18, 12, 5, 5, 0, 0, 0, 0, 0, 5, 0, 16, 16, 20, 24, 
    18, 10, 0, 0, 0, 3, 0, 0, 2, 0, 5, 4, 14, 17, 20, 
    24, 11, 0, 0, 3, 6, 0, 0, 0, 0, 5, 5, 0, 7, 17, 
    24, 14, 3, 2, 3, 0, 0, 0, 4, 0, 0, 0, 0, 2, 4, 
    21, 16, 8, 2, 5, 4, 1, 0, 2, 1, 0, 0, 0, 0, 0, 
    20, 21, 8, 2, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 
    22, 23, 14, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 25, 18, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 26, 15, 7, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=276
    9, 0, 0, 5, 2, 0, 0, 0, 29, 92, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 19, 0, 0, 7, 110, 0, 0, 2, 0, 0, 
    7, 0, 0, 0, 0, 98, 9, 0, 5, 0, 0, 0, 0, 0, 1, 
    81, 0, 0, 39, 0, 40, 47, 42, 0, 0, 0, 0, 0, 34, 0, 
    40, 0, 0, 79, 0, 0, 35, 73, 0, 0, 0, 0, 3, 69, 0, 
    4, 0, 8, 37, 0, 0, 49, 29, 0, 0, 0, 0, 1, 68, 0, 
    6, 0, 45, 0, 6, 0, 51, 0, 22, 0, 0, 0, 0, 22, 32, 
    24, 0, 84, 0, 27, 0, 17, 25, 0, 0, 7, 0, 0, 21, 0, 
    56, 0, 7, 0, 0, 0, 26, 78, 0, 16, 0, 40, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 28, 53, 0, 35, 0, 0, 9, 0, 
    2, 40, 0, 0, 0, 56, 0, 0, 31, 49, 0, 0, 0, 27, 4, 
    0, 51, 0, 0, 14, 29, 0, 0, 20, 72, 0, 0, 0, 25, 23, 
    9, 30, 0, 0, 68, 0, 0, 1, 32, 37, 0, 1, 0, 0, 8, 
    20, 34, 0, 0, 50, 0, 17, 6, 27, 7, 0, 0, 27, 0, 0, 
    16, 15, 0, 0, 19, 34, 43, 0, 43, 0, 0, 0, 11, 0, 0, 
    
    -- channel=277
    0, 154, 26, 0, 0, 15, 0, 14, 0, 0, 116, 14, 1, 3, 0, 
    4, 98, 54, 31, 0, 0, 14, 17, 0, 0, 154, 0, 0, 0, 0, 
    3, 36, 106, 44, 43, 0, 0, 22, 0, 17, 63, 16, 0, 3, 0, 
    0, 82, 102, 0, 62, 0, 0, 0, 11, 95, 0, 59, 0, 0, 18, 
    0, 59, 0, 0, 80, 1, 0, 0, 16, 66, 29, 53, 0, 0, 35, 
    0, 12, 0, 0, 44, 0, 0, 0, 9, 55, 33, 61, 0, 0, 0, 
    0, 3, 0, 9, 0, 18, 0, 39, 0, 26, 34, 57, 0, 0, 0, 
    0, 9, 0, 82, 0, 0, 0, 0, 8, 24, 0, 46, 34, 0, 8, 
    0, 14, 0, 61, 0, 0, 0, 0, 66, 0, 0, 0, 74, 0, 63, 
    0, 13, 9, 0, 13, 0, 0, 0, 0, 29, 0, 0, 26, 0, 33, 
    0, 0, 29, 1, 3, 0, 34, 13, 0, 0, 1, 21, 9, 0, 0, 
    0, 0, 61, 0, 0, 0, 21, 3, 0, 0, 51, 0, 7, 0, 0, 
    0, 0, 50, 0, 0, 22, 17, 0, 0, 0, 29, 0, 0, 0, 0, 
    0, 0, 55, 11, 0, 27, 0, 0, 0, 0, 17, 2, 0, 35, 6, 
    0, 0, 44, 30, 0, 0, 0, 0, 0, 34, 7, 4, 0, 21, 5, 
    
    -- channel=278
    26, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=279
    12, 0, 23, 33, 24, 28, 34, 25, 46, 33, 0, 15, 32, 30, 36, 
    11, 0, 0, 10, 9, 9, 15, 12, 19, 69, 0, 17, 23, 25, 31, 
    12, 0, 0, 1, 0, 41, 5, 0, 22, 17, 0, 0, 12, 12, 18, 
    33, 0, 0, 24, 0, 27, 28, 24, 3, 0, 0, 0, 0, 9, 0, 
    38, 0, 4, 46, 0, 0, 19, 39, 2, 0, 0, 0, 1, 28, 0, 
    11, 0, 12, 31, 0, 0, 24, 19, 2, 0, 0, 0, 0, 35, 3, 
    10, 5, 21, 19, 0, 0, 19, 0, 7, 0, 0, 0, 0, 16, 15, 
    13, 6, 60, 0, 9, 2, 12, 2, 6, 0, 6, 0, 0, 4, 1, 
    30, 0, 33, 0, 8, 3, 2, 38, 0, 22, 16, 35, 0, 5, 0, 
    21, 3, 0, 8, 0, 0, 3, 19, 25, 1, 23, 22, 11, 16, 0, 
    5, 14, 0, 0, 3, 22, 0, 0, 26, 23, 20, 5, 9, 25, 14, 
    0, 29, 0, 0, 5, 27, 0, 3, 13, 47, 0, 11, 9, 24, 28, 
    4, 18, 0, 0, 29, 0, 0, 10, 25, 33, 1, 14, 5, 19, 20, 
    11, 22, 0, 0, 34, 19, 13, 19, 26, 21, 5, 14, 25, 0, 13, 
    13, 22, 0, 0, 11, 17, 33, 22, 35, 7, 11, 13, 24, 5, 10, 
    
    -- channel=280
    0, 93, 22, 0, 0, 11, 0, 0, 0, 0, 69, 0, 0, 0, 0, 
    0, 46, 64, 25, 0, 0, 29, 13, 0, 0, 51, 0, 0, 0, 0, 
    0, 2, 79, 0, 38, 0, 16, 61, 40, 11, 15, 39, 10, 3, 0, 
    0, 0, 0, 0, 73, 0, 0, 0, 0, 59, 25, 50, 11, 11, 55, 
    0, 0, 3, 0, 51, 27, 0, 0, 10, 47, 50, 43, 17, 0, 50, 
    8, 23, 15, 0, 32, 28, 0, 0, 0, 19, 39, 73, 25, 0, 13, 
    9, 18, 7, 10, 0, 17, 0, 30, 0, 17, 32, 62, 37, 0, 0, 
    9, 31, 0, 65, 0, 9, 6, 0, 41, 31, 20, 136, 95, 28, 37, 
    0, 24, 0, 28, 11, 0, 0, 0, 59, 1, 0, 0, 101, 74, 99, 
    0, 4, 14, 6, 35, 53, 37, 0, 0, 9, 0, 8, 0, 0, 49, 
    19, 0, 44, 4, 9, 0, 50, 40, 2, 0, 18, 2, 3, 0, 7, 
    29, 0, 57, 25, 12, 16, 11, 12, 3, 0, 20, 11, 16, 0, 0, 
    19, 9, 56, 21, 0, 42, 36, 25, 9, 0, 26, 11, 28, 23, 0, 
    16, 3, 61, 33, 0, 0, 6, 16, 5, 9, 13, 2, 0, 23, 4, 
    33, 5, 49, 59, 6, 0, 10, 20, 0, 12, 10, 3, 0, 4, 19, 
    
    -- channel=281
    13, 78, 17, 1, 1, 15, 6, 20, 13, 0, 92, 7, 6, 7, 2, 
    15, 49, 20, 29, 13, 0, 1, 10, 0, 0, 92, 4, 2, 3, 0, 
    13, 20, 71, 30, 21, 0, 0, 0, 0, 45, 19, 12, 1, 7, 5, 
    28, 122, 43, 0, 21, 0, 5, 0, 15, 47, 0, 40, 0, 0, 9, 
    2, 31, 0, 0, 35, 0, 0, 0, 11, 32, 11, 23, 0, 0, 11, 
    0, 1, 0, 5, 10, 0, 0, 7, 12, 34, 7, 27, 0, 0, 2, 
    0, 5, 0, 18, 0, 29, 0, 27, 0, 11, 19, 22, 0, 0, 1, 
    0, 1, 0, 41, 0, 0, 0, 0, 11, 0, 0, 0, 12, 0, 16, 
    0, 14, 11, 11, 8, 6, 0, 0, 20, 2, 0, 0, 7, 0, 24, 
    0, 12, 0, 0, 0, 0, 0, 2, 0, 21, 0, 9, 32, 0, 0, 
    0, 0, 21, 2, 1, 0, 9, 0, 0, 0, 22, 12, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 6, 0, 0, 0, 28, 0, 0, 0, 0, 
    0, 0, 24, 0, 0, 17, 0, 0, 0, 0, 12, 0, 0, 1, 0, 
    0, 0, 33, 1, 0, 19, 0, 0, 0, 6, 6, 4, 0, 22, 8, 
    0, 0, 20, 8, 0, 0, 0, 0, 0, 30, 6, 5, 9, 4, 0, 
    
    -- channel=282
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=283
    0, 0, 16, 9, 1, 7, 4, 2, 0, 0, 0, 25, 15, 13, 13, 
    0, 0, 27, 13, 17, 7, 25, 22, 26, 0, 8, 25, 20, 20, 21, 
    0, 0, 14, 0, 43, 10, 10, 22, 23, 0, 24, 31, 29, 27, 23, 
    0, 0, 13, 9, 55, 25, 0, 0, 0, 20, 40, 40, 51, 49, 39, 
    0, 9, 21, 0, 32, 40, 31, 7, 3, 18, 37, 45, 40, 12, 18, 
    20, 24, 27, 0, 38, 44, 24, 0, 1, 10, 31, 49, 42, 5, 1, 
    16, 19, 25, 13, 11, 10, 15, 22, 22, 24, 21, 49, 46, 32, 5, 
    13, 27, 7, 48, 30, 32, 26, 12, 30, 22, 29, 67, 58, 47, 20, 
    4, 12, 23, 39, 34, 35, 18, 15, 23, 3, 25, 0, 31, 33, 41, 
    12, 9, 37, 31, 37, 51, 47, 23, 0, 9, 28, 10, 0, 17, 23, 
    25, 11, 37, 30, 31, 24, 37, 39, 35, 26, 1, 14, 21, 10, 10, 
    26, 9, 38, 48, 48, 40, 30, 32, 31, 2, 7, 19, 27, 8, 0, 
    20, 9, 29, 41, 39, 14, 37, 33, 26, 1, 12, 10, 25, 13, 3, 
    18, 0, 14, 42, 27, 5, 35, 17, 6, 0, 8, 0, 0, 3, 8, 
    12, 0, 3, 49, 30, 25, 17, 14, 0, 0, 2, 2, 0, 3, 13, 
    
    -- channel=284
    0, 58, 10, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 
    0, 32, 52, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 43, 0, 0, 0, 9, 49, 34, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 16, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 10, 5, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 14, 0, 0, 98, 37, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 73, 54, 42, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 16, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 29, 12, 4, 0, 0, 8, 0, 19, 9, 0, 
    0, 0, 8, 0, 0, 0, 0, 7, 4, 0, 0, 0, 0, 5, 0, 
    2, 0, 7, 13, 0, 0, 7, 13, 0, 1, 0, 0, 0, 0, 5, 
    
    -- channel=285
    21, 0, 0, 5, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    21, 0, 0, 9, 0, 0, 0, 0, 4, 34, 0, 0, 0, 0, 0, 
    23, 13, 0, 0, 0, 18, 24, 23, 34, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 4, 0, 7, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 4, 11, 28, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 23, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 1, 1, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 11, 2, 5, 0, 2, 13, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 19, 0, 7, 1, 3, 9, 24, 0, 
    0, 0, 0, 0, 0, 11, 4, 0, 0, 0, 19, 8, 0, 0, 1, 
    0, 0, 0, 0, 0, 10, 0, 5, 8, 19, 9, 0, 0, 16, 10, 
    0, 0, 0, 0, 0, 20, 0, 0, 5, 26, 0, 6, 1, 8, 9, 
    0, 0, 0, 0, 30, 38, 4, 10, 24, 22, 0, 11, 20, 16, 7, 
    0, 0, 0, 0, 3, 0, 10, 18, 26, 17, 2, 9, 20, 0, 1, 
    0, 0, 0, 0, 0, 7, 28, 18, 29, 0, 7, 5, 6, 0, 9, 
    
    -- channel=286
    0, 0, 6, 0, 0, 0, 0, 5, 12, 0, 37, 31, 17, 14, 9, 
    0, 0, 0, 0, 36, 0, 0, 13, 8, 0, 81, 33, 22, 18, 10, 
    0, 0, 21, 18, 48, 0, 0, 0, 0, 12, 55, 27, 29, 34, 32, 
    54, 86, 74, 0, 29, 29, 36, 0, 4, 32, 22, 62, 46, 10, 26, 
    25, 53, 30, 0, 46, 26, 8, 0, 0, 17, 29, 63, 45, 5, 21, 
    22, 24, 11, 10, 32, 10, 0, 0, 28, 36, 24, 55, 41, 17, 13, 
    17, 19, 0, 29, 25, 38, 5, 13, 18, 26, 36, 59, 45, 45, 28, 
    6, 9, 0, 42, 18, 18, 12, 14, 10, 12, 1, 0, 22, 17, 36, 
    5, 12, 29, 39, 40, 61, 47, 3, 4, 0, 12, 3, 0, 0, 19, 
    23, 28, 32, 22, 28, 9, 24, 41, 35, 27, 0, 0, 25, 1, 0, 
    27, 9, 38, 41, 39, 6, 27, 21, 9, 0, 0, 16, 12, 0, 0, 
    23, 6, 44, 32, 18, 0, 39, 26, 12, 0, 19, 0, 13, 0, 0, 
    17, 0, 30, 35, 0, 0, 19, 0, 0, 0, 2, 0, 0, 0, 0, 
    8, 0, 18, 37, 18, 40, 0, 0, 0, 0, 0, 0, 0, 2, 6, 
    0, 0, 0, 34, 22, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=287
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 0, 12, 18, 0, 1, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 5, 1, 9, 11, 0, 0, 0, 0, 15, 0, 15, 24, 0, 
    0, 0, 3, 0, 5, 14, 17, 9, 3, 0, 6, 4, 11, 3, 0, 
    0, 1, 4, 0, 11, 20, 11, 0, 8, 3, 8, 6, 11, 2, 0, 
    0, 0, 0, 0, 0, 0, 18, 3, 17, 10, 7, 5, 9, 6, 0, 
    2, 0, 0, 0, 18, 16, 11, 24, 0, 6, 14, 16, 0, 19, 0, 
    3, 0, 0, 2, 9, 12, 15, 13, 0, 0, 6, 0, 0, 2, 0, 
    0, 0, 6, 6, 10, 24, 17, 3, 1, 0, 0, 0, 0, 0, 0, 
    3, 10, 1, 3, 9, 10, 7, 11, 9, 11, 0, 0, 0, 0, 0, 
    6, 7, 3, 15, 18, 2, 2, 3, 9, 0, 0, 0, 0, 0, 0, 
    5, 1, 0, 13, 18, 0, 4, 0, 0, 0, 0, 0, 4, 0, 0, 
    4, 0, 0, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=288
    36, 43, 29, 5, 2, 34, 58, 94, 58, 17, 17, 3, 43, 54, 31, 
    24, 25, 16, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 6, 
    9, 8, 0, 22, 0, 42, 49, 51, 13, 0, 0, 20, 9, 0, 0, 
    9, 4, 0, 0, 11, 14, 26, 0, 5, 31, 15, 0, 0, 49, 4, 
    2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 18, 37, 103, 
    0, 0, 13, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 
    0, 0, 0, 0, 71, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 24, 7, 0, 0, 7, 8, 54, 155, 170, 147, 168, 150, 45, 0, 
    8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 21, 0, 0, 0, 35, 31, 0, 6, 0, 17, 7, 11, 16, 
    0, 0, 0, 59, 32, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 65, 103, 0, 2, 23, 0, 0, 0, 62, 90, 49, 0, 0, 28, 
    10, 0, 0, 0, 0, 0, 12, 14, 13, 0, 0, 0, 0, 3, 0, 
    0, 0, 5, 0, 0, 0, 14, 10, 2, 0, 0, 0, 13, 0, 24, 
    
    -- channel=289
    12, 5, 12, 19, 11, 8, 8, 3, 9, 22, 17, 16, 9, 0, 6, 
    24, 22, 26, 51, 41, 47, 52, 62, 57, 43, 21, 11, 20, 16, 4, 
    29, 29, 34, 37, 32, 28, 36, 33, 31, 28, 10, 9, 16, 14, 3, 
    29, 29, 32, 61, 43, 65, 72, 75, 65, 62, 35, 17, 15, 2, 2, 
    29, 29, 58, 73, 43, 67, 77, 71, 69, 75, 61, 14, 18, 8, 0, 
    27, 36, 38, 62, 43, 53, 59, 69, 65, 60, 69, 42, 16, 29, 28, 
    16, 35, 23, 37, 37, 56, 71, 51, 54, 65, 48, 40, 43, 54, 30, 
    18, 36, 0, 19, 68, 37, 35, 45, 54, 48, 42, 51, 42, 39, 17, 
    7, 30, 0, 47, 34, 39, 42, 14, 0, 0, 0, 0, 0, 41, 32, 
    21, 41, 11, 25, 27, 26, 25, 43, 45, 42, 51, 43, 44, 48, 25, 
    24, 42, 0, 15, 11, 19, 7, 22, 20, 21, 21, 3, 31, 20, 25, 
    37, 53, 10, 0, 11, 7, 33, 40, 13, 39, 22, 32, 52, 25, 26, 
    44, 18, 0, 21, 21, 2, 1, 1, 1, 0, 22, 26, 22, 3, 11, 
    36, 50, 42, 23, 27, 14, 0, 0, 5, 20, 41, 40, 12, 0, 25, 
    53, 46, 35, 30, 22, 14, 0, 0, 4, 14, 29, 35, 6, 1, 11, 
    
    -- channel=290
    0, 5, 0, 0, 10, 9, 2, 2, 18, 8, 10, 20, 0, 7, 0, 
    4, 5, 0, 0, 17, 30, 41, 46, 53, 54, 28, 30, 18, 0, 35, 
    8, 9, 0, 0, 0, 0, 0, 0, 0, 6, 67, 23, 4, 0, 68, 
    8, 0, 0, 0, 35, 10, 0, 0, 0, 0, 8, 63, 0, 0, 34, 
    14, 0, 0, 0, 16, 7, 0, 0, 0, 0, 0, 55, 30, 0, 0, 
    43, 0, 0, 0, 33, 0, 0, 0, 0, 0, 3, 38, 57, 7, 9, 
    40, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 49, 77, 68, 27, 
    23, 0, 57, 0, 0, 0, 0, 0, 12, 14, 0, 30, 58, 39, 83, 
    0, 0, 58, 0, 9, 14, 0, 0, 0, 0, 0, 0, 0, 0, 114, 
    0, 0, 48, 0, 35, 0, 26, 57, 0, 17, 0, 9, 12, 0, 117, 
    5, 0, 0, 0, 0, 23, 0, 0, 45, 0, 0, 0, 0, 0, 95, 
    0, 0, 38, 0, 0, 17, 66, 0, 96, 9, 0, 31, 0, 37, 114, 
    0, 0, 0, 0, 0, 0, 2, 10, 24, 59, 0, 0, 0, 20, 101, 
    0, 0, 0, 0, 0, 0, 0, 6, 25, 75, 33, 0, 0, 42, 83, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 32, 0, 0, 31, 80, 
    
    -- channel=291
    12, 18, 3, 0, 4, 20, 42, 58, 39, 12, 6, 4, 27, 16, 22, 
    9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 8, 13, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 27, 43, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 10, 0, 0, 0, 0, 34, 41, 58, 76, 92, 72, 44, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 
    0, 41, 14, 0, 0, 0, 0, 0, 0, 37, 65, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=292
    46, 55, 49, 29, 33, 38, 37, 48, 47, 39, 40, 42, 46, 45, 36, 
    45, 46, 33, 0, 0, 0, 0, 0, 0, 16, 26, 49, 43, 34, 45, 
    44, 43, 30, 9, 13, 20, 19, 17, 11, 13, 42, 49, 42, 28, 39, 
    44, 41, 37, 0, 11, 6, 0, 0, 0, 0, 20, 41, 44, 39, 37, 
    45, 37, 2, 0, 5, 0, 0, 0, 0, 0, 0, 36, 50, 51, 72, 
    48, 27, 31, 0, 0, 1, 0, 0, 0, 0, 0, 17, 52, 43, 44, 
    52, 24, 32, 10, 10, 0, 0, 0, 0, 0, 0, 4, 10, 13, 44, 
    47, 13, 48, 26, 0, 13, 7, 0, 0, 0, 0, 0, 0, 17, 49, 
    46, 15, 50, 0, 13, 0, 5, 19, 58, 53, 42, 55, 56, 9, 33, 
    43, 0, 12, 9, 0, 4, 6, 5, 3, 7, 0, 3, 2, 0, 44, 
    41, 0, 22, 9, 8, 1, 32, 6, 25, 21, 20, 50, 1, 23, 37, 
    27, 0, 11, 28, 3, 8, 0, 0, 6, 0, 15, 2, 0, 0, 37, 
    21, 29, 38, 12, 7, 3, 1, 5, 12, 44, 26, 6, 0, 11, 44, 
    26, 9, 8, 3, 3, 0, 10, 10, 13, 9, 9, 0, 0, 17, 32, 
    8, 12, 9, 0, 3, 1, 11, 13, 13, 13, 11, 0, 4, 18, 45, 
    
    -- channel=293
    8, 10, 11, 41, 0, 0, 0, 0, 0, 0, 8, 0, 30, 8, 30, 
    0, 0, 17, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 
    0, 0, 22, 148, 0, 3, 9, 36, 14, 0, 0, 0, 21, 34, 0, 
    0, 8, 16, 113, 0, 0, 49, 0, 0, 0, 28, 0, 9, 36, 15, 
    0, 13, 44, 65, 0, 0, 5, 0, 0, 0, 7, 0, 0, 39, 19, 
    0, 20, 47, 105, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 34, 5, 44, 0, 0, 6, 8, 0, 0, 19, 0, 0, 0, 0, 
    2, 69, 0, 58, 3, 33, 3, 13, 0, 0, 0, 0, 0, 0, 0, 
    25, 92, 0, 62, 0, 0, 0, 48, 18, 10, 68, 39, 0, 0, 0, 
    27, 126, 0, 63, 0, 20, 0, 0, 23, 0, 1, 0, 0, 42, 0, 
    2, 129, 15, 23, 20, 0, 0, 73, 0, 35, 8, 0, 43, 0, 0, 
    8, 150, 0, 10, 79, 0, 0, 33, 0, 0, 0, 0, 90, 0, 0, 
    0, 100, 20, 0, 49, 49, 0, 0, 0, 0, 19, 83, 54, 0, 0, 
    0, 15, 50, 0, 2, 63, 4, 0, 0, 0, 0, 73, 37, 0, 0, 
    3, 9, 40, 35, 0, 25, 11, 1, 0, 0, 0, 13, 52, 0, 0, 
    
    -- channel=294
    230, 222, 232, 183, 188, 180, 189, 203, 233, 245, 235, 240, 219, 199, 192, 
    261, 259, 257, 182, 178, 187, 177, 201, 230, 228, 222, 236, 244, 216, 219, 
    268, 268, 254, 152, 132, 141, 140, 139, 135, 141, 184, 242, 228, 201, 192, 
    267, 268, 231, 180, 166, 213, 206, 195, 186, 178, 175, 226, 229, 195, 167, 
    266, 264, 217, 161, 163, 173, 187, 176, 186, 188, 205, 195, 249, 238, 186, 
    253, 259, 189, 129, 109, 146, 138, 148, 149, 155, 172, 181, 238, 269, 268, 
    218, 209, 164, 135, 115, 138, 159, 118, 131, 161, 127, 142, 207, 240, 274, 
    208, 136, 139, 164, 129, 101, 82, 83, 84, 82, 72, 87, 123, 148, 240, 
    191, 113, 140, 100, 112, 120, 136, 98, 68, 78, 109, 64, 96, 146, 205, 
    214, 113, 125, 54, 84, 83, 81, 114, 172, 147, 157, 150, 172, 114, 150, 
    217, 121, 72, 68, 31, 56, 82, 64, 104, 98, 97, 113, 75, 124, 127, 
    217, 107, 90, 99, 41, 26, 72, 74, 70, 141, 137, 155, 89, 91, 115, 
    202, 138, 75, 147, 78, 18, 13, 19, 25, 142, 185, 161, 36, 47, 107, 
    193, 196, 146, 136, 95, 46, 10, 20, 54, 126, 164, 156, 23, 46, 121, 
    192, 178, 152, 88, 84, 55, 30, 37, 46, 71, 106, 123, 19, 47, 129, 
    
    -- channel=295
    6, 4, 16, 17, 12, 0, 0, 0, 0, 6, 11, 7, 17, 0, 17, 
    3, 2, 18, 31, 3, 0, 0, 0, 0, 0, 12, 4, 12, 24, 2, 
    5, 5, 21, 68, 0, 0, 0, 0, 0, 0, 0, 3, 19, 36, 0, 
    5, 15, 9, 57, 0, 0, 2, 0, 0, 0, 0, 0, 20, 24, 13, 
    6, 18, 18, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 
    1, 28, 30, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 
    4, 37, 17, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    31, 44, 0, 41, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 34, 0, 35, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    27, 47, 0, 22, 0, 5, 0, 0, 20, 0, 0, 0, 0, 9, 0, 
    13, 54, 0, 13, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    6, 60, 0, 0, 12, 0, 0, 36, 0, 14, 0, 0, 48, 0, 0, 
    0, 36, 0, 10, 15, 3, 0, 0, 0, 0, 0, 47, 8, 0, 0, 
    0, 7, 17, 10, 0, 20, 0, 0, 0, 0, 0, 53, 11, 0, 0, 
    0, 0, 10, 1, 0, 4, 0, 0, 0, 0, 0, 23, 4, 0, 0, 
    
    -- channel=296
    9, 12, 11, 0, 0, 8, 23, 38, 18, 0, 0, 0, 18, 21, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 10, 38, 30, 43, 22, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 11, 0, 0, 5, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 48, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 6, 0, 0, 0, 0, 0, 51, 103, 89, 113, 118, 87, 12, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 25, 13, 8, 0, 29, 32, 0, 22, 11, 30, 6, 12, 0, 
    0, 0, 0, 49, 38, 6, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 54, 59, 16, 19, 37, 15, 14, 4, 23, 47, 58, 7, 3, 0, 
    0, 0, 3, 9, 3, 24, 31, 24, 12, 0, 0, 6, 4, 7, 0, 
    0, 0, 14, 0, 4, 12, 27, 26, 16, 3, 0, 0, 24, 11, 0, 
    
    -- channel=297
    16, 16, 13, 18, 18, 8, 9, 6, 12, 21, 24, 24, 23, 24, 34, 
    9, 10, 14, 4, 2, 0, 0, 6, 11, 31, 36, 22, 23, 38, 36, 
    9, 9, 11, 5, 0, 0, 0, 0, 0, 0, 19, 13, 20, 41, 43, 
    9, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 23, 23, 26, 28, 
    10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 6, 
    10, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 9, 
    3, 12, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 16, 
    4, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 
    0, 2, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 2, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 3, 4, 4, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 8, 7, 0, 0, 6, 5, 25, 0, 14, 0, 0, 20, 6, 0, 
    0, 0, 0, 0, 0, 7, 14, 10, 5, 0, 0, 0, 6, 4, 0, 
    0, 0, 0, 0, 0, 10, 12, 7, 0, 0, 1, 13, 13, 0, 0, 
    0, 0, 0, 0, 0, 6, 6, 4, 0, 0, 0, 7, 7, 1, 0, 
    
    -- channel=298
    165, 158, 164, 93, 123, 128, 152, 172, 176, 169, 152, 165, 160, 142, 132, 
    180, 180, 169, 47, 59, 66, 39, 50, 90, 114, 129, 161, 160, 127, 156, 
    179, 178, 161, 51, 84, 98, 91, 84, 64, 46, 123, 175, 139, 106, 114, 
    178, 175, 137, 68, 119, 149, 108, 100, 114, 116, 81, 142, 155, 136, 87, 
    178, 173, 76, 44, 98, 65, 77, 88, 95, 92, 119, 131, 175, 176, 164, 
    164, 155, 117, 37, 30, 71, 56, 53, 52, 68, 69, 83, 168, 179, 179, 
    134, 99, 70, 76, 68, 58, 73, 43, 59, 73, 37, 52, 87, 116, 185, 
    126, 14, 96, 84, 44, 39, 27, 14, 0, 0, 0, 0, 26, 48, 171, 
    122, 34, 86, 0, 69, 54, 82, 77, 105, 106, 127, 103, 110, 85, 128, 
    137, 6, 49, 0, 14, 5, 0, 29, 59, 40, 37, 40, 70, 9, 91, 
    135, 34, 27, 15, 0, 8, 67, 0, 58, 40, 46, 98, 0, 90, 68, 
    118, 0, 46, 78, 0, 0, 0, 0, 8, 58, 85, 60, 0, 6, 55, 
    116, 105, 51, 84, 27, 0, 0, 0, 0, 155, 147, 103, 0, 12, 67, 
    116, 103, 66, 68, 35, 0, 0, 0, 16, 32, 60, 60, 0, 11, 70, 
    98, 94, 80, 9, 26, 4, 0, 3, 6, 19, 33, 54, 0, 12, 98, 
    
    -- channel=299
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 48, 65, 60, 73, 106, 100, 66, 23, 0, 2, 12, 0, 
    0, 0, 2, 2, 0, 0, 0, 0, 0, 2, 0, 0, 8, 30, 16, 
    0, 1, 0, 28, 0, 0, 6, 7, 0, 0, 4, 22, 0, 0, 14, 
    0, 0, 58, 44, 0, 23, 34, 5, 7, 6, 0, 0, 0, 0, 0, 
    8, 28, 0, 17, 28, 0, 3, 31, 35, 18, 41, 19, 0, 0, 0, 
    7, 45, 34, 0, 0, 0, 14, 0, 0, 30, 28, 35, 75, 65, 7, 
    25, 61, 0, 10, 34, 0, 0, 29, 71, 58, 48, 84, 56, 22, 0, 
    0, 0, 1, 75, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 25, 48, 0, 32, 18, 34, 21, 58, 37, 58, 47, 47, 39, 0, 
    0, 0, 0, 0, 6, 3, 0, 5, 4, 0, 0, 0, 0, 0, 0, 
    9, 54, 2, 0, 0, 16, 80, 53, 24, 37, 0, 48, 57, 67, 0, 
    0, 0, 0, 13, 0, 0, 4, 0, 0, 0, 0, 0, 17, 0, 0, 
    0, 20, 1, 20, 2, 0, 0, 0, 0, 61, 44, 53, 1, 0, 0, 
    11, 0, 0, 19, 9, 0, 0, 0, 0, 0, 26, 27, 0, 0, 0, 
    
    -- channel=300
    38, 35, 44, 32, 32, 34, 32, 32, 36, 38, 34, 33, 32, 26, 23, 
    48, 46, 50, 47, 60, 67, 61, 62, 57, 39, 27, 34, 34, 25, 20, 
    51, 51, 51, 55, 86, 99, 97, 100, 99, 81, 37, 41, 36, 19, 11, 
    50, 53, 49, 74, 86, 81, 95, 111, 108, 103, 78, 37, 33, 27, 12, 
    48, 52, 58, 79, 94, 99, 99, 110, 106, 101, 100, 58, 41, 43, 31, 
    41, 51, 47, 85, 77, 93, 101, 100, 99, 99, 97, 76, 55, 50, 51, 
    42, 45, 39, 54, 83, 97, 105, 91, 89, 92, 65, 56, 54, 47, 48, 
    35, 32, 26, 47, 87, 80, 79, 75, 66, 64, 66, 62, 64, 76, 58, 
    39, 36, 34, 41, 68, 56, 61, 60, 47, 44, 54, 44, 59, 75, 55, 
    45, 47, 42, 34, 59, 59, 61, 57, 72, 76, 78, 75, 77, 65, 56, 
    48, 46, 43, 45, 43, 45, 57, 65, 57, 71, 70, 66, 65, 64, 54, 
    65, 54, 39, 54, 45, 37, 48, 44, 40, 43, 58, 61, 39, 58, 43, 
    77, 64, 54, 67, 53, 39, 31, 33, 35, 44, 54, 64, 40, 36, 53, 
    75, 77, 72, 63, 59, 44, 28, 32, 36, 56, 63, 73, 32, 39, 60, 
    83, 82, 76, 58, 56, 45, 35, 38, 43, 51, 60, 65, 35, 40, 60, 
    
    -- channel=301
    64, 67, 57, 35, 36, 55, 69, 91, 80, 58, 55, 51, 64, 68, 56, 
    66, 67, 57, 19, 13, 12, 9, 0, 1, 12, 31, 51, 46, 36, 47, 
    61, 61, 46, 39, 55, 80, 81, 80, 63, 47, 36, 57, 44, 21, 31, 
    61, 56, 48, 26, 72, 70, 75, 63, 72, 82, 66, 27, 43, 52, 34, 
    58, 56, 23, 13, 57, 53, 36, 62, 62, 65, 59, 61, 62, 58, 84, 
    43, 41, 46, 42, 29, 46, 54, 41, 35, 47, 35, 37, 55, 61, 61, 
    41, 9, 13, 34, 79, 61, 43, 49, 53, 42, 32, 31, 17, 15, 52, 
    19, 0, 21, 35, 27, 32, 36, 25, 0, 0, 10, 0, 5, 28, 44, 
    45, 26, 35, 0, 38, 40, 48, 55, 100, 113, 92, 102, 109, 63, 51, 
    41, 17, 0, 15, 14, 14, 13, 21, 17, 21, 9, 11, 12, 14, 50, 
    42, 20, 37, 16, 16, 14, 55, 37, 15, 40, 34, 54, 32, 50, 62, 
    42, 0, 3, 61, 30, 13, 0, 0, 26, 12, 41, 31, 0, 0, 40, 
    45, 63, 76, 32, 26, 22, 8, 11, 23, 76, 81, 46, 12, 21, 69, 
    58, 40, 36, 21, 28, 15, 19, 25, 29, 17, 10, 6, 3, 32, 58, 
    47, 48, 44, 18, 22, 14, 25, 26, 26, 26, 21, 3, 19, 26, 77, 
    
    -- channel=302
    26, 21, 45, 50, 15, 2, 0, 0, 9, 34, 38, 25, 25, 13, 16, 
    40, 38, 70, 93, 65, 53, 55, 78, 68, 33, 32, 27, 39, 53, 0, 
    49, 49, 68, 117, 0, 18, 4, 26, 38, 37, 0, 25, 60, 59, 0, 
    48, 66, 48, 135, 0, 0, 77, 51, 34, 7, 42, 14, 32, 42, 20, 
    45, 69, 96, 102, 11, 40, 70, 38, 39, 34, 51, 0, 16, 44, 0, 
    30, 88, 37, 104, 3, 22, 50, 45, 46, 38, 45, 12, 0, 49, 48, 
    38, 89, 48, 33, 0, 32, 50, 25, 7, 35, 27, 2, 38, 35, 40, 
    54, 87, 0, 74, 49, 32, 23, 46, 29, 15, 33, 25, 0, 20, 0, 
    40, 45, 0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    52, 98, 15, 16, 4, 29, 17, 0, 78, 49, 73, 57, 55, 58, 0, 
    45, 83, 7, 12, 0, 0, 0, 55, 0, 39, 22, 0, 41, 0, 0, 
    61, 124, 0, 0, 22, 0, 9, 37, 0, 15, 8, 43, 57, 36, 0, 
    43, 31, 0, 51, 17, 8, 0, 0, 0, 0, 4, 86, 18, 0, 0, 
    32, 69, 60, 48, 14, 23, 0, 0, 0, 21, 31, 129, 0, 0, 0, 
    55, 42, 61, 41, 12, 3, 0, 0, 0, 0, 9, 56, 0, 0, 0, 
    
    -- channel=303
    58, 57, 57, 39, 40, 52, 61, 68, 60, 53, 46, 48, 61, 42, 46, 
    67, 67, 59, 45, 41, 44, 36, 29, 29, 32, 28, 44, 47, 31, 32, 
    66, 65, 63, 70, 81, 96, 105, 102, 84, 56, 37, 51, 43, 23, 12, 
    66, 63, 62, 76, 77, 95, 102, 100, 105, 106, 68, 29, 53, 41, 19, 
    64, 63, 52, 73, 77, 78, 87, 96, 92, 97, 94, 55, 63, 69, 69, 
    55, 55, 75, 79, 50, 83, 82, 77, 74, 78, 66, 60, 56, 67, 66, 
    48, 41, 35, 68, 96, 85, 91, 79, 77, 75, 57, 41, 29, 37, 62, 
    39, 27, 35, 54, 71, 69, 57, 44, 28, 32, 30, 20, 37, 54, 53, 
    55, 52, 27, 23, 60, 46, 73, 81, 81, 87, 93, 81, 82, 73, 54, 
    62, 45, 12, 40, 27, 43, 31, 37, 57, 48, 49, 47, 46, 50, 52, 
    59, 59, 33, 37, 24, 28, 69, 42, 43, 56, 55, 69, 43, 67, 58, 
    68, 44, 23, 63, 40, 16, 2, 24, 8, 44, 57, 30, 39, 13, 47, 
    77, 98, 61, 49, 53, 24, 12, 15, 24, 58, 79, 66, 25, 30, 58, 
    76, 71, 67, 43, 46, 34, 17, 20, 29, 21, 43, 47, 21, 27, 62, 
    77, 79, 70, 39, 38, 32, 26, 28, 30, 35, 37, 41, 26, 28, 69, 
    
    -- channel=304
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 3, 23, 3, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 28, 123, 119, 52, 112, 71, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 
    0, 0, 0, 0, 0, 1, 74, 0, 26, 0, 0, 65, 0, 26, 27, 
    0, 0, 6, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 
    0, 22, 9, 0, 0, 0, 0, 0, 28, 101, 0, 0, 0, 32, 71, 
    0, 0, 0, 0, 0, 0, 14, 16, 7, 0, 0, 0, 0, 23, 53, 
    0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 20, 91, 
    
    -- channel=305
    8, 18, 12, 14, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 
    2, 4, 0, 3, 9, 10, 22, 16, 0, 0, 7, 5, 5, 7, 0, 
    9, 8, 3, 32, 22, 26, 24, 36, 50, 52, 7, 5, 10, 7, 11, 
    10, 11, 20, 11, 0, 0, 0, 2, 0, 0, 27, 8, 8, 0, 9, 
    6, 5, 18, 9, 0, 11, 5, 0, 0, 3, 0, 0, 0, 16, 16, 
    4, 0, 0, 10, 19, 18, 13, 0, 8, 12, 0, 20, 11, 8, 10, 
    18, 14, 18, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 0, 0, 
    0, 30, 0, 0, 19, 50, 49, 7, 0, 1, 0, 0, 10, 34, 6, 
    1, 0, 1, 29, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 
    8, 16, 0, 8, 6, 21, 41, 0, 33, 45, 38, 43, 12, 32, 15, 
    10, 0, 8, 7, 18, 2, 9, 24, 29, 44, 36, 41, 36, 0, 13, 
    12, 25, 0, 0, 5, 12, 9, 0, 0, 0, 0, 0, 3, 26, 15, 
    8, 1, 16, 0, 3, 5, 0, 0, 8, 0, 0, 0, 0, 0, 19, 
    6, 6, 3, 0, 0, 0, 1, 0, 0, 31, 25, 7, 3, 2, 13, 
    11, 10, 8, 13, 0, 0, 6, 7, 10, 11, 11, 0, 8, 11, 15, 
    
    -- channel=306
    41, 43, 39, 30, 17, 18, 18, 24, 46, 51, 51, 52, 31, 38, 26, 
    58, 58, 51, 20, 15, 18, 32, 43, 47, 50, 47, 53, 55, 42, 45, 
    64, 65, 48, 0, 0, 0, 0, 0, 0, 14, 34, 50, 49, 31, 49, 
    64, 60, 53, 0, 9, 26, 23, 17, 9, 10, 31, 53, 41, 19, 31, 
    64, 56, 43, 0, 5, 29, 14, 14, 19, 28, 13, 35, 52, 29, 17, 
    63, 51, 18, 0, 5, 0, 2, 7, 8, 17, 27, 39, 59, 65, 64, 
    53, 37, 29, 0, 0, 3, 0, 0, 0, 0, 0, 14, 49, 64, 64, 
    33, 16, 9, 0, 5, 0, 0, 0, 0, 0, 0, 0, 7, 23, 56, 
    20, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 61, 
    31, 0, 0, 0, 0, 0, 0, 11, 15, 19, 17, 14, 10, 1, 46, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    33, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 15, 0, 0, 30, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 21, 
    24, 23, 0, 0, 0, 0, 0, 0, 0, 20, 25, 0, 0, 0, 21, 
    24, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=307
    6, 11, 4, 0, 0, 0, 7, 13, 16, 11, 13, 9, 10, 16, 15, 
    4, 5, 2, 0, 0, 0, 0, 0, 0, 11, 11, 8, 7, 16, 18, 
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 15, 6, 5, 12, 18, 
    2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 8, 10, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=308
    2, 0, 13, 52, 0, 0, 0, 0, 0, 0, 4, 0, 26, 0, 23, 
    0, 0, 31, 112, 2, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 
    0, 0, 39, 178, 0, 0, 0, 27, 9, 0, 0, 0, 26, 47, 0, 
    0, 11, 15, 180, 0, 0, 58, 2, 4, 0, 0, 0, 7, 49, 0, 
    0, 21, 72, 115, 0, 0, 30, 0, 0, 0, 21, 0, 0, 41, 0, 
    0, 42, 54, 144, 0, 0, 20, 3, 1, 0, 0, 0, 0, 0, 0, 
    0, 62, 11, 64, 0, 0, 32, 16, 0, 3, 23, 0, 0, 0, 0, 
    13, 95, 0, 82, 17, 28, 13, 40, 6, 0, 20, 0, 0, 0, 0, 
    33, 113, 0, 102, 0, 0, 0, 46, 0, 0, 59, 11, 0, 8, 0, 
    35, 165, 0, 73, 0, 27, 0, 0, 24, 0, 17, 0, 0, 53, 0, 
    6, 177, 5, 34, 22, 0, 0, 86, 0, 40, 8, 0, 67, 0, 0, 
    14, 199, 0, 4, 91, 0, 0, 74, 0, 0, 0, 0, 107, 0, 0, 
    0, 115, 0, 13, 66, 63, 5, 0, 0, 0, 16, 127, 69, 0, 0, 
    0, 33, 70, 29, 14, 85, 4, 0, 0, 0, 0, 134, 53, 0, 0, 
    11, 15, 62, 56, 7, 41, 8, 0, 0, 0, 0, 60, 58, 0, 0, 
    
    -- channel=309
    0, 9, 0, 0, 0, 11, 14, 36, 30, 0, 0, 6, 0, 9, 0, 
    0, 1, 0, 0, 0, 12, 18, 0, 9, 12, 0, 21, 0, 0, 29, 
    0, 0, 0, 0, 34, 14, 19, 0, 3, 27, 81, 13, 0, 0, 52, 
    0, 0, 0, 0, 95, 30, 0, 0, 0, 17, 16, 54, 0, 0, 8, 
    2, 0, 0, 0, 54, 34, 0, 11, 14, 24, 0, 77, 30, 0, 12, 
    29, 0, 0, 0, 48, 14, 0, 2, 0, 19, 10, 43, 77, 0, 0, 
    25, 0, 0, 0, 39, 17, 0, 0, 30, 0, 0, 58, 52, 37, 15, 
    0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 11, 55, 57, 98, 
    0, 0, 64, 0, 38, 27, 7, 0, 32, 63, 0, 14, 78, 15, 126, 
    0, 0, 15, 0, 37, 0, 29, 85, 0, 20, 0, 0, 0, 0, 172, 
    0, 0, 3, 0, 0, 33, 50, 0, 58, 0, 0, 42, 0, 29, 144, 
    0, 0, 38, 2, 0, 24, 55, 0, 125, 0, 3, 24, 0, 10, 178, 
    0, 0, 41, 0, 0, 0, 4, 18, 47, 137, 0, 0, 0, 41, 180, 
    16, 0, 0, 0, 0, 0, 8, 27, 50, 63, 24, 0, 0, 78, 145, 
    0, 0, 0, 0, 0, 0, 5, 12, 22, 27, 37, 0, 0, 57, 168, 
    
    -- channel=310
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 42, 28, 0, 44, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 15, 15, 13, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 26, 20, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 12, 10, 0, 0, 0, 0, 4, 6, 0, 
    
    -- channel=311
    0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 0, 0, 12, 0, 12, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 7, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 0, 
    0, 0, 5, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 3, 
    0, 5, 23, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 28, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 43, 0, 24, 0, 0, 0, 24, 0, 0, 37, 9, 0, 0, 0, 
    13, 48, 0, 32, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 68, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 63, 0, 1, 28, 0, 0, 44, 0, 14, 0, 0, 51, 0, 0, 
    0, 56, 0, 0, 30, 18, 7, 0, 0, 0, 7, 53, 18, 0, 0, 
    0, 0, 13, 8, 0, 36, 7, 0, 0, 0, 0, 44, 27, 0, 0, 
    0, 0, 9, 5, 0, 19, 5, 0, 0, 0, 0, 24, 19, 0, 0, 
    
    -- channel=312
    4, 1, 0, 1, 18, 9, 5, 0, 19, 28, 23, 38, 0, 5, 0, 
    24, 24, 9, 0, 54, 76, 93, 112, 121, 106, 55, 42, 37, 13, 45, 
    34, 35, 14, 0, 11, 0, 0, 0, 0, 32, 98, 29, 12, 11, 84, 
    33, 22, 24, 0, 75, 56, 0, 33, 11, 18, 16, 98, 16, 0, 23, 
    41, 17, 30, 0, 52, 57, 31, 37, 44, 45, 11, 79, 40, 0, 0, 
    70, 20, 0, 0, 73, 26, 8, 39, 42, 40, 71, 78, 90, 33, 34, 
    45, 17, 33, 0, 0, 18, 8, 6, 32, 39, 23, 80, 124, 131, 59, 
    24, 0, 61, 0, 13, 0, 0, 0, 51, 52, 24, 69, 99, 70, 127, 
    0, 0, 36, 12, 25, 39, 9, 0, 0, 0, 0, 0, 0, 6, 141, 
    0, 0, 63, 0, 50, 0, 40, 99, 24, 57, 47, 49, 59, 9, 134, 
    17, 0, 0, 0, 0, 36, 0, 0, 60, 0, 0, 0, 0, 0, 99, 
    23, 0, 55, 0, 0, 1, 91, 0, 105, 38, 1, 56, 0, 56, 135, 
    29, 0, 0, 0, 0, 0, 0, 0, 13, 59, 0, 0, 0, 15, 89, 
    22, 13, 0, 0, 0, 0, 0, 0, 12, 87, 83, 0, 0, 29, 93, 
    25, 9, 0, 0, 1, 0, 0, 0, 0, 12, 45, 0, 0, 16, 81, 
    
    -- channel=313
    0, 7, 0, 0, 0, 6, 11, 16, 0, 0, 0, 0, 2, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 20, 
    0, 0, 0, 0, 37, 15, 22, 7, 0, 0, 44, 0, 0, 0, 20, 
    0, 0, 0, 0, 23, 0, 0, 0, 0, 3, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 18, 4, 0, 39, 
    0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 6, 34, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 56, 0, 0, 1, 4, 0, 0, 0, 0, 0, 16, 9, 37, 
    0, 0, 3, 0, 23, 0, 4, 11, 68, 72, 10, 56, 53, 0, 32, 
    0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 83, 
    0, 0, 0, 0, 0, 26, 58, 0, 54, 0, 9, 59, 0, 34, 52, 
    0, 0, 30, 18, 0, 1, 0, 0, 21, 0, 0, 0, 0, 0, 108, 
    0, 2, 10, 0, 0, 0, 8, 17, 41, 82, 0, 0, 0, 43, 84, 
    0, 0, 0, 0, 0, 0, 21, 25, 20, 0, 6, 0, 0, 42, 74, 
    0, 0, 0, 0, 0, 0, 16, 17, 17, 10, 0, 0, 0, 38, 99, 
    
    -- channel=314
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=315
    38, 35, 42, 25, 32, 35, 40, 36, 54, 52, 44, 50, 26, 27, 12, 
    63, 62, 61, 37, 51, 59, 57, 71, 80, 60, 40, 49, 53, 27, 32, 
    66, 66, 64, 0, 25, 29, 24, 19, 30, 29, 42, 59, 45, 21, 31, 
    65, 65, 48, 24, 60, 82, 60, 60, 53, 55, 47, 58, 41, 21, 25, 
    67, 63, 63, 20, 60, 59, 52, 59, 63, 58, 57, 67, 65, 40, 11, 
    70, 68, 22, 11, 37, 36, 35, 48, 48, 40, 61, 56, 64, 66, 66, 
    61, 55, 38, 3, 28, 47, 53, 32, 44, 67, 27, 40, 74, 80, 70, 
    66, 16, 24, 32, 28, 0, 0, 0, 18, 16, 0, 22, 41, 44, 83, 
    39, 0, 35, 9, 14, 34, 31, 8, 0, 0, 0, 0, 0, 46, 91, 
    44, 0, 40, 0, 29, 0, 11, 28, 48, 35, 40, 36, 56, 10, 51, 
    53, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 1, 4, 7, 51, 
    62, 0, 18, 0, 0, 0, 13, 0, 27, 27, 31, 55, 0, 27, 22, 
    61, 0, 0, 35, 0, 0, 0, 0, 0, 32, 49, 22, 0, 0, 34, 
    52, 57, 18, 33, 7, 0, 0, 0, 0, 53, 42, 18, 0, 0, 38, 
    56, 45, 24, 11, 3, 0, 0, 0, 0, 0, 25, 21, 0, 0, 28, 
    
    -- channel=316
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 46, 60, 82, 85, 55, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 27, 
    0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 
    0, 0, 3, 0, 19, 24, 13, 6, 9, 4, 0, 11, 0, 0, 0, 
    17, 0, 0, 0, 51, 2, 0, 27, 29, 23, 51, 34, 26, 0, 0, 
    8, 5, 22, 0, 0, 0, 0, 0, 9, 20, 4, 42, 76, 75, 1, 
    8, 5, 27, 0, 15, 0, 0, 14, 67, 58, 43, 82, 76, 42, 57, 
    0, 0, 14, 25, 11, 21, 0, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 56, 0, 42, 0, 34, 71, 10, 38, 37, 35, 46, 7, 64, 
    0, 0, 0, 0, 0, 27, 0, 0, 41, 0, 0, 0, 0, 0, 31, 
    0, 0, 38, 0, 0, 11, 93, 20, 79, 22, 0, 43, 0, 61, 67, 
    0, 0, 0, 0, 0, 0, 0, 3, 5, 1, 0, 0, 0, 3, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 63, 57, 0, 0, 14, 34, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 7, 36, 3, 0, 7, 15, 
    
    -- channel=317
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 38, 39, 45, 53, 40, 8, 0, 0, 0, 0, 0, 
    0, 0, 7, 55, 20, 12, 10, 10, 22, 14, 0, 0, 0, 5, 0, 
    0, 0, 5, 70, 5, 6, 31, 39, 29, 9, 0, 1, 0, 0, 0, 
    0, 0, 42, 78, 22, 33, 60, 38, 32, 27, 23, 0, 0, 0, 0, 
    0, 18, 24, 58, 45, 44, 48, 53, 56, 43, 49, 12, 0, 0, 0, 
    7, 48, 42, 46, 0, 36, 50, 41, 29, 34, 37, 21, 26, 25, 0, 
    31, 66, 8, 39, 60, 58, 59, 65, 72, 69, 63, 62, 46, 33, 0, 
    6, 34, 0, 87, 21, 25, 12, 6, 0, 0, 0, 0, 0, 15, 0, 
    15, 59, 39, 40, 39, 47, 47, 35, 48, 51, 62, 55, 54, 61, 0, 
    13, 57, 14, 37, 40, 36, 0, 45, 32, 45, 41, 9, 56, 11, 0, 
    24, 83, 30, 0, 31, 31, 52, 74, 7, 32, 12, 27, 67, 55, 0, 
    29, 17, 0, 35, 35, 30, 27, 24, 16, 0, 0, 28, 43, 17, 0, 
    18, 40, 42, 44, 33, 40, 17, 12, 8, 25, 47, 72, 42, 9, 0, 
    35, 29, 36, 49, 34, 35, 17, 18, 21, 29, 38, 61, 31, 14, 0, 
    
    -- channel=318
    56, 60, 52, 2, 20, 34, 48, 74, 63, 43, 37, 45, 53, 48, 37, 
    57, 59, 37, 0, 0, 0, 0, 0, 0, 0, 12, 48, 37, 10, 45, 
    54, 54, 27, 0, 46, 67, 64, 56, 37, 15, 35, 56, 24, 0, 18, 
    55, 45, 38, 0, 57, 37, 21, 29, 45, 54, 25, 29, 41, 27, 0, 
    54, 44, 0, 0, 34, 15, 0, 28, 28, 30, 32, 48, 55, 55, 91, 
    44, 16, 28, 0, 0, 24, 14, 0, 0, 25, 1, 27, 74, 55, 55, 
    37, 0, 0, 15, 37, 15, 0, 3, 8, 0, 0, 0, 0, 0, 53, 
    2, 0, 32, 0, 0, 20, 17, 0, 0, 0, 0, 0, 0, 8, 65, 
    27, 0, 24, 0, 28, 0, 14, 29, 98, 100, 66, 91, 101, 23, 45, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 
    30, 0, 6, 0, 0, 0, 49, 0, 25, 21, 24, 76, 0, 44, 49, 
    18, 0, 0, 41, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 51, 
    31, 47, 38, 3, 0, 0, 0, 0, 0, 87, 44, 0, 0, 0, 64, 
    40, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 54, 
    18, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 
    
    -- channel=319
    17, 15, 23, 17, 17, 17, 18, 25, 28, 24, 21, 14, 11, 16, 2, 
    28, 27, 36, 38, 47, 49, 47, 50, 50, 29, 10, 18, 18, 15, 5, 
    29, 30, 30, 34, 37, 52, 49, 51, 51, 46, 20, 17, 24, 9, 2, 
    29, 33, 22, 49, 65, 58, 69, 74, 70, 63, 52, 22, 7, 18, 5, 
    27, 33, 46, 49, 62, 68, 66, 72, 72, 67, 63, 38, 23, 12, 3, 
    22, 40, 24, 55, 39, 51, 67, 68, 61, 60, 65, 35, 28, 29, 29, 
    21, 25, 18, 20, 53, 70, 72, 60, 66, 77, 47, 42, 40, 33, 27, 
    24, 13, 0, 44, 50, 26, 33, 49, 44, 32, 45, 45, 26, 42, 31, 
    19, 18, 21, 15, 34, 47, 34, 13, 13, 14, 23, 8, 30, 57, 25, 
    21, 33, 24, 12, 34, 29, 30, 40, 36, 43, 45, 38, 55, 31, 19, 
    24, 26, 18, 19, 21, 13, 13, 48, 5, 29, 25, 11, 34, 31, 23, 
    42, 38, 11, 25, 24, 21, 33, 14, 35, 25, 33, 61, 17, 31, 6, 
    41, 22, 34, 44, 22, 21, 11, 10, 5, 28, 42, 54, 21, 5, 24, 
    50, 47, 42, 44, 33, 21, 6, 11, 23, 31, 30, 49, 9, 16, 24, 
    50, 47, 47, 32, 31, 19, 11, 14, 17, 24, 34, 32, 13, 12, 22, 
    
    
    others => 0);
end gold_package;
