LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 7, 53, 0, 0, 0, 0, 
		0, 0, 0, 13, 0, 0, 0, 
		35, 40, 35, 44, 72, 0, 8, 
		6, 0, 26, 0, 14, 14, 33, 
		0, 24, 7, 70, 0, 0, 0, 
		0, 81, 21, 0, 0, 22, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 99, 43, 19, 59, 
		17, 2, 0, 0, 29, 0, 25, 
		68, 0, 34, 0, 0, 37, 1, 
		0, 39, 66, 23, 18, 0, 0, 
		0, 0, 0, 0, 83, 24, 33, 
		86, 7, 198, 68, 0, 23, 0, 
		0, 116, 0, 0, 0, 13, 0, 
		
		59, 0, 53, 182, 180, 157, 132, 
		95, 142, 134, 18, 0, 0, 42, 
		0, 0, 0, 0, 0, 0, 8, 
		11, 95, 0, 0, 0, 0, 0, 
		0, 0, 29, 11, 66, 106, 139, 
		124, 0, 50, 145, 142, 126, 163, 
		163, 127, 114, 119, 114, 135, 126, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 35, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 33, 
		0, 0, 0, 0, 0, 0, 24, 
		0, 0, 0, 0, 0, 86, 20, 
		0, 0, 0, 106, 0, 0, 5, 
		0, 0, 0, 8, 0, 0, 0, 
		0, 226, 0, 0, 0, 0, 0, 
		
		50, 79, 18, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 43, 0, 
		80, 49, 76, 68, 0, 44, 0, 
		0, 0, 9, 92, 31, 55, 29, 
		79, 0, 0, 0, 0, 0, 0, 
		0, 20, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		128, 143, 117, 89, 33, 0, 52, 
		31, 118, 102, 15, 8, 22, 0, 
		13, 160, 127, 44, 31, 17, 0, 
		3, 42, 53, 38, 62, 24, 9, 
		21, 11, 54, 0, 0, 0, 0, 
		0, 43, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 24, 0, 
		0, 0, 0, 43, 0, 39, 31, 
		99, 0, 0, 115, 0, 104, 88, 
		188, 29, 0, 13, 0, 89, 0, 
		49, 0, 0, 89, 29, 10, 2, 
		0, 0, 48, 0, 24, 0, 0, 
		10, 16, 0, 0, 0, 0, 0, 
		
		71, 91, 80, 47, 43, 68, 47, 
		63, 109, 70, 48, 6, 34, 17, 
		52, 0, 0, 98, 0, 40, 16, 
		66, 68, 0, 0, 0, 0, 8, 
		0, 30, 0, 58, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		71, 61, 74, 71, 0, 0, 30, 
		0, 6, 0, 0, 6, 0, 0, 
		0, 94, 88, 0, 0, 0, 0, 
		0, 0, 102, 42, 66, 51, 29, 
		0, 0, 0, 0, 23, 0, 15, 
		49, 53, 86, 18, 0, 0, 0, 
		0, 69, 26, 0, 0, 0, 0, 
		
		0, 12, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 19, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		1, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		2, 0, 0, 7, 0, 9, 0, 
		46, 0, 0, 0, 0, 0, 0, 
		104, 0, 89, 145, 103, 79, 107, 
		62, 199, 108, 107, 107, 131, 122, 
		
		0, 0, 0, 6, 0, 7, 0, 
		194, 12, 0, 66, 9, 43, 74, 
		8, 126, 0, 52, 175, 98, 0, 
		0, 16, 0, 79, 49, 55, 0, 
		0, 261, 144, 0, 0, 42, 0, 
		0, 25, 267, 0, 73, 0, 0, 
		56, 0, 105, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 4, 0, 
		37, 0, 0, 35, 0, 0, 45, 
		0, 0, 0, 38, 0, 38, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 14, 96, 0, 14, 0, 0, 
		0, 0, 59, 0, 0, 0, 0, 
		64, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 138, 0, 0, 
		0, 38, 17, 0, 16, 0, 0, 
		0, 54, 14, 0, 59, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 35, 0, 47, 0, 61, 0, 
		0, 71, 0, 0, 95, 24, 0, 
		0, 0, 63, 0, 24, 0, 31, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 13, 23, 5, 0, 
		0, 0, 0, 0, 20, 15, 43, 
		12, 0, 0, 0, 0, 3, 0, 
		50, 65, 19, 22, 64, 88, 38, 
		119, 71, 210, 181, 219, 252, 243, 
		252, 142, 243, 222, 250, 273, 276, 
		
		0, 0, 9, 0, 22, 0, 13, 
		0, 46, 0, 0, 147, 0, 0, 
		0, 0, 20, 0, 135, 0, 0, 
		0, 0, 175, 0, 31, 0, 40, 
		30, 37, 0, 0, 0, 0, 57, 
		86, 98, 0, 19, 0, 7, 0, 
		0, 25, 0, 0, 8, 5, 19, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		74, 0, 0, 0, 7, 0, 0, 
		51, 0, 0, 0, 0, 0, 1, 
		45, 63, 0, 12, 0, 0, 0, 
		40, 0, 38, 4, 53, 89, 87, 
		87, 23, 74, 77, 91, 94, 106, 
		
		0, 0, 0, 0, 48, 62, 0, 
		90, 31, 120, 0, 0, 36, 11, 
		0, 22, 0, 14, 0, 0, 0, 
		35, 8, 0, 27, 3, 0, 0, 
		0, 83, 137, 0, 0, 49, 0, 
		0, 0, 0, 84, 0, 0, 7, 
		20, 0, 0, 9, 9, 11, 36, 
		
		200, 217, 142, 132, 80, 21, 129, 
		15, 139, 56, 18, 4, 13, 19, 
		0, 92, 0, 0, 0, 0, 0, 
		0, 48, 56, 21, 21, 3, 13, 
		0, 0, 0, 0, 0, 0, 30, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		39, 34, 11, 53, 7, 0, 24, 
		0, 4, 0, 0, 0, 0, 0, 
		0, 53, 28, 0, 0, 3, 0, 
		0, 14, 0, 61, 0, 11, 0, 
		0, 0, 0, 0, 0, 51, 0, 
		28, 0, 116, 88, 0, 0, 0, 
		0, 99, 8, 0, 0, 0, 0, 
		
		10, 0, 18, 0, 28, 0, 30, 
		162, 33, 21, 0, 113, 0, 0, 
		50, 1, 36, 0, 195, 0, 0, 
		0, 0, 47, 2, 98, 0, 19, 
		9, 180, 0, 0, 0, 0, 0, 
		0, 90, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		98, 110, 105, 105, 77, 61, 79, 
		86, 97, 99, 50, 14, 14, 36, 
		17, 82, 31, 26, 0, 22, 15, 
		0, 72, 22, 17, 2, 0, 17, 
		0, 0, 20, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 17, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		27, 0, 125, 46, 65, 39, 37, 
		141, 40, 124, 98, 77, 101, 78, 
		
		0, 0, 0, 0, 0, 61, 0, 
		103, 33, 99, 48, 0, 0, 0, 
		0, 0, 0, 30, 33, 0, 0, 
		49, 51, 0, 0, 0, 0, 0, 
		0, 86, 114, 67, 22, 0, 14, 
		0, 0, 0, 0, 0, 38, 41, 
		4, 0, 0, 0, 0, 0, 2, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 1, 
		
		0, 0, 0, 0, 18, 57, 23, 
		38, 26, 46, 69, 32, 36, 58, 
		60, 0, 16, 44, 0, 42, 42, 
		32, 46, 0, 0, 24, 10, 39, 
		0, 25, 65, 39, 43, 0, 18, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 7, 9, 16, 30, 0, 0, 
		0, 48, 0, 0, 0, 0, 0, 
		0, 27, 0, 0, 28, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 61, 21, 
		15, 0, 0, 28, 57, 39, 38, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 11, 0, 0, 0, 0, 
		17, 0, 53, 0, 0, 0, 0, 
		77, 0, 0, 23, 0, 0, 0, 
		53, 82, 0, 35, 0, 38, 30, 
		0, 159, 7, 37, 53, 51, 83, 
		
		37, 51, 0, 32, 0, 5, 38, 
		51, 0, 0, 49, 0, 93, 41, 
		124, 12, 0, 79, 0, 100, 11, 
		34, 38, 0, 102, 29, 76, 30, 
		14, 0, 22, 0, 37, 4, 16, 
		15, 0, 56, 18, 24, 0, 1, 
		29, 46, 70, 29, 12, 34, 31, 
		
		13, 19, 31, 18, 41, 34, 9, 
		29, 38, 51, 63, 83, 80, 36, 
		79, 69, 124, 136, 88, 101, 50, 
		93, 82, 102, 90, 70, 65, 57, 
		128, 94, 61, 112, 50, 7, 25, 
		40, 125, 21, 0, 3, 11, 15, 
		0, 18, 0, 0, 0, 0, 0, 
		
		others=>0 );
END gold_package;
