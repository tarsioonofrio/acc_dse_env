library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    4309, -4548, 1922, -1687, 1872, -2230, -4892, -4908, 8348, -4973, -5603, 15533, 2609, 7923, 8185, -989, 951, -10732, -2628, -784, -8448, -3995, -1956, 6940, 1563, 12563, 5468, -3873, -5359, 9306, -3817, -11036,

    -- weights
    -- filter=0 channel=0
    -9, 3, 6, -40, -35, -2, -36, -20, 2,
    -- filter=0 channel=1
    -20, -7, -19, -18, 2, -20, 17, 20, -8,
    -- filter=0 channel=2
    23, 23, 5, -14, 19, -5, 10, -9, -15,
    -- filter=0 channel=3
    7, -17, 13, -18, -17, 31, -5, 7, 20,
    -- filter=0 channel=4
    11, -3, 14, 0, 5, -10, 14, -5, 9,
    -- filter=0 channel=5
    18, 24, 17, 13, -1, 8, 6, -7, -10,
    -- filter=0 channel=6
    34, 15, 29, 6, -3, 20, -5, 26, -5,
    -- filter=0 channel=7
    10, -5, 2, -18, -22, -15, 12, -3, -11,
    -- filter=0 channel=8
    23, 5, 27, 0, 0, 24, -6, 0, 24,
    -- filter=0 channel=9
    11, -5, 7, 23, 16, 13, 10, -4, 11,
    -- filter=0 channel=10
    6, 2, 27, 31, 29, -10, 6, 21, 13,
    -- filter=0 channel=11
    -16, 6, -13, 3, 18, -9, -3, 20, -9,
    -- filter=0 channel=12
    17, -1, 14, 0, 1, 16, -4, 6, 30,
    -- filter=0 channel=13
    0, 14, 8, -22, -13, -12, 0, 3, 6,
    -- filter=0 channel=14
    -4, -2, -14, 6, 9, -5, -14, -1, 18,
    -- filter=0 channel=15
    -6, 2, -15, -14, -11, -3, 7, 1, 10,
    -- filter=1 channel=0
    13, 2, 31, -6, 3, 23, 15, 9, 12,
    -- filter=1 channel=1
    3, -3, 18, -3, -16, -6, -11, 0, 4,
    -- filter=1 channel=2
    -10, 9, 4, -26, -21, -12, -9, -26, -17,
    -- filter=1 channel=3
    12, 13, 11, 0, -19, -16, -5, 8, 20,
    -- filter=1 channel=4
    -29, -22, -29, 4, -13, -30, -24, -6, -5,
    -- filter=1 channel=5
    -16, 23, -13, 9, -8, 0, -8, 0, -12,
    -- filter=1 channel=6
    -28, -6, 3, -5, -21, 18, -1, -6, -11,
    -- filter=1 channel=7
    0, 9, 5, -4, -3, 7, -5, 11, -6,
    -- filter=1 channel=8
    -5, -31, -8, -19, -6, -14, -10, -3, 0,
    -- filter=1 channel=9
    -2, -12, -2, 24, 24, 22, -10, 17, 24,
    -- filter=1 channel=10
    -4, 11, -25, 0, -11, -16, 11, -13, -21,
    -- filter=1 channel=11
    20, -12, -13, 13, 16, 14, 12, 19, 17,
    -- filter=1 channel=12
    -7, 11, 27, 4, -9, 24, -2, 5, 17,
    -- filter=1 channel=13
    -17, -16, 0, -12, -19, 21, 14, 19, 2,
    -- filter=1 channel=14
    -8, -14, -1, -14, 10, -8, -7, 15, 10,
    -- filter=1 channel=15
    -16, 16, 37, -6, 21, 12, 10, 5, -6,
    -- filter=2 channel=0
    3, 7, -11, -18, 8, 19, 15, -10, 0,
    -- filter=2 channel=1
    10, -16, -6, -13, -10, -9, -15, 14, -8,
    -- filter=2 channel=2
    -20, 14, -10, -14, -14, 18, 7, -19, 20,
    -- filter=2 channel=3
    3, -20, -8, 15, 10, 0, -5, -1, -21,
    -- filter=2 channel=4
    4, 8, -1, 6, -7, -10, 12, 17, 9,
    -- filter=2 channel=5
    17, 0, 0, 0, -3, -12, -20, 15, 9,
    -- filter=2 channel=6
    3, -11, -2, -6, -11, 6, 15, 0, -20,
    -- filter=2 channel=7
    11, -17, -12, 3, -7, 7, -4, 20, -20,
    -- filter=2 channel=8
    -15, -11, -20, 4, 19, 2, 9, 4, -4,
    -- filter=2 channel=9
    7, -7, 6, -14, -7, 2, -5, 14, -8,
    -- filter=2 channel=10
    -6, -4, 7, -5, -14, 1, -1, 0, -16,
    -- filter=2 channel=11
    9, -21, 6, -4, -15, -3, 4, 3, 17,
    -- filter=2 channel=12
    -6, -11, -15, -8, -5, 12, 1, 18, 3,
    -- filter=2 channel=13
    -14, -17, -5, -13, -1, 18, -16, -11, -13,
    -- filter=2 channel=14
    -14, -1, -1, -8, -16, -17, 8, -14, 10,
    -- filter=2 channel=15
    3, -15, 14, 6, -19, -15, -12, -7, 0,
    -- filter=3 channel=0
    12, 1, -14, 0, 3, 3, 7, 18, 10,
    -- filter=3 channel=1
    -16, -7, -1, 7, 14, 9, 5, -7, -21,
    -- filter=3 channel=2
    16, 20, -8, -15, -11, -5, 10, 17, 13,
    -- filter=3 channel=3
    -20, -15, 6, -1, -10, 10, -14, 0, 15,
    -- filter=3 channel=4
    -16, -16, -16, 20, -11, 16, -17, 0, 13,
    -- filter=3 channel=5
    0, 10, -12, -13, 15, 0, 5, -6, 3,
    -- filter=3 channel=6
    -1, 20, 5, -20, -20, 0, 20, -1, 18,
    -- filter=3 channel=7
    13, -3, -20, -3, -5, 7, 2, -14, 4,
    -- filter=3 channel=8
    -1, 12, 15, -12, -15, -3, 14, -15, -11,
    -- filter=3 channel=9
    15, 14, -7, 13, -13, 13, -19, 11, -18,
    -- filter=3 channel=10
    20, -20, 2, 13, -3, -20, -19, -6, -2,
    -- filter=3 channel=11
    -17, 10, 0, -8, 5, 0, -19, 9, 9,
    -- filter=3 channel=12
    19, -16, -11, 7, -8, 0, 2, -19, 14,
    -- filter=3 channel=13
    -5, -1, -6, 6, -16, -15, -12, -12, 13,
    -- filter=3 channel=14
    -1, 16, -3, 20, 0, -11, 16, -6, 13,
    -- filter=3 channel=15
    -7, 9, -9, -17, -16, -17, 15, 19, -13,
    -- filter=4 channel=0
    16, 17, 3, 26, -2, 24, 5, 27, 0,
    -- filter=4 channel=1
    0, 0, 5, -9, 14, 0, -6, -9, -14,
    -- filter=4 channel=2
    2, -14, 10, 8, 1, 8, 6, 1, 0,
    -- filter=4 channel=3
    10, -18, -25, -13, 6, 3, 4, -6, -17,
    -- filter=4 channel=4
    -12, -15, 10, -1, -1, 14, 10, 0, 16,
    -- filter=4 channel=5
    1, -4, 4, 10, 12, 20, 5, 11, -2,
    -- filter=4 channel=6
    -14, 24, 12, -14, 19, 17, -13, 24, -1,
    -- filter=4 channel=7
    16, -13, -12, 11, 16, 0, -9, 2, -7,
    -- filter=4 channel=8
    -9, -28, -2, -4, -15, -24, -20, -3, 2,
    -- filter=4 channel=9
    -15, -11, 11, 11, -6, 15, 10, -19, -16,
    -- filter=4 channel=10
    -1, -18, -12, -3, 12, -18, 4, 7, -8,
    -- filter=4 channel=11
    8, 2, -8, 20, -2, 17, 17, -20, 0,
    -- filter=4 channel=12
    5, 6, -22, 12, 9, -13, 12, -6, -6,
    -- filter=4 channel=13
    0, -2, 0, -9, -4, -3, -6, 2, 5,
    -- filter=4 channel=14
    5, 17, 6, -21, 7, -19, -20, 15, -13,
    -- filter=4 channel=15
    34, 28, 36, 15, 19, 27, 17, 0, 35,
    -- filter=5 channel=0
    6, 13, -8, -5, 22, 1, 26, -8, -6,
    -- filter=5 channel=1
    -19, 17, 4, 8, -8, -4, -10, 16, -16,
    -- filter=5 channel=2
    6, 20, 0, -17, -17, 16, 20, 19, -10,
    -- filter=5 channel=3
    -11, -15, 0, -1, 9, 7, 0, -4, -22,
    -- filter=5 channel=4
    -6, -9, -18, 14, -14, -2, -6, 15, 6,
    -- filter=5 channel=5
    -9, 9, 18, -16, -2, 11, -4, -17, -4,
    -- filter=5 channel=6
    -7, -19, 9, -13, 0, 19, -21, -12, 6,
    -- filter=5 channel=7
    -6, 10, -8, -18, -4, -13, 9, 5, -15,
    -- filter=5 channel=8
    -12, 12, 14, 9, 5, 13, 21, 5, -3,
    -- filter=5 channel=9
    14, 10, 4, -2, 19, 0, -16, 12, 6,
    -- filter=5 channel=10
    -21, -6, -17, 8, -16, -4, -6, -15, 2,
    -- filter=5 channel=11
    19, 16, -18, 5, 16, -16, -18, 16, 6,
    -- filter=5 channel=12
    22, 0, -9, 9, 0, 6, 22, -15, -9,
    -- filter=5 channel=13
    12, 7, -10, 13, 26, -17, 4, 25, 11,
    -- filter=5 channel=14
    9, -17, -6, 11, -11, 1, 9, 7, 13,
    -- filter=5 channel=15
    -8, 3, -19, 14, 0, -5, 21, -4, 7,
    -- filter=6 channel=0
    17, 18, -12, -13, -4, -2, -10, 8, -9,
    -- filter=6 channel=1
    -4, 19, -1, 5, 4, 15, -19, 12, 14,
    -- filter=6 channel=2
    -5, -15, 6, 6, 13, 14, 12, -16, 3,
    -- filter=6 channel=3
    10, -20, -12, 19, -16, -12, -14, 3, -14,
    -- filter=6 channel=4
    3, -19, -9, 17, -3, 4, 12, -17, -10,
    -- filter=6 channel=5
    12, -16, 18, -18, -17, 16, -2, 2, 7,
    -- filter=6 channel=6
    -14, -20, -18, 2, 0, -18, 1, -13, -6,
    -- filter=6 channel=7
    -4, 0, -14, -6, -6, -19, 14, -19, 9,
    -- filter=6 channel=8
    2, -2, 7, 5, -9, -4, -18, 7, -12,
    -- filter=6 channel=9
    3, -15, -19, 17, 1, 4, -6, -9, 0,
    -- filter=6 channel=10
    -8, -16, -4, 11, -20, -20, 17, 15, 0,
    -- filter=6 channel=11
    -16, 8, 12, -9, -11, 2, 16, 6, -17,
    -- filter=6 channel=12
    -12, 8, 17, -5, -18, 11, -14, -18, 20,
    -- filter=6 channel=13
    6, 19, -14, -8, -14, 16, -4, 13, 18,
    -- filter=6 channel=14
    4, -7, 11, -8, -18, -12, -19, -10, 0,
    -- filter=6 channel=15
    -3, 0, -3, -9, -8, -7, 10, -7, -13,
    -- filter=7 channel=0
    7, 15, 31, -9, -9, 32, -19, 25, 19,
    -- filter=7 channel=1
    -2, -3, -6, 20, -8, 0, 19, 8, -5,
    -- filter=7 channel=2
    12, 0, 2, -22, -23, -6, 6, -15, -25,
    -- filter=7 channel=3
    19, 29, 9, 15, 17, 32, -7, 20, 19,
    -- filter=7 channel=4
    -6, -19, 4, 9, -24, -16, -13, 9, 18,
    -- filter=7 channel=5
    -17, -18, -11, 0, 5, -4, 0, 17, 7,
    -- filter=7 channel=6
    -15, -13, -10, 13, 4, -19, 1, 20, 9,
    -- filter=7 channel=7
    -14, 11, -7, 5, 0, -11, -10, 18, 9,
    -- filter=7 channel=8
    11, 11, -9, 12, 2, -9, 2, 2, -22,
    -- filter=7 channel=9
    -12, -1, -22, 0, -4, -12, -15, -16, 18,
    -- filter=7 channel=10
    6, 4, 7, 16, -1, 1, 3, -5, -10,
    -- filter=7 channel=11
    -6, 12, 18, -17, -18, -12, -3, 2, 18,
    -- filter=7 channel=12
    24, 12, -7, 30, 11, 29, 0, -7, 19,
    -- filter=7 channel=13
    13, 6, -10, 12, 14, 33, 13, 18, 16,
    -- filter=7 channel=14
    10, 13, 20, -8, 9, -11, 10, 15, 17,
    -- filter=7 channel=15
    1, 22, 20, -6, -18, 15, -6, 16, -1,
    -- filter=8 channel=0
    1, 10, -26, -7, -17, 13, -13, 1, 14,
    -- filter=8 channel=1
    -10, 2, -9, 5, -9, 4, 19, 14, -14,
    -- filter=8 channel=2
    -19, -10, -1, 10, -14, -16, 7, 16, -1,
    -- filter=8 channel=3
    -11, 17, -23, 11, 6, -22, 22, -14, -11,
    -- filter=8 channel=4
    -16, 3, -8, -3, 15, -14, -3, -18, -7,
    -- filter=8 channel=5
    -13, 6, 5, 5, 4, 20, 18, 6, 23,
    -- filter=8 channel=6
    7, -9, 13, 16, -14, 13, 8, 20, 22,
    -- filter=8 channel=7
    -12, -8, -6, 5, 21, 6, -20, 20, -7,
    -- filter=8 channel=8
    21, -12, 19, 13, 19, 14, 10, 23, -4,
    -- filter=8 channel=9
    20, -12, 6, 14, -4, 0, -18, -2, 14,
    -- filter=8 channel=10
    -4, 22, 22, 8, -14, 9, -17, -15, 25,
    -- filter=8 channel=11
    -4, 18, -1, -1, 0, -13, -2, -9, 0,
    -- filter=8 channel=12
    -10, -12, -20, 17, -7, -18, 18, -21, -23,
    -- filter=8 channel=13
    0, 3, 5, 24, -17, -7, 0, -9, 8,
    -- filter=8 channel=14
    0, 4, 18, -1, -2, -5, 9, 11, 2,
    -- filter=8 channel=15
    9, 0, -19, -13, 19, -21, 8, -1, -22,
    -- filter=9 channel=0
    -1, 16, 20, -10, -7, -16, -9, -21, -18,
    -- filter=9 channel=1
    -7, 16, 6, 6, 10, 17, -9, 8, -5,
    -- filter=9 channel=2
    12, -13, 9, -18, 0, -3, 3, 2, -13,
    -- filter=9 channel=3
    9, 2, 7, 16, 9, 4, -21, 8, -10,
    -- filter=9 channel=4
    12, 26, 27, 24, 0, -9, 14, 29, 28,
    -- filter=9 channel=5
    -13, -6, -18, 19, 19, 15, 21, 5, 7,
    -- filter=9 channel=6
    -4, -12, 9, -3, 5, 15, 27, 25, -3,
    -- filter=9 channel=7
    12, -20, -2, -2, -9, -9, 0, -8, -20,
    -- filter=9 channel=8
    -8, 16, 15, 9, 21, -9, -3, -12, 20,
    -- filter=9 channel=9
    -19, 13, -14, -15, 5, 18, 10, -5, 21,
    -- filter=9 channel=10
    5, -4, -9, 11, -6, -3, 19, 1, 4,
    -- filter=9 channel=11
    -12, 19, -19, -17, -16, -9, 6, 4, 12,
    -- filter=9 channel=12
    -9, 18, 3, 12, -8, 2, -16, 15, -8,
    -- filter=9 channel=13
    2, -8, 1, 19, -8, -15, -15, 14, -9,
    -- filter=9 channel=14
    10, 11, -3, 20, 17, -16, 14, 14, 13,
    -- filter=9 channel=15
    -6, 11, -13, 9, 17, 5, 3, 12, -4,
    -- filter=10 channel=0
    23, -4, 10, 30, 20, -4, 16, 0, -16,
    -- filter=10 channel=1
    -2, 9, -16, 1, -11, -20, -12, -12, 17,
    -- filter=10 channel=2
    15, 19, -12, -14, -19, -10, -16, 18, 17,
    -- filter=10 channel=3
    0, -18, -24, -18, 1, -18, 13, -2, -4,
    -- filter=10 channel=4
    4, 1, -13, 23, -8, 19, 0, 16, 11,
    -- filter=10 channel=5
    -1, -15, 9, 20, -14, -7, -15, 18, -3,
    -- filter=10 channel=6
    20, -4, -4, 3, 2, 17, -16, 21, 19,
    -- filter=10 channel=7
    -15, -7, -7, 13, 11, -5, -19, 9, -4,
    -- filter=10 channel=8
    -12, -15, -2, -13, -18, 19, -9, 13, -13,
    -- filter=10 channel=9
    -21, -17, -14, 16, 0, 11, -23, -3, -16,
    -- filter=10 channel=10
    -13, -2, 18, 12, 10, 8, -1, -15, -11,
    -- filter=10 channel=11
    -1, 4, -2, -17, -20, -7, 7, -12, -16,
    -- filter=10 channel=12
    8, -12, -15, 17, -17, 7, 14, 2, -23,
    -- filter=10 channel=13
    6, 21, 8, 15, -13, 18, 14, -19, -14,
    -- filter=10 channel=14
    -8, -19, -9, 12, 2, 14, 4, -9, -3,
    -- filter=10 channel=15
    25, -9, 4, -2, 26, 6, 28, -12, 0,
    -- filter=11 channel=0
    11, 6, -14, -13, -6, -14, -6, -25, 13,
    -- filter=11 channel=1
    -6, -3, -10, -15, -21, 0, 18, 10, -16,
    -- filter=11 channel=2
    -9, 11, -15, 16, -9, -4, -10, 0, -6,
    -- filter=11 channel=3
    6, 0, 19, 16, -7, 17, -5, -13, -5,
    -- filter=11 channel=4
    5, 5, -13, 15, 9, -6, -20, 3, 2,
    -- filter=11 channel=5
    -12, 7, 16, 14, 3, -13, -10, -3, -16,
    -- filter=11 channel=6
    -13, 11, 20, -10, 21, 12, 5, 11, -7,
    -- filter=11 channel=7
    4, 21, 29, 24, 28, 25, 11, 30, 5,
    -- filter=11 channel=8
    22, 19, 6, 13, -6, 6, -6, -1, 28,
    -- filter=11 channel=9
    1, 31, 0, 11, 15, 28, -2, 14, 29,
    -- filter=11 channel=10
    10, 10, 30, 12, -4, 29, -1, -2, 29,
    -- filter=11 channel=11
    12, 15, -5, 10, 5, 1, 4, 17, 17,
    -- filter=11 channel=12
    24, -2, 28, 22, 20, 8, -4, -1, 17,
    -- filter=11 channel=13
    13, -28, -17, -23, -23, -4, -12, -18, -1,
    -- filter=11 channel=14
    15, 3, -13, 13, 1, 12, 0, 9, 17,
    -- filter=11 channel=15
    5, -35, -32, -30, 3, 7, -30, -28, 1,
    -- filter=12 channel=0
    14, -9, -11, -8, 5, -13, -5, 3, 10,
    -- filter=12 channel=1
    10, -2, 15, -10, -2, -9, 19, 16, 14,
    -- filter=12 channel=2
    -7, 12, -18, 13, -8, -6, 11, 11, 5,
    -- filter=12 channel=3
    6, 5, 11, -17, 27, 11, -16, -9, 13,
    -- filter=12 channel=4
    14, -12, 7, 25, -4, 12, 17, 18, 14,
    -- filter=12 channel=5
    17, 17, -8, 5, -1, -6, 14, -2, 0,
    -- filter=12 channel=6
    -18, 0, 11, 23, 2, 2, 24, -2, 11,
    -- filter=12 channel=7
    -16, 19, 2, 16, -14, -23, -22, -1, 11,
    -- filter=12 channel=8
    11, 8, -14, -19, 6, 7, 0, 7, 10,
    -- filter=12 channel=9
    13, -24, -22, -13, -7, -18, -9, -11, 15,
    -- filter=12 channel=10
    -7, -8, 16, 24, 20, 17, 8, 5, -14,
    -- filter=12 channel=11
    20, -5, -17, -10, -2, -18, -19, -16, 8,
    -- filter=12 channel=12
    4, 17, 24, 24, 25, 29, 6, -5, 1,
    -- filter=12 channel=13
    5, 22, 22, 8, 3, 24, -4, 17, -5,
    -- filter=12 channel=14
    -10, -20, -6, 3, -10, -2, 20, -13, -3,
    -- filter=12 channel=15
    8, -7, 18, -2, -27, -21, -7, -25, -24,
    -- filter=13 channel=0
    -3, -6, -17, -7, -25, -21, -25, -31, 0,
    -- filter=13 channel=1
    -20, -9, 16, 0, 12, 15, -19, 19, -7,
    -- filter=13 channel=2
    6, 9, 18, 22, 8, -11, 4, 10, -3,
    -- filter=13 channel=3
    1, -4, 8, 18, -5, 14, 6, 28, 15,
    -- filter=13 channel=4
    3, -28, -28, -19, -18, -8, -31, -8, -28,
    -- filter=13 channel=5
    -17, -2, -5, 11, 10, 7, 11, 4, -23,
    -- filter=13 channel=6
    -32, -23, -36, -31, -27, -38, -14, -11, -8,
    -- filter=13 channel=7
    12, 2, 9, -24, 10, 0, -23, -22, -1,
    -- filter=13 channel=8
    38, 6, 36, 36, 22, 17, 29, 30, 19,
    -- filter=13 channel=9
    -20, -22, 11, -4, -1, -5, -8, -6, -12,
    -- filter=13 channel=10
    10, 23, 0, 5, -2, 23, 4, 22, -1,
    -- filter=13 channel=11
    -13, 0, -16, 9, 20, 16, 0, 9, -18,
    -- filter=13 channel=12
    -7, 16, 21, 9, 24, 36, 24, 27, 32,
    -- filter=13 channel=13
    21, 25, 35, 15, 21, 27, -7, -1, 27,
    -- filter=13 channel=14
    -18, -13, 7, 6, -20, 20, -10, 14, -4,
    -- filter=13 channel=15
    -35, -21, -17, -23, -23, -10, -44, -46, -21,
    -- filter=14 channel=0
    -22, 22, -10, 0, -7, 22, -25, 0, 15,
    -- filter=14 channel=1
    -16, 11, -11, -11, 5, -1, -18, -17, 17,
    -- filter=14 channel=2
    -21, 0, -14, 10, -16, -18, -15, -24, 0,
    -- filter=14 channel=3
    12, 0, -9, 1, -15, -10, -4, 10, 20,
    -- filter=14 channel=4
    -1, -8, 3, -34, -20, -23, -1, 1, -21,
    -- filter=14 channel=5
    15, -1, 6, 3, 24, 12, -12, 8, -1,
    -- filter=14 channel=6
    3, 11, 21, -9, -11, 8, -1, -14, -9,
    -- filter=14 channel=7
    21, 10, 2, 2, 30, 0, 26, -4, 17,
    -- filter=14 channel=8
    -29, -20, -25, -19, -4, -5, -10, -31, -1,
    -- filter=14 channel=9
    17, -2, -12, 28, 27, 16, 8, 15, 3,
    -- filter=14 channel=10
    4, -12, 10, 2, -19, -16, 8, -21, -1,
    -- filter=14 channel=11
    19, 9, -18, 6, -12, 11, 12, -4, 13,
    -- filter=14 channel=12
    21, -5, 32, 1, 7, 25, 21, 2, 22,
    -- filter=14 channel=13
    -26, 11, 19, -25, -21, -8, -30, -3, -1,
    -- filter=14 channel=14
    1, 9, 13, 6, 9, -13, -16, -21, -10,
    -- filter=14 channel=15
    -4, 1, 12, 10, -21, 24, -2, 15, 4,
    -- filter=15 channel=0
    13, 4, -10, 11, 0, 8, -8, -12, -4,
    -- filter=15 channel=1
    15, -18, 17, 16, 1, -15, -20, -3, 3,
    -- filter=15 channel=2
    0, 17, 0, 11, 0, -12, -3, -6, 3,
    -- filter=15 channel=3
    6, 4, 6, 10, 30, -3, 10, -9, -7,
    -- filter=15 channel=4
    15, 19, 15, -11, 8, 8, -8, 14, -6,
    -- filter=15 channel=5
    -6, -22, 3, -17, 1, -2, -23, -22, 2,
    -- filter=15 channel=6
    -18, -24, -17, -7, 0, -14, -23, -5, -25,
    -- filter=15 channel=7
    -15, -22, -26, -3, -8, -4, 0, 11, -11,
    -- filter=15 channel=8
    -5, 13, -7, 19, 31, 2, 22, 20, 22,
    -- filter=15 channel=9
    0, -2, -20, 12, -23, -21, -15, -24, 15,
    -- filter=15 channel=10
    -14, -8, 15, 5, -11, 18, 12, -13, 21,
    -- filter=15 channel=11
    -20, -15, 16, -11, 15, -20, 17, -20, -16,
    -- filter=15 channel=12
    -7, -3, -5, 20, 10, -4, 23, -7, 19,
    -- filter=15 channel=13
    31, 0, 8, 23, 24, -4, 7, -6, -8,
    -- filter=15 channel=14
    15, 8, -11, -8, 0, 4, -21, -14, -12,
    -- filter=15 channel=15
    5, -4, -9, -27, -28, -22, 6, -25, 1,
    -- filter=16 channel=0
    28, 15, 2, 8, 28, 22, 24, 25, -9,
    -- filter=16 channel=1
    15, 0, 12, 7, 12, 19, -14, 18, 15,
    -- filter=16 channel=2
    -16, -1, 1, -5, 13, -14, 0, -24, -18,
    -- filter=16 channel=3
    -16, 7, 0, -11, -19, -3, 0, -4, 9,
    -- filter=16 channel=4
    -31, -1, -12, -3, 6, 9, -26, -3, -23,
    -- filter=16 channel=5
    -2, -1, -10, 0, 14, 13, -12, -3, -12,
    -- filter=16 channel=6
    2, 7, -18, 9, -17, -23, 6, -20, -21,
    -- filter=16 channel=7
    -12, 20, 1, 17, 5, 29, 10, 11, 11,
    -- filter=16 channel=8
    -13, -6, -11, 8, -20, -16, -3, -6, -10,
    -- filter=16 channel=9
    -5, 3, 13, 23, 0, -11, -1, 4, 25,
    -- filter=16 channel=10
    -17, -12, 10, 5, -12, 10, -22, 12, -4,
    -- filter=16 channel=11
    1, -2, 15, 16, 11, -14, -16, 0, 14,
    -- filter=16 channel=12
    -6, -16, 9, -12, 7, 2, 22, 19, 3,
    -- filter=16 channel=13
    -8, -4, 6, -14, 6, -26, -23, 0, -7,
    -- filter=16 channel=14
    9, 5, 21, 18, 4, 3, -16, -14, -13,
    -- filter=16 channel=15
    5, 9, 0, -16, -2, -7, -5, -22, -12,
    -- filter=17 channel=0
    -5, 16, 14, 30, 18, 22, 22, 31, 23,
    -- filter=17 channel=1
    20, -9, 14, -3, 12, -11, -4, 14, -12,
    -- filter=17 channel=2
    -17, 17, -9, -4, -15, -21, 14, 9, -21,
    -- filter=17 channel=3
    35, 28, -20, 22, 22, -5, 36, 25, -21,
    -- filter=17 channel=4
    -15, -30, -21, -21, -1, -12, -21, 11, -9,
    -- filter=17 channel=5
    -31, -23, 10, -21, -18, 9, -7, 18, 17,
    -- filter=17 channel=6
    -21, -13, -15, -22, -22, -7, -18, -11, -17,
    -- filter=17 channel=7
    -8, 2, -10, -1, 0, 11, -14, -17, -3,
    -- filter=17 channel=8
    11, 4, 12, 21, 4, -9, 27, 14, 6,
    -- filter=17 channel=9
    -14, -13, -25, 3, -18, 3, 11, 13, 8,
    -- filter=17 channel=10
    -14, 5, -14, 8, -17, 2, -3, -12, -16,
    -- filter=17 channel=11
    -16, -2, -10, -3, -2, 4, -1, 16, 16,
    -- filter=17 channel=12
    0, 1, -25, 25, 1, 0, 12, 23, -2,
    -- filter=17 channel=13
    39, 34, 21, 27, 0, -1, 27, 32, 8,
    -- filter=17 channel=14
    -3, 3, 11, 16, 3, 2, 10, -7, -17,
    -- filter=17 channel=15
    -16, 2, 34, -9, 9, 24, 6, -16, 1,
    -- filter=18 channel=0
    8, 26, 26, 17, 15, -13, 7, 29, 23,
    -- filter=18 channel=1
    -11, 0, 3, 3, 5, 15, -4, -12, 17,
    -- filter=18 channel=2
    7, 13, -6, -1, -12, 14, 11, -13, -12,
    -- filter=18 channel=3
    6, -23, -10, -18, -16, -14, 3, -24, -26,
    -- filter=18 channel=4
    8, -19, -12, -17, 5, -8, -10, -21, -25,
    -- filter=18 channel=5
    -11, 13, -17, -14, -18, 7, -10, 8, -6,
    -- filter=18 channel=6
    5, -10, 6, 12, -10, -10, -5, 11, -16,
    -- filter=18 channel=7
    14, 23, 13, 19, -4, -3, 4, -8, 14,
    -- filter=18 channel=8
    -23, -8, -18, -27, -3, -21, -12, -5, -30,
    -- filter=18 channel=9
    8, 0, -13, 24, 13, -3, -6, -7, 19,
    -- filter=18 channel=10
    0, -18, 1, -4, 8, -24, -2, 10, 4,
    -- filter=18 channel=11
    -1, -3, 12, 16, -6, 20, -9, -19, -11,
    -- filter=18 channel=12
    22, 18, -8, -3, -14, 10, 3, 17, -2,
    -- filter=18 channel=13
    7, -23, -8, -8, -13, -19, -13, -24, -25,
    -- filter=18 channel=14
    20, -2, -1, 20, 11, 20, -4, 7, -11,
    -- filter=18 channel=15
    26, 9, 19, 6, -1, 23, 20, 21, 15,
    -- filter=19 channel=0
    -10, -12, -1, 0, -8, 11, 20, 13, 10,
    -- filter=19 channel=1
    -4, 0, 0, 16, 17, 3, 6, 19, -12,
    -- filter=19 channel=2
    7, 9, 1, -10, 2, -18, 16, -7, 11,
    -- filter=19 channel=3
    -20, -15, -16, 20, 0, -20, -1, 5, 6,
    -- filter=19 channel=4
    0, 14, -8, -14, -11, -4, -9, 18, -19,
    -- filter=19 channel=5
    17, 6, -19, 4, 12, -18, 13, -7, -9,
    -- filter=19 channel=6
    8, -18, 18, 20, -11, -5, 0, -4, -20,
    -- filter=19 channel=7
    15, 15, 16, -3, -13, -21, -2, 8, -5,
    -- filter=19 channel=8
    0, -21, -2, 10, -15, 19, -10, 13, -2,
    -- filter=19 channel=9
    19, -19, 0, 2, 0, -6, 5, 19, -14,
    -- filter=19 channel=10
    11, -18, 3, 16, 20, 7, -6, -8, -18,
    -- filter=19 channel=11
    -16, -15, 3, -10, -8, -16, 4, -17, -4,
    -- filter=19 channel=12
    17, -11, -12, -12, 8, -19, -21, -20, -3,
    -- filter=19 channel=13
    -1, -5, -16, -13, -5, -14, 6, 21, -21,
    -- filter=19 channel=14
    2, 2, -6, 20, 20, 13, 13, -2, 14,
    -- filter=19 channel=15
    -12, 0, -9, -18, -11, 5, 12, -2, -6,
    -- filter=20 channel=0
    28, 31, 21, 30, 33, 33, -11, 24, 11,
    -- filter=20 channel=1
    20, -3, 9, -1, -3, -17, -1, 5, 3,
    -- filter=20 channel=2
    5, 1, -2, -32, -32, -2, -26, 0, -27,
    -- filter=20 channel=3
    37, 36, 32, 17, 20, -2, -8, -7, -3,
    -- filter=20 channel=4
    -25, -47, -25, -12, -33, -13, -13, -37, -8,
    -- filter=20 channel=5
    8, 2, -6, 12, 6, 18, 2, 10, 27,
    -- filter=20 channel=6
    -12, -23, 8, -30, -14, 13, 6, -20, -14,
    -- filter=20 channel=7
    -5, 17, -4, 18, 21, 22, 25, 32, 22,
    -- filter=20 channel=8
    -12, -2, -46, -31, -22, -10, -24, -25, -10,
    -- filter=20 channel=9
    19, 13, 20, -13, -5, 18, 5, 27, -10,
    -- filter=20 channel=10
    -3, -30, -18, -27, -10, -16, -16, 4, -28,
    -- filter=20 channel=11
    -15, -1, 14, -6, -5, -1, -5, 19, -16,
    -- filter=20 channel=12
    38, 1, 37, 24, 23, 24, 22, 22, 22,
    -- filter=20 channel=13
    -3, 16, -10, -10, -6, 19, -2, 5, -9,
    -- filter=20 channel=14
    4, 7, -8, -12, 3, 18, -9, 20, 18,
    -- filter=20 channel=15
    9, -10, -4, -34, -25, 18, -8, -2, -1,
    -- filter=21 channel=0
    17, 9, 5, 19, 30, 4, 31, -3, 26,
    -- filter=21 channel=1
    -6, 3, -18, -15, -9, 8, -16, 0, 12,
    -- filter=21 channel=2
    20, -5, 16, -20, 6, 7, 0, 19, -6,
    -- filter=21 channel=3
    0, 1, -13, 37, 15, -3, 27, 28, 20,
    -- filter=21 channel=4
    -20, -11, 4, 17, 3, -11, 20, -12, 21,
    -- filter=21 channel=5
    -13, -27, 8, 0, -22, 14, -7, -8, 14,
    -- filter=21 channel=6
    -11, -2, 15, -16, -17, -7, -4, 3, 10,
    -- filter=21 channel=7
    -12, -18, -21, 7, -28, 5, -30, -31, -11,
    -- filter=21 channel=8
    -2, -15, 10, 19, -2, -8, -12, 5, -19,
    -- filter=21 channel=9
    3, -19, -28, -30, -31, -32, -33, -6, -29,
    -- filter=21 channel=10
    8, -20, -22, 0, -12, -6, 1, -13, 6,
    -- filter=21 channel=11
    -2, -17, 19, 2, 11, 8, -7, 5, 5,
    -- filter=21 channel=12
    6, -19, -23, 10, 1, -13, 31, -12, -13,
    -- filter=21 channel=13
    13, 31, 10, 7, 43, 36, 50, 21, 36,
    -- filter=21 channel=14
    -8, 13, 19, 5, -11, 9, -17, 6, -13,
    -- filter=21 channel=15
    8, 14, 10, 0, 23, 36, 21, 32, 36,
    -- filter=22 channel=0
    24, 28, 7, 28, 4, -16, 18, -9, -32,
    -- filter=22 channel=1
    2, 2, -20, -1, 4, -14, 10, -19, 21,
    -- filter=22 channel=2
    8, -3, 2, 23, 17, 18, 28, 24, 7,
    -- filter=22 channel=3
    44, 44, 12, -3, -14, -30, -22, -44, -54,
    -- filter=22 channel=4
    51, 25, 47, 23, 51, 38, 42, 48, 42,
    -- filter=22 channel=5
    24, -8, 0, 20, 8, 21, 2, -7, 16,
    -- filter=22 channel=6
    9, 12, 16, 40, 25, 51, 38, 43, 24,
    -- filter=22 channel=7
    -18, 4, -5, -30, -30, -26, -12, -11, -9,
    -- filter=22 channel=8
    5, -18, -16, -10, -13, -8, -2, 9, 1,
    -- filter=22 channel=9
    -8, -8, 22, 27, 3, 19, 4, 21, 18,
    -- filter=22 channel=10
    12, 20, 8, 21, 17, 27, 5, 7, 14,
    -- filter=22 channel=11
    19, 8, -9, 18, -8, -5, -9, -17, -8,
    -- filter=22 channel=12
    45, 23, 5, 30, 11, 24, -4, -16, -13,
    -- filter=22 channel=13
    7, 43, 38, 23, -2, -11, -6, -29, -36,
    -- filter=22 channel=14
    -9, 2, 0, 6, -15, -5, -19, 17, 19,
    -- filter=22 channel=15
    -4, -2, -9, -15, -20, -27, 5, -15, -31,
    -- filter=23 channel=0
    11, 13, -20, -4, 2, 0, -14, 18, 0,
    -- filter=23 channel=1
    -2, -18, 10, -6, 8, 5, -16, 2, -8,
    -- filter=23 channel=2
    16, -3, -5, -15, 23, -14, 15, 3, 3,
    -- filter=23 channel=3
    9, 0, 15, 1, -19, -13, 0, -11, -17,
    -- filter=23 channel=4
    22, 9, 24, 28, 19, 30, 27, 16, -8,
    -- filter=23 channel=5
    19, 11, -7, -11, 23, 21, -4, -16, 6,
    -- filter=23 channel=6
    -4, -3, 11, 12, 18, -4, 22, -3, 25,
    -- filter=23 channel=7
    8, 9, -14, -18, 18, -13, -20, 12, 19,
    -- filter=23 channel=8
    -6, 14, -21, -23, 4, -10, -24, 17, -18,
    -- filter=23 channel=9
    -13, 6, 5, -4, 6, 16, -5, -12, 0,
    -- filter=23 channel=10
    16, -15, 19, 11, 16, 24, -6, -22, 6,
    -- filter=23 channel=11
    -8, 16, 2, 0, -9, -3, 18, 19, 13,
    -- filter=23 channel=12
    12, 6, -7, -7, -2, 17, 2, -21, -13,
    -- filter=23 channel=13
    15, 22, 23, -7, 15, 9, 17, -16, -9,
    -- filter=23 channel=14
    -5, -20, -20, 12, -20, -2, 16, -15, 17,
    -- filter=23 channel=15
    12, 16, 7, 0, -6, 0, 29, -6, 9,
    -- filter=24 channel=0
    11, 3, 0, 16, -15, 25, -8, 7, -6,
    -- filter=24 channel=1
    15, 14, 15, 11, 3, -6, 12, -15, 8,
    -- filter=24 channel=2
    -12, 0, -7, -5, -30, 0, -5, 11, -10,
    -- filter=24 channel=3
    0, 14, 3, 10, -7, 12, -11, 11, 15,
    -- filter=24 channel=4
    -26, -12, -36, -3, -19, -2, -30, -20, -15,
    -- filter=24 channel=5
    18, -17, 12, 8, 18, 22, 1, 18, -14,
    -- filter=24 channel=6
    5, 5, -19, -3, -7, 4, -14, -23, 0,
    -- filter=24 channel=7
    31, 35, 13, 33, 11, 11, 30, 14, 14,
    -- filter=24 channel=8
    -22, -22, 1, -14, -28, 5, 0, -31, 0,
    -- filter=24 channel=9
    12, 8, 21, 25, 24, 26, 26, 0, 18,
    -- filter=24 channel=10
    1, -12, -3, -15, -7, -15, -24, 3, -18,
    -- filter=24 channel=11
    15, -14, 13, 15, -17, 13, 16, 11, 13,
    -- filter=24 channel=12
    16, -6, 30, -10, 19, 0, -1, 7, -4,
    -- filter=24 channel=13
    -20, -29, -8, 5, 5, -12, -8, -13, -8,
    -- filter=24 channel=14
    10, 0, -21, -19, 19, 18, -13, 13, -1,
    -- filter=24 channel=15
    -8, 11, 12, -6, -2, 11, -19, -9, 18,
    -- filter=25 channel=0
    -8, -5, -5, 5, 0, -11, 9, -6, 16,
    -- filter=25 channel=1
    -10, -11, 1, -6, 6, 5, -6, -4, 6,
    -- filter=25 channel=2
    -10, 1, 24, 12, 26, -6, 23, 25, -6,
    -- filter=25 channel=3
    -8, 3, 0, -8, 5, 6, -1, -10, -10,
    -- filter=25 channel=4
    27, 33, 23, 1, 9, 9, 1, -4, 14,
    -- filter=25 channel=5
    33, 22, 5, 0, 26, 14, 20, 0, 18,
    -- filter=25 channel=6
    20, 33, 24, 3, 30, 32, 33, 26, 1,
    -- filter=25 channel=7
    -31, -25, -31, -10, -15, -13, -9, -1, 1,
    -- filter=25 channel=8
    -11, -19, -21, -17, -19, -14, 8, 10, 1,
    -- filter=25 channel=9
    -6, 0, 3, 12, -3, -13, -28, -28, 9,
    -- filter=25 channel=10
    21, -11, 10, 15, -1, -12, -14, -5, -25,
    -- filter=25 channel=11
    15, -16, -3, -8, 14, 0, 2, -13, 8,
    -- filter=25 channel=12
    -14, -11, 10, -27, -24, 3, 14, -15, -19,
    -- filter=25 channel=13
    13, 32, 0, 27, 11, 25, -3, 25, -2,
    -- filter=25 channel=14
    -6, -10, -2, 3, 2, -1, 0, 10, 10,
    -- filter=25 channel=15
    48, 30, 12, 58, 44, 23, 60, 40, 49,
    -- filter=26 channel=0
    8, -20, -21, 12, 13, 0, 7, -1, -22,
    -- filter=26 channel=1
    2, 7, -19, -9, -11, -4, 7, -13, 1,
    -- filter=26 channel=2
    -3, -15, -19, 9, -17, 13, 11, -5, 15,
    -- filter=26 channel=3
    7, -12, 8, 27, 29, -10, 27, -8, -25,
    -- filter=26 channel=4
    11, 12, 0, 1, 0, -9, 17, -16, -12,
    -- filter=26 channel=5
    -6, -16, 6, -17, -4, -24, -20, 7, -6,
    -- filter=26 channel=6
    -5, 0, -28, -24, -12, -22, -15, 10, -29,
    -- filter=26 channel=7
    -3, 0, 24, -6, -9, -14, 10, -22, -3,
    -- filter=26 channel=8
    36, 30, 30, 44, 37, 51, 41, 49, 31,
    -- filter=26 channel=9
    -25, -19, 20, -6, -4, -10, 16, -13, -7,
    -- filter=26 channel=10
    0, 19, 20, 18, -3, 27, -7, -12, 11,
    -- filter=26 channel=11
    1, 19, 11, 20, 20, -14, 16, 17, -15,
    -- filter=26 channel=12
    -11, -12, -3, 29, -1, -24, 27, -1, -27,
    -- filter=26 channel=13
    0, 24, 12, 2, 25, 17, 16, 21, 13,
    -- filter=26 channel=14
    13, 14, -18, 12, -18, -3, -3, 16, -5,
    -- filter=26 channel=15
    -28, -30, 5, -3, -13, -23, -26, -10, -5,
    -- filter=27 channel=0
    -14, 21, -21, 7, -15, 0, 9, 6, 16,
    -- filter=27 channel=1
    12, -19, -7, -19, -14, -12, -4, 12, 13,
    -- filter=27 channel=2
    8, 3, -5, 12, -12, 8, -16, -12, 4,
    -- filter=27 channel=3
    -14, -4, -19, -5, 18, -14, -15, 18, 7,
    -- filter=27 channel=4
    -20, 12, -9, 12, -21, -8, 17, 9, 14,
    -- filter=27 channel=5
    6, 13, -8, 11, 16, -14, 3, 14, -18,
    -- filter=27 channel=6
    19, 0, 19, 17, -11, -7, -9, 17, -5,
    -- filter=27 channel=7
    2, -10, -7, 6, -20, -13, -10, 8, -5,
    -- filter=27 channel=8
    -19, 3, -19, 13, 11, -10, -5, -21, -3,
    -- filter=27 channel=9
    -21, -12, -3, 15, -3, 6, -11, -4, 3,
    -- filter=27 channel=10
    1, 0, -15, 1, 12, -10, -12, 17, 17,
    -- filter=27 channel=11
    11, -15, -4, 5, 14, 9, -17, 14, -8,
    -- filter=27 channel=12
    -18, -11, -18, 17, 4, 2, -9, 19, 17,
    -- filter=27 channel=13
    0, -20, -1, -18, -19, 1, -21, -2, -17,
    -- filter=27 channel=14
    0, -12, 6, 13, 11, -20, 15, 19, 17,
    -- filter=27 channel=15
    -21, -11, -14, 5, -6, -20, 16, 0, -9,
    -- filter=28 channel=0
    4, -11, 5, 4, 19, -7, -16, 2, 11,
    -- filter=28 channel=1
    -20, -11, -21, 4, -16, -7, 18, -6, 17,
    -- filter=28 channel=2
    -8, -16, -7, 12, 4, 11, 3, -15, -23,
    -- filter=28 channel=3
    8, -7, -6, 20, 6, 16, 7, 19, -12,
    -- filter=28 channel=4
    9, 10, -22, -22, -2, 10, 12, 7, 7,
    -- filter=28 channel=5
    0, 6, -4, -21, 6, 12, -14, 14, 15,
    -- filter=28 channel=6
    3, 3, -5, -6, -17, -1, 13, 17, 5,
    -- filter=28 channel=7
    20, 0, 19, 16, 20, 27, 11, -9, 8,
    -- filter=28 channel=8
    -13, 11, -21, 3, 4, -13, 3, -26, 7,
    -- filter=28 channel=9
    12, 0, 16, -15, -17, 0, -12, -2, -16,
    -- filter=28 channel=10
    0, -22, 3, 7, -19, 11, -14, -12, 2,
    -- filter=28 channel=11
    -6, -11, -10, 20, -15, 3, 8, 9, -1,
    -- filter=28 channel=12
    20, -9, 10, 9, -6, -7, 21, -7, 4,
    -- filter=28 channel=13
    -11, 16, -14, 16, -18, -20, -17, 17, 1,
    -- filter=28 channel=14
    -8, -9, 3, -16, 5, -21, -15, -14, -2,
    -- filter=28 channel=15
    14, 9, 0, -16, 12, -11, -14, -18, 15,
    -- filter=29 channel=0
    16, 17, -17, 4, 11, -22, 10, 18, -10,
    -- filter=29 channel=1
    -4, -5, 7, 5, -14, -16, -4, 13, -7,
    -- filter=29 channel=2
    7, 17, 5, 13, 14, 0, -25, -24, -19,
    -- filter=29 channel=3
    24, 12, -19, 18, -8, -27, 11, 13, -12,
    -- filter=29 channel=4
    6, -16, -11, -3, -11, -20, 0, 1, 12,
    -- filter=29 channel=5
    -6, -14, 12, 4, 0, 5, 18, 15, 18,
    -- filter=29 channel=6
    1, -19, 17, 9, 8, -2, -17, -22, -17,
    -- filter=29 channel=7
    37, 34, 25, 17, 36, 21, 37, 35, 35,
    -- filter=29 channel=8
    3, 19, 24, -1, 29, -4, -4, 16, 0,
    -- filter=29 channel=9
    17, 0, -2, 21, 26, 10, -5, 15, 16,
    -- filter=29 channel=10
    21, -6, 1, -8, 5, 9, -15, 23, 20,
    -- filter=29 channel=11
    -1, 7, -14, 0, 0, 6, 13, 16, 5,
    -- filter=29 channel=12
    -12, 12, 2, -3, 3, 7, 2, 7, 5,
    -- filter=29 channel=13
    -12, -33, 2, -24, 2, -29, -2, -30, -10,
    -- filter=29 channel=14
    2, -13, 13, -16, -17, -18, 3, 6, -9,
    -- filter=29 channel=15
    -11, -11, -33, -13, -30, -3, -14, -10, 6,
    -- filter=30 channel=0
    -20, 16, -19, 17, 12, -10, -12, 7, -5,
    -- filter=30 channel=1
    -2, -21, -9, 6, 9, 3, -15, -13, 16,
    -- filter=30 channel=2
    -13, 7, -1, -14, 10, 0, 18, -16, 4,
    -- filter=30 channel=3
    -2, 0, 5, -13, -13, 13, 17, -1, -8,
    -- filter=30 channel=4
    -20, -9, -20, -5, 17, -12, -9, 15, 19,
    -- filter=30 channel=5
    -20, -10, 17, 17, 1, -7, -3, 14, -1,
    -- filter=30 channel=6
    8, -1, -5, 11, -4, 19, -7, 3, 5,
    -- filter=30 channel=7
    3, -12, 12, 14, -5, -11, 13, -7, 15,
    -- filter=30 channel=8
    -1, 4, 5, 19, 2, -18, -3, 13, -8,
    -- filter=30 channel=9
    14, 4, 2, -15, -16, 16, 4, 5, 2,
    -- filter=30 channel=10
    -16, -4, 10, 8, -15, 18, -19, -10, -20,
    -- filter=30 channel=11
    13, 13, -20, -10, 14, 12, 13, 5, -9,
    -- filter=30 channel=12
    -11, -2, -9, 6, -19, 2, -13, 9, -20,
    -- filter=30 channel=13
    6, 0, 20, -5, -3, 10, 3, -4, -8,
    -- filter=30 channel=14
    14, -8, -11, 3, 12, -20, 1, -12, 18,
    -- filter=30 channel=15
    -10, 13, 0, 2, -12, 6, 8, -2, -16,
    -- filter=31 channel=0
    3, -18, 16, -5, 10, -17, 0, -6, -3,
    -- filter=31 channel=1
    -1, -9, -11, 2, 16, -14, 20, -18, -17,
    -- filter=31 channel=2
    -18, -8, 1, -2, 10, 11, 19, 1, 5,
    -- filter=31 channel=3
    5, 24, -8, 25, 22, -6, 19, 21, 21,
    -- filter=31 channel=4
    9, 7, 12, -20, 8, 15, -22, -16, -12,
    -- filter=31 channel=5
    -25, -26, -24, -25, 8, 2, -12, 13, -11,
    -- filter=31 channel=6
    2, -9, -8, -21, -19, -3, 2, 14, -6,
    -- filter=31 channel=7
    -27, 5, -17, -17, -20, -16, -15, 0, 1,
    -- filter=31 channel=8
    10, 14, -6, 23, 23, 1, 12, 9, 24,
    -- filter=31 channel=9
    -18, 5, -27, -32, -22, -18, -10, -22, 9,
    -- filter=31 channel=10
    -15, 3, -9, 10, 18, -15, -1, -20, 3,
    -- filter=31 channel=11
    9, -1, 14, -20, 5, -18, 4, 12, -7,
    -- filter=31 channel=12
    -8, 9, 7, 12, -2, 8, -10, 0, 3,
    -- filter=31 channel=13
    30, -6, 25, 13, 0, 31, 17, 0, 21,
    -- filter=31 channel=14
    -7, -16, 14, 6, -4, 6, -13, 0, -11,
    -- filter=31 channel=15
    -6, -5, 1, 0, -21, -16, -32, 2, 5,

    -- ifmap
    -- channel=0
    241, 239, 243, 248, 245, 251, 252, 252, 248, 239, 237, 247, 259, 270, 273, 267, 252, 232, 216, 194, 183, 181, 185, 196, 202, 209, 213, 213, 208, 193, 
    243, 245, 247, 250, 251, 257, 258, 257, 250, 241, 240, 259, 264, 262, 260, 252, 228, 204, 169, 153, 141, 137, 138, 144, 165, 182, 202, 212, 211, 200, 
    244, 251, 255, 253, 254, 257, 261, 258, 252, 246, 249, 285, 259, 235, 223, 205, 178, 142, 120, 114, 105, 101, 100, 109, 119, 150, 175, 195, 206, 203, 
    224, 232, 246, 256, 257, 260, 262, 260, 253, 230, 246, 260, 219, 183, 162, 138, 121, 90, 87, 95, 95, 86, 82, 75, 82, 102, 127, 163, 194, 205, 
    174, 184, 194, 233, 258, 265, 265, 264, 261, 234, 252, 240, 188, 154, 125, 94, 70, 61, 85, 113, 113, 98, 86, 76, 80, 70, 85, 120, 168, 197, 
    145, 127, 143, 207, 255, 265, 263, 260, 255, 234, 215, 186, 162, 135, 85, 63, 60, 63, 90, 129, 140, 117, 88, 89, 77, 54, 44, 81, 142, 188, 
    141, 83, 90, 203, 258, 263, 257, 252, 233, 226, 183, 160, 161, 136, 83, 61, 63, 58, 87, 126, 148, 122, 95, 89, 74, 54, 35, 48, 107, 170, 
    148, 85, 99, 206, 256, 250, 245, 237, 254, 235, 186, 155, 170, 141, 96, 67, 64, 57, 69, 116, 156, 133, 107, 87, 72, 58, 44, 39, 71, 132, 
    161, 79, 144, 229, 253, 228, 213, 190, 249, 231, 184, 166, 178, 148, 98, 77, 55, 60, 51, 105, 170, 149, 118, 81, 70, 72, 55, 38, 39, 92, 
    160, 92, 165, 249, 263, 229, 171, 160, 210, 249, 204, 185, 185, 159, 113, 85, 65, 52, 42, 127, 186, 156, 126, 77, 74, 78, 71, 49, 32, 57, 
    143, 90, 168, 251, 261, 245, 177, 145, 174, 224, 193, 180, 207, 187, 140, 101, 84, 60, 44, 161, 193, 163, 118, 71, 74, 78, 70, 54, 42, 54, 
    144, 84, 162, 238, 237, 248, 211, 131, 135, 200, 182, 194, 231, 222, 159, 119, 103, 60, 65, 184, 198, 153, 102, 63, 63, 74, 71, 70, 66, 80, 
    147, 89, 168, 207, 203, 230, 226, 145, 126, 169, 166, 194, 226, 216, 164, 134, 123, 64, 80, 180, 190, 140, 103, 77, 65, 73, 78, 89, 94, 110, 
    152, 114, 182, 170, 160, 192, 227, 166, 130, 152, 182, 223, 238, 187, 157, 136, 121, 75, 95, 173, 173, 134, 91, 64, 56, 67, 90, 110, 125, 133, 
    161, 136, 186, 165, 131, 139, 211, 171, 134, 108, 174, 217, 186, 148, 129, 133, 124, 98, 114, 176, 166, 142, 113, 74, 56, 71, 100, 131, 144, 156, 
    174, 147, 178, 177, 117, 103, 162, 188, 146, 111, 163, 199, 165, 130, 107, 113, 121, 118, 140, 150, 131, 130, 101, 49, 38, 63, 101, 144, 159, 185, 
    183, 151, 171, 190, 129, 90, 121, 179, 144, 127, 137, 131, 153, 129, 110, 110, 104, 128, 175, 148, 126, 122, 84, 49, 41, 75, 113, 156, 187, 213, 
    192, 162, 167, 187, 144, 84, 92, 150, 146, 133, 120, 91, 131, 117, 130, 121, 94, 121, 154, 112, 107, 97, 51, 29, 50, 102, 148, 194, 219, 228, 
    193, 183, 173, 181, 160, 97, 87, 126, 150, 118, 73, 87, 117, 130, 174, 150, 99, 107, 109, 97, 74, 37, 15, 0, 46, 103, 169, 216, 224, 216, 
    176, 201, 181, 178, 165, 102, 83, 147, 185, 173, 104, 109, 122, 155, 197, 178, 124, 101, 96, 68, 38, 10, 0, 0, 30, 74, 132, 159, 155, 143, 
    145, 201, 184, 182, 174, 119, 102, 204, 220, 167, 120, 79, 85, 127, 144, 133, 99, 65, 46, 19, 0, 0, 0, 0, 0, 12, 52, 72, 63, 51, 
    86, 154, 168, 183, 181, 131, 145, 249, 252, 186, 91, 52, 58, 71, 72, 67, 48, 31, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 80, 115, 157, 176, 135, 198, 259, 242, 163, 62, 19, 15, 16, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 60, 121, 160, 160, 230, 253, 191, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 72, 104, 159, 239, 240, 109, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 53, 134, 237, 204, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 94, 178, 145, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 103, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    41, 45, 39, 41, 45, 47, 44, 43, 44, 46, 39, 40, 48, 48, 50, 49, 44, 33, 23, 12, 10, 14, 19, 26, 32, 37, 39, 41, 41, 36, 
    43, 54, 47, 46, 49, 47, 45, 46, 46, 52, 42, 42, 48, 42, 44, 46, 32, 23, 8, 3, 0, 0, 3, 4, 12, 18, 29, 39, 41, 39, 
    43, 54, 54, 50, 51, 45, 44, 45, 49, 59, 32, 37, 40, 33, 25, 20, 9, 5, 4, 4, 0, 0, 1, 4, 3, 11, 16, 29, 36, 37, 
    28, 34, 41, 46, 50, 47, 44, 46, 50, 56, 10, 0, 2, 8, 0, 0, 3, 7, 11, 0, 0, 0, 0, 0, 0, 2, 7, 18, 29, 37, 
    0, 1, 9, 30, 48, 51, 47, 49, 53, 63, 24, 0, 0, 5, 1, 0, 8, 25, 12, 0, 0, 0, 0, 0, 0, 0, 2, 15, 20, 32, 
    0, 0, 12, 27, 44, 50, 47, 44, 42, 42, 30, 9, 4, 3, 7, 5, 4, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 16, 19, 25, 
    0, 0, 28, 44, 43, 46, 46, 42, 28, 34, 25, 24, 13, 0, 0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 17, 
    0, 0, 18, 28, 39, 40, 48, 45, 42, 42, 45, 24, 1, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 
    0, 0, 6, 0, 27, 33, 47, 24, 6, 0, 34, 12, 0, 0, 0, 0, 0, 0, 19, 20, 0, 0, 0, 1, 0, 0, 0, 0, 14, 18, 
    0, 0, 0, 0, 22, 43, 49, 25, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 32, 17, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 
    0, 0, 0, 0, 13, 50, 53, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 37, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 40, 42, 59, 4, 0, 0, 13, 0, 0, 0, 0, 0, 16, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 3, 0, 0, 0, 26, 32, 45, 15, 0, 2, 16, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 13, 25, 41, 24, 14, 13, 0, 0, 0, 0, 0, 0, 8, 18, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 6, 
    0, 1, 0, 0, 0, 0, 11, 23, 34, 8, 0, 0, 0, 0, 0, 0, 0, 23, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 
    0, 0, 0, 0, 0, 0, 0, 3, 35, 10, 0, 0, 0, 0, 0, 0, 0, 9, 18, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 18, 0, 0, 0, 0, 0, 0, 0, 0, 21, 9, 0, 0, 0, 0, 2, 14, 6, 21, 36, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 10, 40, 41, 38, 41, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 22, 20, 18, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 27, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    72, 79, 84, 78, 76, 79, 80, 75, 71, 77, 84, 82, 76, 71, 68, 65, 66, 67, 66, 64, 60, 59, 61, 64, 68, 63, 58, 52, 47, 44, 
    67, 71, 76, 77, 79, 82, 81, 79, 79, 91, 105, 94, 76, 69, 70, 71, 65, 56, 60, 66, 64, 56, 49, 50, 56, 59, 58, 56, 52, 48, 
    68, 72, 76, 73, 76, 82, 80, 77, 84, 128, 169, 128, 84, 76, 72, 59, 43, 58, 90, 106, 103, 82, 66, 51, 50, 57, 60, 61, 58, 52, 
    72, 73, 75, 73, 74, 79, 77, 74, 81, 134, 174, 135, 83, 57, 44, 29, 43, 86, 126, 151, 155, 139, 105, 88, 63, 39, 47, 63, 67, 58, 
    61, 47, 62, 76, 75, 75, 76, 73, 72, 83, 121, 133, 89, 50, 46, 55, 58, 95, 157, 185, 175, 153, 142, 125, 80, 45, 35, 57, 73, 64, 
    57, 24, 56, 85, 78, 72, 75, 73, 69, 68, 79, 110, 118, 91, 72, 76, 76, 109, 175, 197, 168, 145, 139, 122, 94, 54, 23, 39, 69, 70, 
    96, 54, 75, 97, 82, 72, 78, 88, 83, 73, 94, 139, 153, 125, 96, 95, 93, 96, 146, 192, 171, 130, 108, 105, 91, 63, 30, 18, 52, 74, 
    153, 134, 147, 128, 91, 76, 99, 159, 180, 154, 156, 177, 176, 141, 103, 98, 92, 70, 103, 178, 188, 140, 104, 98, 96, 76, 42, 10, 25, 63, 
    210, 196, 212, 176, 105, 74, 131, 244, 300, 240, 194, 206, 195, 158, 117, 91, 72, 63, 110, 180, 207, 178, 121, 98, 104, 96, 67, 17, 0, 40, 
    232, 242, 251, 208, 127, 78, 110, 223, 318, 293, 241, 238, 217, 172, 130, 102, 72, 63, 151, 227, 227, 186, 128, 108, 113, 108, 89, 54, 14, 18, 
    214, 243, 278, 224, 139, 93, 61, 147, 275, 270, 230, 257, 255, 188, 152, 133, 89, 90, 188, 256, 233, 179, 128, 103, 115, 118, 103, 84, 55, 28, 
    214, 248, 270, 206, 136, 101, 67, 94, 188, 216, 221, 276, 295, 231, 172, 158, 120, 113, 201, 267, 232, 167, 121, 94, 95, 110, 121, 114, 93, 59, 
    231, 260, 253, 180, 128, 105, 75, 70, 135, 207, 236, 270, 289, 250, 197, 168, 136, 132, 213, 265, 224, 170, 128, 101, 99, 118, 138, 135, 111, 80, 
    248, 269, 271, 182, 116, 114, 93, 73, 125, 219, 290, 294, 261, 241, 206, 164, 132, 139, 207, 251, 224, 172, 121, 102, 111, 126, 145, 140, 106, 86, 
    269, 277, 298, 214, 132, 137, 131, 99, 111, 215, 299, 283, 223, 185, 164, 158, 139, 130, 182, 231, 211, 165, 128, 104, 112, 131, 133, 117, 99, 87, 
    293, 293, 317, 249, 160, 158, 175, 121, 114, 172, 206, 232, 192, 144, 141, 135, 134, 136, 129, 149, 188, 168, 105, 71, 79, 104, 110, 104, 98, 85, 
    318, 307, 324, 283, 185, 170, 204, 175, 129, 113, 140, 162, 154, 148, 145, 129, 146, 136, 100, 121, 147, 118, 74, 53, 62, 87, 109, 109, 97, 88, 
    332, 316, 323, 303, 214, 162, 196, 209, 168, 115, 116, 139, 145, 178, 185, 143, 137, 161, 154, 116, 81, 74, 52, 46, 73, 86, 110, 110, 96, 89, 
    325, 317, 316, 305, 238, 176, 202, 229, 200, 128, 91, 120, 170, 233, 246, 179, 128, 134, 131, 101, 66, 39, 31, 55, 83, 96, 102, 100, 87, 80, 
    315, 311, 304, 296, 239, 191, 254, 294, 239, 192, 156, 179, 243, 280, 292, 244, 155, 105, 77, 67, 69, 54, 61, 79, 95, 119, 116, 107, 95, 89, 
    311, 316, 302, 286, 232, 219, 321, 409, 358, 270, 223, 224, 249, 273, 281, 243, 179, 115, 77, 76, 87, 104, 112, 118, 122, 136, 146, 145, 130, 126, 
    287, 317, 309, 298, 266, 277, 355, 428, 417, 297, 201, 192, 202, 209, 210, 193, 167, 147, 128, 120, 123, 135, 150, 160, 164, 173, 184, 180, 175, 173, 
    232, 284, 306, 305, 288, 316, 388, 410, 332, 244, 188, 157, 157, 156, 158, 163, 154, 143, 141, 148, 157, 158, 165, 179, 190, 190, 192, 194, 191, 186, 
    183, 221, 270, 275, 288, 354, 405, 357, 263, 202, 167, 154, 151, 146, 144, 143, 144, 146, 148, 156, 167, 172, 181, 195, 205, 202, 200, 201, 203, 215, 
    185, 171, 200, 241, 292, 369, 386, 300, 218, 181, 168, 164, 158, 152, 150, 148, 148, 152, 157, 164, 178, 189, 199, 203, 200, 200, 202, 217, 239, 254, 
    201, 173, 163, 199, 279, 372, 366, 271, 193, 168, 172, 168, 160, 154, 153, 152, 156, 160, 167, 176, 186, 198, 202, 199, 192, 190, 210, 244, 251, 237, 
    206, 186, 172, 167, 226, 331, 336, 241, 179, 166, 175, 181, 170, 159, 155, 154, 159, 167, 176, 181, 183, 193, 199, 197, 190, 202, 229, 235, 214, 198, 
    209, 192, 186, 173, 169, 237, 267, 200, 161, 159, 168, 180, 184, 173, 162, 162, 171, 179, 182, 186, 186, 181, 181, 193, 212, 235, 240, 228, 196, 173, 
    207, 192, 189, 183, 164, 161, 193, 172, 134, 137, 150, 161, 169, 171, 171, 175, 182, 192, 200, 197, 185, 176, 179, 204, 243, 267, 266, 236, 185, 152, 
    213, 189, 185, 183, 176, 157, 150, 146, 127, 123, 127, 133, 140, 145, 147, 158, 180, 205, 217, 203, 185, 176, 181, 211, 257, 283, 267, 219, 185, 154, 
    
    -- channel=4
    25, 23, 27, 24, 11, 7, 11, 11, 11, 12, 14, 18, 20, 23, 24, 20, 16, 24, 44, 63, 71, 69, 59, 46, 29, 13, 13, 16, 15, 11, 
    19, 13, 18, 17, 9, 6, 10, 11, 5, 0, 0, 0, 18, 24, 19, 17, 31, 54, 60, 52, 51, 67, 80, 86, 83, 58, 28, 13, 8, 2, 
    6, 0, 8, 14, 9, 13, 17, 18, 7, 0, 0, 0, 2, 22, 41, 84, 115, 78, 12, 0, 0, 0, 0, 28, 45, 60, 52, 27, 16, 13, 
    22, 27, 28, 28, 20, 23, 26, 24, 17, 0, 27, 69, 69, 90, 131, 137, 100, 26, 0, 0, 0, 0, 0, 0, 0, 29, 64, 45, 20, 12, 
    74, 122, 104, 47, 16, 13, 18, 13, 14, 34, 112, 173, 90, 62, 70, 48, 0, 0, 0, 0, 0, 10, 0, 0, 0, 28, 46, 47, 28, 13, 
    59, 90, 70, 39, 20, 17, 14, 9, 13, 39, 61, 47, 0, 0, 0, 0, 0, 0, 0, 0, 2, 30, 21, 17, 35, 31, 15, 25, 37, 30, 
    0, 0, 0, 0, 17, 19, 9, 0, 9, 34, 7, 0, 0, 0, 0, 0, 0, 0, 24, 40, 22, 15, 35, 53, 43, 10, 10, 16, 32, 31, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 26, 15, 12, 35, 42, 23, 31, 28, 0, 0, 18, 8, 0, 0, 5, 34, 51, 
    0, 0, 0, 0, 16, 27, 0, 0, 0, 0, 0, 0, 15, 26, 0, 0, 29, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 52, 
    36, 0, 0, 14, 25, 16, 24, 42, 79, 83, 23, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 15, 38, 12, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 38, 34, 4, 24, 50, 142, 155, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 68, 70, 20, 8, 15, 0, 0, 0, 0, 
    40, 0, 2, 101, 92, 28, 26, 0, 35, 104, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 74, 58, 16, 21, 27, 0, 0, 0, 0, 
    10, 0, 0, 106, 98, 47, 40, 8, 13, 35, 0, 0, 50, 76, 0, 0, 26, 0, 0, 20, 66, 28, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 58, 20, 24, 35, 0, 0, 0, 0, 0, 68, 129, 69, 38, 34, 0, 0, 34, 54, 40, 33, 9, 0, 0, 0, 0, 10, 0, 
    0, 0, 1, 16, 0, 0, 10, 0, 0, 0, 0, 94, 102, 91, 82, 80, 51, 0, 0, 38, 48, 17, 32, 26, 8, 10, 26, 52, 25, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 39, 132, 235, 188, 74, 56, 42, 9, 0, 40, 127, 95, 48, 45, 44, 36, 45, 40, 20, 0, 0, 
    0, 0, 0, 32, 16, 0, 0, 0, 0, 30, 129, 103, 54, 0, 0, 0, 0, 0, 5, 58, 83, 130, 124, 78, 36, 14, 0, 0, 0, 0, 
    22, 0, 1, 26, 22, 0, 10, 40, 0, 0, 30, 15, 0, 0, 0, 0, 0, 11, 0, 0, 7, 121, 99, 2, 0, 0, 0, 0, 0, 15, 
    40, 4, 5, 19, 31, 0, 0, 0, 42, 58, 5, 0, 0, 0, 0, 0, 0, 59, 115, 111, 111, 85, 41, 0, 0, 0, 0, 8, 36, 38, 
    36, 12, 8, 27, 65, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 139, 100, 5, 0, 0, 0, 8, 36, 74, 76, 72, 
    13, 18, 6, 26, 58, 0, 0, 0, 0, 0, 0, 0, 0, 31, 106, 111, 72, 31, 2, 0, 0, 0, 0, 0, 0, 0, 33, 55, 49, 38, 
    51, 69, 11, 4, 0, 0, 0, 0, 59, 109, 106, 140, 184, 226, 238, 212, 150, 83, 19, 0, 0, 0, 0, 0, 0, 0, 1, 6, 2, 0, 
    102, 158, 74, 41, 12, 0, 0, 27, 198, 264, 193, 100, 94, 101, 93, 82, 49, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 101, 112, 100, 33, 0, 0, 148, 249, 184, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 64, 109, 9, 0, 26, 202, 200, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 6, 0, 0, 0, 
    0, 0, 11, 54, 19, 0, 90, 174, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 26, 0, 0, 0, 11, 
    1, 0, 0, 1, 30, 89, 177, 162, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 19, 1, 0, 0, 0, 56, 95, 
    0, 0, 0, 0, 21, 122, 250, 184, 64, 35, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 53, 49, 
    0, 0, 0, 0, 0, 39, 134, 136, 36, 32, 32, 39, 43, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    11, 0, 0, 0, 0, 0, 10, 32, 11, 0, 0, 18, 38, 56, 57, 33, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 25, 0, 
    
    -- channel=5
    117, 117, 112, 108, 111, 109, 109, 108, 108, 106, 106, 111, 118, 121, 120, 116, 110, 110, 108, 109, 110, 111, 113, 106, 103, 102, 104, 107, 103, 98, 
    116, 119, 115, 109, 109, 109, 109, 108, 104, 86, 84, 93, 108, 115, 112, 105, 107, 96, 96, 85, 86, 97, 107, 118, 115, 113, 107, 104, 100, 96, 
    106, 113, 114, 112, 110, 113, 111, 113, 108, 67, 55, 51, 88, 104, 110, 119, 110, 89, 63, 35, 27, 35, 60, 73, 98, 108, 111, 106, 103, 98, 
    101, 112, 119, 118, 117, 118, 117, 117, 120, 127, 97, 80, 101, 121, 120, 117, 95, 73, 41, 20, 9, 13, 16, 31, 57, 85, 110, 109, 102, 96, 
    112, 127, 140, 129, 118, 114, 114, 115, 119, 146, 132, 108, 90, 85, 81, 72, 61, 51, 37, 27, 28, 31, 28, 34, 32, 64, 96, 111, 105, 96, 
    70, 96, 127, 131, 121, 118, 114, 110, 109, 118, 105, 80, 51, 29, 30, 31, 44, 56, 47, 32, 34, 44, 55, 46, 45, 46, 76, 104, 111, 103, 
    12, 22, 67, 93, 113, 116, 110, 91, 95, 80, 75, 53, 30, 26, 37, 40, 44, 74, 80, 59, 35, 46, 64, 60, 50, 40, 60, 94, 110, 108, 
    0, 0, 22, 56, 95, 110, 77, 39, 0, 1, 20, 37, 27, 34, 43, 53, 57, 72, 87, 74, 34, 30, 42, 51, 42, 31, 37, 77, 109, 114, 
    0, 0, 11, 53, 87, 113, 75, 41, 0, 0, 2, 31, 29, 25, 39, 38, 59, 55, 58, 45, 14, 20, 24, 35, 41, 32, 29, 47, 92, 116, 
    4, 22, 18, 49, 82, 100, 126, 99, 66, 30, 33, 23, 22, 22, 28, 33, 44, 37, 41, 19, 8, 30, 34, 49, 40, 36, 26, 28, 52, 95, 
    17, 35, 35, 46, 84, 90, 118, 112, 110, 74, 61, 36, 10, 12, 20, 21, 20, 24, 54, 22, 30, 39, 45, 57, 53, 47, 30, 23, 29, 63, 
    6, 31, 42, 57, 104, 104, 91, 92, 95, 64, 65, 39, 7, 0, 17, 24, 12, 27, 56, 34, 37, 40, 47, 55, 62, 53, 40, 24, 27, 45, 
    0, 25, 21, 52, 105, 116, 93, 93, 84, 49, 43, 43, 36, 22, 25, 34, 23, 45, 55, 36, 23, 25, 30, 33, 43, 40, 32, 26, 40, 49, 
    3, 26, 0, 23, 65, 103, 83, 77, 66, 38, 9, 21, 30, 59, 54, 44, 35, 60, 64, 38, 34, 35, 41, 41, 38, 38, 40, 48, 56, 70, 
    1, 18, 0, 0, 20, 68, 55, 82, 57, 78, 62, 40, 52, 66, 71, 60, 53, 64, 78, 49, 35, 30, 39, 51, 54, 57, 68, 72, 74, 82, 
    0, 10, 0, 0, 18, 40, 42, 51, 72, 109, 112, 100, 88, 66, 67, 51, 44, 81, 104, 93, 73, 48, 42, 65, 74, 71, 73, 69, 79, 80, 
    0, 4, 7, 0, 12, 34, 41, 15, 57, 88, 87, 86, 52, 40, 36, 32, 44, 62, 55, 88, 95, 76, 78, 72, 81, 78, 72, 72, 85, 90, 
    6, 5, 11, 0, 0, 31, 52, 27, 24, 47, 54, 71, 33, 24, 2, 15, 54, 60, 25, 41, 61, 75, 72, 47, 49, 60, 72, 80, 90, 98, 
    26, 12, 15, 3, 0, 14, 18, 32, 32, 38, 63, 55, 35, 25, 0, 0, 48, 85, 95, 78, 68, 73, 56, 56, 46, 69, 81, 89, 93, 98, 
    40, 14, 21, 18, 12, 15, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 53, 82, 80, 56, 30, 17, 25, 32, 63, 73, 78, 80, 75, 
    37, 11, 20, 17, 6, 4, 8, 0, 0, 0, 0, 1, 27, 38, 42, 26, 20, 25, 19, 14, 7, 0, 0, 0, 8, 22, 35, 37, 32, 31, 
    44, 27, 17, 0, 0, 0, 4, 0, 0, 0, 40, 80, 91, 100, 93, 65, 48, 30, 9, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    65, 63, 42, 25, 0, 12, 3, 24, 37, 41, 52, 46, 44, 45, 43, 28, 17, 13, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 62, 66, 46, 22, 34, 23, 36, 24, 28, 6, 0, 0, 0, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 60, 44, 34, 27, 30, 15, 23, 10, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 43, 49, 44, 16, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 72, 72, 37, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 
    0, 0, 0, 0, 54, 91, 62, 33, 23, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 4, 48, 38, 31, 15, 20, 24, 21, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 7, 7, 3, 7, 11, 14, 24, 28, 30, 23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    86, 89, 88, 80, 79, 76, 75, 75, 77, 79, 78, 80, 88, 94, 93, 89, 83, 88, 96, 107, 109, 108, 104, 91, 81, 72, 72, 75, 71, 64, 
    82, 87, 88, 80, 78, 75, 77, 73, 68, 48, 42, 52, 77, 89, 85, 81, 94, 96, 98, 80, 78, 89, 107, 121, 113, 100, 80, 69, 63, 58, 
    74, 77, 79, 83, 81, 83, 82, 83, 74, 9, 0, 0, 54, 82, 102, 129, 138, 97, 39, 0, 0, 0, 26, 54, 83, 87, 88, 77, 70, 63, 
    82, 90, 94, 91, 88, 90, 90, 88, 90, 85, 96, 88, 101, 133, 155, 158, 100, 44, 0, 0, 0, 0, 0, 0, 19, 66, 96, 85, 71, 61, 
    125, 137, 140, 103, 83, 84, 83, 82, 90, 156, 167, 133, 97, 91, 73, 45, 17, 7, 0, 0, 0, 8, 0, 0, 2, 46, 73, 84, 76, 62, 
    80, 94, 99, 90, 83, 86, 82, 81, 85, 116, 108, 65, 17, 0, 0, 0, 0, 13, 12, 7, 16, 25, 33, 32, 24, 22, 50, 75, 86, 75, 
    0, 0, 0, 27, 72, 87, 80, 62, 76, 70, 45, 4, 0, 0, 2, 8, 17, 53, 68, 58, 23, 25, 56, 55, 35, 5, 24, 66, 85, 78, 
    0, 0, 0, 0, 49, 79, 42, 0, 0, 0, 0, 0, 6, 21, 22, 32, 39, 69, 81, 63, 15, 6, 17, 25, 11, 0, 0, 44, 83, 96, 
    0, 0, 0, 2, 46, 92, 34, 0, 0, 0, 0, 15, 20, 5, 10, 11, 48, 29, 13, 3, 0, 0, 0, 1, 3, 0, 0, 13, 65, 98, 
    0, 0, 0, 10, 35, 77, 115, 129, 111, 44, 26, 7, 4, 0, 5, 0, 19, 0, 0, 0, 0, 16, 21, 23, 11, 2, 0, 0, 9, 64, 
    8, 20, 13, 15, 44, 56, 133, 149, 163, 104, 72, 19, 0, 0, 0, 0, 0, 0, 0, 0, 30, 45, 38, 37, 27, 21, 0, 0, 0, 17, 
    0, 1, 32, 54, 92, 74, 80, 90, 119, 84, 53, 5, 0, 0, 0, 0, 0, 0, 18, 32, 46, 39, 31, 36, 47, 35, 7, 0, 0, 0, 
    0, 0, 26, 56, 88, 89, 76, 86, 94, 28, 7, 20, 48, 26, 0, 7, 2, 6, 31, 38, 22, 7, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 1, 0, 9, 31, 72, 60, 53, 41, 0, 0, 9, 47, 74, 47, 44, 21, 20, 45, 43, 24, 14, 28, 16, 2, 0, 0, 15, 18, 14, 
    0, 3, 0, 0, 0, 37, 21, 39, 22, 58, 55, 82, 79, 77, 88, 64, 29, 20, 57, 44, 36, 18, 19, 26, 29, 39, 53, 55, 34, 27, 
    0, 0, 0, 0, 0, 10, 9, 22, 36, 129, 185, 165, 122, 69, 65, 42, 14, 37, 111, 131, 87, 36, 30, 59, 68, 68, 63, 33, 27, 36, 
    0, 0, 1, 0, 0, 0, 15, 0, 25, 101, 122, 100, 37, 2, 5, 2, 0, 34, 55, 79, 93, 106, 97, 68, 64, 35, 17, 4, 28, 51, 
    2, 0, 6, 0, 0, 5, 43, 9, 2, 29, 22, 53, 0, 0, 0, 0, 17, 33, 0, 6, 66, 88, 69, 12, 0, 0, 4, 29, 55, 70, 
    33, 4, 8, 0, 0, 0, 0, 8, 6, 34, 45, 44, 4, 0, 0, 0, 17, 77, 111, 108, 91, 72, 35, 20, 0, 16, 43, 71, 81, 87, 
    48, 8, 13, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 107, 108, 50, 0, 0, 0, 0, 42, 71, 88, 86, 83, 
    39, 4, 10, 22, 7, 0, 0, 0, 0, 0, 0, 0, 19, 64, 78, 54, 21, 20, 2, 0, 0, 0, 0, 0, 0, 7, 26, 26, 22, 18, 
    64, 39, 12, 0, 0, 0, 0, 0, 0, 35, 87, 135, 169, 186, 175, 134, 78, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    99, 98, 58, 25, 0, 0, 0, 59, 134, 132, 93, 68, 65, 64, 57, 28, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 75, 86, 78, 6, 0, 26, 115, 113, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 74, 61, 9, 0, 67, 95, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 39, 35, 50, 70, 29, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 78, 116, 104, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 30, 
    0, 0, 0, 0, 69, 141, 139, 64, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 67, 63, 38, 6, 5, 12, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 21, 23, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    153, 150, 143, 142, 148, 152, 152, 153, 152, 145, 139, 143, 153, 157, 158, 158, 152, 146, 138, 131, 126, 127, 130, 132, 135, 139, 142, 146, 147, 148, 
    160, 155, 144, 140, 148, 153, 153, 154, 154, 140, 134, 139, 149, 154, 151, 145, 137, 124, 119, 114, 110, 113, 114, 116, 123, 135, 144, 150, 152, 151, 
    157, 155, 149, 143, 147, 153, 152, 153, 152, 140, 136, 128, 136, 141, 130, 118, 107, 103, 110, 102, 99, 96, 101, 102, 110, 130, 143, 147, 150, 150, 
    141, 143, 146, 150, 151, 153, 152, 154, 154, 146, 127, 107, 120, 119, 103, 93, 100, 108, 97, 87, 89, 95, 93, 97, 107, 109, 129, 142, 145, 145, 
    115, 124, 147, 161, 158, 154, 155, 157, 156, 126, 109, 122, 116, 101, 102, 117, 111, 95, 87, 84, 85, 86, 92, 99, 92, 101, 121, 135, 141, 139, 
    98, 104, 151, 173, 163, 156, 156, 151, 148, 136, 120, 120, 120, 111, 106, 108, 102, 95, 94, 86, 80, 87, 95, 90, 96, 105, 108, 120, 135, 140, 
    96, 107, 135, 158, 160, 156, 151, 140, 133, 122, 123, 117, 105, 98, 95, 99, 100, 93, 90, 90, 87, 88, 87, 90, 98, 104, 112, 110, 127, 144, 
    83, 104, 125, 133, 151, 154, 137, 123, 113, 106, 108, 93, 79, 83, 85, 93, 99, 89, 81, 95, 94, 87, 86, 95, 102, 104, 106, 108, 120, 140, 
    81, 85, 101, 130, 144, 145, 124, 109, 88, 76, 55, 64, 67, 80, 88, 87, 92, 96, 97, 91, 86, 95, 89, 89, 99, 104, 106, 102, 104, 127, 
    69, 82, 83, 125, 145, 141, 105, 65, 47, 53, 50, 59, 67, 78, 87, 87, 100, 96, 104, 91, 75, 84, 83, 93, 97, 97, 101, 105, 101, 110, 
    57, 65, 86, 119, 141, 143, 95, 41, 62, 63, 58, 65, 79, 76, 89, 96, 97, 97, 98, 76, 65, 78, 87, 91, 96, 103, 96, 99, 102, 110, 
    57, 64, 77, 99, 135, 146, 121, 67, 65, 67, 75, 79, 84, 84, 89, 94, 97, 87, 78, 68, 74, 82, 93, 91, 90, 97, 99, 100, 104, 119, 
    64, 64, 60, 82, 132, 150, 134, 89, 78, 91, 91, 66, 71, 79, 86, 83, 90, 83, 73, 72, 75, 86, 92, 91, 94, 100, 101, 99, 109, 128, 
    60, 55, 63, 83, 109, 140, 138, 108, 96, 94, 82, 56, 51, 79, 90, 80, 86, 91, 78, 72, 81, 92, 88, 89, 98, 95, 97, 105, 114, 139, 
    53, 45, 63, 83, 86, 115, 129, 132, 104, 85, 76, 58, 56, 77, 75, 88, 110, 102, 86, 83, 82, 80, 91, 92, 92, 92, 96, 110, 129, 146, 
    44, 38, 55, 76, 79, 90, 108, 115, 103, 84, 41, 70, 92, 84, 91, 90, 106, 116, 99, 79, 95, 98, 89, 86, 86, 89, 99, 119, 139, 140, 
    43, 36, 47, 71, 72, 71, 95, 106, 101, 75, 67, 90, 99, 101, 97, 89, 111, 109, 83, 97, 107, 86, 86, 94, 100, 115, 129, 136, 139, 138, 
    53, 43, 48, 70, 77, 60, 73, 91, 90, 82, 87, 103, 91, 97, 90, 81, 94, 111, 111, 98, 73, 89, 103, 95, 112, 125, 138, 137, 135, 142, 
    63, 55, 55, 65, 74, 60, 59, 76, 88, 89, 76, 84, 84, 90, 84, 76, 80, 99, 97, 85, 83, 95, 97, 95, 105, 121, 129, 131, 134, 140, 
    73, 61, 58, 62, 72, 67, 70, 68, 56, 85, 90, 79, 87, 65, 61, 76, 74, 77, 78, 82, 99, 96, 89, 82, 79, 96, 100, 105, 107, 108, 
    71, 61, 58, 57, 66, 72, 80, 81, 70, 65, 78, 68, 49, 35, 44, 56, 70, 76, 74, 88, 93, 93, 81, 66, 68, 70, 80, 91, 87, 87, 
    57, 60, 54, 57, 76, 82, 65, 43, 62, 48, 35, 42, 33, 33, 38, 43, 59, 79, 83, 79, 75, 68, 62, 58, 58, 62, 70, 69, 67, 67, 
    45, 62, 57, 63, 76, 72, 47, 32, 19, 31, 62, 54, 50, 52, 54, 63, 70, 70, 69, 68, 68, 62, 58, 58, 59, 59, 57, 59, 60, 58, 
    46, 59, 63, 57, 64, 73, 47, 27, 25, 63, 71, 66, 63, 63, 64, 65, 68, 68, 68, 67, 64, 63, 61, 60, 60, 58, 55, 54, 52, 57, 
    61, 57, 52, 65, 71, 60, 36, 27, 52, 70, 62, 60, 58, 60, 63, 67, 70, 71, 70, 65, 63, 63, 61, 58, 54, 54, 51, 52, 59, 62, 
    62, 62, 51, 58, 63, 48, 37, 49, 73, 64, 61, 59, 60, 64, 64, 65, 65, 65, 62, 60, 59, 59, 54, 50, 52, 51, 52, 60, 58, 45, 
    59, 62, 57, 47, 41, 44, 54, 65, 76, 65, 60, 65, 63, 64, 63, 60, 58, 57, 57, 54, 52, 55, 57, 57, 55, 55, 58, 48, 42, 44, 
    57, 58, 55, 49, 34, 36, 66, 71, 77, 72, 65, 64, 67, 65, 60, 58, 57, 57, 54, 54, 58, 57, 56, 60, 63, 60, 45, 37, 52, 63, 
    52, 54, 52, 52, 50, 40, 66, 88, 73, 72, 69, 67, 67, 67, 67, 64, 59, 55, 57, 58, 58, 61, 62, 66, 63, 52, 43, 52, 61, 62, 
    58, 54, 51, 53, 64, 66, 67, 79, 77, 74, 69, 65, 68, 71, 71, 65, 62, 63, 64, 59, 59, 66, 66, 63, 55, 49, 42, 45, 60, 67, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 47, 63, 53, 23, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 49, 56, 39, 44, 60, 32, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 27, 14, 22, 0, 0, 4, 55, 35, 12, 33, 72, 75, 1, 0, 0, 0, 
    99, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 42, 19, 37, 0, 0, 0, 44, 42, 8, 16, 61, 75, 49, 0, 0, 0, 
    137, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 63, 52, 26, 41, 20, 0, 0, 15, 55, 37, 20, 35, 65, 72, 13, 0, 0, 
    124, 25, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 31, 56, 59, 47, 55, 26, 0, 0, 1, 53, 69, 25, 20, 51, 73, 68, 0, 0, 
    98, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 43, 50, 51, 53, 79, 15, 0, 0, 24, 54, 79, 20, 9, 43, 68, 85, 32, 0, 
    117, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 21, 70, 31, 46, 96, 5, 0, 0, 55, 64, 79, 23, 0, 31, 57, 77, 59, 0, 
    125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 38, 20, 95, 0, 0, 0, 79, 74, 70, 33, 8, 7, 34, 60, 53, 9, 
    109, 0, 52, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 34, 28, 82, 0, 0, 0, 79, 73, 73, 49, 25, 3, 12, 44, 37, 0, 
    91, 0, 75, 131, 0, 0, 0, 0, 0, 0, 0, 2, 38, 25, 13, 33, 67, 0, 0, 0, 65, 66, 70, 41, 14, 3, 0, 22, 6, 0, 
    87, 0, 55, 165, 25, 0, 0, 0, 0, 0, 0, 35, 74, 20, 0, 13, 33, 0, 0, 0, 41, 63, 74, 47, 0, 0, 0, 0, 0, 0, 
    97, 0, 29, 160, 105, 0, 0, 1, 0, 0, 0, 0, 49, 5, 5, 15, 0, 0, 0, 0, 0, 55, 81, 45, 1, 0, 0, 0, 0, 0, 
    101, 28, 24, 131, 159, 0, 0, 16, 2, 0, 0, 0, 1, 0, 22, 46, 0, 0, 0, 0, 0, 42, 70, 41, 0, 0, 0, 0, 0, 0, 
    77, 49, 29, 96, 170, 40, 0, 10, 31, 47, 0, 0, 0, 0, 35, 106, 0, 0, 0, 15, 22, 45, 61, 24, 0, 0, 0, 0, 0, 0, 
    26, 45, 24, 64, 154, 85, 0, 33, 52, 76, 10, 0, 0, 0, 33, 145, 33, 0, 0, 26, 71, 69, 48, 18, 0, 0, 0, 0, 0, 0, 
    0, 38, 11, 48, 140, 77, 0, 45, 134, 102, 51, 0, 0, 0, 35, 138, 108, 32, 41, 53, 79, 91, 77, 66, 15, 0, 0, 0, 0, 0, 
    0, 46, 14, 52, 136, 34, 0, 0, 151, 157, 90, 20, 1, 3, 48, 118, 124, 103, 106, 109, 106, 108, 121, 125, 113, 75, 57, 72, 88, 86, 
    0, 43, 25, 55, 112, 0, 0, 0, 103, 204, 139, 68, 62, 68, 83, 129, 144, 130, 146, 147, 149, 147, 157, 172, 182, 174, 165, 172, 186, 191, 
    47, 34, 13, 52, 56, 0, 0, 21, 162, 216, 184, 138, 135, 140, 140, 160, 174, 166, 170, 172, 180, 185, 188, 193, 199, 204, 197, 201, 213, 214, 
    176, 77, 10, 50, 1, 0, 0, 130, 223, 218, 186, 170, 175, 174, 172, 176, 185, 187, 189, 191, 198, 202, 200, 198, 199, 206, 207, 214, 216, 208, 
    257, 169, 62, 38, 0, 0, 27, 220, 241, 191, 182, 184, 189, 183, 178, 180, 187, 189, 192, 198, 203, 208, 205, 206, 204, 207, 209, 211, 209, 207, 
    276, 229, 155, 68, 0, 0, 114, 260, 226, 178, 180, 190, 198, 186, 178, 181, 186, 191, 194, 205, 210, 206, 212, 222, 228, 223, 208, 206, 221, 215, 
    276, 250, 215, 151, 0, 0, 138, 266, 190, 183, 176, 186, 205, 194, 186, 183, 186, 191, 198, 213, 222, 214, 217, 230, 238, 227, 220, 232, 249, 219, 
    281, 255, 235, 211, 113, 0, 126, 239, 178, 176, 169, 171, 191, 200, 196, 187, 188, 196, 205, 213, 227, 227, 219, 213, 215, 221, 245, 272, 286, 227, 
    280, 250, 237, 229, 197, 124, 131, 216, 193, 178, 169, 170, 174, 182, 184, 176, 182, 189, 203, 221, 228, 224, 208, 183, 176, 208, 260, 298, 293, 237, 
    265, 244, 227, 228, 213, 197, 172, 197, 208, 189, 182, 185, 181, 179, 165, 151, 155, 164, 187, 220, 222, 212, 188, 152, 142, 186, 262, 298, 270, 245, 
    
    -- channel=9
    141, 138, 133, 131, 134, 134, 135, 135, 138, 132, 123, 127, 138, 143, 147, 146, 139, 133, 126, 121, 117, 118, 120, 117, 117, 119, 126, 134, 136, 133, 
    146, 141, 135, 134, 136, 135, 135, 135, 133, 118, 110, 117, 133, 137, 133, 126, 123, 118, 120, 112, 108, 110, 114, 118, 117, 121, 125, 129, 131, 131, 
    138, 131, 127, 130, 134, 136, 135, 137, 134, 104, 82, 80, 113, 120, 116, 116, 118, 112, 95, 71, 62, 68, 86, 98, 113, 122, 125, 125, 127, 128, 
    120, 117, 122, 131, 139, 141, 141, 142, 143, 124, 96, 92, 114, 120, 120, 127, 122, 98, 65, 50, 45, 47, 52, 63, 81, 102, 121, 124, 124, 126, 
    118, 124, 139, 139, 139, 140, 140, 142, 147, 157, 154, 147, 127, 121, 120, 111, 88, 71, 62, 59, 61, 67, 67, 67, 71, 97, 114, 121, 120, 119, 
    102, 126, 148, 142, 136, 139, 138, 136, 137, 137, 127, 116, 92, 73, 69, 70, 74, 74, 69, 62, 70, 82, 83, 78, 84, 87, 100, 115, 121, 122, 
    61, 72, 93, 113, 134, 141, 134, 119, 118, 113, 104, 81, 62, 61, 68, 73, 78, 88, 88, 81, 71, 77, 88, 93, 93, 87, 94, 107, 121, 125, 
    35, 35, 43, 75, 120, 134, 112, 77, 50, 51, 56, 54, 52, 68, 78, 87, 89, 95, 104, 99, 72, 68, 80, 89, 85, 76, 80, 101, 120, 128, 
    24, 24, 28, 72, 113, 135, 98, 43, 0, 0, 11, 46, 56, 65, 73, 75, 92, 92, 85, 70, 54, 57, 58, 70, 77, 72, 72, 82, 107, 128, 
    43, 40, 35, 77, 113, 132, 123, 84, 50, 37, 43, 45, 51, 56, 68, 73, 85, 77, 63, 40, 34, 58, 68, 77, 74, 75, 73, 71, 81, 109, 
    48, 55, 52, 71, 105, 120, 132, 122, 112, 81, 68, 54, 44, 49, 65, 67, 70, 63, 55, 37, 52, 73, 83, 86, 83, 81, 69, 63, 63, 88, 
    47, 53, 55, 76, 114, 121, 120, 102, 99, 93, 86, 59, 41, 39, 53, 60, 58, 52, 57, 56, 70, 79, 83, 83, 88, 90, 79, 64, 64, 81, 
    37, 39, 47, 82, 117, 125, 122, 104, 96, 82, 60, 43, 50, 49, 53, 63, 68, 63, 60, 61, 63, 71, 73, 75, 83, 81, 71, 63, 73, 89, 
    31, 36, 41, 63, 86, 115, 114, 103, 95, 69, 37, 38, 62, 85, 73, 70, 76, 80, 76, 71, 70, 66, 68, 70, 69, 66, 68, 78, 95, 113, 
    24, 28, 34, 44, 53, 85, 86, 95, 80, 76, 44, 44, 69, 89, 98, 95, 87, 85, 97, 88, 78, 76, 89, 89, 83, 80, 86, 102, 116, 121, 
    17, 21, 26, 31, 42, 62, 74, 88, 93, 103, 110, 129, 119, 98, 101, 87, 83, 92, 103, 105, 97, 75, 71, 86, 92, 94, 102, 107, 109, 109, 
    17, 19, 30, 35, 47, 55, 63, 59, 76, 94, 114, 121, 101, 87, 79, 70, 71, 82, 102, 127, 115, 103, 111, 108, 109, 107, 110, 107, 112, 121, 
    35, 28, 37, 39, 43, 48, 64, 56, 55, 74, 86, 89, 63, 55, 45, 54, 73, 83, 65, 62, 83, 114, 111, 85, 84, 89, 103, 108, 120, 131, 
    55, 40, 45, 45, 43, 43, 52, 61, 54, 61, 71, 78, 66, 47, 27, 38, 70, 98, 101, 90, 95, 100, 88, 74, 59, 74, 91, 104, 113, 118, 
    60, 39, 46, 50, 50, 43, 24, 7, 24, 50, 55, 36, 25, 8, 14, 21, 35, 82, 116, 121, 105, 79, 63, 57, 56, 73, 71, 79, 83, 81, 
    48, 30, 39, 48, 55, 49, 26, 0, 0, 0, 0, 0, 6, 19, 38, 36, 31, 47, 60, 62, 50, 34, 20, 18, 29, 48, 61, 66, 64, 63, 
    44, 35, 31, 34, 32, 18, 8, 6, 17, 13, 42, 77, 90, 99, 103, 91, 79, 67, 46, 26, 25, 30, 33, 31, 35, 40, 45, 45, 44, 42, 
    70, 65, 45, 37, 24, 20, 12, 33, 63, 89, 99, 88, 86, 87, 88, 77, 63, 56, 52, 46, 44, 41, 41, 38, 35, 35, 38, 39, 35, 30, 
    62, 82, 73, 63, 50, 42, 28, 54, 76, 80, 53, 39, 35, 36, 43, 45, 48, 52, 51, 47, 44, 40, 34, 29, 24, 25, 24, 24, 22, 19, 
    27, 51, 71, 68, 45, 25, 36, 65, 83, 61, 40, 38, 39, 43, 48, 50, 49, 47, 42, 37, 31, 27, 24, 24, 27, 34, 29, 23, 14, 6, 
    27, 35, 52, 61, 45, 32, 45, 61, 64, 43, 39, 40, 43, 45, 44, 42, 40, 36, 34, 33, 29, 27, 26, 32, 42, 44, 36, 22, 14, 22, 
    29, 29, 29, 42, 58, 63, 68, 58, 54, 40, 39, 38, 35, 39, 42, 42, 39, 36, 34, 34, 37, 43, 44, 41, 39, 30, 20, 16, 39, 59, 
    26, 28, 26, 30, 60, 92, 102, 82, 69, 55, 47, 40, 35, 31, 34, 38, 38, 35, 34, 36, 38, 41, 45, 43, 30, 13, 9, 27, 52, 57, 
    25, 30, 29, 28, 43, 77, 98, 91, 69, 69, 66, 61, 56, 47, 40, 32, 27, 24, 26, 30, 35, 43, 43, 33, 14, 3, 6, 20, 26, 41, 
    32, 31, 32, 34, 37, 47, 58, 63, 56, 57, 60, 65, 72, 70, 66, 59, 49, 37, 27, 26, 34, 41, 36, 28, 17, 13, 17, 29, 38, 43, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 4, 7, 13, 11, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 23, 12, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 38, 37, 32, 6, 0, 0, 0, 0, 0, 0, 3, 13, 0, 0, 0, 
    0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 19, 1, 4, 25, 30, 17, 15, 3, 0, 0, 17, 13, 7, 9, 20, 21, 13, 0, 0, 
    6, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 15, 15, 0, 0, 15, 27, 23, 32, 38, 27, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 24, 24, 37, 28, 0, 0, 25, 38, 40, 32, 33, 26, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 32, 39, 42, 40, 32, 0, 0, 0, 23, 28, 21, 17, 23, 29, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 37, 38, 27, 0, 0, 0, 0, 9, 15, 14, 19, 19, 25, 29, 
    0, 15, 0, 0, 0, 0, 0, 38, 6, 0, 0, 0, 0, 0, 2, 5, 25, 26, 8, 0, 0, 0, 3, 25, 22, 12, 16, 19, 15, 13, 
    6, 30, 0, 0, 0, 0, 0, 37, 59, 6, 0, 0, 0, 0, 0, 1, 0, 4, 2, 0, 0, 5, 22, 31, 29, 29, 21, 19, 7, 0, 
    2, 18, 0, 0, 0, 0, 0, 6, 31, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 27, 32, 36, 39, 29, 12, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 24, 2, 0, 0, 0, 0, 0, 0, 7, 20, 8, 0, 0, 1, 4, 16, 22, 17, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 21, 10, 9, 11, 17, 16, 3, 0, 6, 23, 29, 27, 9, 3, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 1, 26, 32, 29, 15, 1, 3, 7, 6, 0, 13, 31, 40, 29, 15, 12, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 38, 42, 66, 57, 30, 35, 23, 4, 0, 8, 51, 51, 11, 18, 46, 56, 49, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 9, 0, 0, 12, 52, 44, 10, 1, 0, 3, 6, 0, 0, 11, 40, 51, 59, 64, 50, 29, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 28, 3, 0, 0, 9, 28, 0, 0, 0, 0, 9, 10, 0, 0, 2, 55, 70, 45, 9, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 1, 12, 0, 0, 17, 12, 25, 5, 0, 0, 0, 0, 29, 51, 57, 60, 65, 66, 57, 15, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 1, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 85, 83, 56, 34, 38, 28, 17, 3, 4, 7, 15, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 35, 39, 30, 30, 32, 41, 41, 39, 35, 34, 49, 52, 47, 46, 48, 52, 
    60, 19, 0, 0, 0, 0, 0, 0, 0, 9, 50, 94, 113, 120, 127, 121, 96, 77, 66, 51, 49, 57, 69, 75, 77, 76, 76, 73, 75, 75, 
    104, 98, 46, 3, 0, 0, 0, 0, 30, 89, 111, 97, 97, 98, 98, 100, 91, 81, 84, 85, 82, 83, 86, 85, 79, 74, 77, 80, 82, 84, 
    90, 103, 92, 49, 4, 0, 0, 2, 70, 108, 82, 68, 67, 67, 71, 77, 84, 85, 87, 90, 88, 85, 81, 75, 68, 69, 73, 76, 73, 66, 
    78, 85, 93, 83, 28, 0, 0, 27, 90, 97, 75, 72, 77, 80, 78, 79, 82, 81, 81, 83, 81, 75, 70, 75, 81, 90, 95, 88, 66, 54, 
    91, 87, 86, 83, 63, 11, 0, 30, 78, 73, 78, 76, 76, 83, 82, 78, 77, 77, 78, 82, 86, 90, 88, 87, 97, 106, 101, 84, 72, 83, 
    97, 93, 85, 80, 81, 83, 57, 51, 80, 74, 74, 72, 66, 67, 76, 84, 87, 85, 83, 88, 92, 97, 103, 102, 99, 92, 85, 86, 104, 120, 
    86, 98, 93, 84, 88, 109, 131, 101, 99, 101, 95, 83, 74, 65, 65, 72, 73, 75, 79, 85, 91, 95, 100, 99, 84, 69, 69, 82, 99, 107, 
    83, 95, 99, 87, 84, 90, 111, 116, 95, 105, 107, 106, 107, 96, 83, 73, 68, 64, 61, 65, 77, 89, 89, 80, 62, 50, 52, 77, 88, 91, 
    87, 87, 96, 93, 85, 81, 83, 94, 90, 95, 98, 100, 108, 110, 112, 106, 94, 80, 68, 64, 72, 80, 79, 74, 61, 60, 68, 87, 99, 98, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    75, 76, 71, 65, 69, 69, 68, 65, 64, 67, 72, 75, 73, 68, 65, 61, 61, 71, 76, 78, 80, 81, 81, 73, 68, 62, 57, 53, 48, 45, 
    69, 71, 67, 62, 69, 69, 69, 65, 64, 61, 67, 68, 68, 65, 63, 61, 68, 68, 77, 76, 77, 82, 85, 88, 86, 78, 65, 57, 50, 46, 
    62, 68, 66, 63, 68, 73, 69, 69, 72, 77, 82, 58, 61, 71, 76, 80, 72, 67, 76, 70, 65, 60, 66, 68, 82, 87, 81, 70, 60, 52, 
    70, 82, 79, 70, 71, 73, 69, 69, 80, 138, 139, 83, 76, 90, 85, 73, 61, 84, 96, 98, 89, 77, 62, 57, 68, 75, 90, 86, 69, 54, 
    85, 99, 106, 87, 73, 67, 65, 65, 76, 137, 136, 105, 75, 62, 57, 52, 61, 98, 122, 126, 120, 108, 90, 88, 60, 60, 83, 98, 81, 59, 
    58, 68, 111, 110, 80, 67, 64, 62, 68, 86, 87, 84, 65, 36, 42, 54, 73, 117, 149, 136, 114, 106, 116, 99, 69, 50, 64, 95, 96, 71, 
    25, 31, 91, 103, 82, 69, 68, 63, 68, 60, 76, 96, 86, 63, 74, 82, 84, 125, 167, 153, 104, 96, 108, 94, 73, 48, 51, 80, 99, 84, 
    36, 60, 108, 94, 77, 73, 70, 74, 52, 42, 85, 124, 105, 82, 81, 92, 89, 101, 145, 160, 112, 83, 78, 82, 70, 51, 35, 56, 94, 99, 
    80, 127, 144, 112, 79, 79, 103, 158, 118, 89, 106, 138, 112, 82, 77, 75, 76, 68, 120, 146, 116, 91, 68, 74, 80, 66, 39, 29, 69, 102, 
    132, 187, 175, 124, 82, 67, 146, 235, 234, 162, 146, 141, 112, 88, 77, 67, 57, 58, 138, 156, 131, 113, 79, 92, 93, 80, 53, 26, 39, 78, 
    150, 208, 202, 133, 92, 57, 104, 192, 250, 185, 165, 165, 125, 92, 79, 76, 40, 71, 190, 181, 152, 116, 86, 100, 106, 96, 69, 45, 36, 53, 
    136, 207, 207, 141, 114, 75, 45, 123, 192, 155, 164, 195, 155, 101, 93, 96, 49, 99, 213, 190, 150, 105, 87, 93, 107, 102, 90, 69, 58, 44, 
    136, 212, 177, 123, 125, 101, 43, 94, 145, 139, 170, 211, 195, 139, 119, 115, 70, 131, 211, 187, 133, 97, 81, 78, 89, 98, 103, 88, 81, 56, 
    153, 216, 152, 101, 108, 117, 56, 74, 116, 160, 187, 200, 178, 171, 150, 120, 77, 142, 206, 175, 135, 110, 90, 83, 92, 107, 117, 105, 83, 69, 
    167, 209, 161, 98, 94, 127, 76, 89, 109, 203, 247, 198, 154, 156, 147, 120, 93, 133, 183, 163, 135, 104, 85, 93, 110, 124, 129, 103, 78, 75, 
    176, 208, 192, 113, 108, 136, 112, 86, 114, 217, 239, 196, 158, 126, 124, 111, 98, 137, 164, 160, 151, 112, 76, 85, 110, 119, 110, 84, 82, 75, 
    187, 213, 216, 135, 113, 144, 154, 85, 110, 146, 148, 146, 108, 103, 101, 97, 116, 126, 84, 121, 156, 115, 78, 73, 92, 102, 90, 76, 79, 68, 
    206, 214, 223, 160, 110, 141, 174, 131, 106, 85, 98, 126, 96, 117, 96, 86, 136, 131, 71, 90, 97, 78, 61, 50, 67, 84, 90, 86, 79, 74, 
    219, 213, 220, 181, 117, 127, 157, 158, 133, 81, 99, 118, 122, 163, 121, 78, 120, 147, 140, 112, 73, 62, 51, 77, 86, 104, 104, 92, 83, 81, 
    232, 207, 214, 193, 131, 133, 165, 141, 101, 65, 92, 98, 150, 189, 155, 97, 88, 105, 111, 92, 70, 50, 51, 88, 107, 137, 133, 118, 111, 107, 
    245, 208, 211, 188, 126, 142, 233, 199, 118, 84, 114, 160, 213, 232, 217, 163, 120, 88, 55, 57, 68, 70, 83, 94, 120, 141, 146, 135, 125, 124, 
    266, 234, 218, 181, 120, 170, 275, 281, 241, 183, 182, 222, 241, 244, 231, 186, 154, 119, 93, 89, 104, 119, 131, 133, 142, 150, 160, 149, 140, 140, 
    268, 268, 250, 212, 165, 237, 288, 297, 251, 182, 172, 167, 164, 163, 160, 144, 135, 127, 128, 132, 138, 140, 145, 147, 149, 152, 158, 155, 153, 150, 
    206, 249, 269, 228, 208, 285, 302, 262, 174, 144, 130, 123, 120, 118, 123, 125, 129, 128, 132, 139, 143, 144, 145, 154, 156, 155, 154, 154, 151, 151, 
    155, 194, 238, 215, 240, 300, 288, 189, 141, 138, 134, 135, 131, 129, 129, 127, 127, 127, 132, 138, 142, 147, 155, 167, 169, 171, 168, 166, 170, 181, 
    155, 159, 184, 205, 277, 326, 250, 138, 130, 135, 141, 138, 131, 130, 129, 126, 127, 131, 137, 146, 156, 166, 172, 170, 170, 168, 174, 189, 205, 208, 
    159, 152, 151, 183, 283, 338, 238, 138, 137, 138, 143, 138, 127, 127, 131, 133, 136, 139, 146, 152, 159, 173, 176, 166, 156, 155, 185, 205, 204, 192, 
    158, 154, 152, 157, 233, 300, 232, 156, 151, 150, 157, 151, 140, 131, 126, 128, 135, 141, 148, 150, 153, 160, 161, 158, 153, 169, 186, 183, 161, 160, 
    155, 154, 157, 149, 164, 211, 179, 151, 134, 145, 159, 163, 163, 149, 140, 137, 140, 141, 143, 146, 145, 146, 147, 158, 172, 188, 178, 165, 129, 143, 
    157, 151, 153, 152, 144, 147, 138, 128, 117, 126, 135, 141, 152, 154, 158, 160, 161, 164, 163, 149, 139, 139, 148, 175, 204, 209, 187, 159, 137, 138, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 53, 3, 0, 0, 0, 0, 0, 4, 42, 49, 46, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 67, 74, 53, 32, 25, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 75, 73, 40, 28, 25, 9, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 33, 9, 0, 0, 11, 30, 59, 66, 41, 18, 7, 0, 0, 0, 0, 0, 0, 
    59, 13, 4, 20, 0, 0, 0, 0, 10, 29, 21, 53, 78, 52, 16, 0, 1, 0, 0, 30, 60, 43, 13, 0, 0, 0, 0, 0, 0, 0, 
    100, 74, 82, 70, 0, 0, 0, 58, 157, 162, 113, 96, 101, 55, 27, 2, 0, 0, 0, 30, 76, 68, 38, 0, 0, 0, 0, 0, 0, 0, 
    129, 105, 126, 92, 6, 0, 6, 85, 193, 202, 145, 110, 113, 77, 30, 11, 0, 0, 0, 78, 126, 94, 53, 11, 2, 7, 0, 0, 0, 0, 
    134, 104, 142, 112, 22, 0, 0, 26, 118, 173, 123, 107, 123, 98, 40, 15, 0, 0, 24, 127, 149, 89, 40, 7, 7, 13, 5, 0, 0, 0, 
    123, 97, 158, 123, 21, 0, 0, 0, 52, 98, 81, 105, 144, 127, 68, 43, 25, 11, 51, 141, 137, 76, 29, 5, 3, 0, 4, 5, 0, 0, 
    128, 112, 158, 112, 11, 0, 0, 0, 8, 56, 83, 150, 174, 145, 88, 68, 43, 27, 67, 143, 121, 61, 28, 1, 0, 0, 11, 24, 11, 0, 
    146, 132, 156, 110, 21, 0, 0, 0, 0, 48, 104, 186, 169, 126, 101, 71, 35, 26, 67, 122, 120, 79, 44, 15, 2, 18, 32, 33, 0, 0, 
    169, 151, 162, 126, 55, 15, 6, 0, 0, 71, 173, 198, 155, 89, 67, 47, 22, 8, 43, 93, 89, 61, 26, 6, 5, 25, 34, 6, 0, 0, 
    193, 176, 184, 152, 99, 40, 47, 23, 9, 48, 124, 118, 79, 39, 29, 26, 5, 20, 42, 46, 50, 71, 38, 0, 0, 1, 1, 0, 0, 0, 
    209, 196, 198, 168, 117, 65, 67, 60, 41, 33, 35, 28, 23, 11, 24, 34, 18, 22, 2, 0, 26, 38, 3, 0, 0, 0, 0, 0, 0, 0, 
    206, 199, 197, 176, 132, 83, 82, 94, 62, 38, 11, 13, 34, 32, 58, 67, 36, 32, 32, 26, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    180, 190, 183, 175, 140, 88, 67, 115, 114, 54, 25, 5, 34, 74, 111, 92, 53, 36, 49, 36, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    158, 187, 173, 173, 150, 94, 78, 122, 135, 64, 22, 31, 84, 143, 169, 134, 74, 33, 3, 0, 0, 0, 0, 0, 10, 32, 32, 25, 16, 6, 
    157, 199, 178, 167, 132, 78, 120, 217, 223, 183, 138, 139, 178, 208, 207, 176, 123, 55, 4, 0, 0, 7, 29, 47, 57, 65, 69, 67, 59, 52, 
    168, 204, 190, 172, 134, 114, 175, 278, 308, 254, 176, 138, 143, 150, 142, 118, 92, 62, 43, 39, 48, 59, 72, 82, 85, 89, 96, 95, 89, 86, 
    154, 174, 183, 196, 162, 158, 226, 306, 274, 179, 97, 67, 67, 67, 66, 64, 65, 63, 58, 63, 73, 75, 79, 85, 90, 95, 95, 97, 97, 91, 
    113, 127, 150, 166, 151, 170, 262, 294, 206, 110, 74, 67, 71, 69, 64, 60, 59, 56, 56, 62, 71, 78, 80, 93, 103, 109, 107, 109, 105, 104, 
    110, 101, 117, 122, 140, 200, 282, 240, 137, 75, 79, 82, 79, 70, 63, 58, 54, 55, 60, 68, 78, 88, 101, 114, 120, 119, 114, 112, 125, 145, 
    117, 96, 91, 107, 139, 220, 271, 194, 94, 74, 80, 81, 78, 68, 65, 63, 64, 69, 74, 85, 98, 108, 115, 118, 112, 101, 101, 127, 161, 165, 
    118, 102, 94, 101, 144, 197, 237, 169, 84, 74, 80, 81, 78, 73, 70, 71, 73, 79, 88, 92, 97, 103, 108, 107, 97, 94, 123, 156, 158, 122, 
    124, 105, 102, 100, 117, 153, 157, 124, 72, 70, 78, 85, 88, 84, 75, 68, 74, 84, 92, 94, 96, 96, 91, 86, 91, 117, 143, 147, 118, 86, 
    129, 105, 101, 102, 91, 94, 83, 69, 49, 46, 60, 76, 83, 83, 80, 81, 87, 92, 98, 102, 96, 84, 77, 83, 109, 146, 168, 155, 109, 83, 
    124, 105, 96, 98, 90, 77, 64, 52, 44, 36, 41, 47, 53, 62, 64, 69, 82, 98, 114, 115, 97, 82, 79, 96, 137, 172, 182, 148, 101, 73, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    322, 332, 335, 337, 339, 343, 343, 341, 338, 329, 326, 335, 352, 366, 369, 362, 342, 309, 277, 249, 236, 238, 253, 270, 283, 294, 304, 307, 298, 279, 
    330, 344, 347, 346, 344, 348, 347, 348, 343, 339, 337, 341, 348, 358, 361, 346, 302, 249, 205, 178, 166, 166, 177, 195, 220, 251, 285, 304, 302, 287, 
    337, 354, 361, 356, 352, 350, 351, 349, 345, 353, 353, 351, 333, 322, 302, 263, 208, 180, 159, 146, 131, 131, 137, 140, 162, 197, 240, 276, 291, 287, 
    305, 313, 335, 347, 352, 350, 352, 351, 343, 324, 290, 284, 263, 229, 188, 155, 148, 135, 128, 110, 100, 102, 109, 124, 124, 143, 177, 230, 270, 285, 
    215, 206, 250, 319, 353, 360, 359, 360, 348, 284, 240, 206, 197, 166, 137, 124, 124, 114, 108, 95, 80, 70, 88, 91, 92, 91, 125, 184, 246, 281, 
    143, 130, 186, 282, 347, 364, 365, 359, 341, 290, 247, 215, 197, 172, 137, 115, 98, 92, 97, 105, 96, 85, 77, 76, 71, 64, 90, 145, 211, 264, 
    139, 122, 188, 278, 335, 356, 354, 345, 308, 265, 234, 213, 185, 145, 100, 80, 72, 68, 77, 96, 116, 107, 81, 75, 63, 67, 72, 111, 177, 242, 
    129, 130, 182, 275, 326, 337, 336, 338, 316, 285, 236, 188, 156, 117, 88, 66, 58, 52, 73, 97, 123, 121, 106, 89, 82, 80, 83, 92, 136, 197, 
    102, 98, 163, 241, 307, 304, 296, 272, 286, 250, 215, 162, 140, 122, 101, 79, 55, 71, 101, 130, 147, 134, 120, 101, 91, 88, 87, 87, 105, 151, 
    67, 48, 128, 221, 302, 298, 230, 141, 130, 157, 168, 164, 152, 143, 109, 98, 69, 89, 125, 151, 151, 114, 100, 86, 83, 85, 84, 88, 97, 129, 
    37, 28, 93, 206, 299, 325, 217, 123, 69, 114, 140, 166, 170, 158, 134, 108, 96, 106, 114, 130, 112, 90, 79, 68, 75, 73, 80, 83, 100, 125, 
    44, 40, 74, 162, 256, 325, 275, 174, 106, 119, 152, 168, 174, 169, 148, 121, 103, 105, 91, 105, 88, 85, 73, 64, 59, 63, 72, 84, 102, 141, 
    69, 58, 65, 119, 205, 294, 291, 195, 131, 151, 168, 158, 125, 125, 132, 115, 94, 75, 82, 90, 93, 93, 86, 75, 70, 80, 83, 93, 108, 157, 
    80, 68, 76, 94, 166, 242, 270, 207, 159, 161, 174, 141, 98, 79, 99, 96, 94, 81, 82, 90, 97, 89, 74, 71, 75, 86, 94, 102, 131, 188, 
    78, 74, 87, 83, 126, 174, 231, 205, 167, 133, 122, 92, 87, 71, 72, 83, 101, 117, 119, 114, 96, 93, 75, 60, 57, 64, 84, 118, 178, 231, 
    74, 70, 78, 75, 82, 112, 173, 178, 163, 77, 39, 40, 48, 82, 74, 79, 112, 145, 123, 92, 86, 95, 83, 55, 43, 55, 96, 169, 229, 266, 
    66, 54, 54, 67, 52, 73, 102, 168, 150, 96, 63, 77, 112, 126, 103, 85, 115, 146, 159, 121, 79, 56, 50, 44, 54, 98, 166, 241, 280, 296, 
    59, 46, 42, 62, 57, 54, 58, 105, 126, 123, 116, 105, 142, 148, 130, 92, 86, 128, 178, 142, 90, 57, 45, 69, 103, 169, 230, 271, 290, 293, 
    60, 57, 51, 61, 60, 52, 54, 69, 91, 92, 99, 95, 121, 140, 137, 101, 84, 86, 82, 61, 46, 38, 40, 44, 100, 178, 247, 271, 275, 268, 
    59, 75, 70, 61, 52, 49, 87, 111, 124, 122, 100, 133, 130, 128, 123, 107, 94, 82, 34, 7, 5, 18, 31, 7, 34, 72, 123, 139, 139, 128, 
    31, 71, 77, 61, 52, 70, 102, 155, 163, 157, 110, 75, 40, 26, 15, 13, 27, 36, 38, 13, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 11, 55, 68, 89, 119, 115, 114, 70, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 82, 106, 115, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 50, 82, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 77, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
