library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 1, 0, 
    26, 0, 33, 30, 0, 75, 4, 
    148, 0, 56, 79, 0, 116, 0, 
    192, 61, 56, 120, 52, 88, 0, 
    160, 68, 148, 53, 85, 54, 45, 
    188, 45, 160, 134, 0, 0, 0, 
    45, 250, 36, 0, 0, 0, 21, 
    
    -- channel=1
    0, 61, 0, 0, 0, 0, 41, 
    0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 178, 0, 
    0, 0, 0, 60, 104, 0, 0, 
    0, 0, 62, 8, 10, 10, 0, 
    
    -- channel=2
    0, 0, 17, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 
    0, 0, 11, 9, 0, 0, 53, 
    0, 0, 0, 0, 0, 0, 29, 
    0, 0, 0, 32, 0, 11, 0, 
    0, 0, 0, 0, 12, 52, 64, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    49, 96, 0, 0, 122, 25, 28, 
    17, 154, 92, 0, 73, 0, 0, 
    0, 0, 0, 0, 51, 0, 34, 
    0, 0, 0, 0, 0, 0, 50, 
    0, 5, 59, 14, 0, 37, 109, 
    0, 0, 0, 0, 203, 289, 242, 
    41, 0, 63, 183, 253, 238, 158, 
    
    -- channel=4
    0, 14, 7, 0, 68, 26, 0, 
    54, 86, 98, 0, 112, 4, 0, 
    0, 24, 106, 3, 158, 0, 30, 
    0, 59, 111, 0, 107, 0, 51, 
    35, 121, 59, 41, 0, 5, 60, 
    2, 117, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    68, 16, 87, 85, 146, 54, 68, 
    229, 179, 144, 44, 265, 0, 87, 
    94, 224, 105, 0, 521, 32, 27, 
    63, 243, 250, 0, 252, 0, 46, 
    46, 391, 180, 74, 71, 48, 133, 
    184, 364, 4, 0, 0, 5, 0, 
    167, 82, 0, 0, 0, 7, 52, 
    
    -- channel=6
    48, 35, 23, 159, 126, 81, 114, 
    99, 110, 66, 0, 52, 0, 106, 
    0, 277, 0, 0, 17, 0, 0, 
    0, 40, 84, 0, 50, 0, 0, 
    0, 0, 69, 0, 153, 133, 122, 
    117, 70, 173, 73, 0, 4, 0, 
    73, 179, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    41, 43, 0, 0, 0, 6, 0, 
    206, 152, 210, 166, 166, 208, 187, 
    299, 221, 284, 228, 263, 291, 339, 
    
    -- channel=8
    189, 227, 133, 122, 119, 56, 127, 
    0, 146, 22, 0, 3, 0, 0, 
    0, 14, 23, 0, 0, 0, 0, 
    0, 0, 50, 0, 0, 0, 90, 
    0, 0, 0, 0, 0, 12, 90, 
    0, 0, 0, 3, 0, 8, 0, 
    0, 0, 0, 19, 30, 20, 0, 
    
    -- channel=9
    0, 0, 41, 53, 133, 89, 35, 
    163, 102, 117, 127, 191, 156, 128, 
    208, 213, 245, 268, 289, 235, 141, 
    246, 180, 85, 222, 218, 214, 75, 
    229, 425, 188, 131, 160, 176, 64, 
    186, 320, 390, 109, 127, 64, 69, 
    97, 126, 94, 41, 9, 42, 34, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 47, 10, 41, 37, 0, 
    0, 0, 0, 59, 146, 35, 0, 
    78, 0, 39, 26, 101, 0, 0, 
    134, 106, 113, 0, 0, 0, 0, 
    0, 132, 0, 25, 0, 0, 7, 
    69, 43, 0, 17, 34, 27, 68, 
    
    -- channel=11
    66, 0, 72, 172, 265, 174, 114, 
    149, 133, 189, 75, 0, 0, 54, 
    0, 0, 0, 4, 0, 0, 32, 
    30, 100, 0, 0, 0, 0, 0, 
    0, 112, 127, 42, 68, 201, 75, 
    93, 0, 0, 103, 126, 49, 122, 
    62, 61, 92, 18, 12, 0, 32, 
    
    -- channel=12
    0, 6, 0, 0, 25, 28, 0, 
    0, 8, 101, 0, 0, 22, 19, 
    0, 0, 0, 0, 0, 0, 42, 
    0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 138, 0, 
    0, 0, 0, 144, 155, 126, 142, 
    46, 0, 0, 47, 75, 64, 0, 
    
    -- channel=13
    0, 26, 15, 17, 0, 32, 0, 
    15, 0, 45, 82, 0, 126, 93, 
    130, 16, 120, 213, 18, 163, 89, 
    201, 99, 30, 145, 33, 119, 35, 
    271, 108, 111, 124, 74, 43, 20, 
    140, 117, 79, 71, 0, 0, 8, 
    72, 193, 0, 0, 0, 0, 31, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    6, 0, 0, 173, 124, 75, 98, 
    92, 32, 72, 15, 26, 50, 70, 
    70, 126, 42, 46, 85, 104, 0, 
    53, 41, 24, 83, 57, 94, 0, 
    45, 96, 96, 28, 162, 129, 102, 
    189, 140, 292, 119, 32, 0, 0, 
    64, 205, 54, 19, 2, 23, 58, 
    
    -- channel=16
    170, 191, 134, 136, 79, 109, 147, 
    151, 173, 139, 151, 72, 120, 108, 
    114, 107, 45, 138, 57, 127, 83, 
    39, 174, 46, 118, 83, 103, 133, 
    0, 40, 61, 0, 54, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    20, 81, 12, 0, 0, 0, 0, 
    73, 0, 0, 2, 72, 19, 24, 
    40, 50, 0, 7, 223, 41, 3, 
    0, 0, 0, 0, 58, 0, 73, 
    0, 98, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 19, 0, 
    58, 0, 0, 80, 1, 4, 69, 
    0, 0, 0, 142, 131, 45, 123, 
    83, 97, 0, 0, 0, 0, 0, 
    0, 251, 47, 49, 15, 33, 0, 
    0, 0, 0, 0, 113, 121, 113, 
    61, 0, 0, 47, 57, 39, 102, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    178, 163, 187, 165, 136, 68, 158, 
    80, 189, 137, 60, 51, 0, 33, 
    0, 151, 84, 0, 50, 0, 0, 
    0, 98, 80, 0, 17, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    49, 28, 7, 62, 11, 0, 37, 
    46, 14, 45, 0, 91, 27, 49, 
    0, 211, 57, 0, 87, 5, 0, 
    0, 8, 175, 77, 158, 49, 23, 
    29, 29, 34, 0, 131, 67, 0, 
    139, 112, 157, 113, 0, 0, 0, 
    98, 304, 13, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 
    53, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 52, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 74, 0, 0, 0, 0, 
    
    -- channel=23
    17, 134, 52, 0, 0, 49, 0, 
    0, 6, 69, 82, 0, 106, 0, 
    97, 0, 0, 165, 0, 85, 33, 
    213, 0, 0, 0, 0, 0, 0, 
    123, 0, 35, 55, 0, 0, 0, 
    0, 0, 0, 0, 179, 201, 215, 
    0, 0, 114, 190, 217, 173, 210, 
    
    -- channel=24
    363, 339, 298, 304, 100, 74, 235, 
    94, 267, 90, 63, 0, 75, 89, 
    72, 267, 67, 24, 0, 92, 0, 
    0, 9, 0, 84, 22, 114, 48, 
    0, 0, 29, 0, 84, 23, 30, 
    7, 0, 183, 51, 8, 0, 0, 
    0, 40, 65, 28, 12, 40, 2, 
    
    -- channel=25
    93, 70, 122, 68, 46, 95, 103, 
    203, 111, 140, 73, 92, 57, 104, 
    171, 161, 178, 57, 167, 70, 37, 
    115, 167, 192, 0, 144, 28, 55, 
    58, 127, 172, 158, 118, 50, 172, 
    167, 285, 120, 43, 0, 41, 34, 
    123, 182, 0, 0, 6, 7, 47, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 19, 19, 108, 20, 
    88, 0, 112, 223, 347, 442, 447, 
    371, 127, 310, 415, 452, 480, 474, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    91, 0, 145, 65, 0, 0, 33, 
    179, 0, 0, 0, 0, 0, 12, 
    239, 114, 0, 147, 0, 0, 15, 
    118, 0, 0, 36, 125, 144, 175, 
    0, 139, 90, 142, 154, 139, 171, 
    
    -- channel=28
    15, 1, 41, 33, 80, 50, 41, 
    27, 34, 72, 96, 93, 60, 84, 
    0, 60, 53, 49, 77, 57, 84, 
    0, 80, 68, 22, 59, 55, 79, 
    0, 26, 58, 29, 80, 60, 52, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 
    41, 33, 86, 0, 10, 0, 0, 
    0, 0, 30, 0, 0, 0, 50, 
    0, 0, 0, 18, 0, 0, 0, 
    0, 234, 92, 0, 0, 141, 82, 
    0, 0, 0, 27, 71, 62, 73, 
    
    -- channel=30
    177, 162, 210, 287, 198, 216, 209, 
    185, 197, 257, 206, 8, 121, 85, 
    144, 148, 63, 197, 0, 172, 46, 
    167, 183, 67, 181, 0, 84, 9, 
    63, 62, 141, 56, 145, 40, 38, 
    0, 0, 70, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 2, 66, 20, 
    50, 0, 0, 8, 0, 81, 38, 
    78, 18, 0, 151, 0, 47, 19, 
    59, 0, 7, 0, 144, 102, 0, 
    58, 0, 173, 140, 47, 28, 40, 
    59, 91, 105, 102, 70, 117, 39, 
    
    
    others => 0);
end gold_package;
