library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    339, 337, 348, 352, 355, 322, 362, 390, 368, 304, 254, 262, 281, 302, 312, 
    353, 356, 360, 363, 357, 294, 317, 310, 241, 141, 76, 96, 152, 248, 302, 
    244, 288, 365, 373, 377, 295, 209, 136, 86, 49, 20, 27, 49, 126, 241, 
    79, 153, 340, 365, 315, 226, 127, 60, 46, 64, 64, 60, 40, 50, 177, 
    1, 64, 285, 279, 133, 99, 62, 46, 37, 57, 61, 53, 48, 39, 101, 
    0, 23, 257, 258, 61, 65, 66, 61, 41, 55, 49, 39, 44, 35, 31, 
    0, 1, 183, 288, 126, 99, 70, 64, 38, 44, 30, 31, 33, 34, 54, 
    0, 0, 50, 193, 149, 75, 46, 52, 63, 102, 53, 34, 27, 61, 153, 
    0, 0, 0, 39, 121, 64, 75, 66, 61, 145, 87, 51, 50, 126, 251, 
    4, 0, 0, 0, 16, 58, 55, 36, 37, 88, 48, 17, 43, 219, 280, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
