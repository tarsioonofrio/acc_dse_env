library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    145, 219, 247, 
    330, 242, 157, 
    230, 201, 143, 
    
    -- channel=1
    203, 101, 44, 
    207, 95, 66, 
    44, 67, 0, 
    
    -- channel=2
    96, 0, 173, 
    36, 73, 54, 
    0, 0, 0, 
    
    -- channel=3
    463, 333, 345, 
    389, 326, 255, 
    55, 0, 0, 
    
    -- channel=4
    94, 0, 0, 
    0, 0, 0, 
    0, 0, 108, 
    
    -- channel=5
    11, 36, 11, 
    176, 12, 79, 
    0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 
    2, 0, 0, 
    340, 488, 518, 
    
    -- channel=8
    60, 143, 110, 
    440, 183, 143, 
    58, 0, 0, 
    
    -- channel=9
    219, 257, 296, 
    231, 147, 65, 
    182, 159, 281, 
    
    -- channel=10
    0, 0, 0, 
    0, 0, 0, 
    0, 131, 100, 
    
    -- channel=11
    178, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=12
    105, 0, 0, 
    0, 0, 16, 
    0, 155, 281, 
    
    -- channel=13
    191, 178, 210, 
    151, 253, 210, 
    65, 52, 76, 
    
    -- channel=14
    0, 0, 0, 
    0, 0, 15, 
    0, 0, 0, 
    
    -- channel=15
    355, 276, 220, 
    0, 0, 33, 
    0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 
    32, 0, 0, 
    0, 140, 119, 
    
    -- channel=17
    24, 0, 48, 
    401, 192, 179, 
    400, 227, 164, 
    
    -- channel=18
    46, 131, 63, 
    0, 94, 199, 
    208, 204, 183, 
    
    -- channel=19
    224, 0, 0, 
    0, 0, 0, 
    0, 173, 162, 
    
    -- channel=20
    61, 38, 20, 
    0, 0, 0, 
    85, 22, 232, 
    
    -- channel=21
    0, 43, 28, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=23
    0, 0, 17, 
    0, 9, 41, 
    44, 0, 6, 
    
    -- channel=24
    26, 248, 109, 
    0, 80, 53, 
    0, 0, 0, 
    
    -- channel=25
    66, 22, 91, 
    67, 196, 244, 
    139, 58, 51, 
    
    -- channel=26
    190, 258, 303, 
    448, 408, 291, 
    453, 356, 311, 
    
    -- channel=27
    246, 131, 197, 
    288, 213, 205, 
    370, 159, 167, 
    
    -- channel=28
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=29
    124, 0, 5, 
    320, 118, 61, 
    280, 446, 340, 
    
    -- channel=30
    110, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
