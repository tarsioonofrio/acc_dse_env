-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        INPUT_SIZE : integer := 8;
        ADDRESS_SIZE    : integer := 12;
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(ADDRESS_SIZE-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(2-1 downto 0);
    signal bram_addr     : std_logic_vector(10-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(10-1 downto 0);
          

    MEM_IFMAP_LAYER0_ENTITY0 : if BRAM_NAME = "ifmap_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009e009f00a500a600a0009c00a2009f009e009f00a100a000a100a600a900aa",
            INIT_01 => X"00a700a200a000a0009c0095009600940095008f008c008d008f0089007e0074",
            INIT_02 => X"00980097009f00a600a200a000a400a200a3009c009b009f00a300aa00ab00ab",
            INIT_03 => X"00a900a0009a00970091008b008c008d009500930091008e008f0088007d0077",
            INIT_04 => X"00970097009e00a700a000a300a500a500a300a2009e009d00a100a600a700a9",
            INIT_05 => X"00aa009f00910079006e00620065007200780086008f008c008e008b00820078",
            INIT_06 => X"009b009b00a000ae00a700a700a900a900a500a500a700bf00b1009d00a200a4",
            INIT_07 => X"009e0095006800670062005c0050004a0056005300710084008c008c0088007f",
            INIT_08 => X"009b009c00a100aa00a900a300a900a600a400a400ad00f600c300970092008e",
            INIT_09 => X"006f004e005500710070006a0061005d004a0054005500690080008a00850081",
            INIT_0A => X"009400850082009300a100a500a700a700a300a500a300b4009d008000610042",
            INIT_0B => X"0045004200590076007a00770072005e0063005b003a0043006c008c008a0086",
            INIT_0C => X"007f006d002f0058009900aa00a800aa00a900a600a400930081007f00640044",
            INIT_0D => X"004e0048005300840092007c0069006b00730055003f002e004f0084008d0086",
            INIT_0E => X"00830063002a0046008f00a700a500a800ab00a1008c00780082009000740058",
            INIT_0F => X"005b0055004d007c00a300880066006a00640055003600310039006b008a0088",
            INIT_10 => X"00aa00670036007c009900a100a300a600a500ae0071007d009d009c00790056",
            INIT_11 => X"0052005400500051008a00920071005700530056004700380028004a00850089",
            INIT_12 => X"00b40086005e009a00ae009e009c009900cf00ed00cf009c00ae0094007d005d",
            INIT_13 => X"0056004a003b004c0089008f0085006a005600570054004b00320028005f0084",
            INIT_14 => X"00b7006c008e00a500b1009b009f007a00d500ed00dc00a400b7009c007d0078",
            INIT_15 => X"004e0050002d005b00af009d009b006b005700670058004e003b0029003b0068",
            INIT_16 => X"00bc0064008700aa00bb00a600ad0086007500c200c700aa00b900bd00860075",
            INIT_17 => X"006600540026007d00d200a00092005d0053005e0068005500490037003e004c",
            INIT_18 => X"00bd005a007f00af00ae00a600b2009f006100a800a8008900ba00d800a0007b",
            INIT_19 => X"007800730032009600c2009b007b005b00540054005f005600540049004f0049",
            INIT_1A => X"00bd005d009800b90077008800ad00a700670093009100a700bd00e200b4008d",
            INIT_1B => X"007e00750047009a00ba00950072005700500048005000630064005a0061005e",
            INIT_1C => X"00c2006c00a800ba00690063009c00a700640073008a00c600be00ac0091009a",
            INIT_1D => X"009200670047009800b300890082006e0055005b005f006d0073006400610075",
            INIT_1E => X"00c5008400ac00b80082004e008c009b00730082008f00e600f2009100870083",
            INIT_1F => X"0079006c005f009000a800980070005700470057006900700078006700790088",
            INIT_20 => X"00cb009200a800bf00a8004e007e008a008a0060009a00ad00a2008c00710071",
            INIT_21 => X"00650069007000ab009c00940087006d004e004f005e0065006b007d00970090",
            INIT_22 => X"00d600a300a400b700b0005e0060009c0094006a008100760072007400660073",
            INIT_23 => X"0056006500900076004400800085004b003c003a004700660074008f0096008c",
            INIT_24 => X"00d400b200a700ad00b0007c0056008d009900870068004d0086007c00810093",
            INIT_25 => X"0055005c009600840075006b004b0040002c004100560085009b00a0009a0097",
            INIT_26 => X"00c700bb00ab00ae00b1009000560077007a0089009000460081006c009100b8",
            INIT_27 => X"00740049008300890086005900330034002f005a007900a300ab00a4009e0095",
            INIT_28 => X"00a500c300b300b100b500980063008300ab0067005d0050005d007a00b200bf",
            INIT_29 => X"0096006400590057003c002e00260018002e003c006c009000900080007f0078",
            INIT_2A => X"007500c300b100b200b5008a0053009600f500db00850086009500b000be00c2",
            INIT_2B => X"00a8007d006e003d002300220031003a003d003a00450048004e0045003b0037",
            INIT_2C => X"004f00af00ae00b000b1008c006d00d300fd00fc00d0007c0072007c0074007a",
            INIT_2D => X"006800440044003c003400320033003800380033002b0033003b0030002b002a",
            INIT_2E => X"00290060009000a800b200a500a500f600fd00e3006e003c0035003100310030",
            INIT_2F => X"002d002a002e002a0026002e002e002b002a002e002e0032003700350033002d",
            INIT_30 => X"001d001d003b008300a6008400c200fe00f1008d003d00320032003300310032",
            INIT_31 => X"002f002a00270022002300270026002a002d0038003e003b00380032002e0033",
            INIT_32 => X"0030001e002200490080008000d7010000bb00420036003200340034002e002d",
            INIT_33 => X"002b00290024002700280028002b002e003b003e0040003b0036003200460053",
            INIT_34 => X"00340023001f00290042008000e000f0007c003a003100380036002c002c002f",
            INIT_35 => X"002e002b002b002c002c002d0036003a0036002e002b0024003300490055004c",
            INIT_36 => X"00320023001d0023002c004e00ca00d30061004100360030003a00300028002d",
            INIT_37 => X"002f0030002f002e0033002700270030002f0027001c002800430043002e0033",
            INIT_38 => X"00320023002000210029002e006800aa0040003600340035003d003a0036002d",
            INIT_39 => X"002a0029002e0031002e002a0028002700250028002c003f002f001f000f0033",
            INIT_3A => X"0044002a001f00260025002b002a00470031001f001b002600310038003a0035",
            INIT_3B => X"0038003c003900350032002d00270021002a003e004f004900380026000d0028",
            INIT_3C => X"003d00310023002b0027002a002c0028002a001b0017001e001b001d0024002f",
            INIT_3D => X"0038003e0042004b00450031002b002b003c0055006d005d003c001a001d0014",
            INIT_3E => X"00360038002d002b00280028002800260024001a0016001d0019001d00130012",
            INIT_3F => X"0020002f003d004a004200350034002d00430059006900590030001800220015",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY1 : if BRAM_NAME = "ifmap_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0070006f007400760070006d00730071006f00710074006f006f007500750077",
            INIT_01 => X"00750071006f0070006d006b006b006a006b0065006200610061005f005b0055",
            INIT_02 => X"0070006e0072007400700071007500720074006e006f006e0071007700750073",
            INIT_03 => X"0073006f00700073006e00680066006400690066006600610062005f005b0058",
            INIT_04 => X"006e006d006f006f006a007300750075007300730072006d006f007300720071",
            INIT_05 => X"00740072006f0060005a004e004d0055005600600067006300630062005f0059",
            INIT_06 => X"006b006e006d0070006e00750078007700730075007b00920082006f00730072",
            INIT_07 => X"0070006f00500057005a005a004b003f0046003e00550062006600650063005e",
            INIT_08 => X"006b007200730072007200710078007400710074008000d6009c0072006f006c",
            INIT_09 => X"0050003500450067006e00720066005e0048004e0049005300600065005e005d",
            INIT_0A => X"006d0068006400700073007100740073006f00740076008a007a0066004b0032",
            INIT_0B => X"003a0038005300710079007a007400600064005b003a003a005400690062005f",
            INIT_0C => X"0064005f0025004a0075007600730076007500740078006b0062006c00570043",
            INIT_0D => X"0053004b00540082008e007600630066006f00530047002f003d00620063005d",
            INIT_0E => X"00730060002b0040006f00750072007400770071006d005e006e0083006a0057",
            INIT_0F => X"005f0058004d00760099007c005d0062005d0051003c0035002f005300670061",
            INIT_10 => X"00a10069003a0079007c00710075007a0079008700590069008d008f006f0050",
            INIT_11 => X"00510055004e0047007d00870067004f004d0052004900390023003b006a0067",
            INIT_12 => X"00b0008b0064009a009500740074007600b400d600b4008300990083006e0055",
            INIT_13 => X"0054004a00390044007d0085007c0062005100550055004c0031001e004b0067",
            INIT_14 => X"00b70074009700a9009c00700076005900c500e000bf0087009f0089006c006f",
            INIT_15 => X"004c0050002c005500a5009300930064005300660058004f003b0024002e0051",
            INIT_16 => X"00bf006c009000af00a70078007b005d005f00b600ab008e00a100ab0077006b",
            INIT_17 => X"006200540026007900c90098008b00590050005d00680057004b003500370038",
            INIT_18 => X"00c20060008600b4009c007b007b006d0044009a0090007200a600ca00950071",
            INIT_19 => X"007200720032009300bb00950076005800530054005f005700570049004a0037",
            INIT_1A => X"00c0005f009a00bc006e006a007c007400480084007d009500ae00d800ac0083",
            INIT_1B => X"007500720047009800b50090006e005500500049005000640065005800590049",
            INIT_1C => X"00c4006b00a700ba006d00590077007a004a006a007b00b900b400a5008c008f",
            INIT_1D => X"008800640047009800af00850080006d0056005d0060006e007400600055005f",
            INIT_1E => X"00c5008100a700b2008900530078007d005e0078008300dd00ec008a00820079",
            INIT_1F => X"0070006800580086009f0093006c0055004800580068006d006e005600600068",
            INIT_20 => X"00cb009200a400b600aa0056007d007e00790050008f00a300980084006a006a",
            INIT_21 => X"00650065005a008f008a008d00820069004c004f005d005b00530058006c0068",
            INIT_22 => X"00d700a600a700b800b60066006000950089005d0074006900660069005b006e",
            INIT_23 => X"005b00670080006000380078007e0045003800380046005d005e00700074006e",
            INIT_24 => X"00d300b800af00b500b800830058008b00940080005a00400079006f0075008f",
            INIT_25 => X"005c0060008b0075006d00630044003b0029003e00450069007700780073006f",
            INIT_26 => X"00c000bd00b000b300b60095005a0079007c00880086003b00760061008600b0",
            INIT_27 => X"0076004b0077007c00810056003100330031005a005b007600790071006f006b",
            INIT_28 => X"009c00c100b200ad00b5009d0067008700af0069005a004d005a007600ad00b6",
            INIT_29 => X"00940064004e004d003d0034002e0021003900470064007d007b006d00710069",
            INIT_2A => X"007800c800b200a900b300900057009900f700de008c008d009c00b600c400c0",
            INIT_2B => X"00ac0085006d003e0031003600460051005500540063006500680060005c005a",
            INIT_2C => X"006900c500b700ac00b10092007000d300fc00fd00e0008f0084008d00850085",
            INIT_2D => X"007c005d00570052005400540055005d005e005b00600068006c00610061005f",
            INIT_2E => X"0059008900a800ae00b600aa00a600f500fb00e7008800580050004c004b0048",
            INIT_2F => X"004f0051005100520056005a005900570059005d005e00600060005e005f005a",
            INIT_30 => X"005b00570066009900b3008800bd00fa00f5009f005e00540054005500530054",
            INIT_31 => X"005600540052004f0053005600550059005c00670067006500660063005e0067",
            INIT_32 => X"006f005e0055006a0094008800d500fd00c6005d005b0058005a005a00530052",
            INIT_33 => X"005200510050005300560059005c005f006c006e006d006c006c0069007b0089",
            INIT_34 => X"0072006300560053005f009100e500f5008f005c0057005e005c005200520053",
            INIT_35 => X"0054005300560058005a0061006a006e00690061005f005b006c0082008a007d",
            INIT_36 => X"006e0062005900560053006a00db00e4007e0068005e00570061005700500052",
            INIT_37 => X"00540057005900590061005c005d00660065005d005500650081007e00620060",
            INIT_38 => X"006c0061005c005800580054008500c500640061005e005f0067006400600053",
            INIT_39 => X"004f00500058005c005c005f005d005c005a005d0066007d006e005a003c005d",
            INIT_3A => X"007c00640058005b00570059004f006b0059004d00470052005d00640066005c",
            INIT_3B => X"005e006300630061005f005e00580053005b0070008400830074006100400055",
            INIT_3C => X"007400660055005b005a005c00580051005500480043004a0047004900500056",
            INIT_3D => X"005f0065006d00770071005f0058005800690082009c00910073005200520040",
            INIT_3E => X"006b0069005900560059005c00570051004f00450042004900450049003f003a",
            INIT_3F => X"0046005700680077006f0060005f0057006d0083009200870063004d00540043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY1;


    MEM_IFMAP_LAYER0_ENTITY2 : if BRAM_NAME = "ifmap_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0031002f00330035002e0029002f002d002c00290029003400310029002d002c",
            INIT_01 => X"002800260027002b002c002d002d002b002c0027002b00290026002400240021",
            INIT_02 => X"00330028002d00380031002b002f002d002e0026002900360034002900280021",
            INIT_03 => X"001e00210029003200350037003400300032002e002d00260022001f00200022",
            INIT_04 => X"002f002100240030002a002c002d002d002b002b003000390033002600250023",
            INIT_05 => X"0027002f0036003100340032002f003200300037003300270023002200220021",
            INIT_06 => X"00280020001f002c002b002e00300030002c002d0039005f004b0029002f0036",
            INIT_07 => X"003a0043002f0041004c00540042003200340027002d002e002b002700270024",
            INIT_08 => X"002900300031002f002b0028002f002c0029002a003b00a4006b0038003c0047",
            INIT_09 => X"0032001f00380062006f00760069005d00430046002f002d0030002e00240024",
            INIT_0A => X"0036004000390035002c00270029002900250027002a0055004e003a002b001f",
            INIT_0B => X"002b002d004c006e0078007a0074006000610056002f00250031003a002c0028",
            INIT_0C => X"003900500011001c0030002b0028002b002a002500270034003b004b00460039",
            INIT_0D => X"00480040004a00790084006c005a005e0067004d004500270024003a00300027",
            INIT_0E => X"005a005c002600290038002a002400270031003300330031004d006b005d004f",
            INIT_0F => X"005800520045006b008c0070005100580054004a003a00310020003200330027",
            INIT_10 => X"00900069003b00710052002b002900320042005f003b004e007900800065004a",
            INIT_11 => X"004d00520049003d0070007b005d00460045004c00430035001b0023003b002d",
            INIT_12 => X"00a3008f0069009500700033002f003c009200c600a600770091007d006b004f",
            INIT_13 => X"004f00470035003a0070007a00720059004a004e004e0047002b000f002c0039",
            INIT_14 => X"00af007a009e00a8007a00320033002f00b300e200bc0083009b008400680068",
            INIT_15 => X"0045004d0028004d009a0089008a005c004d0060004f0049003b0021001f002e",
            INIT_16 => X"00bd0074009900b20088003b0037002c005000bc00a400850097009f006a005f",
            INIT_17 => X"0059004f0022007100c0008e00820052004b0058005e0051004e00370030001a",
            INIT_18 => X"00c20069009000b9008500440035002f002c0098007e005e009400b700810062",
            INIT_19 => X"0069006d002f008c00b2008c006f0053004f0050005500510059004900400018",
            INIT_1A => X"00c1006700a300c000620042003a0032002700780067007f009b00c8009d0075",
            INIT_1B => X"006b006d0044009300ae008800680050004c00460048005e0063005100450022",
            INIT_1C => X"00c4007000ac00bc006d0043003e003700220058006700a900a9009f008c0086",
            INIT_1D => X"007d005f0046009500aa007f007a00690053005b005a0068006f00500035002f",
            INIT_1E => X"00c5008800ae00b5008e004d0058004d0034005d007400d300e6008900820070",
            INIT_1F => X"0065005f004b00760092008a006500500044005700630063005d003600300030",
            INIT_20 => X"00cc00a000b200bc00ac005a007e0071005200250085009b008d00750058005a",
            INIT_21 => X"005c0057003a0068006d007e007600610048004d005e00520037002d0037002e",
            INIT_22 => X"00d700b400b800c200ba006900660091006f003d0069005f0059005900490062",
            INIT_23 => X"0058005f00660040002000690073003d003300350041004e0040004400400036",
            INIT_24 => X"00cd00c000bd00c100bc00850060008f008d006f00500037006c006000640085",
            INIT_25 => X"005d005d0078005d005c0056003a00340027003c0028003b003e0036002d002e",
            INIT_26 => X"00b400bb00b500b900b800980063008400820087007e0033006c0056007b00a8",
            INIT_27 => X"00760049006700690076004e002c00320034005d003c0044004000340032002e",
            INIT_28 => X"009200bb00af00ac00b400a0006f009200b9006f005700490056007400ad00b1",
            INIT_29 => X"009400650042003f003900360033002900450053004b0052004c003d0045003f",
            INIT_2A => X"007c00c800b000a800b30093005b009f00fa00e10090009300a400c000d000c5",
            INIT_2B => X"00b5008f006d003e003a004400570066006e006f007a00770078007000700073",
            INIT_2C => X"008500d500c000b100b60096007100d100f700fc00e8009d009500a2009c0098",
            INIT_2D => X"0094007700680065006f006e0073007d008300820087008d008e008400890084",
            INIT_2E => X"008700a800bc00bc00c000ae00a400ed00f100e40099006f00690069006b0065",
            INIT_2F => X"0073007800710074007d007d007e00800084008b0089008900870086008b0085",
            INIT_30 => X"008d0082008600b000bf008900b500f200f500af007f00760077007900780074",
            INIT_31 => X"00750075007300710078007d007d008200860091008e008e00920090008c0095",
            INIT_32 => X"00a2008c007c008800a7008f00d100f900cd00760080007d007f007f00790073",
            INIT_33 => X"0071007000710075007b00830086008a0096009800930095009a009800a700b6",
            INIT_34 => X"00a500930082007a007e00a400ea00f700990072007b00830081007700770077",
            INIT_35 => X"00770077007b007f0083008d0096009a0096008d008c008a009e00b200b600a9",
            INIT_36 => X"00a20095008a0085007e008a00e900ea008c007e0081007c0085007b00740077",
            INIT_37 => X"007a007e00820084008c008a008b00940093008b0085009900b600b0008e008b",
            INIT_38 => X"00a10093008f008d008a007d009f00d30077007900800082008b008700830078",
            INIT_39 => X"00760078008200870088008b008a00880087008a009700b200a4008c00670088",
            INIT_3A => X"00b1009400890092008b00840071008500720069006900750080008700890080",
            INIT_3B => X"00830089008b008a008900880083007d0085009a00b300b500a80092006c007f",
            INIT_3C => X"00a800940084008f008b0086007d0070007300680066006d006a006c00730078",
            INIT_3D => X"008000870090009c00980086007f007f009000aa00c500be00a40082007e006b",
            INIT_3E => X"00a000950084008600860084007b0073007200690065006c0068006c00620059",
            INIT_3F => X"0064007600890098009100830082007b009100a700b600af0091007c0081006e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY2;


    MEM_IFMAP_LAYER0_ENTITY3 : if BRAM_NAME = "ifmap_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00eb00e700e800e800e800e800e800e800e800e800e900e900e900e900e900e9",
            INIT_01 => X"00e900e800e700e600e800e800e800e900e800e900e800e800e800e900e900e8",
            INIT_02 => X"00ee00eb00eb00eb00eb00eb00eb00eb00eb00eb00ec00ec00ec00ec00ec00ec",
            INIT_03 => X"00ed00ec00ec00ea00ea00ea00eb00ec00ec00ec00eb00eb00eb00ec00ec00eb",
            INIT_04 => X"00ed00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00eb00eb",
            INIT_05 => X"00ec00ec00eb00ea00e300e700e700ea00ea00ea00ea00ea00ea00eb00eb00ea",
            INIT_06 => X"00ee00eb00eb00eb00eb00eb00eb00eb00ea00ea00ea00ea00ea00ea00eb00eb",
            INIT_07 => X"00e900e800e400df00ba00d100cf00e400ec00ea00ea00ea00ea00eb00eb00eb",
            INIT_08 => X"00ed00ea00eb00eb00eb00eb00eb00eb00ea00ea00eb00eb00ea00ea00eb00eb",
            INIT_09 => X"00ec00e900db00cb00a300c300d600e600ed00eb00eb00eb00eb00ec00ec00ec",
            INIT_0A => X"00ef00ec00ec00ec00ec00ec00eb00eb00ea00eb00ed00ed00ea00e800eb00e5",
            INIT_0B => X"00d000c200b900ae00a500b800cf00e200ec00ec00ec00ec00ec00ed00ed00ed",
            INIT_0C => X"00e400e400e800e700ea00ed00ed00ec00ed00ed00ef00ef00e100e000e900dd",
            INIT_0D => X"00b700a1009f009a0090008f009c00c600e900ec00eb00eb00eb00ec00ed00ef",
            INIT_0E => X"00d400e000e600e300e500ea00ed00ee00ef00ef00ef00f000c900db00e900d6",
            INIT_0F => X"00c100b900b800ad00a5009f00a200ba00e500ea00e900e900ea00ec00ed00ee",
            INIT_10 => X"00d800dd00e100e100e300e700ec00ee00ee00ee00ed00ef00c500dc00e900e6",
            INIT_11 => X"00d100d100db00d000d100d200d900da00e100e400e400e600e600eb00ed00ee",
            INIT_12 => X"00760077007c008800ac00e100eb00ed00ec00eb00eb00e900d600e200e800ec",
            INIT_13 => X"00e400e300e700e100e100d900c900b900ac00a700a700ba00df00eb00ec00ee",
            INIT_14 => X"006d0067006c006f009200de00e300e500ec00ea00e700e600e500e700e800e6",
            INIT_15 => X"00e700e700e500df00bf00a400920089008600800079009500d800ea00eb00ed",
            INIT_16 => X"00c300bc00c700c800d100df00d500d300d800dc00db00d200d100d300d800dc",
            INIT_17 => X"00e100e200e100da00b700af00b500b200ba00aa008e00b900db00e700ea00ec",
            INIT_18 => X"00c100bf00ca00d600df00d600cb00ab00b100cf00ae0062005d0065006f007a",
            INIT_19 => X"0089009900ca00df00da00dc00df00d900dd00d400c400de00db00dd00e800eb",
            INIT_1A => X"0071006f0071007d008a00aa00bf00be00d000d8009e0036002d003100350042",
            INIT_1B => X"0066009f00dd00ea00e900e300df00cf00ca00d300d400c700b300bc00d300dd",
            INIT_1C => X"003d0045003f0044007b008b009700c300d600ce00a30067005f0065008a00b5",
            INIT_1D => X"00cf00dd00db00cd00b7009e00930083007d0082008800850080008a00b600c5",
            INIT_1E => X"0028003a0055007f00840060007700a300ad00b800b600b500b700c600da00c8",
            INIT_1F => X"00ae009f0091008400740062005e00630069006b007a008a0096009d00bc00b9",
            INIT_20 => X"000d001a008600ce008a0076008d00ac00b500cf00dc00e400e000e600e200b0",
            INIT_21 => X"0090008a008e0091009a00950095009a009d00a000ad00bb00be00b200a5009d",
            INIT_22 => X"0005003a00c800e100c500c700d400e200e500e900e800e600d100df00dd00d2",
            INIT_23 => X"00c600b400c100bc00bd00c200c000b800ac00ab00a10090008800830080008a",
            INIT_24 => X"0027009100be00ba00b800c000c200c200c200bf00c000be00b100b4009a0093",
            INIT_25 => X"0091009c0092007100720084007e006f005c005b005d005e0069007900810081",
            INIT_26 => X"007a00a2008f008900830080007f008200830080007f00810081007c00680064",
            INIT_27 => X"006600760070005e005e005e0057005300500053005d0065006c007300790082",
            INIT_28 => X"0049004c004d0050005400570057005a005e0066006b00710073007600760078",
            INIT_29 => X"0073006e006a0064005f0055004f00500050004d00500052005c0071007d0088",
            INIT_2A => X"000d0003000900120012001500140016001a0022002a00300034003c00420046",
            INIT_2B => X"004700480043003c003700350035003900390039004800570068007800820089",
            INIT_2C => X"0024000b00080020002400160008000300010000000000000006000500010003",
            INIT_2D => X"000d00180015001500150016001e0027003900550071007b0074007a00860099",
            INIT_2E => X"0023001a000d001b004700460031001b000f00050002000000110039001f000a",
            INIT_2F => X"000400040007000e00190029003e0056007a00900084007200750084009200ac",
            INIT_30 => X"0010000d00040003002d00410036002400120004000200000007007600a10083",
            INIT_31 => X"007000690069006d0076008a009a0097007f0069006a00780081008e00a400b8",
            INIT_32 => X"0028000c00000000000c001e0020001500070002000200030000004400b600cd",
            INIT_33 => X"00c400c200c300bb00ac0096007b0067005f0068007a00810084009800ab00b9",
            INIT_34 => X"0045001a000100010004000c0012000c000400020002000400010020009900cb",
            INIT_35 => X"00c300bf00b3009b0077005b0051005e0075007d007d0081009000a200ad00b8",
            INIT_36 => X"0053002f00010002000200050007000400010001000100030001001b008e00cd",
            INIT_37 => X"00c600a900790055004a0055006600790080007a00790084009300a500b000ba",
            INIT_38 => X"005c003600060003000200010001000100010001000100010000000f0066009d",
            INIT_39 => X"0075004a0038004a00630073007a007c007b007d00800088009400a200b100bc",
            INIT_3A => X"0057002b0013000b0008000500020002000300030003000200000004002a0047",
            INIT_3B => X"003500390050007100840086007b007400780083008b008f009c00a900b600bc",
            INIT_3C => X"0052002e0024001f001b00160011001000120013001400130013001700250040",
            INIT_3D => X"0057006800740080008b008300750073007b0083008b0094009f00ae00b900bb",
            INIT_3E => X"0055003e003a00370033002f002e00300031003300350037003b004400510068",
            INIT_3F => X"0074007f0085007f007f00760072007a00810088008d0095009e00a800b400ba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY3;


    MEM_IFMAP_LAYER0_ENTITY4 : if BRAM_NAME = "ifmap_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00eb00e700e800e800e800e800e800e800e800e800e900e900e900e900e900e8",
            INIT_01 => X"00e700e700e900e900e800e700e800e900e900e900e800e800e800e900e900e8",
            INIT_02 => X"00ee00eb00eb00eb00eb00eb00eb00eb00eb00eb00ec00ec00ec00ec00ec00ec",
            INIT_03 => X"00ea00ea00ec00ec00eb00ea00ec00ec00ec00ec00eb00eb00eb00ec00ec00eb",
            INIT_04 => X"00ed00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00eb00ea",
            INIT_05 => X"00e900ea00eb00eb00e600eb00e900ea00ea00ea00ea00ea00ea00eb00eb00ea",
            INIT_06 => X"00ee00eb00eb00eb00eb00eb00eb00eb00ea00ea00ea00ea00ea00ea00eb00eb",
            INIT_07 => X"00e900e800e600e200c000d800d200e400eb00ea00ea00ea00ea00eb00eb00eb",
            INIT_08 => X"00ed00ea00eb00eb00eb00eb00eb00eb00ea00ea00eb00eb00ea00ea00eb00eb",
            INIT_09 => X"00ee00ed00e100d200ac00cd00da00e500eb00eb00eb00eb00ec00ec00ec00ec",
            INIT_0A => X"00ef00eb00eb00eb00eb00eb00ec00eb00ea00eb00ec00ec00eb00e900ed00e7",
            INIT_0B => X"00d800cd00c600bc00b300c400d700e400eb00ec00ec00ec00ec00ed00ed00ed",
            INIT_0C => X"00e500e300e600e400e800ec00ed00ed00eb00eb00ec00ed00e500e400ed00e2",
            INIT_0D => X"00c500b400b400b000a3009f00a900ce00ee00ed00ec00eb00ec00ee00ed00ed",
            INIT_0E => X"00dc00e600ea00e800ea00ed00ee00ed00ed00ed00ec00ee00cc00de00ec00da",
            INIT_0F => X"00cc00c900c900bf00b600ae00b000c700ef00ef00ee00ee00ef00ef00ef00ee",
            INIT_10 => X"00ea00ec00ee00ef00f000ee00ed00ec00ec00ec00ed00ef00c600dd00ea00e7",
            INIT_11 => X"00d500d800e400da00dd00e000e900eb00f000ee00ef00f000f000f000f000ee",
            INIT_12 => X"008c008a008e009b00bc00ea00ec00ea00e900eb00ed00ed00d800e400ea00ed",
            INIT_13 => X"00e600e600ec00e800ed00e900db00cc00bd00b300b400c700eb00f100f000f0",
            INIT_14 => X"00820079007d007f009f00e500e400e200e800ea00ec00ed00ea00eb00ed00eb",
            INIT_15 => X"00ec00ed00ed00e800ce00b800a5009c0095008c008500a200e400f100f000f0",
            INIT_16 => X"00d400ca00d300d300d900e300d500d100d500de00e200dd00db00dd00e100e5",
            INIT_17 => X"00ea00ec00ed00e700cc00c600c800c200c500b2009700c300e600f000f100f0",
            INIT_18 => X"00cf00ca00d300d900e100db00d000ae00b400d500b80070007200790081008a",
            INIT_19 => X"009800a700d800ec00e800e900ea00e200e400db00cb00e600e300e600ef00f1",
            INIT_1A => X"0082007d007d0083009100b600c900c700db00e600ac00470046004900490054",
            INIT_1B => X"007200a800e300ef00ed00e700e400d300d000da00db00ce00ba00c500dd00e7",
            INIT_1C => X"00510056004f0055008d009b009d00c800e400df00b4007900700075009700c0",
            INIT_1D => X"00d400de00db00cb00ba00a6009a008a0085008b0092008e0089009900c500d4",
            INIT_1E => X"00350046006200900097006b0073009e00b400c200c200c100c200d100e400d2",
            INIT_1F => X"00b500a500960088007d006f006a006f007600790087009700a400ae00ce00cb",
            INIT_20 => X"000f001d008c00d80096007b008500a200b500d100e000ea00ea00f100ee00bd",
            INIT_21 => X"009f009a009e00a300ab00a500a500ab00ae00b100be00cc00cf00c400b700af",
            INIT_22 => X"0005003e00cf00e800cd00cf00d400e000e600ec00ee00ee00dd00ee00ee00e4",
            INIT_23 => X"00d900c800d800d500d400d600d400cc00c100bf00b500a5009c0092008f009a",
            INIT_24 => X"002d009b00cc00c400c500d300d300d000ce00cb00cf00cf00c100c600b000a9",
            INIT_25 => X"00a100ab00a300850089009d009600870073007000720074007d0085008d008e",
            INIT_26 => X"008700b300a0009a0098009800960096009600930093009500950091007e007a",
            INIT_27 => X"007800860080006d007000750070006700610067006f00750079007d00850090",
            INIT_28 => X"0057005a005a005d0062006600660069006f0077007c00830089008800840085",
            INIT_29 => X"00880085007f0077006d00650061005c005e0064006400620068007700870095",
            INIT_2A => X"0019000b0010001a001a00190019001e0024002b0033003b0045004b004d004f",
            INIT_2B => X"005700580051004800430044004500450047004e005900640071007c00880092",
            INIT_2C => X"002e0010000d002c002d0019000b00080004000200020004000d001200130017",
            INIT_2D => X"001d00260021001f0026002c0032003a0046005a0073007b0073007b008b00a0",
            INIT_2E => X"0029001b00130029005100460032001f000f0005000200000011004000320024",
            INIT_2F => X"001e001e001e0023002b003700470061007c008300780069006f0086009800b3",
            INIT_30 => X"000f000a000a000c002c0034002b0021001200040002000100080075009e0080",
            INIT_31 => X"0070006900670069006b0073007e007e006a0056005e00740082009300ac00c2",
            INIT_32 => X"0028000a000300040006000c000c000a00060001000100020000003a00800082",
            INIT_33 => X"007f007b00770071006e0060004b00420047005d00760084008d00a200b600c5",
            INIT_34 => X"004d001d00010001000100020003000200010000000000000001000c002d002f",
            INIT_35 => X"002e003000320031002a00260030004d006e007e00800087009900b000bb00c6",
            INIT_36 => X"005e003400010001000000010001000000000000000000000002000300190020",
            INIT_37 => X"001900190019001d00290042005c0071007c007e007f008b009d00b300bf00c9",
            INIT_38 => X"0066003c0007000200020003000300020001000000000001000300010013001f",
            INIT_39 => X"0011000d001b003a005a0073007e007c007b008200870091009f00b000c000ca",
            INIT_3A => X"006300330017000c000a000b000a0007000400040004000300060005000d0015",
            INIT_3B => X"001b0032004d00620071007e007e007d0080008a0094009a00a800b800c500ca",
            INIT_3C => X"00600039002c0023001e001c001a00170015001500160017001b001f00280037",
            INIT_3D => X"00460058006600700079007a007a007f0085008b009500a000ac00bd00c800ca",
            INIT_3E => X"0065004b0043003d003800350035003700370038003a003e0043004700540060",
            INIT_3F => X"0067006d00740079007f007c007d008300880091009800a200ab00b700c300c8",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY4;


    MEM_IFMAP_LAYER0_ENTITY5 : if BRAM_NAME = "ifmap_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00eb00e700e800e800e800e800e800e800e800e800e900e900e900e900e900e9",
            INIT_01 => X"00e900e900e900e800ea00ea00e800e600e700e900e800e800e800e900e900e8",
            INIT_02 => X"00ee00eb00eb00eb00eb00eb00eb00eb00eb00eb00ec00ec00ec00ec00ec00ec",
            INIT_03 => X"00e900e900ea00ea00ed00ee00ed00eb00ea00ec00eb00eb00eb00ec00ec00eb",
            INIT_04 => X"00ed00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00ea00eb00ea",
            INIT_05 => X"00e700e700ea00ec00e900ee00eb00ea00ea00ea00ea00ea00ea00eb00eb00ea",
            INIT_06 => X"00ee00eb00eb00eb00eb00eb00eb00eb00ea00ea00ea00ea00ea00ea00eb00ea",
            INIT_07 => X"00e600e700e800e700c500db00d500e600eb00ea00ea00ea00ea00eb00eb00eb",
            INIT_08 => X"00ed00ea00eb00eb00eb00eb00eb00eb00ea00ea00eb00eb00ea00ea00eb00eb",
            INIT_09 => X"00ec00ed00e600db00b300d000dd00e800ed00eb00eb00eb00ec00ec00ec00ec",
            INIT_0A => X"00ee00eb00eb00eb00eb00eb00eb00eb00ea00eb00ec00ec00ec00ea00ed00e8",
            INIT_0B => X"00da00d200cf00c800bd00ca00dc00e800ed00eb00eb00eb00ec00ed00ed00ed",
            INIT_0C => X"00e500e400e700e600e900ec00eb00eb00ec00ec00ed00ee00e600e500ee00e4",
            INIT_0D => X"00cc00be00bf00be00b100ab00b100d300ef00ea00e900eb00ec00ed00ed00ee",
            INIT_0E => X"00de00e900ee00ea00ea00ec00eb00ec00ee00ee00ed00ef00cb00dd00eb00da",
            INIT_0F => X"00d200d200d300cb00c400bb00b900cc00f000ee00ed00ee00ee00ee00ee00ee",
            INIT_10 => X"00f100f300f600f300f000ed00eb00eb00ed00ed00ed00ef00c400da00e700e5",
            INIT_11 => X"00d900de00eb00e300ea00eb00f000f100f300f000f000f000ef00ef00ef00ee",
            INIT_12 => X"00950094009900a100bf00e900e900e800ea00eb00ec00eb00d600e200e800ec",
            INIT_13 => X"00e800eb00f100ef00f700f300e200d300c300ba00b900c900eb00ef00ef00ef",
            INIT_14 => X"008d00850089008900a500e700e100e000e900ea00ea00eb00eb00ec00ee00ec",
            INIT_15 => X"00ee00f000f100ee00d500bf00ac00a3009f0099008f00a600e500ef00ee00ef",
            INIT_16 => X"00e000d700e000df00e300e700d300ce00d600de00e100db00df00e100e600e9",
            INIT_17 => X"00ed00ef00f100ed00d000cb00cf00ca00d300c400a400ca00e900ee00ef00ef",
            INIT_18 => X"00de00d900e000ea00f100e300d000ae00b700d600bc0079007e0084008b0093",
            INIT_19 => X"00a100ae00dc00ed00eb00ee00f000e900ed00e500d400ed00ea00e900f200f2",
            INIT_1A => X"00980093008d009700a500c100cd00cc00e200ea00b7005c005b005b005a0062",
            INIT_1B => X"008100b300e900f100f100ed00e900d900d400dc00df00d600c400cd00e300ea",
            INIT_1C => X"006c007200640066009b00a400a400cf00ea00e400be008a0083008700a800cf",
            INIT_1D => X"00df00e800e300d400c300ae00a30093008c009000980097009300a000cb00d8",
            INIT_1E => X"004d005e00740099009c006e007600a100b600c500c600c800ca00d900ec00d9",
            INIT_1F => X"00ba00ac009f0095008a007b0076007b00800082009100a100ae00b800d500d0",
            INIT_20 => X"0023002f009700dc0096007b008600a200b400d300e100e900e800f000ee00be",
            INIT_21 => X"00a300a200aa00b100bb00b600b600bb00bd00bf00cc00d900da00d000c100b7",
            INIT_22 => X"0018004f00d900ef00d400d300da00e500ed00f600f500ef00dc00ef00f100ea",
            INIT_23 => X"00e400d600e600e500e700ea00e800e000d400d100c500b300a900a1009e00a5",
            INIT_24 => X"004700b300de00d800d900e500e600e300e300e400e400dd00cf00d700c100bc",
            INIT_25 => X"00b800c300ba009c00a100b400ad009e008a008700850083008c0097009e009c",
            INIT_26 => X"00a100cf00c200bd00bb00be00c000c100c000be00bd00bd00bc00ba00a3009a",
            INIT_27 => X"009a00aa00a30091009400990090008800820086008b008d009000920094009c",
            INIT_28 => X"006d0071007a007f0086008e00930096009800a000a500ac00b500ba00b400af",
            INIT_29 => X"00ac00a800a3009b0094008b0084007f008100850081007a007e008a0092009c",
            INIT_2A => X"002900190023003000340038003a003d003e0046004d0057006a0079007e007e",
            INIT_2B => X"007f007e00780070006a0068006700660069006e0073007700800088008d0095",
            INIT_2C => X"0037001400130035003a0029001e00180011000f000f0014002a0038003c003e",
            INIT_2D => X"00470051004d004c004e004f0053005a00650076008a008a007d00800089009e",
            INIT_2E => X"002d001a001200290054004c003900250015000b000700070023005b004e003e",
            INIT_2F => X"003c003e003f0045004a00530063007b009200950087007200740085009200af",
            INIT_30 => X"001100090008000b002e0039002f00230014000700040003000f008600b30094",
            INIT_31 => X"0083007d007c007f007e00850090008d0074005b006100740081009000a500be",
            INIT_32 => X"0023000700030004000700110011000c00070003000200030002004000920094",
            INIT_33 => X"0090008d00890081007a006a00530045004600580071007e0087009e00b000c2",
            INIT_34 => X"0040001500010002000000050009000500020000000000010001000b003b0044",
            INIT_35 => X"004300450043003b0031002a002e00470066007400780080009300ab00b700c4",
            INIT_36 => X"0052002b00010002000000020005000200000000000000000000000200260036",
            INIT_37 => X"002e002b0024002200270038005200690073007300760083009600ae00bb00c7",
            INIT_38 => X"005d0032000300010000000100030002000100000000000100020000001c002f",
            INIT_39 => X"0017000c0016003700510063006f007000710077007e0089009700ab00bc00c9",
            INIT_3A => X"00590025000b00040002000400040002000100010001000200060002000d0018",
            INIT_3B => X"00190029003e0052006500710070006f0073007e0089009100a100b300c100c9",
            INIT_3C => X"0052002400160011000f000f000d000c000c000d000e000f00140015001b002d",
            INIT_3D => X"00430051005500580069006e006b00700077007f008a009700a400b700c400c8",
            INIT_3E => X"0053003000260025002300210022002600280029002c002e002d0030003b004a",
            INIT_3F => X"0053005c00610061006b006a006c0075007b0085008d009900a300b200bf00c7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY5;


    MEM_IFMAP_LAYER0_ENTITY6 : if BRAM_NAME = "ifmap_layer0_entity6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009e009e008b008400a600b600bb00c100c700cd00d100ce00da00df00e300e6",
            INIT_01 => X"00d500e200e700eb00ec00e800ea00ea00ec00e200e600ee00e800e400ed00ee",
            INIT_02 => X"00aa00ac0097008900ae00c100c500c700ce00d700d900d200e100e700e900ed",
            INIT_03 => X"00db00e400e800f200f500ea00ec00f200f100e400eb00f300e900e800f600f6",
            INIT_04 => X"00ae00b0009d008e00b500c900ce00c700d100df00da00d400e000e600e600ef",
            INIT_05 => X"00dd00e400e900ef00e800d500ec00f300f500e700ee00f800ed00e600fa00f5",
            INIT_06 => X"00b400b200a0009300ba00cb00d400cf00d600e400dd00d600dc00e700df00f0",
            INIT_07 => X"00e000e400e900e400b100ac00e600f300f800e800ee00fa00ee00e400f900f4",
            INIT_08 => X"00ba00b900a5009300bd00cc00d900cf00d300e700de00d600da00e700d300eb",
            INIT_09 => X"00e200e000e800d4009f00a800e000ed00f700e700eb00f600e800ea00f800f2",
            INIT_0A => X"00c100be00aa008e00bf00cb00db00d300d700ea00dd00d600d600e400c700cd",
            INIT_0B => X"00cf00ce00eb00c10070009e00de00e600f500e500e200f100e400e700f300eb",
            INIT_0C => X"00c400bf00ac008500bf00ca00de00d900df00eb00da00d600d700e300bc00b0",
            INIT_0D => X"00bb00ba00cd00bb0078008900ac00b700db00df00d800eb00e200e100f000eb",
            INIT_0E => X"00cc00c500ae008c00cb00da00e000e000e800ed00dc00dc00dc00dd00c900cd",
            INIT_0F => X"00ac008a006400530047003e0041003c006800b600d100e400da00d400ef00ec",
            INIT_10 => X"00af00aa009d008900b000ba00af00c500d100d400ce00d200d400c900c100c1",
            INIT_11 => X"008e00690059005b00540053005e0045004e007900a200b700ae00a300cf00c3",
            INIT_12 => X"00720073007100680069006b006f0080008b00920097009b009d009300970096",
            INIT_13 => X"00760064006300630055005600560053008b0080009a00990076006d0084007b",
            INIT_14 => X"0042004c004b00440053005a0054005a005d006a00660067006a006b0072006c",
            INIT_15 => X"005a005a005b005500480042005f00720080006e009300c7007d0067005c005e",
            INIT_16 => X"00350041004b004d006f006a00550046005d0071005f005d006c0073006b0061",
            INIT_17 => X"0062005f00620061005a0055009500bb00b30092007000cc009a005f00570055",
            INIT_18 => X"003a0056005e004a00640064004d005500780085007f006c0069006e00620057",
            INIT_19 => X"005100510057005f005f007000aa00c300d000c1007f00ad00b200500055004f",
            INIT_1A => X"004a00590057004b0052004400470050005900670076006f0065006a00690062",
            INIT_1B => X"006000620062006d0072008e00b400b800bf00c000a0008400aa0050003c0043",
            INIT_1C => X"004d004f0052004e004f004800460056006d0079008100850089008800870083",
            INIT_1D => X"0092009400920096009400a300b300b500b900b000aa0065005a00490037003b",
            INIT_1E => X"0060005e006a0068006d00830084008a00900098009b009a009b009b009e0094",
            INIT_1F => X"0096009d009c009200770082009200a900b100a800a700690045006200560048",
            INIT_20 => X"006a006500730083008100870090008f00920096009a009a009a009900970090",
            INIT_21 => X"00820086008b007f005e00750092009f00a700a300a20084009000c0009a0069",
            INIT_22 => X"005f006c0076006d005f005d0081009100950097009600900086007e007a007b",
            INIT_23 => X"007a0085009b00940083009300a2009c009d009700990095009f00a4009d0094",
            INIT_24 => X"00660059004900460056006f007b008c008f0081007800750078007e0085008d",
            INIT_25 => X"0096008e0099009f0097009d00a500a100990098009a009000830079007d0095",
            INIT_26 => X"0056003d0047006e0080008a0082007b0076006c00760084008f0098009c0099",
            INIT_27 => X"009500890091009a0099009a00a000a400980090007d0069005c004b00560084",
            INIT_28 => X"00680067006b007200730074007b007600740086008d0090008f008d00850075",
            INIT_29 => X"00620059008200960097009a0098009100750060005a00500041004700490041",
            INIT_2A => X"0063006b006f006f00720077007d007e0075007d007d008100830082005b003d",
            INIT_2B => X"0039003800730094008b00820072005f005600530049003a003c004b0033001b",
            INIT_2C => X"003e006800740072007400750066005b00540051004e0070008500820060004c",
            INIT_2D => X"00530056006b006c00600058005300510046003d0033002d0034002e001e0018",
            INIT_2E => X"00390060006a0069006b006800410035003b00400044006e0087008500730062",
            INIT_2F => X"0058004f004e00500051005000460037002c0031002d00290022001e001b0018",
            INIT_30 => X"0041005a00680069006d006d004f0049005500580062006a0062005300440041",
            INIT_31 => X"0046004a00510052004800330029002c003d0037002700230020001e001b0019",
            INIT_32 => X"00430057006900670066006300580051004c0045003b0039003a003f00420046",
            INIT_33 => X"00480044003e0036002e002f0031002c0038002e001e001c001d00190018001e",
            INIT_34 => X"0036003a0041003a00370032002d002c002e00330037003a003e0040003e003a",
            INIT_35 => X"003300260025003000310030002a002600290020001b001c001b0019001c001f",
            INIT_36 => X"001e001d001a001b001f0020002100270031003400350033002e002800260028",
            INIT_37 => X"0026002c004200370029002500240025001f001b001a001b001c001e00210017",
            INIT_38 => X"0021001f001b001c001c001e001f002000230021001e001e002200270029002d",
            INIT_39 => X"002a003400490031001e002300260020001b001a001b001d001e0026001a000d",
            INIT_3A => X"001f001e001a001a00190019001a001b001d002000250028002a00290028002a",
            INIT_3B => X"0027002e00400026001c0024001e001d001a0019001b001c0021002500090004",
            INIT_3C => X"0017001b0019001c001e002000220025002700270028002700260023001e0021",
            INIT_3D => X"001c002400390024001e001d001d001d001800180017001b0024001300040005",
            INIT_3E => X"001c001e0020002200210022002300250026002600240022001e0018000f000c",
            INIT_3F => X"00080013002d00200019001b001b001c00180015001400220019000500040007",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY6;


    MEM_IFMAP_LAYER0_ENTITY7 : if BRAM_NAME = "ifmap_layer0_entity7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00be00bb00a6009e00c100d000d300d800db00dd00de00da00e500e800eb00ed",
            INIT_01 => X"00dc00e900ee00ef00f100ef00f100f100f200e700eb00f300ed00e700ef00f1",
            INIT_02 => X"00c800c700b000a000c700d900da00da00df00e500e500db00e900ee00ef00f3",
            INIT_03 => X"00e100ea00ee00f500f700ed00ef00f500f500e900ef00f800ec00e800f600f7",
            INIT_04 => X"00c900c800b300a200c900dc00df00d600dd00e900e200db00e500ea00ea00f4",
            INIT_05 => X"00e200e900ee00f300eb00d600ea00f100f700e900f000fa00ee00e500f900f4",
            INIT_06 => X"00cb00c700b300a400c900d900e100d900df00eb00e300d900dd00e800e200f4",
            INIT_07 => X"00e400e700ed00eb00b800af00e400f100f800e800ee00fa00ed00e300f700f2",
            INIT_08 => X"00cf00cc00b500a100c900d600e100d500d700ed00e200d700d900e500d400ec",
            INIT_09 => X"00e300e100ec00e100aa00ae00e000ec00f700e700eb00f600e700e700f500ef",
            INIT_0A => X"00d000cd00b7009a00c900d400e200d700da00ee00df00d700d700e500c700cd",
            INIT_0B => X"00d100d000ef00cc007c00a700e300e900f600e500e100ef00e200e600f100e8",
            INIT_0C => X"00cc00c700b3008b00c200cb00dd00d500db00e900d800d400d800e600bc00b0",
            INIT_0D => X"00be00c000d400c00081009700b700be00e000e000d600e500db00de00eb00e0",
            INIT_0E => X"00cd00c600af008a00c000cb00ce00cc00d400df00d000d200d500d800c700ce",
            INIT_0F => X"00b200950071005d0055005000500045006c00b700ce00de00d000c500dd00d4",
            INIT_10 => X"00ad00a8009a008500a500ac00a000b300be00c200bd00c300c700bf00c100c6",
            INIT_11 => X"00980079006b006c00680068006e004f0052007a009f00af00a3009500be00af",
            INIT_12 => X"0073007400720069006d006e0070007f00870088008c00930097008f009e00a1",
            INIT_13 => X"0086007700780078006c006c0066005c008f008000970091006e006a00820078",
            INIT_14 => X"004e00570056005200630069006100640065006d006a006f007200760084007f",
            INIT_15 => X"006d006d006e006b00600057006c00770084006f009000bf0078006f00660068",
            INIT_16 => X"004a0055005f00620080007a0062005100680081007100730084008b0086007b",
            INIT_17 => X"007800730074007700710068009e00bd00b70094006d00c50095006700630063",
            INIT_18 => X"0051006b0071005d00750073005d0066008900980095008300820088007d0071",
            INIT_19 => X"006c006c0072007b0076007f00af00c200ce00bd007600a200a7005000620065",
            INIT_1A => X"0061006e006a005d0062005400590064006e007b008a0086007e00830082007c",
            INIT_1B => X"007b007f007e00870086009900b500b400b800b70097007a00a0004d00480059",
            INIT_1C => X"0066006500660061005f00580058006b0082008e0097009e00a300a400a1009d",
            INIT_1D => X"00ab00ad00aa00a900a200a900b100ae00b000a800a4006200570046003f004b",
            INIT_1E => X"007b0076007f007c007e0094009800a000a700af00b300b400b700b800b900ae",
            INIT_1F => X"00ad00b200af00a000800085008e00a100a900a200a6006c0046005f00590052",
            INIT_20 => X"0085007d008a00980094009a00a600a700aa00ae00b300b600b900b900b500ab",
            INIT_21 => X"00980098009a008b006600780090009b00a500a200a30088009100bb0099006c",
            INIT_22 => X"007c0085008d008300740072009800aa00af00af00b000ad00a700a0009a0097",
            INIT_23 => X"0090009600a800a0008c009800a5009e00a3009b009c0097009e009e00980093",
            INIT_24 => X"008100710060005d006e0087009400a400a9009f0096009200940099009f00a5",
            INIT_25 => X"00aa00a000a800ac00a100a400a800a400a0009e009e009200840079007d0096",
            INIT_26 => X"0070005500600087009b00a5009c0093008e008d009700a000a700ad00ae00ab",
            INIT_27 => X"00a7009b00a200a800a300a100a300a6009e00970082006f00620052005c008a",
            INIT_28 => X"008500840087008f008f008f0096008e008a00a100a900ab00a900a500970086",
            INIT_29 => X"0074006b009400a400a300a3009f00980080006c0066005b004b004e00500048",
            INIT_2A => X"0084008c0090008f0090009300970096008b00920094009a009f009c006e004e",
            INIT_2B => X"004b004a008400a30099008f007e006d00670064005a004c004b005200390021",
            INIT_2C => X"005e0089009400920092009100810073006a006600630087009d009a0072005d",
            INIT_2D => X"00650068007d007c0071006a006600650058004f0045003f004300350025001f",
            INIT_2E => X"0056007d0086008600890085005c004d00520059005c00830099009600840073",
            INIT_2F => X"006a00610060006100630065005f004f003c0040003c0039002f00260022001f",
            INIT_30 => X"005a0074008100830089008a006a0061006c0074007c007e0071005f00540053",
            INIT_31 => X"0059005c00620064005c004a00430045004a00420033002e002b002600230020",
            INIT_32 => X"005c00700082007f007c0078006e00660061005a0050004c004b00500054005b",
            INIT_33 => X"005f005900510049004100410043003d0045003a002a0028002a002800230025",
            INIT_34 => X"004c004f0056004e004a00450040003f00410046004a004d0051005200510050",
            INIT_35 => X"0049003b003700440043003f003600320036002d002800280029002800270025",
            INIT_36 => X"002d002b0028002a003100340035003a00440047004800460041003b003a003b",
            INIT_37 => X"0038003f0055004900390033002f002f002c0028002700280029002a002a001d",
            INIT_38 => X"002b002800240026002c00300031003200350034003100310035003b003e003d",
            INIT_39 => X"00370045005e0042002c002e002f0028002700270028002a0029002e00200012",
            INIT_3A => X"0028002700230024002700290029002b002e00330038003a003d003d003c0037",
            INIT_3B => X"002e003c005500360028002e00250024002600260028002a002b0028000d0007",
            INIT_3C => X"0022002600240028002c002f0031003300360039003b0039003900370033002b",
            INIT_3D => X"001f0030004e003200290025002300230025002500240029002d001400060007",
            INIT_3E => X"0029002b002d002f0030003000300031003200330031002d00280022001a0011",
            INIT_3F => X"0008001b003f002c0021002200220023002300220022002c001f000600050008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY7;


    MEM_IFMAP_LAYER0_ENTITY8 : if BRAM_NAME = "ifmap_layer0_entity8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00de00da00c200ba00de00ec00ee00f100f300f500f400eb00f000f100f200f5",
            INIT_01 => X"00e300f000f500f800f900f300f300f300f500eb00ef00f700f100ea00f300f6",
            INIT_02 => X"00e500e200c900b800df00f000f000ee00f300f700f500e800f300f500f500f8",
            INIT_03 => X"00e600ef00f300fb00fb00ee00ee00f400f800ec00f300fc00f000ec00fa00fb",
            INIT_04 => X"00e100de00c700b500db00ee00ef00e400eb00f400ec00e400eb00ef00ee00f7",
            INIT_05 => X"00e500ec00f100f600ec00d700e800ef00f800eb00f200fc00f100e800fb00f7",
            INIT_06 => X"00de00d800c200b300d600e400eb00e100e500ef00e600dd00e100ec00e600f7",
            INIT_07 => X"00e600ea00f000ee00ba00b000e500f100f800e900ef00fb00ee00e400f800f3",
            INIT_08 => X"00df00d900c100ac00d200dd00e700d900da00eb00e100d700db00e800d600ee",
            INIT_09 => X"00e500e300ee00e400b000b200e500ef00f700e700ea00f500e700e800f600f0",
            INIT_0A => X"00dc00d500bf00a400ce00d500e100d500d600e600da00d600d600e300c800ce",
            INIT_0B => X"00d000ce00ed00cf008200ad00e600e900f400e100db00e800dd00e700f200e6",
            INIT_0C => X"00d400ca00b9009600c400c900d900d000d300db00d000d300d400dd00b900af",
            INIT_0D => X"00bb00bd00d200c50089009d00b800bb00dd00dc00ce00da00d100db00e700d8",
            INIT_0E => X"00d300c900b3009300c500cc00ce00cb00d000d200c600cd00ce00ce00c000cb",
            INIT_0F => X"00b3009b007a006a0064005e00580049006f00b700ca00d700c600b900ce00c1",
            INIT_10 => X"00b300ad00a0008c00aa00af00a100b300bb00b800b400bd00c300b900ba00c4",
            INIT_11 => X"009f008900800080007e007e0080005a0058007c009e00ac009c008900b0009f",
            INIT_12 => X"007b007e007b0070007200720072008000860086008900900098009200a000a7",
            INIT_13 => X"0093008b0090008c0082008300780068009500830096008d006a006900800075",
            INIT_14 => X"0059006600620058006b00730068006a006b007600710073007b008600970092",
            INIT_15 => X"0080007f007f0078006f0068007a00800086006e008b00b600720075006d0070",
            INIT_16 => X"00580068006e006a008e00890071005e00740092007f007d009400a500a50097",
            INIT_17 => X"008e0082007f007f007b007200a500bf00b4008e006400b8008c006d006c006c",
            INIT_18 => X"006400820084006800810082006d0076009a00ab00a80097009b00a5009a008b",
            INIT_19 => X"0082007d0081008c0086008900b300c100cb00b90070009800a000540069006d",
            INIT_1A => X"00780086007e006a00710065006c00790083009100a1009f009900a1009e0095",
            INIT_1B => X"009200930091009b009600a100b600b100b500b500940076009d0050004e0060",
            INIT_1C => X"007f0080007d00720074007100730086009f00a800b000b800be00bf00be00b9",
            INIT_1D => X"00c500c400be00b800ac00ad00af00a800ab00a500a300630057004700430051",
            INIT_1E => X"00970095009a0091009900b300b800c100c900cd00cf00d000d100d200d400c8",
            INIT_1F => X"00c600c900c300ab00860087008b009b00a500a100a800710049005c005a0056",
            INIT_20 => X"00a5009f00a700b000af00b900c600c900cd00d000d200d200d200d000c900be",
            INIT_21 => X"00aa00aa00a90094006c007a008e009900a700a500a7008e009300b50098006f",
            INIT_22 => X"009d00aa00ae009d008d008f00b600ca00d000d300d100ca00bf00b500a700a2",
            INIT_23 => X"009b00a000b200a90093009d00a700a000a900a200a1009c009e009600960094",
            INIT_24 => X"00a2009400800079008a00a400b100c200c700bc00b200ab00aa00ac00ac00b0",
            INIT_25 => X"00b400a800b000b500aa00ad00af00ac00a800a500a3009600850076007d0099",
            INIT_26 => X"008f0075007f00a600bc00c500ba00b000a900a300ab00b200b900be00bf00ba",
            INIT_27 => X"00b400a500ac00b100ad00ac00af00b200a4009c008800740067005700620090",
            INIT_28 => X"00a600a500a800b000b000ae00b300aa00a400b800be00bd00b900b500a80096",
            INIT_29 => X"00810076009d00ad00ad00ad00ab00a200850070006a005f005000540056004e",
            INIT_2A => X"00a500ac00b100af00ae00b000b300b000a400ab00ab00ad00af00ab007e005e",
            INIT_2B => X"00580055008e00ac00a2009800880075006c0068005e0050004f0058003f0027",
            INIT_2C => X"007c00a600b200af00af00ad009a008b0082007e007a009a00ae00a90083006c",
            INIT_2D => X"007200720086008500790071006d006c005f0056004b00450049003b002b0026",
            INIT_2E => X"006f009600a0009f00a3009e00740064006800700073009700ac00a800950083",
            INIT_2F => X"0077006b006a006a006a006c0064005400450049004400410037002c00280025",
            INIT_30 => X"0071008a0097009a00a100a20080007700810088009000920084007200650062",
            INIT_31 => X"00650067006d006c006300500048004b0055004d003d003a0034002d00290027",
            INIT_32 => X"00740088009a00970094008f0084007c00760067005b00570056005b00630065",
            INIT_33 => X"00650063005e005200480048004a0045004e00440034003200330030002f0030",
            INIT_34 => X"00600064006a0063005c0056005200510052004f005100540057005b005e0058",
            INIT_35 => X"004d00440044004c004a00480040003b003f0036003100320031003000340030",
            INIT_36 => X"003b003900360037003c003d003e0044004e004f004f004d0048004400450042",
            INIT_37 => X"003d0047006100520041003c0038003900350031003000310032003200320023",
            INIT_38 => X"00320030002c002d0031003500350037003a003b00380038003c004200470044",
            INIT_39 => X"003b004b0068004b00350038003a003300310030003100330032003500250014",
            INIT_3A => X"002d002c00280029002c002e002e003000330039003f0041004400440044003d",
            INIT_3B => X"00320042005d003f003100380030002f002f002f003100330034002e000e0005",
            INIT_3C => X"0027002b0029002d003200360038003b003e0040004200400040003d003a0031",
            INIT_3D => X"002400350055003b00320030002f002f002e002e002d00320036001800030003",
            INIT_3E => X"002f003200340036003800380038003a003a003700350032002d0027001e0014",
            INIT_3F => X"000b002100480036002c002d002d002e002c002c002b00340025000800030007",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY8;


    MEM_IFMAP_LAYER0_ENTITY9 : if BRAM_NAME = "ifmap_layer0_entity9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009b00a700b000be00b100a600a800a600aa00b300bb00bb00bb00bb00b800b8",
            INIT_01 => X"00b600b400b800ba00bb00bb00bc00bd00bb00bb00bc00c300c900c900ca00c0",
            INIT_02 => X"009900a300ab00bb00b3009b009a009f009f00a500ab00af00a900ab00a200a5",
            INIT_03 => X"00aa00a400a600a500a700ad00a900a800a900ad00be00ca00cc00ca00cb00bd",
            INIT_04 => X"009b00a000a800b800bb00ae00b000bc00b600b300b100be00c000c200bc00b9",
            INIT_05 => X"00c100c200c100c200c300c500c100bf00bf00c500ce00cf00d000ce00cc00bd",
            INIT_06 => X"0097009d00a600b100b400b900c700c500b600cc00cd00c600d200c500c400cb",
            INIT_07 => X"00cd00cf00d200cb00cf00d200c500cc00d000c600cc00c900d100cf00ce00c0",
            INIT_08 => X"0097009e00a800ae00b100b500bf00c400b700c200bd00b900c400b900b900ca",
            INIT_09 => X"00c700c700c800c000c300c700be00bc00c900c700c900c400ce00cc00cf00c4",
            INIT_0A => X"0094009c00a700ae00ab00ae00c400c300c000be00bd00b800bb00bd00bd00bf",
            INIT_0B => X"00be00c300bb00c600c000bc00c000c100cd00ce00cb00d100d400d000d100c4",
            INIT_0C => X"0094009900a500ae00a800b000cb00c300bc00bc00bb00be00b600c200c500c3",
            INIT_0D => X"00c400c100c800cd00c600c500c500c900c500c800c600c300c500cb00cf00c3",
            INIT_0E => X"0099009b00a300ac00ac00bc00c700d100c400be00bd00bf00c100bc00bb00c4",
            INIT_0F => X"00ca00c200c400ce00c200c900c400c800b500bb00c800c900c800c400c700bd",
            INIT_10 => X"00a0009f00a300ac00ae00b000b000be00b400af00b000b000b500aa00ac00b6",
            INIT_11 => X"00bb00b200b500bb00b100bc00b400bb00c700c400bc00bc00c500c000c200b8",
            INIT_12 => X"00ab00a700a200ac00aa00ab00b400b0009b009c0096009c009600920099009e",
            INIT_13 => X"00a600a600a4009d009d00a2009c00a600c800c700bc00bd00c500c100c200b6",
            INIT_14 => X"00af00b400a800b000ad00b100b600ae009c00a0009f009a009f00a300a800ad",
            INIT_15 => X"00aa00a400a000a200a000a800a700ac00c200c300c400c400c500bf00c100b7",
            INIT_16 => X"00b500bb00b200bb00b700aa00ae00b600b300b300b400b500b800bb00c100c1",
            INIT_17 => X"00c100c000bc00b900b800ba00c000c000bb00bc00c000bd00be00bf00c400ba",
            INIT_18 => X"00b900be00ba00ab00990084009500c100c600bf00ba00bc00bf00c100c300c4",
            INIT_19 => X"00c300c000be00bc00bc00be00c000bf00bf00c100c300c500ca00ca00cc00c1",
            INIT_1A => X"00ba00c200bc009e00840074005e006d009100b100c200c200bf00c100c400c7",
            INIT_1B => X"00c700c700c800c600c400c400c700c600c500c400c400c400c600c500c600b9",
            INIT_1C => X"00ba00c500c400c600c200b8008d005c00540068008e00b300c300c900cc00cc",
            INIT_1D => X"00cc00cc00cc00c700c200c200c200bf00bd00be00be00be00bf00be00c000b5",
            INIT_1E => X"00b800c700c600c800c500c800c900b100750054005d008000ad00ca00d000cd",
            INIT_1F => X"00ca00c800c700c700c300c400c500c300c100c300c200bf00bf00bd00be00b2",
            INIT_20 => X"00b900c900cb00d000cd00ce00d000d600af005c004c005b0069008c00b500cb",
            INIT_21 => X"00ce00ca00c500c200c100c200c200c200c200c300c100bf00c100be00be00b4",
            INIT_22 => X"00bb00cc00cf00d600d400d400d300d000cb007c004700570054005400630084",
            INIT_23 => X"00a700be00cb00cb00c300c000c500c400c200c200c000bf00c100bf00c000b7",
            INIT_24 => X"00be00cf00cf00d600d400d300d300d000d30089004800570053005400560053",
            INIT_25 => X"0059006b0083009b00a300b600cb00cc00ca00c600c200bf00c100c000bf00b6",
            INIT_26 => X"00bf00d200d100d700d500d400d400d500cc0071002f003a003f004c0057005d",
            INIT_27 => X"005a00500046003e003a004d007a009f00b400c200c900c800c800c400c400b9",
            INIT_28 => X"00bf00d000cf00d300d100d200d100d4009d00650041002500330044004a0058",
            INIT_29 => X"005b0056005500490037002e003e0048004e006b0085009e00b800c300c400ba",
            INIT_2A => X"00ba00ca00cb00d100cf00ce00d100c80095008c00970064002d003500320060",
            INIT_2B => X"009c00a00080004800620070005900420043008300a600a300ad00b700bc00b2",
            INIT_2C => X"00b900c900ca00d200d200d000d100d100d200d300d700bd00900092009400a8",
            INIT_2D => X"00ca00ce00c0009a00a300b200b1009f009c00b200bf00c200c400c100bc00b0",
            INIT_2E => X"00b000bc00c000c400c000bc00b900b700b600b200b300ad00aa00aa00ab00ad",
            INIT_2F => X"00a900a000a100a700a500a100a500aa00aa00a000980096009d00a300a4009c",
            INIT_30 => X"00720063006e006b00660061005e005d0058005500580050004d004e00530065",
            INIT_31 => X"0071006c006a006b006c006e006f0071007500770078007700780079007a007c",
            INIT_32 => X"007a006d007100750073007000720071006f0070006f006d006e006d006e006c",
            INIT_33 => X"007300700069006b006c006a00650068006a006b006d006d00670066005e0065",
            INIT_34 => X"00780061006b0070006d00680062005e005e005d005800560052004f0050004e",
            INIT_35 => X"0050004f00480045004300420041004100400041004200400043003f0035004d",
            INIT_36 => X"005b00370041004500420042003f003d00420040003c00390039003c003d003f",
            INIT_37 => X"003f00420040003a00380039003b003c003a00390038003900340031004b005c",
            INIT_38 => X"005d003c00420044004300430040004100450041003e003b003b003b003c003d",
            INIT_39 => X"0040003f003a003800370037003800380039003a003800350041005d00610051",
            INIT_3A => X"00590039003d00390039003b0039003b003c003a00380036003c003d003b003d",
            INIT_3B => X"0041003d003a0039003c003c003d003d0042003e0039004600610059003b0043",
            INIT_3C => X"0059003c003f003e003e003e003e003f003e003d0041005200540051004e0051",
            INIT_3D => X"005800540055005300500043004200400034003800560067004c0039003d004b",
            INIT_3E => X"005c003c003d003c003f00420043004100420043004100480049004900480046",
            INIT_3F => X"0049004a004b004b004b00400040003e00410056005800400039003c00400049",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY9;


    MEM_IFMAP_LAYER0_ENTITY10 : if BRAM_NAME = "ifmap_layer0_entity10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009c00b000b300c000b900ab00ad00ad00af00b300b600b800b900b800b600b5",
            INIT_01 => X"00b300b300b700b900ba00ba00bb00bd00bb00bb00bc00c300c500c400ca00b7",
            INIT_02 => X"009b00b300b800c300be00a2009f00a400a300a500a900b000ab00ae00a400a7",
            INIT_03 => X"00ac00a600a800a600a900af00ab00a900aa00ae00bf00cc00ce00d000d700be",
            INIT_04 => X"009a00b200b900c400cb00c100b200a800a000af00be00c400c300c500be00bc",
            INIT_05 => X"00c400c300c200c300c400c600c100bf00c000c400cd00cd00ce00d000d700bf",
            INIT_06 => X"009a00b200bc00c300ca00c500bc0080006c0098009a009b009e009500950094",
            INIT_07 => X"00a700a100a300ad00a800a300ae009f00bc00d000cc00ce00cc00cd00d400bc",
            INIT_08 => X"009a00b100bb00bf00c600c400bd007e0080008b006a006b0073007800760071",
            INIT_09 => X"007700720072007e007600700088007000a000cb00c900ce00ce00cd00d600be",
            INIT_0A => X"009700ae00bb00bd00c500c800b7009300a900a8009100a500aa00920095009d",
            INIT_0B => X"00b400b200b000bd00b000b300bc00b100c400d000cf00d000d000d100d800be",
            INIT_0C => X"009800ac00b900bd00c200c6009300600095009700900098009800790080008b",
            INIT_0D => X"009c009700aa00a2009600ad009600a4009c00a600cc00d200d300cf00d400bc",
            INIT_0E => X"009b00ac00b600bb00c200b500770065007b008300830078009200870087007f",
            INIT_0F => X"007b007b0083007b006d0084007b009f007b008400bf00c700c900c900d000ba",
            INIT_10 => X"00a100af00b400b900c000ba00ab00af00a200a500ac00a600af00ac00ad00aa",
            INIT_11 => X"00ac00b200b200af00a300ac00b200be00ac00b000c800cd00c800c900d100b9",
            INIT_12 => X"00ac00b700b400ba00be00c000c200b700a000a500a200a3009f009e00a400a2",
            INIT_13 => X"00a700ae00ac00a200a000a300a500b600c800c600ca00cd00ca00ca00d000b8",
            INIT_14 => X"00b100c400ba00be00c000c100c100b700a300a700a5009f00a400a600aa00ac",
            INIT_15 => X"00a800a600a600ab00a800ad00ab00b200c700c600c700c700c800c800d000b8",
            INIT_16 => X"00b700cc00c300c800c900bb00be00c600c200c100c100c100c100c200c600c6",
            INIT_17 => X"00c600c300c300c600c500c400c400c500c900cb00c900c900ca00c800d100bb",
            INIT_18 => X"00b900cd00c600b200a6008d009a00c400ca00ca00c700c500c500c700c900ca",
            INIT_19 => X"00c900c700c600c400c400c600c700c600c700ca00cb00ce00cf00ce00d400bd",
            INIT_1A => X"00ba00d000c800a50090007c005f006b008f00b300c700c700c500c600c900cc",
            INIT_1B => X"00cc00cd00ce00cc00c900c900cd00cd00cc00cb00cb00cb00ca00ca00cf00b7",
            INIT_1C => X"00ba00d400d000cc00ce00c1008f005b00510065008e00b500c600cc00cf00cf",
            INIT_1D => X"00cf00cf00cf00ca00c500c500c600c500c500c500c500c500c400c500cc00b5",
            INIT_1E => X"00b800d600d200ce00d100d400cf00b300740053005d008000ae00cb00d200ce",
            INIT_1F => X"00cc00ca00ca00c900c600c700c900c900c800ca00c900c700c600c600cb00b4",
            INIT_20 => X"00ba00d700d600d500d600d600d400d900af005b004900560065008a00b500cc",
            INIT_21 => X"00d000cb00c700c600c700c900c900c800c800ca00c900c900ca00c800cc00b6",
            INIT_22 => X"00bb00d800d800d900db00d900d600d300cc007b00440052004f005100610082",
            INIT_23 => X"00a500bc00c900ca00c400c100c700c600c600c700c800c800c900c700cc00b6",
            INIT_24 => X"00bc00d900d500d600d800d800d600d200d4008800460053004e00500050004d",
            INIT_25 => X"00530066007e0097009f00b200c900cc00cb00c900c800c600c700c500c900b4",
            INIT_26 => X"00bb00da00d600d500d700d800d700d800cc0070002d0037003a0045004d0051",
            INIT_27 => X"0050004d0046003e003b004f007c00a000b500c400cd00cd00cb00c800ca00b4",
            INIT_28 => X"00bc00d800d200d100d300d600d400d4009a005f003a00210030003e0041004d",
            INIT_29 => X"00520054005400480038002f003f0048004e006b0084009e00b500c100ca00b6",
            INIT_2A => X"00b800d200ce00cf00d100d300d400c800910085008f0061002d0032002e005a",
            INIT_2B => X"0096009e007f004700610070005800410043008200a500a200a800b500c500b0",
            INIT_2C => X"00b700d200cd00d000d300d400d500d200d100d100d400bf00940093009300a6",
            INIT_2D => X"00c800d000c3009d00a600b500b400a2009f00b400c100c500c300c100c700b1",
            INIT_2E => X"00ae00c400c300c200c200be00bb00b900b800b500b700b500b200b000ae00ad",
            INIT_2F => X"00aa00a400a600ac00aa00a600aa00b000af00a5009d009b009d00a300af009e",
            INIT_30 => X"0070006c007000690067006400610060005c005a005e00570054005300570067",
            INIT_31 => X"00730070006f00700071007300740076007a007b007c007b0079007a0084007c",
            INIT_32 => X"00750073007100700071006f00710071006f0070006f006e006e006d006e006b",
            INIT_33 => X"00730073006c006e006f006d0068006b006d006e007000700064005f00620065",
            INIT_34 => X"007100660069006a006a00660061005d005f005e005900550052004e004f004e",
            INIT_35 => X"0050004f0047004400430041004100410041004200420041003c003700470064",
            INIT_36 => X"0054003c0041004000400040003e003c00420040003d00380039003c003d003f",
            INIT_37 => X"004000430041003b0038003a003b003c003a0039003800380038004800750080",
            INIT_38 => X"0053003b003f003e003f0041003d003f0043003e003c0039003a003a003c003d",
            INIT_39 => X"004100440040003e003d003c003e003d003a003a003d0041005b008800890063",
            INIT_3A => X"004f0035003d00390037003b003a003c003d003c00390037003c003e003d003f",
            INIT_3B => X"0043003f003c003b003e003e0040003f003e003c0047006e008e0077004f004a",
            INIT_3C => X"0052003a00420041003f003e003e003e003f003e0041004f004f004c004a004d",
            INIT_3D => X"005400500050004e004c003f003e004100420056007c008d0066004200400045",
            INIT_3E => X"004e0034003a003a003a003a003b0039003a003b003a00450047004700460045",
            INIT_3F => X"004800480049004a0049003f003f0044005a0080008000580042003f00410044",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY10;


    MEM_IFMAP_LAYER0_ENTITY11 : if BRAM_NAME = "ifmap_layer0_entity11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009500bb00c100cd00ca00b700b500b400b600bd00c100c000c000c000bd00bd",
            INIT_01 => X"00ba00b900bd00c000c100c100c000be00bb00bb00bc00c300ca00d100d400ab",
            INIT_02 => X"009d00cc00d700e300e000be00b300b300b300bb00c300c300bb00be00b400b7",
            INIT_03 => X"00bc00b700b800b700b900bf00bc00bc00be00c200d300e000df00de00e300b7",
            INIT_04 => X"009900c900d500db00df00d500c400b800b100c300d300d400d000d200cc00ca",
            INIT_05 => X"00d100d100d000d100d200d400d000d000d000d500de00df00da00d700e000b8",
            INIT_06 => X"00a600cf00d300de00e200dc00c900830077009e00a600b100b200a700a600ab",
            INIT_07 => X"00b700b200b200ba00b900ba00b400a500cf00e400dc00dd00e000df00e600ba",
            INIT_08 => X"00a700cb00ca00da00e000e100d6008e00990098007800810081007e007c0083",
            INIT_09 => X"008600840082008a00880088008d007b00ba00e300da00d900de00dc00e300b9",
            INIT_0A => X"00a400c900cb00d900dc00da00d100a500c400b5009c00b400b300a000a300ac",
            INIT_0B => X"00bf00c100be00c900bf00c000c600be00d400e100e100e100df00e100e800bc",
            INIT_0C => X"00a400c600c800d900d900d600ac0068009e00a500a600af00a50090009700a0",
            INIT_0D => X"00b200ad00bd00b600aa00b700ad00b900a600b200dc00e200dd00e000e700bc",
            INIT_0E => X"00a900c900c700d800da00cb0092006f00860095009d0090009b008f008f0090",
            INIT_0F => X"0093008e0094008e007f008d008e00b00089009500d100dc00d900dc00e400ba",
            INIT_10 => X"00b100ce00c700d900db00cd00c100c500b800b700bb00b800c000ba00bb00bd",
            INIT_11 => X"00c000c200c200bf00b200ba00bc00c800c100c600d600db00db00dd00e400b9",
            INIT_12 => X"00ba00d400c500d600d700d600dc00d200b900bb00b600ba00b600b400b900ba",
            INIT_13 => X"00c100c600c300b800b500b600b600c600de00de00dd00df00df00de00e300b7",
            INIT_14 => X"00bc00de00c800d800d700d400d600cc00b500b800b600b000b500b800bc00bf",
            INIT_15 => X"00bd00ba00b800b900b600b800ba00c900df00dd00dc00db00db00dc00e300b8",
            INIT_16 => X"00bf00e200cf00e000dc00d100d700de00d900d700d600d700d900db00df00df",
            INIT_17 => X"00df00dd00db00da00d800d600d900db00db00db00d900d600d700db00e300ba",
            INIT_18 => X"00bc00dc00d400ce00b5009900ac00d900e200e100dd00dc00de00df00e100e2",
            INIT_19 => X"00e100dd00dc00da00d900db00dc00da00d900dc00de00e000e000e000e600bb",
            INIT_1A => X"00bd00df00d600c1009d007e00630073009d00c600dd00dd00da00dc00df00e2",
            INIT_1B => X"00e200e000e100df00dc00dd00e000e000df00de00de00de00dd00dd00e200b7",
            INIT_1C => X"00bd00e200de00e900dc00c40092005a0054007100a100ca00da00e000e300e4",
            INIT_1D => X"00e200e100e000dc00d700d700d800d900d800d800d800d800d700da00e100b6",
            INIT_1E => X"00bb00e500e000ea00e100e100da00b300730058006a009100c000dd00e400e1",
            INIT_1F => X"00df00db00da00d900d600d600d900db00db00dd00dc00da00d900dc00e200b7",
            INIT_20 => X"00be00e900de00e900e400e200e000e100b500620050005b006a009200c000d9",
            INIT_21 => X"00e000e100dd00da00d900da00da00d900da00dd00dd00dd00dd00dc00e300bc",
            INIT_22 => X"00bf00ea00dd00e900e700e300e200dd00d500820049004f004b005000640088",
            INIT_23 => X"00ad00c800d700dc00d900d900df00de00dd00dd00db00db00da00db00e300bd",
            INIT_24 => X"00bd00e800d900e400e300e100e200dc00dd0090004a0050004a004c004e004c",
            INIT_25 => X"00530064008100a100b000c900e100e200df00dc00d900d700d700d900e100bb",
            INIT_26 => X"00bb00e800d700e100e000e100e300e200d5007700320038003b0045004d0052",
            INIT_27 => X"005000480042003f0041005b008500a200b800cc00da00df00dd00dd00e300bc",
            INIT_28 => X"00b700e700de00df00df00e600e400e100a20062003c0027003500430044004e",
            INIT_29 => X"005100520053004800390031003f0043004b006d008b00a800c600d700df00c3",
            INIT_2A => X"00b000e200e200de00de00e200e200d4009b008b0096006a003500390033005e",
            INIT_2B => X"009a00a10082004900630072005a00430045008600ab00a900b700c500d000be",
            INIT_2C => X"00af00e100e100df00df00de00de00de00de00e000e400cc009f009f00a000b3",
            INIT_2D => X"00d600dc00cf00a900b200c100c000ad00ab00c300d200d600d800d100d200bd",
            INIT_2E => X"00a600d400d700d100ce00cc00c900c700c700c300c500c200c000c100c200c4",
            INIT_2F => X"00c400c200c400ca00c800c400c800cd00ce00c500c000bf00c500c500c900b5",
            INIT_30 => X"006500780082007800760070006b006a006500620066006300620065006c0080",
            INIT_31 => X"0090009200920093009400960098009e00a400a600a800a800a800a500a70092",
            INIT_32 => X"006f008200860086008a008800890088008400860083007e007f008000830083",
            INIT_33 => X"008a0086007f008100810080007c007e00810082008400840077007300730060",
            INIT_34 => X"0068007100780078007a0076006c00640060005b005500590058005500570056",
            INIT_35 => X"0056004f0046004300420041003f003c003b003c003c003b00360032003f004b",
            INIT_36 => X"003d0037003d0039003a003f003b003600380033002f002f0030003200310032",
            INIT_37 => X"003300370035002f002d002e0032003700360034003400340030003a00680068",
            INIT_38 => X"0044003d0041003c003e003d00370039003d00380037003a003b003800380036",
            INIT_39 => X"0039003b0037003400330033003400340033003500370039004b00710078004b",
            INIT_3A => X"003e0034003b0035003900390034003600360032003000320039003800340035",
            INIT_3B => X"0039003600340033003600370035003000320034003d005f007c0065003e0032",
            INIT_3C => X"003e0035003a0037003b003d003c003c00390037003a004b004c004800440045",
            INIT_3D => X"004b004a004b00490046003a0037003500330045006b007f005b003a00360033",
            INIT_3E => X"004000330033002e0033003800390035003400330032003e0040003e003c0039",
            INIT_3F => X"003c003e00400040004000350034003700460067006900480035003200340032",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY11;


    MEM_IFMAP_LAYER0_ENTITY12 : if BRAM_NAME = "ifmap_layer0_entity12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"004100460030001e00170028002c002d002d0028000a000f002c003500330030",
            INIT_01 => X"0041005a005d005b005f0051003c00370070006f00290044004d003300360043",
            INIT_02 => X"0045004f003c001e002900410031003100310023000700190041004500370031",
            INIT_03 => X"004d005500530050005700510037003b00830079001f002f003800360041003d",
            INIT_04 => X"00490054004800290040004a0032003600360020000b0024003c0043002f0027",
            INIT_05 => X"004b004d003b003e005300550030003f008b0080001700290046004e00490030",
            INIT_06 => X"0058004b00500036005000440037003f003a001c00110025002b003300280027",
            INIT_07 => X"00550062004b00460056005400320044008e0089002f004b0064005d00410026",
            INIT_08 => X"005f0059006f00420051003d003d0044003e0016000f0016001f00230033003f",
            INIT_09 => X"0048004b00480047004d00530033004e0095009c005700570063005f004b0058",
            INIT_0A => X"005200530052004d0047003a00400039003b00140011001c0032003d00470047",
            INIT_0B => X"0045004300440038002900530046004e009c00ac00620059005e006f00700063",
            INIT_0C => X"004500400020003b0048004a0049003100310012001d003e005200550056003f",
            INIT_0D => X"00220034005f002b0019005e0055004e00a600b4006d006b006c00830056002f",
            INIT_0E => X"003b0035001900460051004e0050003d0028000a0035005e00570058004b0019",
            INIT_0F => X"000d002d005c00390032006500590062009000b30078007c007c008000340018",
            INIT_10 => X"0044002f0031006600770059003f004f00420022005100600059005a0029000e",
            INIT_11 => X"0034005c00430047006f0071006e00730088009c0079007f007c0073001f0016",
            INIT_12 => X"004d0035003700720080007b00410037004f0052006f006e006a004500140025",
            INIT_13 => X"005c006900530061007600780073005c00900093007d007f0077005f000e0017",
            INIT_14 => X"0055003a003600700081008400640031002700540068006d007d005d003f0053",
            INIT_15 => X"0061005e0068006e006d007f0055003900980096007b007c0072005d000c0015",
            INIT_16 => X"006c00350032006b007e00830080004b0033005b0055006b008a006e00810093",
            INIT_17 => X"008400780071007700750073005a005d00a0008d0071007d00790065000e0009",
            INIT_18 => X"0060002a002b005c006a0080008200770078007b007200890094006e00690084",
            INIT_19 => X"0092008700800086008c0078007e0077009800910063006a0082006300120028",
            INIT_1A => X"00610042003b00590064006f008500880093008c00960091008e00880083007f",
            INIT_1B => X"007d007b008800930097008e009c008800920090006d00700082005c00320053",
            INIT_1C => X"00690048004b005f0068005e00850085008f0087008000850093009600a00098",
            INIT_1D => X"0091009000840087008a008a00a200a500a3007f007e00770076005f003b004d",
            INIT_1E => X"005e00440044005b00650062007b0083009300c1008a004f007c0093009300a2",
            INIT_1F => X"00b400ab0098009000900079009400b300b400a00080007b0070003f001a0054",
            INIT_20 => X"0058004f004a0059006e007800780081007800b800c000570072009c00a400a6",
            INIT_21 => X"009a00a100b700b600bb00ad0094008f00b500c3008e007c006b002c00290076",
            INIT_22 => X"005b00590067006000740064006f006a0072008000bb00a8008c009900ac00ac",
            INIT_23 => X"00a700a4009d00a300a100a500ab009c00a1009100a70072006a004a002a005e",
            INIT_24 => X"006500610078007a0072004e005f005b0073006e008100cc00a7008900a00099",
            INIT_25 => X"00b300ba00aa00b200b3009c00a200a5009c008c006800480054005900460072",
            INIT_26 => X"006e006b007a0060005a004c00480064006d007f0057008c00bd009f00a600b4",
            INIT_27 => X"00ae00ad00be00bc00a2009900a200a100990095004b004a0042003e0070008a",
            INIT_28 => X"0077006a0059004e00590047003c0067004b005f00720042007f00b500ae00be",
            INIT_29 => X"00ba00ab00b800c100a400a000ab00a50092008b0068005c004d005e00700073",
            INIT_2A => X"007e005e003a0067006a004c0048005f005e004100780063005b00a100c400bc",
            INIT_2B => X"00b600c100a700a700aa00a0009a00a10091008a006e005100690088006d0064",
            INIT_2C => X"006f0052004600680071005e004500540074006d0055007d007f009b00ba00c8",
            INIT_2D => X"00bb00bb00b1009d009400a200a400a600a20095007900610078007300610061",
            INIT_2E => X"0065005c008c00b40097007b0055004c0067007c005a0054009200af00ad00c8",
            INIT_2F => X"00bc00ad00ad009f009f00ac00a300ad00a4008b008300830070005f00640060",
            INIT_30 => X"0077009000c000d100c2009d007f006c006a005e006a006f007c00af00b000c5",
            INIT_31 => X"00b800aa00b000a5009c00c500af00a300930083007a006500640060006b0066",
            INIT_32 => X"006e0074008a00a900c500c400a0008800810063005c008a0092009f00b400a9",
            INIT_33 => X"008e008d00af00b200a600bc00b30097008f009a0070003a005b006500660049",
            INIT_34 => X"005b0057004a006b00a500b900bf00a300860080006a00660076008400920074",
            INIT_35 => X"004d006300a100b600b7009f00ad00a7009c0087005e002b005b005c0044004d",
            INIT_36 => X"0051005f0032002c005f009400a600bb00ae0090007e0072006800720077006b",
            INIT_37 => X"00510052009d00b600a900b200a900960098006c002c003f0061004500500056",
            INIT_38 => X"005a005f00340015001c006d009200b000ca00b5008e007f0078007700720082",
            INIT_39 => X"00810076009000a9009f00ad00b4009800770044002c00550033007200a7006a",
            INIT_3A => X"005f005b00390034001800310077009c00bb00cb00ba009b008d008500740075",
            INIT_3B => X"006d0077008b0099009f00a7009c007d00650041004400400037009000aa007a",
            INIT_3C => X"005e004b00200049002e002100360073009600b000c300c200b1009b00880092",
            INIT_3D => X"008b0065005e00770065005f0060006900830076006b006d0080008f009a006a",
            INIT_3E => X"004e00230018004c00410028001b003b00780088009600b000c000b700a500ba",
            INIT_3F => X"00cf00aa006b0056004200550070008c00a90095008900890096008f009a0080",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY12;


    MEM_IFMAP_LAYER0_ENTITY13 : if BRAM_NAME = "ifmap_layer0_entity13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"004400510040002e00210039004b005000530046001400220047004b00460042",
            INIT_01 => X"00570078007c0079007e006c0054005200880081003b005b00600043004c0057",
            INIT_02 => X"00500066004a002f0038005c005400540058003e00120030005d005c004d0049",
            INIT_03 => X"006b0075006f006a0075006c004d00530097008b002d004100470042005a0051",
            INIT_04 => X"005f006d00580038005400690056005a005c00350014003c005900580042003c",
            INIT_05 => X"00670066004e00540072007200420056009e008f00230037005400620062003b",
            INIT_06 => X"0074006400640049006d006600580060005e002d001a00380041004300360037",
            INIT_07 => X"006a007500610062007600720045005b00a000960040005d0078007e005e0032",
            INIT_08 => X"007800680080005d0072005e005a005e005d0027001a0024002f003700490056",
            INIT_09 => X"00690071006b00650067006d004a006700a200ac00700074008100840067006c",
            INIT_0A => X"0069006600620062005f0059005b004e00580023001b002b004d005d006a006c",
            INIT_0B => X"006700650064004e0039006e0062006600a700ba0082007f0081009000840078",
            INIT_0C => X"005e00600030004f005a0064005d003f004a001d0026005a007e008100820063",
            INIT_0D => X"003a0047007300390025007b0071006a00b700c1008d008c008900a00065003b",
            INIT_0E => X"00560054002f006900670061005e0047003800140049008b008a008c00720029",
            INIT_0F => X"001a00410073004f003b007d0078008c00b000c3009600940090009b003f0018",
            INIT_10 => X"0062004e004a008c009500720050005c0047002c0071009000880086003f0017",
            INIT_11 => X"0045007c005e00560070008b009b00a500aa00b1009600960092008e00290016",
            INIT_12 => X"00740051004e009400a3009b005400450051005a0089008e008a005d00210038",
            INIT_13 => X"007c008f007300800097009c009c008100a700ad0098009a0094007900160018",
            INIT_14 => X"0078004f0049009100a500a6007f004100360072008e007f007e005d0047006c",
            INIT_15 => X"00870085009200a1009c00a50075005700a900af0097009c0091007400130017",
            INIT_16 => X"007b00450042008a00a100a800a5005f004b008c008a0070006d0066008800a2",
            INIT_17 => X"0099009a00970087007c00850076008800bd00aa0092009d009400770014000b",
            INIT_18 => X"006a0039003c0079008700a400ad009800900093007f00760073005c0066008b",
            INIT_19 => X"008d008a008500740078006b0077008800b000ae0087009100a10072001a002b",
            INIT_1A => X"00740055004e0074007f008c00ac00ab0099007c00820078007700760071006e",
            INIT_1B => X"0069006c0077007d0083007a00810075009000a2008d009a00a600700041005f",
            INIT_1C => X"00840060006300780082007200a500a8008b006b00680070007c0081008e0084",
            INIT_1D => X"007a0077006b006f00730076008d0090008e007b0092009f009d00700048005e",
            INIT_1E => X"0079005a005d0076007f007c009700a6009900ab00790045006b007c007b008b",
            INIT_1F => X"009b009000800077007a0067008300a7009f008c008000a00095004b00220068",
            INIT_20 => X"007000640064007e008d0098009500a3008a00a300a6004700640085008b008d",
            INIT_21 => X"0081008800a0009e00a30097007d007e00a900b1007a008f008f003d0033008b",
            INIT_22 => X"00700070008300810093007c00900089008f007900a80099007a007f00920093",
            INIT_23 => X"008d008b0084008a0086008f00990086009100820092007a00860064003a006f",
            INIT_24 => X"007900760095008e008d0061007b0076008f007e007900bb0091006e00880082",
            INIT_25 => X"009a00a10094009a00970086009600910086007b006100570067007700610086",
            INIT_26 => X"008800870097006f007a0065005d007d008600990060007d00a90088009200a0",
            INIT_27 => X"0096009400a600a7008d00800090009100840082004b005e00530057009500a9",
            INIT_28 => X"0094008c0070005e007900680054008200660074008d004a007600a3009b00aa",
            INIT_29 => X"00a50095009d00a70092008900930091007f007c006d007100600077009c00a1",
            INIT_2A => X"009800770048007d00810065006300790078005b009a007d005d009600b500a9",
            INIT_2B => X"00a200ad0091008f008f00870081008b007d007800750066008100ab009a0099",
            INIT_2C => X"008800680052007b00880076006200730096008d007500940081009500ad00b3",
            INIT_2D => X"00a500a8009f008f007e008b008c008d00880085007a006d009800a400960095",
            INIT_2E => X"007d006f009600bf00ac009e0079006f0091009900730069009400a1009a00ac",
            INIT_2F => X"00a1009b009c008d008900930088008f0089008c007b0086009c0095009e0095",
            INIT_30 => X"009500a200c800dc00d100bd00aa00930091007a007d0088008b009f009600a4",
            INIT_31 => X"009b009b009f008e008500a900930088007f007e006b0072009a008f00a0009c",
            INIT_32 => X"008b0089009d00be00d500d700bf00b000a90084007500a300ad0097009a008f",
            INIT_33 => X"007c008100990098009100a30095007c007700830060004a0091009500970078",
            INIT_34 => X"0073006f0061008600bf00cf00d300c100b100ad0091007f0090008f00860068",
            INIT_35 => X"0049005c008b009b00a1008a0094008e008300750055003c00920091006f006d",
            INIT_36 => X"006a007200410040007800b200c300d500ca00b900ad0099008e0096008d007d",
            INIT_37 => X"006c0060008e009a009000a10095007f00830062003100610093006c00760075",
            INIT_38 => X"00740070003e00260029008700b400c700d400cc00b700b200ab00a4009e00a1",
            INIT_39 => X"009d008b0087008d00870099009c007e00670042003b007c0054008800c50083",
            INIT_3A => X"007f007b004f004e00250042009500bf00d000db00d600c200b800b400a5009f",
            INIT_3B => X"0087007d007b0083008a009300870072006c004f0055005b004e00ac00c9008f",
            INIT_3C => X"007d00680034006b00430030004e009700bd00cb00d900da00cd00c300b400b6",
            INIT_3D => X"00a50074005e007a006100590059006f0096008a00820086009f00b500bc0081",
            INIT_3E => X"00660033002800730060003a0029004e00a000b500b900cf00da00d200c400ce",
            INIT_3F => X"00d600b4007c007100560066008400a000ba00a700a700a700b400b300b9009c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY13;


    MEM_IFMAP_LAYER0_ENTITY14 : if BRAM_NAME = "ifmap_layer0_entity14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00320040002e001e0016002400370039003b0036000c0012002b002c00310032",
            INIT_01 => X"003a004d0051004d0053004e003800390061005d001f003a0041002900350042",
            INIT_02 => X"003a00510039001d0023003d003b003c0040002f0007001b0038003e003b002f",
            INIT_03 => X"0044004a004a0044004e00510033003c006f006000150027002d002c00450042",
            INIT_04 => X"004800570046002300350048003c004100450026000700230034004100300021",
            INIT_05 => X"0043004200320037004d0052002d003e0074006300100026003f004b004d0033",
            INIT_06 => X"005e004c0050002f004700480041004a0048001e000c0022002800340023001e",
            INIT_07 => X"004b0057004400450051004d002e00430077006b002a0049005f006000440022",
            INIT_08 => X"0061004f006a003c004b00440048004c00490018000c0011001c00250033003b",
            INIT_09 => X"0048004f004b004700470049002d004d0080008100520055005e006100490050",
            INIT_0A => X"0052004d004b0043003d0045004d003d00430013000d0016002c003b00470049",
            INIT_0B => X"004800480049003500220049003e004d008800930060005b005c006e0068005c",
            INIT_0C => X"0048004600190033003e004f004f00320038000f001800360049004b004d003e",
            INIT_0D => X"002200330060002a001600580048004a009500a10068006c006b00830051002b",
            INIT_0E => X"003f003b00150046004d0048004b003a00290008002f0051004b004b003e0012",
            INIT_0F => X"0006002700590040002a005e00480053008300a2007200780076008500340015",
            INIT_10 => X"004900350031006800790058003900460033001700470053004e004f00220007",
            INIT_11 => X"00280051003c003e00500063005b005d0073008d007800790079007c00210014",
            INIT_12 => X"0056003a003800760083007f00400033003b004000610063005e003a000d001c",
            INIT_13 => X"0053005d0049005000620069005f004a007400840077007e007f0065000d0017",
            INIT_14 => X"005b003b0035007400840087006700300020004b006000610066004a00320049",
            INIT_15 => X"005a0052005900610062006c004700310077007c0077008a007b005b000a0014",
            INIT_16 => X"00650033002f006e0081008700870048002e00540052004f005e005600750087",
            INIT_17 => X"00780066005d005e005c0058004a0058008400730076008d0077005b000b0007",
            INIT_18 => X"0058002800280060006b0083008b0077006b006600570059005f004a0051006c",
            INIT_19 => X"0076006e0064005d006600550057005f007c007800650071007b0059000f0020",
            INIT_1A => X"005f003f0037005c0064006e008b0089007b00610065005c005a005800560056",
            INIT_1B => X"005500580064006c0072006c006e005f006d0075006b0073008000580031004c",
            INIT_1C => X"006a0045004700600068005600860087007400570051005800600060006e006a",
            INIT_1D => X"0062005f0057005c0061006b007f0080007a005e00740077007a005c00350046",
            INIT_1E => X"006000400040005c0067005f0079008500810096006400330058006500620071",
            INIT_1F => X"008300770065005f0060005300710098009400780062007c00760039000d0048",
            INIT_20 => X"0057004c0047005a0073007c00780082006e008e0096003a0054007400770078",
            INIT_21 => X"006c0071008500860089007e0067006e009f00a3006300720075002a0021006b",
            INIT_22 => X"005600580064005d0075006300750069006e0066009b008b006b006f00810081",
            INIT_23 => X"007c0077006d007600710076007c007100830075008300630069004800270057",
            INIT_24 => X"005f006000780073006d004700630056006c0063006a00b00082005e007b0075",
            INIT_25 => X"0089008d008100880083006f007800790075006b00500043004800510043006e",
            INIT_26 => X"006d0070007d0057005800480047005e00640079004900730098007600870094",
            INIT_27 => X"0085008200940095007d00710079007a00720071003a004e003d00380073008a",
            INIT_28 => X"007700740059004300580048003c006600480057006d003700650092008d009c",
            INIT_29 => X"00980088008c00980086007b007f007c006d0069005d0062004d0062007a0077",
            INIT_2A => X"007e00610032005d00600046004b0060005a003b007600610049008300a20097",
            INIT_2B => X"009600a30084007f007d0076006e007500690066005e004f006b008e0070006a",
            INIT_2C => X"0070005100370059005c004e004500590077006b00530076006b007d0097009c",
            INIT_2D => X"0094009b0094007e006c007b0078007500720066005400560081007900630069",
            INIT_2E => X"006200560078009a0077005f0045004e0073007e0057004e007d008b00840096",
            INIT_2F => X"008d008e0092007e007900840076007b007300580052006f00790065006a0067",
            INIT_30 => X"0074008800a700b6009f00770060005c0066005a0066006f007000880083008f",
            INIT_31 => X"0086008e009600800075009c0084007700660059004e0053006a00600071006c",
            INIT_32 => X"006c006d0071009200a6009e007b0069006600520055008c0091007e0086007b",
            INIT_33 => X"00680073008a008900830096008a006a0061006f004a002d006000650069004b",
            INIT_34 => X"0058005500370056008b00970097007e0068006800570057006f006e006e0052",
            INIT_35 => X"0035004b0079008c009100780081007a00740062003e00200061006200410040",
            INIT_36 => X"0052005c00220020004b00750086009c008d006d006200570052005a005b005f",
            INIT_37 => X"005200460079008b0081008f0080006b0071004e001d003f0063004700470042",
            INIT_38 => X"005a00560023000d000f004e0072009400a2008b006f00620061005b00560071",
            INIT_39 => X"0078006a0073007e007600870087006a004f002a0026005b002c006000990053",
            INIT_3A => X"005c0056002d0025000d001f0057007a009600ad009e007a00750072005d005c",
            INIT_3B => X"004d005500670071007e00850073005b004e0032003b003c002a006c00860062",
            INIT_3C => X"005200470018003800240017002300540076009200a500a500960082006f0079",
            INIT_3D => X"006c0042003f0062004e0045004600560075006c0060006200780074007b0059",
            INIT_3E => X"0041001b001100400034001d000f0025005900640074009600aa00980088009c",
            INIT_3F => X"00a600790045004a002f00470066007f009c008b008300820093008800920075",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY14;


    MEM_IFMAP_LAYER0_ENTITY15 : if BRAM_NAME = "ifmap_layer0_entity15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00b3008b004d0058008d009d009c0097009c009e009000970097008800790076",
            INIT_01 => X"007e006c0054005400620062005e0053005a00560054006000750057004c004d",
            INIT_02 => X"00b8008500800092009f009f009e00a700a500a20099009a009600960088007d",
            INIT_03 => X"0081006d005a0052005d0062005e0058004e004c005b006a00760062005b005a",
            INIT_04 => X"00b4009800b000aa00a40098009b00a400a200aa00a2009f009c00970092008c",
            INIT_05 => X"0092007c00580047005500620067006b0065006d006f006f006f0065005d005f",
            INIT_06 => X"00af00ae00b800b500a8009800a400a300a600b300a700a800ae00a2009f00a4",
            INIT_07 => X"009700890059003a0048005a0063006b00750080007d007900690061006d006f",
            INIT_08 => X"00af00ae00a700ac00a200a100b000af00b200b200b300b400b000a800a000a4",
            INIT_09 => X"00ad009c007800450042005a0063005e0069007c007f007b0070006800710074",
            INIT_0A => X"00b500ae009000aa00a900a600b000b300b400b400b400b500b000ae009f0096",
            INIT_0B => X"00b500af009b00740060007d0083007000750078007a0079007900780076007c",
            INIT_0C => X"00c0009c008a00b200af00ae00b000af00b800b400ba00b800bb00bb00ad0099",
            INIT_0D => X"00a600ad00ad00a7009600950094007900730075006d006f0078007a007b0080",
            INIT_0E => X"00b9007d009c00ab00ad00af00af00b800bc00b700c100c200bd00b900b800a6",
            INIT_0F => X"00a400ac00b100b000aa0089008f007a006b006e0060006700750076007b007d",
            INIT_10 => X"009b0095009f00a000ac00ad00b200b400bb00ba00ba00bf00bb00af00ac00a0",
            INIT_11 => X"009a009700a600b000b7009b00a6008500680068007000770076007a007a007d",
            INIT_12 => X"009a0098009300a900b200b200b700aa00b000bc00c600c100ae00a700a500a9",
            INIT_13 => X"009d008c009200a900b300a000ab008d005f0068007500770074007b0076007d",
            INIT_14 => X"00860070009f00b100ae00b800b800ba00ba00c200bf00b0009b009e00a700bb",
            INIT_15 => X"00ae00930086009700a0009c009b007c004a006600690066006b0075007b007f",
            INIT_16 => X"0041005b00ae009d009300b100bf00be00bc00b000ac00b000b800ae009400a3",
            INIT_17 => X"00b0009a0085009500980095008300500042006100670066006700710078007d",
            INIT_18 => X"0015005c00bf00b100bc00ca00bd00b600b3009c00a500bc00c800ae00980072",
            INIT_19 => X"005f007f00780089009700880072004e00400049005900620062007100750076",
            INIT_1A => X"002c006300a800ad00c800c300bc00bb00a5009500b400c200b900a800a8009a",
            INIT_1B => X"006b00920091008a009c007f0064004800390040005300600062006a006c006f",
            INIT_1C => X"006900760075009f00c400be00b400bb00ad00ad00c600c100ab00a500b400bc",
            INIT_1D => X"00ae00bb00ad00b300a0008000690048004300450057006c0063006400610066",
            INIT_1E => X"008a00710068009d00c600c400b400a800b400bf00cb00cd00d200bf00c400c8",
            INIT_1F => X"00c000bb00bc00be00a800990071005000460040006000870078005a005a0062",
            INIT_20 => X"0096008a0073009300be00bb00b0009600ab00c700d300c600d300c200be00cb",
            INIT_21 => X"00bf00ba00b800bd00be00a600640046002f0038006a008f0095005c004a005e",
            INIT_22 => X"009b009b009200a500bd00c000bf0091009c00d200a9009500c000c200b200a8",
            INIT_23 => X"00a900b500aa00a7009a00750043002b002200310068008f009c006a003f0050",
            INIT_24 => X"00a500a2008a00a600c400be00ba0089007400c9009d00a900d200b60080008f",
            INIT_25 => X"007c0093007f006100520038002f0033002b00400069009d009d007b00390041",
            INIT_26 => X"00a900960078009e00be00be00be0098003c009900bc00b900c300a5009000ce",
            INIT_27 => X"00b100890065003d00370033004700500037004a006e00a000b0008e00360032",
            INIT_28 => X"00aa00a0009600a600ba00bc00ba009a00200031007e0092009b008c008c00c0",
            INIT_29 => X"00cc009c0061003e0049004900520057003a003e006b00a600bc00a700480033",
            INIT_2A => X"00b200ab0097009c00b500b200a3007c0024001d00280037004e006300650082",
            INIT_2B => X"0090007b005f003700340033003c0055004e004d0066009900bb00b100590037",
            INIT_2C => X"00b500ab0092009800a900a700950069004f005e0042002e002f0047005c0078",
            INIT_2D => X"005a00370038002900230022001e0037005200560061007700ad00ae006a003c",
            INIT_2E => X"00b1009c009e00a3009c00a000940089008f00760066006b006e006d007d0067",
            INIT_2F => X"002f0011001000130018001c000e0013002b004100600063008c00ad00850043",
            INIT_30 => X"009e008b00a700b60097008c00ab00c000ac0074008500880092008d007f0065",
            INIT_31 => X"004100250020001900180011000a000f001400420061004e00620094009c0069",
            INIT_32 => X"00a000a400ae00ab009e0088009400b100b8009300a90097007f008b008e007d",
            INIT_33 => X"0067004d003f002b002100180011001a001f003e004800320048005a00780088",
            INIT_34 => X"00a000a300a700a700b100a8008c007800ab008f00760082007b009c00a60091",
            INIT_35 => X"007c0069005b004e004c00420038004300460041004100490064007b0051006a",
            INIT_36 => X"009c009f008c009300b400aa0099007b008b009c0073007e0083009e00a800a2",
            INIT_37 => X"007f0077007b00780070006800690077007400690068006d007a0086005c0068",
            INIT_38 => X"00a4009e007b008b00ad009c008d008c008d0079008200a10097009d00a600a8",
            INIT_39 => X"0090008a008f008400810085008a0094008f0089008600840078006400730093",
            INIT_3A => X"008e0095009000a800a700a1009e009e00a50090009700a900a100a0009e00a2",
            INIT_3B => X"009900910089007f008d00950096009e009f00960094008f007b0077008b009f",
            INIT_3C => X"009800a600b300b900a700a700aa00a800a700a400ad00b200a9009d00890085",
            INIT_3D => X"0092008f008c0088008c00970098009d00a6009c009900900085008300900099",
            INIT_3E => X"009f00b200b700ab008b007d0091009f00a2008b0095009c009e009800830073",
            INIT_3F => X"0084008e0094008f0090009d009c00a100a7009f0094009c009c009600990098",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY15;


    MEM_IFMAP_LAYER0_ENTITY16 : if BRAM_NAME = "ifmap_layer0_entity16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"007600600031003b0060005f00540053005f00610053005a005c0052004b004f",
            INIT_01 => X"005b0050003b00320037003800380033003c00380033003a004c0035002f002f",
            INIT_02 => X"0082005800590069006c0060005d006800650062005a005b00540057004f0048",
            INIT_03 => X"00520048003d00320037003800370033002b002800350041004b003d003a0039",
            INIT_04 => X"008400680081007a006c0059005f006a006200690062005e00550050004f004c",
            INIT_05 => X"0055004c0036002a0033003a003f0042003c0042004300420043003e00380039",
            INIT_06 => X"0081007f008800840070005a0068006900650071006500660067005a0057005d",
            INIT_07 => X"004f004e0033001f002a00330039003e0046004d004b004a003c003700430045",
            INIT_08 => X"0080007f0079007f006d006300720072006f006f00700071006c00630059005c",
            INIT_09 => X"005e0059004e002c002700340038002e00350043004700490042003b00450047",
            INIT_0A => X"008900830068007f0076006a007100740073007500740071006d0069005a0054",
            INIT_0B => X"006a00680067004f003a004d0052003d003e003f00430046004900480046004b",
            INIT_0C => X"0098007700660087007a00750073006f0079007b007c0070007300710066005c",
            INIT_0D => X"00640065006d006e005c0057005b0043003e00400038003b00450048004a004e",
            INIT_0E => X"009300590078007e00780076007200790080007a007c00730073006d006c0064",
            INIT_0F => X"00650068006d006a0066004b00570048003b003c002e0035004200440049004b",
            INIT_10 => X"0076006f0078007200770074007500770080007a006f006d007300670061005e",
            INIT_11 => X"005e005900610064006d005f00720059003e003a00400047004600480048004b",
            INIT_12 => X"0077007100690078007c007a007b006f0076007b007d00790076006d0065006f",
            INIT_13 => X"0069005500520060006a0064007a0067003d003e004700490047004b0044004b",
            INIT_14 => X"006400480072007e0078007f007c007e007f00810080007b0079007700780090",
            INIT_15 => X"00830063004f0058005f0061006c005b002e003e003d003b004000460049004c",
            INIT_16 => X"00220034007f0069005d007a00840083008100730078008c00a6009700740085",
            INIT_17 => X"008d006e005600610060005c00560031002a003c003e003c003e00420045004a",
            INIT_18 => X"00040040008e007d008c009a008c0084007f006b007b009c00b2009300770053",
            INIT_19 => X"0040005b00530064006f005c004d00310029002f00370039003b004300420044",
            INIT_1A => X"00180048007a007b009c0096008f008d0077006a008f00a00097008100800077",
            INIT_1B => X"004d00740073006d007b005a0044002d0023002b00330037003b003e003a003e",
            INIT_1C => X"00450052004a0070009600910086008f0083008400a1009c007d007200850097",
            INIT_1D => X"009100a0009200980081005d004b002f002f003000380044003c003c00360039",
            INIT_1E => X"00570041003b0070009800960086007d008f009b00a700a5009b0084008f00a0",
            INIT_1F => X"00a2009e009f00a100890078005400390033002b0040005f0051003700360039",
            INIT_20 => X"0058004e004000660090008d0081006c008b00a500af009d009e00860086009f",
            INIT_21 => X"009a009400930098009a008700490031001e0023004b0067006f003d002c0039",
            INIT_22 => X"0056005700570074008f009300910069008000b30085006c0091008b007a0079",
            INIT_23 => X"007d0087007c007900720058002a00180013001d00490066007500500027002e",
            INIT_24 => X"005c005c004d0076009c009900910062005c00aa0074007a00a50083004b0062",
            INIT_25 => X"004c0061005500400036001b0011001b001a002800450075007f006400240028",
            INIT_26 => X"005e0054003c006e009c00a3009b00730027007c00940089009500710057009c",
            INIT_27 => X"00780050003d0027002700180022002e001f002d004500780099007b00220020",
            INIT_28 => X"0061005d00590072009600a200980075000d001d00640074007300560049007c",
            INIT_29 => X"0086005b002f001b00310032003100320019001e0042007d00a2009600380020",
            INIT_2A => X"006a006800570063008d009600810057000f000b00160025003600390029003e",
            INIT_2B => X"005300480036001a00200023002200330028002b003e0070009b009e004a001f",
            INIT_2C => X"00700068004f005a007b008900730042002f004200280017001b0026002c0045",
            INIT_2D => X"0036001f0026001d00190016000f001f00310033003a004e008600940057001f",
            INIT_2E => X"006d005800590060006900810073005e006100470036003c0042003e004b003c",
            INIT_2F => X"001a000a0009000e00110013000b000c0017001f003a003b005e008800690023",
            INIT_30 => X"005b00460060007000600068008900930075003a00450043004a0045003f0035",
            INIT_31 => X"002900190013000d000c0009000d0012000c0024003e00270034006800790047",
            INIT_32 => X"005b005c006200620061005600690086008e006b007c006100440049004e0049",
            INIT_33 => X"003e002b0026001c0016000e000b00140014002a003000140025003800580064",
            INIT_34 => X"005b005e006100620071006f005b004c0084006e005000510047005f00630054",
            INIT_35 => X"0048003d003800330035002b0020002b002e0028002500280040005a00300042",
            INIT_36 => X"00570060005000520071006d00620048005c007300450046004a005e00600058",
            INIT_37 => X"00450047004c004a0042003c003d004b00490040003f0041004c005e0036003a",
            INIT_38 => X"006000610043004c0069005a004e005000570048004c00620057005c005d005a",
            INIT_39 => X"004f00540055004600420048004d0057005300520050004f004300350046005e",
            INIT_3A => X"00490054005100650061005b0058005b00690059005b00630059005d005d005a",
            INIT_3B => X"005800550049003c004900520054005b005d0056005700550043004400570064",
            INIT_3C => X"00530060006a00710060005f0060005f00660069006d0068005b005a0052004a",
            INIT_3D => X"0052004e004d004a004d00550057005c00640059005a0054004e004d0057005a",
            INIT_3E => X"005c006b0071006800520042004d005c005f0051005b005a0058005b004d003d",
            INIT_3F => X"0046004d005600520053005c005b00600065005c0057005b005c005a005b0057",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY16;


    MEM_IFMAP_LAYER0_ENTITY17 : if BRAM_NAME = "ifmap_layer0_entity17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0053003d001a002400410043003a0036003f00410034003b003e0035002e0034",
            INIT_01 => X"00470041002b0027002f002f002d0026002f002d002a00320045002e00290029",
            INIT_02 => X"00610035003a0046004600430044004d0044004100380039003400390032002e",
            INIT_03 => X"003c0034002b0026002f002f002c00280020001e002b00380043003500330031",
            INIT_04 => X"00640047005c0051004400390044004e00400047003f003b0034003000310030",
            INIT_05 => X"003b00320021001e002b003000350038003300380039003800390035002f0031",
            INIT_06 => X"0060005f0061005900490037004900480041004e00420042004300370036003f",
            INIT_07 => X"002f002e001a001200220029002f0035003d00440040003e0030002d003a003c",
            INIT_08 => X"005c0061005400570049003f004c004b004a004a004b004b0043003b0035003b",
            INIT_09 => X"003b00340033001e001f0029002e0027002e003b003d003d00340030003a003c",
            INIT_0A => X"006500660047005900510046004c004c004c0051004e00470044004300350031",
            INIT_0B => X"0043004100480039002b003e00420032003800360038003a003c003d003c0041",
            INIT_0C => X"0078005900490063005300500051004b0051005700550042004c004f00430035",
            INIT_0D => X"003c0040004a004d004100400041002f00350036002d0030003a003d003f0042",
            INIT_0E => X"0075003b005b005b00510051004f00540057005600560048004d004c004a003f",
            INIT_0F => X"00420049004c00490047002f0038002f002c00310023002a00370039003e0040",
            INIT_10 => X"005c0054005b00510053004f005000500058005300490046005100480043003d",
            INIT_11 => X"0043004100460046004f0040004f003c002c002d0034003b003a003d003d0040",
            INIT_12 => X"00610058004c005a005b005600530047004f00520054005300580053004d0055",
            INIT_13 => X"0051003e00390046005000480059004b002b0031003a003c003a003f00390040",
            INIT_14 => X"00510030005600620059005b00520054005b005400500050005e00650067007e",
            INIT_15 => X"006b004900370043004b004c0051004400200031002f002d0033003a003e0041",
            INIT_16 => X"0014001f0063004d00400056005a005a005f00450045005f008f008800670079",
            INIT_17 => X"00760052003f00500052004d00420021002100300030002e00300036003b003f",
            INIT_18 => X"000000320070005c006e007a006900620060004800540077009d007d005f0049",
            INIT_19 => X"00340047004100540060004f0041002a0025002500290029002d00380039003a",
            INIT_1A => X"0014003c0061005c007d00780070006f0059004c006e0080007f00640062006c",
            INIT_1B => X"004400630062005b006a004c003a00290021002300250026002e003400320035",
            INIT_1C => X"003b0046003a0058007b0075006a0073006600670082007d005f005000660089",
            INIT_1D => X"0083008c007e0084006f004e0040002a002b0028002a0032002f0032002e0031",
            INIT_1E => X"004900350032005e007e007c006c00620072007d008a0088007b00620071008c",
            INIT_1F => X"008f0089008a008c0075006900490033002f00230032004d0043002d002d0032",
            INIT_20 => X"00480041003a00560077007500690053006e0089009300820082006b006d0087",
            INIT_21 => X"0084007f007e008300870077003d002a001a001b003c00550061003300240033",
            INIT_22 => X"00470048005100660078007c007a005000630097006a0054007c00790065005c",
            INIT_23 => X"0063007300680065005e0048001f0011000e0015003a005500680046001f0029",
            INIT_24 => X"004f004e0044006400860088007d004b00470093005b0061008e007100370048",
            INIT_25 => X"0035004f00450032002a0014000d00160014002300370060006f005b001e0023",
            INIT_26 => X"005100480032005800870099008a005d001f006f007f0071007c005c0047008d",
            INIT_27 => X"0067004100330021002400190024002c001a002b0036006000890073001e001a",
            INIT_28 => X"00530052004f005f0082009600860062000a0017005600630065004c00420074",
            INIT_29 => X"007a004e00270017002e002f002f002e0014001b0034006700920089002f0019",
            INIT_2A => X"005c005c004e0053007b0087006e0046000c00080010001d002f003400250038",
            INIT_2B => X"00460039002b00120019001c001d002c002100260031005e008c008d003d0018",
            INIT_2C => X"0061005d0046004e006b0076006000300025003a002200130013001f0026003b",
            INIT_2D => X"00270013001b001200110011000a0018002a002c003000400078008000460018",
            INIT_2E => X"005e004d00520058005b006b005f004b004a003700300039003a003500430033",
            INIT_2F => X"0010000400030008000e001300070006001100170030002f005100730057001b",
            INIT_30 => X"004b003b00570069005300520075007e005500220039003e0042003d0039002e",
            INIT_31 => X"002400170012000d000f000e000c000e0007001c0036001e002800550068003e",
            INIT_32 => X"004d004d005100560055004500570070006f004f0064004f003b00430045003a",
            INIT_33 => X"00330026002000150011000c0006000e000f00220029000f001f002e004c005a",
            INIT_34 => X"004f00510052005500650060004a0039006d0057003a003e003d0058005a0044",
            INIT_35 => X"003b0035002f002a002c0023001800230026001d001b001f0039005200270038",
            INIT_36 => X"004c0057004a004a0066005f00530039004d00630037003a003f00540057004d",
            INIT_37 => X"0039003c00430044003b00310031003f003c003100300033003f0054002d002f",
            INIT_38 => X"0055005a00400045005e004e00410044004c003c0042005a004a004e00530051",
            INIT_39 => X"00430047004c0040003b0039003e0048004400420040003e00320029003d0053",
            INIT_3A => X"003d004b0049005c00570051004e0050005d004c00500059004a004c004e0050",
            INIT_3B => X"004a0045003e0035004000420044004b004d00480048004400320038004e0059",
            INIT_3C => X"00460051005a0064005600550057005500560057005d005a004a0046003f003c",
            INIT_3D => X"0042003c003e003e004100460047004c0055004d004e0047003e0041004d004f",
            INIT_3E => X"004f005d005f005900460039004600510053004000470047004a004c003d002f",
            INIT_3F => X"0038003f004800460045004c004b00500056004f0049004e004f004c004f0049",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY17;


    MEM_IFMAP_LAYER0_ENTITY18 : if BRAM_NAME = "ifmap_layer0_entity18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00a000b900d100d900e600f600f900f600f800f300e600dd00da00dd00d800c7",
            INIT_01 => X"00bc00bb00b800b400a600900079008b006a00660066004f005e0065005b005e",
            INIT_02 => X"00e100ef00f200e600e800f500f300eb00ed00e600d800cd00c900cb00c800ba",
            INIT_03 => X"00af00ab00a1007f008e008d007a00870076005200250034005f006b00610064",
            INIT_04 => X"00fc00f900f100dc00d900e200df00d600d500cf00c300b800b300b600b300a7",
            INIT_05 => X"009f0098009400810080008c0080007200570028000400260063007300690069",
            INIT_06 => X"00e900e100de00d300d300cb00c800c000bb00b700ae00a400a000a500a00099",
            INIT_07 => X"0091008d008c008a007d007d007f0069003b0025001a0037007000780070006d",
            INIT_08 => X"00cf00c300cf00c900be00b400b300ab00a3009f00990092009100970093008d",
            INIT_09 => X"00870088008300870081007a0084005a003a003d00300056007500780072006d",
            INIT_0A => X"00b600ab00aa00a20099009c009f00970090008d008c008a008b008d008a008a",
            INIT_0B => X"0087008c0086008a008c008900660045004b003e00430074008100800070006e",
            INIT_0C => X"008d00880088008600880086008c008500870089008b008d008f0092008e0091",
            INIT_0D => X"00910091008a008f008e006b002f00210048004b006c007f00840084006f0070",
            INIT_0E => X"0076007d0080008100880083008a00840088008c009000930096009e009a0099",
            INIT_0F => X"009200950093009400800042000d0011005000750080007a007b008000720070",
            INIT_10 => X"0073007e00840085008b0087008f0089008b0091009500980094009a00a300aa",
            INIT_11 => X"009e00a2009d00940073002c000e001e0069008b0088007e0077007a0074006f",
            INIT_12 => X"0076008000880088008d00880091008d008d0093009a00a5009d009a00a200a7",
            INIT_13 => X"009b00930091008a00630038002e0037006d007c007a007e007300740075006e",
            INIT_14 => X"007d0084008b0089008e00880090008c008b0090009600990083008b00900098",
            INIT_15 => X"00a600ba00d300d60080005c0045002a0055005f006300730070006f0071006b",
            INIT_16 => X"00850089008e008a008d0088008e008a0089008f00880084008e00b600c900cb",
            INIT_17 => X"00d200ce00cf00c000a200bd0092002a001b002800670072006d006a006c0068",
            INIT_18 => X"008c008b008f008b008f008c008a008900870085009000a400ab00a000890073",
            INIT_19 => X"006a005d004b003b006f00dc00c9005f000d0007003e00740063006500690064",
            INIT_1A => X"0090008a008f008c009200920082008700820091008c006e005e005c00310013",
            INIT_1B => X"001d003200190012007800d100d2009d0026000600130044004500520063005f",
            INIT_1C => X"0091008b0092008e0090008e007900800085007f0054004400560052002e0016",
            INIT_1D => X"00130032001e004100af00c900cd00cb006600100012001600230038004f0058",
            INIT_1E => X"008f008b00940090008a0084008b00830075004200480056006a004e00280022",
            INIT_1F => X"00240046007300b600cb00c500cd00c3006c003d002500120018004f00640053",
            INIT_20 => X"008e008b00930090008500720084007900510059003c0045005500440053009b",
            INIT_21 => X"00c000db00ed00eb00d700d700d300720030005d003500140041008b008f0054",
            INIT_22 => X"008f008d008e008900740045003a00430051004b001d001c00240019008c00f2",
            INIT_23 => X"00ec00eb00e300dc00db00df0095003a00390054004e004e008500a100a7005b",
            INIT_24 => X"008f008c00880086008d0047002d00340043002100170016002f0029009b00d9",
            INIT_25 => X"00c700be00bf00d000dc00df00ad0067005d0073008700950098009400a50059",
            INIT_26 => X"008f008c007e00b500bd004c0021002b003900150010001700390042009e00c2",
            INIT_27 => X"00b600b300c400c900c200ce00de00b30097009c009500970096009200880042",
            INIT_28 => X"008c0085009a00ea00b5005a0026002a0034000b000b000b0014003100a000ba",
            INIT_29 => X"00b000b900b900730045005a00a100c400b700aa00a0009900930088004d0026",
            INIT_2A => X"0082008000a300a3008b006a002d002e001c00030009000f001e003600a200b4",
            INIT_2B => X"00ac00be00710015001400150030009500bb00ab008e00850080004300150027",
            INIT_2C => X"007c00840067001a0048006c0034003000120007000b003b005a006300a500b0",
            INIT_2D => X"00b100a9002a001d002f0026000e00460095008800750075003c000e00150030",
            INIT_2E => X"0079007c0049001e003b00720044001f000d000e00180048004f006c00bb00bb",
            INIT_2F => X"00bf008b001b002b001e001b001c001b006c0084007b005900160015002a003b",
            INIT_30 => X"006d00660047003f003c0071004d001c0010001f003000470046008800bd00b3",
            INIT_31 => X"00b40074001f003600350029001b000e00480085007c003c001200220032003b",
            INIT_32 => X"00570051003d003c003a0069004b00150014002e004c00600061009100a400a3",
            INIT_33 => X"00aa00710020003900470031002500110029006c00600021000c001d00280032",
            INIT_34 => X"004900490040003c0039005f0057002f003d0062008900a500a900b000b700b6",
            INIT_35 => X"00b6007c002200360060005c0033001b00110046003b000c00060012001d0028",
            INIT_36 => X"004900490045004e004100590045002f0034003c004a0056005b006000620060",
            INIT_37 => X"006200530020003c003b003e001d001400040011000a00030007000a00110021",
            INIT_38 => X"004b005300480036002d0027000f0004000300020005000700070008000a000b",
            INIT_39 => X"000b000d000800420043002f0038000f00020002000100030006000a000f0020",
            INIT_3A => X"005000590051002f0015000a00100019000e000a000e000e000e000e000e000c",
            INIT_3B => X"000a000900060017003e0048002a000700030004000500050007000b00150021",
            INIT_3C => X"0049004f00490037002e002f003b003a001a00110019001c001f0020001d001c",
            INIT_3D => X"001800150010000c00140016000800060008000700080008000b000f001b001f",
            INIT_3E => X"00450048004c004e005800530048003800200026002b002a002f003300320031",
            INIT_3F => X"002c0026001e001c002200220013000c000e0010000f000d0012001a001e001d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY18;


    MEM_IFMAP_LAYER0_ENTITY19 : if BRAM_NAME = "ifmap_layer0_entity19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"002500310039003a0042004e0050005100560052004900420041004300430038",
            INIT_01 => X"0032003200400073003400380032002700160022002e0024001d001200150013",
            INIT_02 => X"00430048004d00440043004a004800420044004000390034003200360037002e",
            INIT_03 => X"0029002a0027002900280023001e00210022002e001e001b001c001500160012",
            INIT_04 => X"004800440048003e003a003d003800310030002d002b00280026002a002b0026",
            INIT_05 => X"00220023001e001c00230021001f002200300022000d000e0015001400130011",
            INIT_06 => X"00380036003d003c003e0030002b00240023002300220020001f002100220020",
            INIT_07 => X"001d001e001b001d0020001c001d0025002a0012000b000f0016001300100011",
            INIT_08 => X"003900390042003b003400240020001b001c001d001c001a001a001a001c001e",
            INIT_09 => X"001c001c001c001c001c00300043002a00190012000d0019001b001f00130011",
            INIT_0A => X"003b003a002f0021001a001a0019001600170019001a001900180018001b001f",
            INIT_0B => X"001d001e0021001e0021005d005e003c0029001b001e002c002b002d00180013",
            INIT_0C => X"0022001c001700140016001700160015001600160019001a00180019001d0023",
            INIT_0D => X"0020001f0023001e003300590037002500380028002b002d0024001e00170015",
            INIT_0E => X"0011001100100012001600170016001600180017001a001b0019001b001d0027",
            INIT_0F => X"0028002d00330030004100400012000b00220025001f00200019001600160015",
            INIT_10 => X"0011001200120012001500160017001700190018001c001e002500380033003b",
            INIT_11 => X"003b003a00370036003d002800110010001a00190018001b001a001700150014",
            INIT_12 => X"001300120012001200150014001600180018001900200031003e004c00390034",
            INIT_13 => X"0031002e0032003a003800310030002c00290023001900190019001800140014",
            INIT_14 => X"00140012001300120015001500150017001900190024003500310042003e004a",
            INIT_15 => X"0068008900a600b8007c0068004b00210038003d002600190018001900120013",
            INIT_16 => X"001500120014001300180018001600180019001d001f00300055009700b200be",
            INIT_17 => X"00cd00cd00ca00c500b200d00098001600180025004600280015001600110011",
            INIT_18 => X"0014001400160015001800180019001a00190020004200700090009b008c0075",
            INIT_19 => X"006400580047003d007500e800d5004e000f000a00320046001a001500110010",
            INIT_1A => X"0014001600190016001700170019001a001a00480067005b0050005600340012",
            INIT_1B => X"00110022000f0010007c00dd00e0009b002400070016003b0021001300120010",
            INIT_1C => X"00180017001b0016001800190013001500370055003a0029003d004e00320018",
            INIT_1D => X"000b002b001e004900bf00d800d100cd0067000e00100017001b001600140012",
            INIT_1E => X"001a0016001a001700190025003c0034004c00340038003b0050004d002e0026",
            INIT_1F => X"00230049007c00c400df00d800d900d2007600390015000e001f0047003e0011",
            INIT_20 => X"0019001400190017002100350060005c0049005d003e004200510047005a00a2",
            INIT_21 => X"00c400df00f500f500e300e400de00790025003b001100090048008c00750013",
            INIT_22 => X"001900150018001a0028002c00350045005800520025002900310020009400fb",
            INIT_23 => X"00f600f200e900e200e100e2008b001f000b001900280043008500a200970022",
            INIT_24 => X"0016001300160026005d0046002e0036004b00260018001b0038003100a300e3",
            INIT_25 => X"00d600cd00cb00da00e500e400a3004a0039005a008000950097009600a00033",
            INIT_26 => X"0013000f0026007c00af005a0024002a003f0017000b00150040004f00aa00d0",
            INIT_27 => X"00c700c500d300d600ce00d900e300b1009800a800a700a2009a00970088002a",
            INIT_28 => X"0012000a006500dc00be006f002f002e0039000a0009000e001f004200b100cc",
            INIT_29 => X"00c200ca00c6007c004f006600ac00d300c800b800b100a9009c008c004a0011",
            INIT_2A => X"000e0014008400a50096008000370034001e0003000a0016002d004800b400c6",
            INIT_2B => X"00be00cd007b0019001a001e003800a300ca00b8009e009300880044000d0011",
            INIT_2C => X"000a00230053002100530082003e00350013000700100048006c007500b700c2",
            INIT_2D => X"00c300b7002f001e0031002b0014004f00a10094008400810040000a00090018",
            INIT_2E => X"000a00210037002300460088004e0024000f0011002200580061007e00cd00cd",
            INIT_2F => X"00d000980020002b0020001f0020001f00750091008a00630017000c00190021",
            INIT_30 => X"000a001500360041004700880057002100150027003f00570056009a00cf00c5",
            INIT_31 => X"00c60081002500380037002c001c000f004d0093008b0043000e0014001c001f",
            INIT_32 => X"0007000e002f003e004500800056001c001e003c005e006f006f00a200b600b4",
            INIT_33 => X"00bc007f0029003c004b00350023000f002c007a006f00260007000d00100016",
            INIT_34 => X"000b00110027003b004600750068003d00510079009f00b700b900c300c900c7",
            INIT_35 => X"00c60088002a003c006600620034001c0015004f0045001000030007000c0016",
            INIT_36 => X"00130014001d0043004900670055003c00450050005b0064006800710071006d",
            INIT_37 => X"006d00590025004100400042001f001700080014000e000500060006000b0018",
            INIT_38 => X"0017001c001d0025002c002c00160007000a000a000c000c000d001000110010",
            INIT_39 => X"000f000f000900430044003000380010000400030003000400060009000e0019",
            INIT_3A => X"002100250027002000170012001900200017001500170017001700150013000f",
            INIT_3B => X"000b000a00070018003e00470029000800040005000500060009000e0018001d",
            INIT_3C => X"0023002500290032003c00430051004d002c0024002d00300031002c00270023",
            INIT_3D => X"001d001b0015001000170019000a0009000b0009000a000b000e0014001f001e",
            INIT_3E => X"002a002a003b0057006d006f006600520037003e00450047004a004800460043",
            INIT_3F => X"003b0033002b0029002f002c0018001200140016001500130016001c0020001e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY19;


    MEM_IFMAP_LAYER0_ENTITY20 : if BRAM_NAME = "ifmap_layer0_entity20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000d000b000e000a0009000a0005000200030003000100020004000600050000",
            INIT_01 => X"000100000023005600160017001d0008000d001b0027001d0013000800060005",
            INIT_02 => X"000d000c000a0004000700080003000000040002000100010002000400040001",
            INIT_03 => X"000100010010001300070006000600070021002e001700160013000800040006",
            INIT_04 => X"0007000400030000000400040001000000040004000400040004000600050003",
            INIT_05 => X"00040003000c0009000400070006000a00280023000d000c000f000600030006",
            INIT_06 => X"000100030008000b001200040003000300050006000800070008000900060006",
            INIT_07 => X"00070005000a00090004000a00100017001e00160011000e000f000600050008",
            INIT_08 => X"000c0013001d001a001700060007000800070008000900080009000a00070008",
            INIT_09 => X"0009000700080007000800250040002700100010000e0015000e000f000d0009",
            INIT_0A => X"0018001e0016000c0009000600090008000500050009000a000b000a00070009",
            INIT_0B => X"000a000b000b000700140055005d003b0022000e001300200017001b00100009",
            INIT_0C => X"000c000b000a000700080008000a000700060005000a000e000d000c000a000c",
            INIT_0D => X"0009000e000e000700250056003c00280035001c001c001c0014001000060007",
            INIT_0E => X"0003000600060007000b000a000c000900090008000c000e000e001200100013",
            INIT_0F => X"00100015001a00160031003e0014000a001e001a0010000d0009000800040007",
            INIT_10 => X"0007000a00090008000b000a000e000b000d000c000e000f0013002400220028",
            INIT_11 => X"00240020002200220033002b000f00090014000c0009000a0008000800080008",
            INIT_12 => X"000c000c000b0008000c000a000e000d000e000e001400220027003100280026",
            INIT_13 => X"0020001b002700320036003b0034002600230015000b000c00060009000b000a",
            INIT_14 => X"000c000b000b0009000c000a000d000d000d0010001b0028002000320032003f",
            INIT_15 => X"0058007700a100b4007900710054002200320031001d00110009000a000c000a",
            INIT_16 => X"0009000a000e000b000e000c000d000c000c001200180027004d009300af00ba",
            INIT_17 => X"00c800c800d200ca00b100d5009e001c0013002200460025000a0009000b0009",
            INIT_18 => X"0008000a000f000d0010000e000d000e000c0018003e006c008e00a20093007d",
            INIT_19 => X"006e005e0054004a007e00f100d70054000c0009003400490019000d00090008",
            INIT_1A => X"000b000b000f000e00110010000c000e001400440067005d0056005f003d0019",
            INIT_1B => X"0016002300110017008900eb00eb00a7002a0007001700420028001100090007",
            INIT_1C => X"000f000d0012000e00100012000b001200360053003b002e004400530037001b",
            INIT_1D => X"000c0027001c004c00c800e800e700e0007300160013001a001f0016000d0008",
            INIT_1E => X"0010000d0013000e000e001e00390037004f00350039003c0052004e00320029",
            INIT_1F => X"00230047007c00c800e700e600ec00dd007e0044001a000e00200049003f0009",
            INIT_20 => X"0011000e001300110018002f005d005c004f0062003c003d004c0047005e00a6",
            INIT_21 => X"00c600e200fa00fc00ed00f000e7007c002a004a001c000c004c0095007e0011",
            INIT_22 => X"00120010001200150024002a003800480060005800240024002d0022009a0100",
            INIT_23 => X"00fa00f900f400ed00ed00ee009600270015002e003b004d008e00ae00a30026",
            INIT_24 => X"0011001000100022005c0049003c00420054002c001c0021003e003700ae00f0",
            INIT_25 => X"00e100d900d900e700ef00ee00b100560045006a009200a400a400a100a90037",
            INIT_26 => X"000d000a0020007d00b40062003500380048001c000e001b0049005900b900e0",
            INIT_27 => X"00d500d500e400e300d700e100f200c000a500b400b500b000a6009f008d002a",
            INIT_28 => X"000c0007006500e500c9007b003e00390041000f0009000f0026004f00bf00da",
            INIT_29 => X"00d000db00d8008a0058006d00b800e400da00c900bf00b500a60093004d000e",
            INIT_2A => X"000d0018008b00b300a2008d0045003d00230004000b001b0036005600c200d4",
            INIT_2B => X"00cc00db0088002400200022004000b100dd00cc00ad009f00900049000f000d",
            INIT_2C => X"00090027005b00310060008f004c003e00150007001500510079008300c500d0",
            INIT_2D => X"00d100c1003800260037002e0019005900b200a90095008d0048000e00080014",
            INIT_2E => X"00050022003b003000530095005c002d000f0013002a0064006f008c00db00db",
            INIT_2F => X"00de00a0002600330025002300240027008200a4009b006e001d000c0016001e",
            INIT_30 => X"00070017003a004d005400940065002a0016002b004a0065006400a800dd00d3",
            INIT_31 => X"00d40089002b0040003f003400230015005600a2009a004e001300120018001c",
            INIT_32 => X"000900150037004c0052008c0065002500210043006c007f007e00b000c300c2",
            INIT_33 => X"00c900870030004600560041002e001500320083007b0031000b000a000b0014",
            INIT_34 => X"000b001700310049005700840078004b005d008600b100c800c800cf00d400d5",
            INIT_35 => X"00d60094003500480071006e0040002200180055004c001600070009000d0016",
            INIT_36 => X"000f00160025004e00570073006000480052005d006900720077007d007e007b",
            INIT_37 => X"007c00660030004c004b004e0029001b00090018001000060008000a000f0019",
            INIT_38 => X"0015001f0023002b003200300019000c000e000e0011001100140018001a0019",
            INIT_39 => X"00180014000d004a004e003b00410012000300050004000300050009000d001a",
            INIT_3A => X"00210028002c0025001e0017001e0025001c0019001c001c001b001800170013",
            INIT_3B => X"000f00090006001c00470053002f000800020005000500040006000b0015001c",
            INIT_3C => X"002500290030003b0049004f005c00590038002f0038003b00390030002b0028",
            INIT_3D => X"0023001b00150015002100250010000800080009000a000a000d0012001d001c",
            INIT_3E => X"002c00310046006500800080007600630047004e00540055005700530051004f",
            INIT_3F => X"0047003c00310031003a00380020001300130018001800150019001f0022001c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY20;


    MEM_IFMAP_LAYER0_ENTITY21 : if BRAM_NAME = "ifmap_layer0_entity21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"005300520051004d00510055005b005c005c005f0065005c005700520050004c",
            INIT_01 => X"00440041003f003e003c00380034002f002a0025002300220024001d00190015",
            INIT_02 => X"005400530053004d00500054005a005d005a0058005f006100580052004e004c",
            INIT_03 => X"0047004400400042003d00360034002e002a0026002400230024001e001d001f",
            INIT_04 => X"005200510050004b004b00540058004c005200560057006300650058004d004c",
            INIT_05 => X"0049004400400040003a00370034002d002b00280029002c0031003000310035",
            INIT_06 => X"005300510050004e004a005700500032005500610057005b0068006600580050",
            INIT_07 => X"00490040003f003f003b00380039003a003d003f004400470049004700450045",
            INIT_08 => X"004f004f004f004f004a0053004c003700530054004b004b004e0059005a0057",
            INIT_09 => X"0053004200430046004e005000540057005700560059005900580054004f0049",
            INIT_0A => X"004c004a004b004d00490049004600460046004500470049004b004e004e0051",
            INIT_0B => X"005a00590060006200640068006600680063005f0061005e0057005000490042",
            INIT_0C => X"004a004800470049004a003e002b00330044004000440047004b004a0051005e",
            INIT_0D => X"00600062006e0072006600640068006d0063005b00550050004c004900460043",
            INIT_0E => X"00470048004700480047003a002a002900390036003a003f0041004700520060",
            INIT_0F => X"0069005e005d00670067006a006c0061005d005b0054005000500050004f004d",
            INIT_10 => X"00490049004b0052005800670057002e003800380045005200510057005a0057",
            INIT_11 => X"00620063005e005b00610066006a0066005e00630061005c00590059005b005f",
            INIT_12 => X"0056005f006d007b0088009900680033003c003b004900610065006c0066005a",
            INIT_13 => X"005f00610061005d005d00630069006e00670069006c006c006d006e006e006e",
            INIT_14 => X"007f008b0096009d00a000a200570032004300380035005800650070006b005a",
            INIT_15 => X"005e0060005e00600060005f0060006500680071007d007e007b007700740070",
            INIT_16 => X"0098009d009f00a200a0009f005a002c00480045003a00560067005a0061005c",
            INIT_17 => X"005a0060005f005e006300620057005c0061007000830083007f00790074006c",
            INIT_18 => X"009b009e00a0009d009800940072003000440058005e0067007300600058005d",
            INIT_19 => X"005900650062005e00630065005400550069006e007d0084007f0076006b005f",
            INIT_1A => X"00940094009500920090008e00880050002f0048005e006800720071005c005e",
            INIT_1B => X"005d00670061005d0060006100550052006b006b006f0079007000640057004d",
            INIT_1C => X"00860087008a008c008e009300970089005d00490032003e0059005e005a0062",
            INIT_1D => X"0066006900670061005e005e00560053005f0065005c0066005f0052004a004b",
            INIT_1E => X"00830086008b00900098009f009a0098009e00760035003900670064005f0066",
            INIT_1F => X"006e0074006f006a0061005b00570055005400620055005300530055005a005f",
            INIT_20 => X"00870090009800a000a400a100890073009d00910080006e007b007a00680067",
            INIT_21 => X"0069006d006c00680061005a00580057004f005c00570055006500690069005e",
            INIT_22 => X"0094009a009f00a400aa00b300b0007f00b000c5009d00980071009100800067",
            INIT_23 => X"00670065006800660061005f005b0059004f0056005b005b006d006800560046",
            INIT_24 => X"009b00a400b200c500dd00ee00f800c4009c00c800b000b8006c008e0089006a",
            INIT_25 => X"006400630064006500650063005f005900500051005c00530058005200490047",
            INIT_26 => X"00bf00d600eb00f900fd00f600fb00f400a0009e00ac00c300710072008b006e",
            INIT_27 => X"0062006200610063006700680066005c0053004e00550049004b0050004a0048",
            INIT_28 => X"00f500fc00fd00fe00f300bb00ba00c9009100800097009c0074006a00800072",
            INIT_29 => X"0068006700650067006c006e0069005c0052004c00540055004e0053004d0049",
            INIT_2A => X"00fb00fc00fc010000e9007e006b0072006900730078006e0063006300680067",
            INIT_2B => X"006d006e006b006b0070006e00600056004e004c005a0068005b00520052004f",
            INIT_2C => X"00f800f800f600eb00c8007c00720076005d00570053004f00500056004b0044",
            INIT_2D => X"005f0064006200610062006100610061005b0057005b006f006e005500520052",
            INIT_2E => X"00eb00d600b50096008a0088008500840064003d0039003c004300590060003a",
            INIT_2F => X"0033004500470050005e006500680065005d0057005e006d0077006200510051",
            INIT_30 => X"00990082007a0078007c007a006f0067006a005a0039003400450066006a0053",
            INIT_31 => X"00400047004d0055006400670066006d006a0057005d006300710073005c0050",
            INIT_32 => X"006d006f0072006d006500610066006d0075007800670055005d0065005f0059",
            INIT_33 => X"004a004b0052005a0072007700690066006f006b005e006200650075006b004f",
            INIT_34 => X"00690062005d005b0063006a006f0071007000680061005f0050004c0054005c",
            INIT_35 => X"00510048004f00590075007b0069005e006000670067006500600069006f005a",
            INIT_36 => X"00570057005e0065006c006e006b0064005b005100560068005d0049004c005c",
            INIT_37 => X"0058004d004f004f005b0064005d00560057005c006100600060006000660065",
            INIT_38 => X"005a0060006700690065005f00560050005100550060006a006200550060005d",
            INIT_39 => X"00580051004f004c0047004c0054005b005c00560053005a00620060005b0060",
            INIT_3A => X"00640063005f00560050004f004f004f005200530062006c0063006000610059",
            INIT_3B => X"005c0054004f0051004c004a00520059005a005500520056005d005c00530053",
            INIT_3C => X"0057004e00490047004d0057005900530051004f0061006a006400670059005c",
            INIT_3D => X"00600057005800590052004f005400530056005a0056005300560056004f0049",
            INIT_3E => X"003e003f004600490054005600530051004e004a005e006b005f0068005b0058",
            INIT_3F => X"005b00580058005900550050005500530054005900560050004c004d004c0048",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY21;


    MEM_IFMAP_LAYER0_ENTITY22 : if BRAM_NAME = "ifmap_layer0_entity22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"005e005e005d0059005a005a0060006000610066006e0065005e005800550052",
            INIT_01 => X"004e004b0049004800450041003d00380033002e0029002700280022001d0019",
            INIT_02 => X"0060005f005f005900590059005f006200610060006a006b0060005900550052",
            INIT_03 => X"004f004b004700490044003d003b00350031002c0027002500260020001f001f",
            INIT_04 => X"005e005c005c00570054005a005d0051005900600063006e0070006200560054",
            INIT_05 => X"004f004900440046003f003a00360030002e002b0029002b002f002e00300031",
            INIT_06 => X"005f005d005c005a0053005d00560039005d006b00630068007400720065005a",
            INIT_07 => X"004e004300420042003e003800380039003c003e0041004200430041003f003d",
            INIT_08 => X"005c005b005b005b005300590052003e005c005f00580058005c006800690064",
            INIT_09 => X"005b0046004500480050004d005000530053005100510050004f004b0046003f",
            INIT_0A => X"00580056005700590052004f004c004d0050005200550057005a005e005e005f",
            INIT_0B => X"0063005e006200630064006400600062005d005800580053004c0045003e0037",
            INIT_0C => X"00550054005200540051003d002a00370053005700580059005b0057005d0065",
            INIT_0D => X"00620064007000730069006700670067005b0050004e004a0044003f00390036",
            INIT_0E => X"0052005300520054004c00370026002c004c00550052005100500053005b0063",
            INIT_0F => X"006700600061006c006d00720071005e0052004d004d004b004700440040003b",
            INIT_10 => X"005100520054005b005e00680055003100490054005b0063006100640065005e",
            INIT_11 => X"0065006800650062006a006f00720067005700550052004e004a004600470048",
            INIT_12 => X"005c006500730080008e009d00680036004b0054005d00710075007c00750065",
            INIT_13 => X"0067006a006b00670068006e007400760064005a005500540055005500550052",
            INIT_14 => X"0082008e009900a000a600aa005900350050004d0046006800770082007f006b",
            INIT_15 => X"006a006c0069006a006a0069006e00720069006200620060005e005b00590055",
            INIT_16 => X"009a009f00a200a400a700a9005d002e00510056004a0067007b0070007a0072",
            INIT_17 => X"006a006d006a0067006b00690067006e00660061006500630060005e005a0055",
            INIT_18 => X"009d009f00a1009e009e009f0075003000490065006c00780087007800740075",
            INIT_19 => X"006b0073006c00660069006a0064006900700060006000650062005d0055004c",
            INIT_1A => X"0099009800970093009300930087004c002c0049006700750083008500730071",
            INIT_1B => X"006c00770071006b006a006a0065006400750069005d0062005d0055004a0040",
            INIT_1C => X"008f008e008e008e008f00940095008300540041003500460063006b0068006d",
            INIT_1D => X"0072007c007d0075006e006c00650062006c006f0058005a005500480041003f",
            INIT_1E => X"008c008d008e0091009900a0009900930097006f0034003a006a00680065006e",
            INIT_1F => X"007b0089008700800073006c006800650063006f0059004e004a0048004a004d",
            INIT_20 => X"008f0095009b009f00a400a000880072009b008f007a0068007600770066006c",
            INIT_21 => X"00780084008500800075006d006b006a0061006c00620056005a0054004f0044",
            INIT_22 => X"009a009d009f00a100a700b100b0008100b300c70097008e00680089007b006c",
            INIT_23 => X"0079007e00830080007700730070006e00630069006a005e005c004a00340027",
            INIT_24 => X"009d00a400b000c100da00ec00f700c700a300ce00ad00b10065008800860071",
            INIT_25 => X"0077007e00820081007d007a0076007100680067006a0050003e002c00250027",
            INIT_26 => X"00c000d400e800f600fa00f200fa00f700a900aa00ae00c1006e0070008b0078",
            INIT_27 => X"0076007e008000800080007f007e0074006c00660060003e002a00250027002b",
            INIT_28 => X"00f500fb00fa00fb00f100ba00be00d200a10092009c00a0007d00730087007a",
            INIT_29 => X"0078007f00810080007f007f007d0074006a006200570042002d002a00290029",
            INIT_2A => X"00fb00fb00fb00fe00ea008300740082007f008a0082007c007a00770072006b",
            INIT_2B => X"007600800082007f007d0077006f006c0063005a00520050003d002f002c0029",
            INIT_2C => X"00fc00fc00f900ef00cb0080007b0083006f006c00660067006a006900510044",
            INIT_2D => X"0066007500780074006e006b0070007300680059004b005400510034002d002d",
            INIT_2E => X"00f500df00bf00a0009000890089008a006d004b00510057005a00660063003a",
            INIT_2F => X"003a0056005f0065006d0074007a00740061004d0046005000590042002f002f",
            INIT_30 => X"00a5008d008600840082007b00700069006b005e004a00470053006e006f0056",
            INIT_31 => X"0048005a0066006c0076007b007b007c006c00490042004400520054003d0030",
            INIT_32 => X"00750078007a0075006a00610065006a00700073006a0057005c006800680061",
            INIT_33 => X"0054005f006c00720086008e0082007a007700640045004000450057004f0032",
            INIT_34 => X"006c00660060005e0065006b006e006b0067005d0056005100420048005d0068",
            INIT_35 => X"005e005f006b0071008900940085007a0072006b005100420040004b0055003f",
            INIT_36 => X"00580057005d0063006b006c006500570049003c00410053004a003f004e005e",
            INIT_37 => X"00590057005f005d0069007b007a0072006d0068004e003b003c003f004a004b",
            INIT_38 => X"005d005f0061005f005b00540045003800320031004200550053004900550048",
            INIT_39 => X"003e003e0043004400450058006400680065005a0040003300350036003a0045",
            INIT_3A => X"0060005b00510044003b003700340030002f002e004000520052004f004d0039",
            INIT_3B => X"003500320034003a003a003f0047004a004800410034002e0030003100300036",
            INIT_3C => X"0049003c0031002b002c0030003400300030002c003a0049004b004f003e0035",
            INIT_3D => X"0032002e003400390034002f0033002f002f0031002e002a002b002d002b002a",
            INIT_3E => X"0029002500270025002a00290029002d002f002b003600470043004c003b002e",
            INIT_3F => X"002b002a002d0030002f002d0031002d002b002d002a00270025002800280026",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY22;


    MEM_IFMAP_LAYER0_ENTITY23 : if BRAM_NAME = "ifmap_layer0_entity23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"005500540053004f00500052005d005f005a0055004f0048004b004e0054004f",
            INIT_01 => X"0044003e003c003d003c003b00380033002e0029002500230024001e00190015",
            INIT_02 => X"005600550055004f004e0050005a005d00540049004600470044004500470048",
            INIT_03 => X"00460043003e003e003800350034002e00290025002200200021001b001a001b",
            INIT_04 => X"005400530052004e004900500056004800460041003800430048003f0036003c",
            INIT_05 => X"00420041003d003a0030002f002d00260024002100220025002a0029002a002c",
            INIT_06 => X"005500530052005000480052004d002b00430045003200340041003f0032002f",
            INIT_07 => X"0032003400390036002d002b002b002c002f00320038003b003c003b00380037",
            INIT_08 => X"00520051005100510048004c0046002c003d00330022001d001f002700260023",
            INIT_09 => X"0029002b0039003b003d003d00410044004400420047004800470043003e0038",
            INIT_0A => X"004d004c004c004f00470042003e0038002c0021001a001700160014000f000e",
            INIT_0B => X"001f0035004f005400530052004e0050004c0048004d004b0044003c0035002e",
            INIT_0C => X"0049004700460048004700370020002000260018001400130012000b000e0015",
            INIT_0D => X"001800290046005900560050004f0052004b004800480043003b0034002d002a",
            INIT_0E => X"004400450044004500430033001c00110017000c000a000b0009000b00110018",
            INIT_0F => X"001c00160021003f004d004f004d00400041004900480042003c0036002f002b",
            INIT_10 => X"004400450047004e0052005d004600130012000c001900250020002100210014",
            INIT_11 => X"001600180019002100310038003c003b003b004b0049003f0039003400340035",
            INIT_12 => X"00500059006700750080008d005500160015000f002100380039003d0035001c",
            INIT_13 => X"001500160016001400180023002d003a003d00480046004100410040003f003d",
            INIT_14 => X"00770083008e00950098009800470018001e001100150031003c0044003f0021",
            INIT_15 => X"0019001b00150011000f0014001c002b00370046004d004a0049004700440041",
            INIT_16 => X"008f00940096009900990099004f0017002800220019002e003d003000370027",
            INIT_17 => X"001d0024001f0015001300150012001f002a003b004c004d004d004c004a0045",
            INIT_18 => X"009200950097009400920092006b0020002b00370034003b00470034002c0029",
            INIT_19 => X"00220032002c001e001a001c00120019002e0032004500510051004f00490042",
            INIT_1A => X"0090008f008f008b008a0089007e0040001a002e003d00410046004000280024",
            INIT_1B => X"00240036003300280021001d00120013002f0033003c004e004f004a00400037",
            INIT_1C => X"0085008400860086008600880089007700470031001b0021002e002a00200022",
            INIT_1D => X"00280039003d00320027001c0011001100240033003000410046003e00360032",
            INIT_1E => X"007d007f00810085008c0091008800810084005a001e001e0040003300270027",
            INIT_1F => X"003100450045003d002c001c00140013001900300029002d00350039003c003d",
            INIT_20 => X"007d0084008b0091009500910075005a00800072006200500057004d00310028",
            INIT_21 => X"002e003f0044003c002d001f001900170015002a002b002d00400042003e0032",
            INIT_22 => X"0088008c00900093009a00a4009e0068009500a6007a007700500067004b0029",
            INIT_23 => X"002d00380041003c00300028001f001b00150023002f00320041003900230014",
            INIT_24 => X"0090009700a400b600d200e600eb00b2008500ab008a0095004d00670055002d",
            INIT_25 => X"002b0038003f003c003500300027001d0017001d002f00270027001f00160015",
            INIT_26 => X"00b700cd00e100f000f800f200f200e6008d00840084009f0053004d00560031",
            INIT_27 => X"002a0037003c003a00390037002f00210019001a0027001c0019001d001c001b",
            INIT_28 => X"00f100f800f700f900ec00b000ab00b50078006200720076004d003c00470034",
            INIT_29 => X"002e00360039003a003b0039003000200018001700250025001c0020001f001a",
            INIT_2A => X"00f800f900f900fd00e0006a005300550047004e005100410030002e00340031",
            INIT_2B => X"0033003700360039003d00330024001b00150016002700360028001f001f001c",
            INIT_2C => X"00f700f800f500eb00c2006d0060005e0041003500230019001c002b002d0020",
            INIT_2D => X"002e0033002f002f0030002d002b00290022001e0024003a00390021001d001e",
            INIT_2E => X"00ec00d700b6009800880081007a007400510023000d00090014003400490022",
            INIT_2F => X"0011001c001a0020002f003b003b00310023001a00220034003f002c001c001d",
            INIT_30 => X"009a0082007a0078007b00760068005c005a0046001f0012001d003d00450034",
            INIT_31 => X"0022002400240028003a00470041003d00300017001f00280038003c0027001c",
            INIT_32 => X"0069006b006d0068005f0058005b005d006000620056003e00380038002f0031",
            INIT_33 => X"00280025002a0030004c005b004800390036002c001d0023002a003d0037001d",
            INIT_34 => X"005f00590053005100560058005b0058005300490044003e00280023002c0034",
            INIT_35 => X"0028001e002700310051005f004700320029002a0025002300220030003a0028",
            INIT_36 => X"004b0049004f005500570053004c004000330027002a003b0032002200290031",
            INIT_37 => X"0026001e0024002700370045003c002d002600260022001d0020002400300033",
            INIT_38 => X"004c004e004f004d00440039002c0021001d001e002e003d0037002900320026",
            INIT_39 => X"001d001a001d001e001d0025002e0030002e002500190018001e00200024002f",
            INIT_3A => X"0050004a0040003200260020001e001b001b001b002d003c0035002f002c001d",
            INIT_3B => X"001c00170017001c00190018002000250023001d00150015001a001e001c0022",
            INIT_3C => X"003a002d0021001a001a001d0021001c001b001800270033003100320021001c",
            INIT_3D => X"001b00150019001d00180015001900170017001a001600120015001a00190017",
            INIT_3E => X"001b001700180015001a001900180019001a001600210030002a003300230018",
            INIT_3F => X"001500140015001800170017001d00190018001b001600120011001600180016",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY23;


    MEM_IFMAP_LAYER0_ENTITY24 : if BRAM_NAME = "ifmap_layer0_entity24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"001700130015004100a400bc00b700b200aa00ac00ba00ba00b800b700b600b7",
            INIT_01 => X"00b400a4007f005c006b006e009900c200c300c900c500c600c900c800c700c5",
            INIT_02 => X"001700130015002e009900ca00bf00b200a4009e00a900b700ba00b800b400b2",
            INIT_03 => X"00b400ad008a0056004a006a00b400ce00cf00d500d000ce00cf00cd00cc00ca",
            INIT_04 => X"001700140017001f007f00c800b900a8009f009e009a00a200b200b200b300b2",
            INIT_05 => X"00b500be00b6007d0047007200c500d100d500d800d500d300d400d300d000ce",
            INIT_06 => X"0017001500180017006300bd00af00a000a800a800a6009500aa00ba00bf00c3",
            INIT_07 => X"00c300c800bc008d0063009200d200d600d500d400d400d500d900d900d700d6",
            INIT_08 => X"0019001700170015004800aa00a5009700af00b700b9009b0092009d00a900bc",
            INIT_09 => X"00c500c400b2008d007900ac00d300db00dd00d900d900d900d600d400d100ce",
            INIT_0A => X"001a001b001a00170031008f00a4009a00a900c200c800a60082007d00800097",
            INIT_0B => X"00a500a50094008f009300b600bc00c900d400d900d500db00dc00d700d700d3",
            INIT_0C => X"001e001a001b00190025007d00b400ab00a900c500ca00b3008b0071007a0082",
            INIT_0D => X"00770085007a008c00b900cb00bf00c900d700da00d700db00dc00da00dc00e0",
            INIT_0E => X"005e0030001f0024006400af00c100a800a300c000c600c300ae0091008e0084",
            INIT_0F => X"006a0079007a008b00c000d100bd00d500f200ed00ef00e800d000d500de00e5",
            INIT_10 => X"00b4009e0072007a00b100be00be00a0008500ad00c500c800c200b900a70092",
            INIT_11 => X"008100810085008d00b100c900bd00dc00f100eb00e800d500bd00c700e100ea",
            INIT_12 => X"00c500c000b200ba00c100c300c5009d008000a300b900bf00c100c300b20097",
            INIT_13 => X"007200810083008600aa00c200d000ea00ec00f000eb00c900b900bb00d000eb",
            INIT_14 => X"00ca00c400bb00c000c800cd00c50097009500af00b800bd00c100bb00a80088",
            INIT_15 => X"007500800080008100a700b500cd00f000f300f300ee00ce00ba00bb00c100dd",
            INIT_16 => X"00cd00cd00c500c000cb00d000c200a000a800bf00c100bf00c100ac00920077",
            INIT_17 => X"007c008e0085008700a700b000bf00ea00f300f100ec00d700ba00b800b900c4",
            INIT_18 => X"00ce00cc00c800c100c500c700bf00b400ac00b300b700ad00ae00ae00980083",
            INIT_19 => X"008d00a6008e009a00a900ac00bf00e600f000f100ef00e400c800ba00b800c0",
            INIT_1A => X"00d200ca00c600bf00c900b400b100ca00ab009a008e008e00a800a80093009c",
            INIT_1B => X"00af00a9009600a4009e00a000c500e600f100f100f400f200e200bf00c300d7",
            INIT_1C => X"00d300c900c700c000cf00aa00a100d700bd00ba00ad00ac00be00b10089007f",
            INIT_1D => X"00b400ae009600a000af00b000c100ec00f500f200f300fb00ef00c900d400e1",
            INIT_1E => X"00d300c400c500c100d100b5009a00d900ce00c500c300b900aa00ad00a60098",
            INIT_1F => X"00a300b800a6009800c000b500af00cc00ee00f300f400f700df00d500e200e2",
            INIT_20 => X"00d600c200b400b500c500c4009b00c600d600c000ae00b700ad00a100ae00b2",
            INIT_21 => X"008000a400bd009300a700b4009c0076009d00d700ef00eb00ce00d600ea00e4",
            INIT_22 => X"00d700c600a600a300b400ca00be00b900cf00d200cd00d600c100ae00b000ad",
            INIT_23 => X"0081008900bf009900a300c800ab00870074009000b800c100bb00d200ef00eb",
            INIT_24 => X"00d800cd00ae00a400b900cb00d200c200bf00d300da00e200e100cb00be00b3",
            INIT_25 => X"0097007900a8009e00a700c200aa00ac009a0083009900a900a200b800de00ec",
            INIT_26 => X"00d800d000c000b400c500ca00d100d200ba00bd00c500cc00d100d500cf00b5",
            INIT_27 => X"00b20095009200af00b700ae009c00ab00a3009400a900b400a600a000ac00cc",
            INIT_28 => X"00da00d500ca00b600bf00cb00c900ca00ca00c300c100c000b200c600cf00c7",
            INIT_29 => X"00d300cb00a600bb00b1009b009300a600a700ab00b600af009c009c009f00a7",
            INIT_2A => X"00d900d700d100ba00b300c800d000c800d100d700d200ba00a100b600c400c2",
            INIT_2B => X"00cb00cf00be00b9009b008e009b00a600ac00b300ad009f0096009e009e008f",
            INIT_2C => X"00d600d500d600c000a900c500da00d900d700d900d400c300aa00b300c300bf",
            INIT_2D => X"00be00c000c000aa0084008e00a700aa00aa00b300ad009d009d00930086007d",
            INIT_2E => X"00d500d100d300ca00a800c100d800de00df00de00d300cd00c200c200c900c6",
            INIT_2F => X"00c600c400bc00990086009b00ab00a700a600bd00b200a500a3008e00850089",
            INIT_30 => X"00d300ce00ce00ca00af00bf00d300d500d600d800c600ab00c200ce00c900c9",
            INIT_31 => X"00c800c500b100960090009e00a7009d009f00b500b000a80098009600950090",
            INIT_32 => X"00d200cc00c900c100b500bc00d000d200cd00ce00a0007a00b100d000c600c2",
            INIT_33 => X"00c100b800a60096008b009c00a00099009b00a0009f009b00980098008c0083",
            INIT_34 => X"00d200ca00c600bb00ae00b200cd00d600d100cb00a4008300b400ca00bb00b6",
            INIT_35 => X"00b600a9009d008b00860099009a00900097008d0083008d009d009b00960093",
            INIT_36 => X"00d200c800c200b500a800a800c400d700d400c700bd00b800cb00b900ad00ac",
            INIT_37 => X"00a3009b00930076008300940091008d00900084007f0085009500a300a2009c",
            INIT_38 => X"00d000c200bd00b400a2009e00bd00d300d300c500c200c700bf00ac00a300a4",
            INIT_39 => X"009e00930082006d008900900090009100900084007c0086009700a2009f0093",
            INIT_3A => X"00c200b100b000b5009f008f00b300cd00d000c700c200be00b500a5009c00a1",
            INIT_3B => X"009500880070007200890085008a00920092008300830090009600950094008d",
            INIT_3C => X"00ac009d00a500b200a70085009c00c700ce00c700c700c200a000850084008b",
            INIT_3D => X"008c007e006b007e00820081008a0095008d008c0091008e0088008c00950098",
            INIT_3E => X"009700860090009b009e007d008200b700c500bf00b700a500800067005e0069",
            INIT_3F => X"007700700075007c0079007d008b008f008b008c0081007d00840095009b0096",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY24;


    MEM_IFMAP_LAYER0_ENTITY25 : if BRAM_NAME = "ifmap_layer0_entity25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"001300150010002f008300930093008e008700890090008e008d008c008c008f",
            INIT_01 => X"008c007e00600049005f005d008200a4009b009c009b009d009e009b00980097",
            INIT_02 => X"001400140011001f007a00a1009b0092008a0088008b00950098009600920097",
            INIT_03 => X"009f00960075004900410058009c00af00a800a900ab00ad00ac00a800a400a3",
            INIT_04 => X"0014001400140015006600a20097008c008d00950088008b009a00990098009f",
            INIT_05 => X"00a600ab00a1006d003a006100b100b700b300b200b100b200b100ad00a900a6",
            INIT_06 => X"0014001400150011004f0099008c0082009700a4009d0087009900a600a900b0",
            INIT_07 => X"00b000af00a100760052008500c400c300bd00b700b400b300b300b100ad00ab",
            INIT_08 => X"00150014001500130038008900820077009c00b200b300920084008b009400a7",
            INIT_09 => X"00af00a900980078006d00a700ce00d200d100c900c300bf00ba00b600b100ac",
            INIT_0A => X"00160016001700160026007300820078009200b900c3009e0076006c006b0084",
            INIT_0B => X"0092008f00810084008f00b700be00c700cf00d100cc00d100d100ca00c700c2",
            INIT_0C => X"0018001300150014001e007100a10094009700ba00c200aa0080006200690071",
            INIT_0D => X"00680074006b008000b200ca00c000c500ce00cf00d100d700d800d600d700da",
            INIT_0E => X"005800290018001d006000ae00ba009c009500b500bd00ba00a4008400810076",
            INIT_0F => X"005c006b006c007c00b400cc00bb00ce00e600e000e700e400cd00d300dc00e2",
            INIT_10 => X"00b10099006d007500af00bd00b70093007800a100bc00c000b800ad009a0083",
            INIT_11 => X"007300730077007f00a600c500bc00d800e900e200e300d300bc00c600e000e8",
            INIT_12 => X"00c200bc00af00b600bf00c200be00900073009800b100b600b700b600a4008a",
            INIT_13 => X"006600760077007b00a000bd00d000e900e800eb00ea00cb00bb00bd00d100eb",
            INIT_14 => X"00c700c000b700bb00c600cd00bf008a008800a500b000b500b800af009a007c",
            INIT_15 => X"006b007600770078009e00b000cd00f000f300f400f200d400c000c000c600e0",
            INIT_16 => X"00c900c900c100bb00c900d100bc0092009b00b600b900b700b7009f0084006b",
            INIT_17 => X"00730085007c007e009e00aa00bd00eb00f600f600f200de00c200c000c000ca",
            INIT_18 => X"00cb00c900c500bd00c400c600b700a5009f00aa00b000a500a400a2008a0078",
            INIT_19 => X"0085009f0087009200a100a500bd00e700f400f800f700ea00d000c300c100c7",
            INIT_1A => X"00d000ca00c400b900c100a7009c00b900a100910087008700a1009e0089008f",
            INIT_1B => X"00a400a4009500a20099009d00c300e400f200f700f900f500e800c700cc00de",
            INIT_1C => X"00d200cc00c500b600bf008e007d00c100b500b100a600a700b800aa00820072",
            INIT_1D => X"00a500aa0098009e00ab00ae00bd00e700f200f400f500fb00f200cf00dd00e9",
            INIT_1E => X"00d400c800c500b900bd0091007000c000c700be00bd00b400a400a700a00089",
            INIT_1F => X"009200b000a2009100b800b100a800c300e800f100f500f900e400dd00ec00eb",
            INIT_20 => X"00d800c700b600ae00b0009b006e00ad00d000ba00a800b200a8009b00a700a4",
            INIT_21 => X"006e009600b10086009a00ab00900068009100d100ee00ed00d200dd00f300ed",
            INIT_22 => X"00db00ce00a9009e00a300a7009500a200ca00cd00c800d100bc00a800aa00a1",
            INIT_23 => X"0070007800ad0087009300ba009b00730062008400b200bc00b900d400f300ef",
            INIT_24 => X"00dd00d600b300a100af00b500b300b100bd00cf00d400dd00dc00c500b800ab",
            INIT_25 => X"008b00670095008c009700b10094009300830070008a009c009700b100d900ea",
            INIT_26 => X"00df00da00c600b200c200c200be00c800ba00b800bf00c700cb00d000c800b1",
            INIT_27 => X"00ab0087007f009e00a8009b0083008f0089007e0094009f00930090009e00c5",
            INIT_28 => X"00e100dd00d000b700bf00c700be00c200c600bc00be00ba00ab00c100c600bf",
            INIT_29 => X"00cf00bf009400a900a00087007b008d008e0095009f009800870088008c009a",
            INIT_2A => X"00de00dd00d600be00b300c300c800be00c600cd00d100b2009700b300b600b5",
            INIT_2B => X"00c500c400ae00a50086007c00890093009900a10099008b0083008b008b007d",
            INIT_2C => X"00db00da00db00c600aa00bf00d200cf00cb00ce00cf00b4009c00ae00b400b0",
            INIT_2D => X"00b600b500b00096006f007d00960098009800a1009a008a008a00800073006a",
            INIT_2E => X"00da00d600d900cf00aa00bc00d200d500d400d300c700b600ae00ba00ba00b5",
            INIT_2F => X"00ba00b600ab008500720089009a0095009400ab009f00920090007b00730076",
            INIT_30 => X"00d800d400d400d100b300bd00cf00cd00cd00cd00b1008a00a700c300bb00b6",
            INIT_31 => X"00b900b5009e0082007d008d0096008c008d00a3009d0095008500830082007c",
            INIT_32 => X"00d700d200d000c800bb00be00ce00cc00c600c400830050009100c200b800ae",
            INIT_33 => X"00ae00a5009300830078008b008f00880089008e008c00880085008500790070",
            INIT_34 => X"00d700d000cd00c200b500b700cd00d100cc00c200810051008e00ba00ab00a1",
            INIT_35 => X"00a1009500890078007300870089007e0085007b0070007a008a008800830080",
            INIT_36 => X"00d600cd00c800bc00b000af00c600d400d000c000a0008e00aa00a8009b0095",
            INIT_37 => X"008d0085007f0064007100830080007b007e0072006c00720082009000900089",
            INIT_38 => X"00d200c400c000b700a900a600c000d200d100c000b600b400ab0099008d008c",
            INIT_39 => X"0086007d006f005c0078007e007e007f007e00720069007400850090008d0081",
            INIT_3A => X"00c400b300b300b900a6009700b500cc00cd00c200ba00b300a6009200850088",
            INIT_3B => X"007e0072005d00610078007300780080008000710071007e008400830082007b",
            INIT_3C => X"00b100a100aa00b800ae008c009c00c300c900c100bf00b600910071006c0073",
            INIT_3D => X"0076006a0059006e0072007000780083007b007a007f007c0075007a00820086",
            INIT_3E => X"009d008c009700a100a60082008000b100bf00b700af009a0070005300470053",
            INIT_3F => X"0063005e0065006e006c006c0079007e0079007a006f006b0073008400890084",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY25;


    MEM_IFMAP_LAYER0_ENTITY26 : if BRAM_NAME = "ifmap_layer0_entity26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0017001c0013002800710073006d007400710067006a0069006900690069006b",
            INIT_01 => X"006a0063004c003a0054005600720089007c007d007c007d007f007d007a0078",
            INIT_02 => X"0018001b0014001a006a00820076007c007d0072006d00750078007600720079",
            INIT_03 => X"00850083006a0044003e0051008c0096008a008c008900880088008500810080",
            INIT_04 => X"0018001a00170012005800830074007b008b008d007400740081007f007d0084",
            INIT_05 => X"008e009a0098006900370059009f009e009700970092008e008e008b00880084",
            INIT_06 => X"00180019001900120045007c006a0073009c00a6009200780089009400950097",
            INIT_07 => X"0096009c0094006d004a007a00b100a900a1009d00980095009600940091008e",
            INIT_08 => X"00190018001900170033006d0060006800a100b800b2008d007c008000860093",
            INIT_09 => X"009700960089006c0060009800b700b500b300ae00a800a400a0009c00980093",
            INIT_0A => X"001a001a001b001c00230059005f0066009600c100c7009f0074006600620076",
            INIT_0B => X"008200830077007a008400a700a600aa00b200b700b300b700b700b100af00a9",
            INIT_0C => X"001a00160019001a001d005c0080007b009300c300c700ab007e005e0063006a",
            INIT_0D => X"0060006d0065007a00ac00c000aa00b000c300c400c500ca00c500bf00bf00c2",
            INIT_0E => X"004d0021001100190058009a009b007e008c00be00c100b900a30081007b0071",
            INIT_0F => X"005800670068007900b100c600a500bd00e400db00e000da00ba00bb00c400cd",
            INIT_10 => X"0095008000560060009b00a700990077006f00a800bf00bf00b700aa0094007f",
            INIT_11 => X"007000700074007c00a300bb00a200c100df00d500cf00bb009d00a600c400d2",
            INIT_12 => X"00a1009e0092009b00a700a9009f00750068009b00b300b500b600b4009f0087",
            INIT_13 => X"0064007400750079009e00b200b200cc00d800d600cb00a70093009600b000cf",
            INIT_14 => X"00aa00a5009e00a500af00b000a00070007b00a400b100b400b600ac00950079",
            INIT_15 => X"006a007400750076009c00a600af00d100de00d800cd00a900910093009f00ba",
            INIT_16 => X"00ac00ae00a900a600b000b0009d007a008d00b100b900b600b6009d007f0068",
            INIT_17 => X"00730084007b007d009f00a400a300ce00e000d900cd00b50092008e0093009c",
            INIT_18 => X"00a700a700a500a000a500a40099008f009100a300ae00a400a3009f00850076",
            INIT_19 => X"0086009f0087009200a300a300a800cd00df00dc00d600c700a3009000900098",
            INIT_1A => X"00a900a200a0009b00a30088008300a40092008800840085009f009e00870092",
            INIT_1B => X"00a700a20090009e0098009800b000cb00d700d800dd00da00c5009f00a200b6",
            INIT_1C => X"00ae00a400a2009d00a80078006d00b200a600a700a100a300b600ab00840078",
            INIT_1D => X"00a900a3008c009500a600a400aa00cc00d300d500da00e400d600b000bb00c7",
            INIT_1E => X"00af00a000a1009f00aa0084006800b700bc00b600b800b000a200a800a3008d",
            INIT_1F => X"009100a50092008500af00a5009600a900ca00d400d900dd00c400ba00c700c7",
            INIT_20 => X"00b3009f0092009400a10097006d00a800c700b500a400ae00a5009c00aa00a6",
            INIT_21 => X"00690088009f0077008f009e007e0050007600b700d100cd00af00b700c900c5",
            INIT_22 => X"00b500a400850083009500a50097009f00c200c700c400cd00b900a800ac00a2",
            INIT_23 => X"00680069009b0077008600ad0088005c004b006f0098009e009800b000cb00c8",
            INIT_24 => X"00b700ac008e0085009f00b000b100aa00b100c500cf00d900d900c600bb00aa",
            INIT_25 => X"0083005a0085007e008b00a20082007e006f006000760084007c009200b800c7",
            INIT_26 => X"00b900b000a1009500af00b700b600bc00aa00aa00b900c200c900d000ca00af",
            INIT_27 => X"00a4007b00710091009d008c0071007b007700700086008e007f0079008400a6",
            INIT_28 => X"00bd00b700ad009b00ab00ba00b100b200b400ac00b200b100a400bc00c300bd",
            INIT_29 => X"00c900b60088009d00930078006a007c0080008a0094008a00780077007a0082",
            INIT_2A => X"00bd00bc00b700a1009e00b700bb00b000b800bf00c000a4008b00a600ad00b1",
            INIT_2B => X"00c000bc00a200960076006b00790085008e0096008d007d0075007c007d006c",
            INIT_2C => X"00ba00ba00bb00a6009400b400c700c500c100c300c000a80091009f00a900aa",
            INIT_2D => X"00af00ac00a30086005d006c0086008b008d0097008e007c007c00720065005b",
            INIT_2E => X"00ba00b500b700ac008f00b000c900cf00ce00cb00bd00af00a500ab00ae00ac",
            INIT_2F => X"00b200ab009e007500610078008a0088008a00a1009200840082006d00640068",
            INIT_30 => X"00b800b200af00a9009200aa00c600ca00c800c500ab008800a100b400ab00aa",
            INIT_31 => X"00ad00a800900073006c007c0086007e0082009900910087007700750074006f",
            INIT_32 => X"00b800b000a8009d009300a200c000c800bf00b900810052008d00b300a6009f",
            INIT_33 => X"009f0096008400740069007a007f007a007f00840080007a00770077006b0062",
            INIT_34 => X"00b800ac00a300940086009200ba00ca00c000b200820058008c00ac00980090",
            INIT_35 => X"00910084007a00690064007700790070007a00710064006c007c007a00750072",
            INIT_36 => X"00b700a9009e008e007e008400b200cc00c300af009d009000a4009800870083",
            INIT_37 => X"007c0074006f0054006100730071006d00720066005f0064007400820082007b",
            INIT_38 => X"00b100a10099008e0077007a00b200cc00c500b400aa00a8009d0087007a007b",
            INIT_39 => X"0077006d005e004b0068006f0070007100700064005c006600770082007e0073",
            INIT_3A => X"00a30090008d00910074006b00a900c800c200b700ac00a30096008100730079",
            INIT_3B => X"00700064004e005100680065006a00720072006300630070007600750074006e",
            INIT_3C => X"008e007e0083008f007c005f009100c000be00b700b200a800820062005c0065",
            INIT_3D => X"0068005c004b005f00630061006a0074006d006c0071006e0067006c00740077",
            INIT_3E => X"007b00680070007800740057007600ae00b500ae00a4008d0063004500390046",
            INIT_3F => X"0057005100580060005d005e006b0070006b006c0061005d00650076007b0076",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY26;


    MEM_IFMAP_LAYER0_ENTITY27 : if BRAM_NAME = "ifmap_layer0_entity27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00d900d200cd00c700da00d600cf00bd00bb00ae00a600a90096009a008c008f",
            INIT_01 => X"00a700bf00db00df00db00d700e200e100db00be00af00bb00c800aa00a100a2",
            INIT_02 => X"00de00dd00dc00d700d800e100d300b300b400c000be00bc00c700ce00d100db",
            INIT_03 => X"00e500eb00ec00ec00e900e200e100e500e700d400d000cd00d800b700ba00c8",
            INIT_04 => X"00ea00e900e700e800e900ef00d900ad00a400b400ad00b700be00bc00d400e0",
            INIT_05 => X"00da00eb00e300e100e500df00d600e100ea00e800e600d800d100ca00d000d3",
            INIT_06 => X"00f500f400f400f200f400f300e4009e0092009d0083009f0091008800a2009f",
            INIT_07 => X"00a900cb00c300d300d100cb00d000e200e600e900e400d500c700db00e000d4",
            INIT_08 => X"00f500f300f400f400f500f100cf00750063006c0059006b0064005b0064005c",
            INIT_09 => X"0066007c007c009500b600b900ca00e900e100e200e300cd00c200d500e200de",
            INIT_0A => X"00f500f400f400f300f500ed00d8007e0048005a005b006600650067006b0063",
            INIT_0B => X"00590059005b005d007e00be00d800eb00e700df00d800c400ae00bd00d900ec",
            INIT_0C => X"00f500f300f300f400f100db00d9009e0050007200840097008c0084008f008a",
            INIT_0D => X"0082007a00720078006e009b00dd00e900eb00e000c600c000a700ab00cc00eb",
            INIT_0E => X"00f400f300f300f600e300c700d700990051009200bb00ca00cf009e00830083",
            INIT_0F => X"0081008d00830084009f0084009f00d700e500d700d400d100c500ab00b200dd",
            INIT_10 => X"00f400f300f400f500e300ce00da0082005100820080008100b800910074007d",
            INIT_11 => X"007c0089008e007d00990093009000c600d600db00e900dc00b800a400a900c9",
            INIT_12 => X"00f300f300f400f200e400be00a8006e005300860077006e008f008000730078",
            INIT_13 => X"007d00830092007d0095009b008c00c400e900f000f000e900c800c800d700dc",
            INIT_14 => X"00ef00f100f400f500dc00850082005f004e00740074006c006d006b006d006c",
            INIT_15 => X"007300780078007300880096008f00a700d000e400f500f300f400f500f500f4",
            INIT_16 => X"00de00e900f200f400d800a900a50059003d0043005b0064005f005f00620060",
            INIT_17 => X"0060005f005a0061006900790081007e009b00d800f800f300f400f400f400f4",
            INIT_18 => X"00d000df00ec00e300bf00b700b500640037003800580065006f006300560054",
            INIT_19 => X"00520054005d0071006d00620070008100ae00e200f500f400f400f400f400f4",
            INIT_1A => X"00c800cc00db00c300aa009a009c006600680063006c006600730075005e0055",
            INIT_1B => X"005a006a007a008c00800068006c007c009600b300c300d400ef00f500f400f4",
            INIT_1C => X"00c800d200cf00a900a400940093008a0081005c006a005d0059005d0054004d",
            INIT_1D => X"004c005100510051004f004a004b00520065007b008c008f00bf00f400f400f4",
            INIT_1E => X"00d200e200c400770070009600ba00c0006c004d004d0037002d002f003c003f",
            INIT_1F => X"003b003f003b003600310032003d00400047004b005b0067008700e100f600f4",
            INIT_20 => X"00c700c100b40060005d009100c000a100560049005c00620068004f004f0047",
            INIT_21 => X"0025001c001e001b003400320016001c00180035005b0068008000ce00f700f3",
            INIT_22 => X"00d300c700c200710078009d009f00470044005a0074007c0095007900800066",
            INIT_23 => X"004e00620070006400940093005c0063005e006c0087008e009c00b700f200f5",
            INIT_24 => X"00dc00ca00b70066006e00a50084001e00390062006b00530052006500810064",
            INIT_25 => X"009900ae009e009f00ac00a800a200a300a000af009c00770072008700e400f7",
            INIT_26 => X"00db00cf00bc00620053008d006f002a003a0048004c003e003500380040005d",
            INIT_27 => X"00a0007c005b00650074006b006700670063009b007e00430051007600d900f8",
            INIT_28 => X"00d900d200c7006500380058005d003c0038002e003f0046003c003600400041",
            INIT_29 => X"006300720069006700640060005d00610066006f006400490052007200d400f9",
            INIT_2A => X"00d100cd00ca0075005300460051004400320023002b00330044004d0057003f",
            INIT_2B => X"003400470052004800400043003e005d0058003c0053006c0070006c00cc00fa",
            INIT_2C => X"00cd00ca00c50068005d006f00470049003f002900260022004b0063008e004f",
            INIT_2D => X"001e005600930076006300720066009900b2003f004a008d0077005a00c300f6",
            INIT_2E => X"00c600c200b900570031006c00610063005f0033002700240028003200570037",
            INIT_2F => X"0020004f0097007f007a00880074009c009f00370035004a003e004e00c200f0",
            INIT_30 => X"00b600b400a9004d0025003b006c0090006a003c002b0020001d001c001e0021",
            INIT_31 => X"0027002a003a0058006a0079007a00750043002f003300320033005000ba00e1",
            INIT_32 => X"00a800a500a4007d005b0060006f008d0060004a00370024001e001e001d001f",
            INIT_33 => X"00230018004000ae00cd00cb00b300b500570026002b00300042005b00ae00d3",
            INIT_34 => X"00a200a300af00b400980076006c008d005b0053004e0030001900180019001d",
            INIT_35 => X"00270026004700a400b800b100a900a60051001e001e0031004e005f00a900ce",
            INIT_36 => X"009a00ac00b300a6009200750067009200570055005200360020001e00210025",
            INIT_37 => X"0036004d00560065006b0079008e0089003c001e00210036004e005b00a500c7",
            INIT_38 => X"00a600a9009e0094008f008500670071004f0051004b003c002a0027002a002c",
            INIT_39 => X"003000360041004d005a006e0083008b0035001d002600360046005b00a900c4",
            INIT_3A => X"00a200970093008d00890085006b004e0048004e0046003c0032002a002e0030",
            INIT_3B => X"00310033003b0042004c0059006500710045001d00230034003f006200ae00ba",
            INIT_3C => X"0094008d008e008c008f008c006a003c0042004a00420037003900340036003a",
            INIT_3D => X"003a003a00410046004900500057005d004d002500260037004a008300b300b4",
            INIT_3E => X"0090009500a000a2009e0092007e003d00390039003a00430046004500490048",
            INIT_3F => X"0044004900590062005e0061006300610052004500400047007700a400b600ba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY27;


    MEM_IFMAP_LAYER0_ENTITY28 : if BRAM_NAME = "ifmap_layer0_entity28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00d700d000d000ca00d700d100ca00b900b800a8009800a0009d00a7009a009d",
            INIT_01 => X"00b500cb00e100e100de00db00e500e400dd00c500b800c400d000b800b000a5",
            INIT_02 => X"00e200e000e100d900d500dd00cc00ab00b400bd00b200b100c400cd00d000e0",
            INIT_03 => X"00ec00f000f200f300ee00e500e400e700e700d600d400d200de00be00bf00c5",
            INIT_04 => X"00eb00ea00ea00eb00ea00ef00d600a600a600b100a800b100b800b700ce00df",
            INIT_05 => X"00dc00ec00e300e800eb00e400d900e000e900e900e600dd00d900ce00d100d2",
            INIT_06 => X"00f500f400f400f300f400f400e300990092009b0082009f0090008a00a200a0",
            INIT_07 => X"00ac00cd00c200dc00de00d300d300e000e600e900e500db00cf00df00e200d4",
            INIT_08 => X"00f500f400f400f400f500f000cd00700062006d005b006d0065005c0064005c",
            INIT_09 => X"0068007d007c009a00c200c200c900e300dc00de00e300d300cb00dc00e800e1",
            INIT_0A => X"00f500f400f400f300f600eb00d4007b0047005d005f00690067006a006e0066",
            INIT_0B => X"005b0059005b005d008100c500d900e600dd00da00d600c600b400c500e200ed",
            INIT_0C => X"00f500f300f300f400f000d600d5009c004f00770089009a0090008b009b0096",
            INIT_0D => X"008e00800079007e007200a000e100e900e900da00c000ba00a500b000d400ec",
            INIT_0E => X"00f400f300f300f700e200c100d300960051009800bc00c800cd00a5008d0090",
            INIT_0F => X"008e0096008d008f00a7008c00a300d600e000d100d300d200c700ae00af00dc",
            INIT_10 => X"00f400f300f400f500e100ca00d8007f005100860084008700b90097007c0087",
            INIT_11 => X"008600910096008800a4009e008e00c000cf00d800e700d700b1009e009c00c4",
            INIT_12 => X"00f200f200f400f200e300bd00a8006e0053008c0080007600930087007c0081",
            INIT_13 => X"0085008b00970086009e00a4009100c100e500ef00ef00e600c100be00cc00d7",
            INIT_14 => X"00e800ef00f300f400da00810080005e004f007a007a00700071007000730073",
            INIT_15 => X"007c0080007f007e0090009e009900aa00ce00e300f600f400f300f300f500f4",
            INIT_16 => X"00cd00e300f200f200d300a1009f0058003c0045005e00660062006100670066",
            INIT_17 => X"00680064005f00670071007f00890080009900d700f800f300f400f400f400f4",
            INIT_18 => X"00bc00d500e400dc00b400aa00ad006300370039005a00660072006700580055",
            INIT_19 => X"00550055005d0073007000650076008600b000e100f500f400f400f400f400f4",
            INIT_1A => X"00b800bc00ca00b500980086008d006300670066006f00670076007800600056",
            INIT_1B => X"005c006b007d00920084006a006e007f009800b300c300d200ee00f500f400f4",
            INIT_1C => X"00b600c200bd00980092007b007f007e007c005d0069005e005a005d0055004f",
            INIT_1D => X"004e0053005400550051004b004c00530065007a008a008a00bc00f400f400f4",
            INIT_1E => X"00bd00cc00a700650065007d00a900ae0067004d004f0036002b002f003b003e",
            INIT_1F => X"003b003e00390034002f0030003d00400046004a005a0061008000df00f600f4",
            INIT_20 => X"00ae00a4009700540052007c00ac0092005300490057005a0064004b004c0044",
            INIT_21 => X"00210017001a00170030002f001400190015003200560064007800ca00f700f3",
            INIT_22 => X"00c000b400b3006800680087008e004000410057006c007800950076007d0062",
            INIT_23 => X"00460059006a00600090009000590060005a00670082008b009700b200f100f4",
            INIT_24 => X"00d100bd00ab005e006200920076001c0036005f0067004f005300640080005f",
            INIT_25 => X"009200aa009b009e00ab00a800a000a1009e00ac009b0077006f008000e200f7",
            INIT_26 => X"00d000c100b0005b004c007f00640028003500440049003900320035003d0059",
            INIT_27 => X"009c007700570062007100680063006400600098007a003f004d007000d600f8",
            INIT_28 => X"00ca00c300be005f0033004e0053003800330027003c004400390033003b003d",
            INIT_29 => X"005f006e006600650063005f005c00600064006c00600046004f006c00d000f9",
            INIT_2A => X"00c200c000c0006e004c003e0049003f002e001d00280030004100480053003b",
            INIT_2B => X"00300043004d0043003c0040003b005800520036004e0069006b006500c900f9",
            INIT_2C => X"00c300be00bb00610055006300410043003a00260023002000480060008d004c",
            INIT_2D => X"0019004f008c0071005e006d0061009200ab003a0045008a0074005300c000f4",
            INIT_2E => X"00bd00b700b00052002c00630059005e005a0030002400210026002f00550034",
            INIT_2F => X"001c004a0091007b0077008600710097009c003300320047003b004700c000ee",
            INIT_30 => X"00ae00ad00a30048002200360065008b0066003a0028001e001a0019001a001e",
            INIT_31 => X"00250026003500560068007500760072003e002b0030002e002f004b00b800df",
            INIT_32 => X"00a200a0009e00780057005900670088005c004800340022001c001b001b001d",
            INIT_33 => X"00200015003d00af00cf00ca00b100b4005400220028002c003e005700ab00d1",
            INIT_34 => X"009c009c00a800b0009300700066008800560051004b002d001600160017001a",
            INIT_35 => X"00230022004500a400b900b100a900a5004e0019001a002d004b005c00a700cc",
            INIT_36 => X"009500a700ad00a1008d00710063008e00530053004f0033001d001c001f0022",
            INIT_37 => X"003200480051006100660074008a00850037001b001d0032004c005900a400c6",
            INIT_38 => X"00a400a6009b0090008b00820063006c004c0050004800380026002400270029",
            INIT_39 => X"002d0033003d004800540067007c00830031001a002100320045005900a900c3",
            INIT_3A => X"00a000940092008d00870082006600490045004d00420038002f0028002b002d",
            INIT_3B => X"002e00300036003d00460054005e006a0040001a001f0030003d006200af00ba",
            INIT_3C => X"0093008d008e008c008f008b006800390040004a003f00340037003100330036",
            INIT_3D => X"00360036003d00420044004a0051005700480021002300340048008400b600b5",
            INIT_3E => X"0092009600a100a3009d0091007c003a00370038003900410043004200460045",
            INIT_3F => X"004300480057005f005c005f0060005e00510044003e0046007600a300b600b9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY28;


    MEM_IFMAP_LAYER0_ENTITY29 : if BRAM_NAME = "ifmap_layer0_entity29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00d100ca00bf00b600d100d100c600af00ab00a5009d00a00095009a008d008f",
            INIT_01 => X"00a400bc00d600db00d100ca00d900d600d000b100a100ad00b7009d00950095",
            INIT_02 => X"00d400d400d200cd00cf00db00c800a300a500b600b800b600c200c900cd00d7",
            INIT_03 => X"00df00e300e300e400dd00d400d300d700df00cd00c300bb00c600aa00ad00ba",
            INIT_04 => X"00e600e500e300e200e300ec00d300a4009f00ad00b700b800bc00bf00cf00e0",
            INIT_05 => X"00db00e500e000d600d600d000c800d300de00e000db00c500b900bc00c500c6",
            INIT_06 => X"00f500f400f400f100f200f100e300af00a800b000a100bb00ae00a000b800b6",
            INIT_07 => X"00b900d500d000ca00b900ba00c400d400d700dc00d500bb00a900c500d400c8",
            INIT_08 => X"00f500f300f400f400f500f100cd0084008b00a1008a00a7009f008b009b008d",
            INIT_09 => X"008e00a6009900a400a900a900c400e000d100d100d400b100a000b800cc00d2",
            INIT_0A => X"00f500f400f400f300f600ee00d700810071009c00a000aa00aa00aa00b100a7",
            INIT_0B => X"009d009d0098008f009400b300cd00e400da00ce00c100aa009300a000c000df",
            INIT_0C => X"00f500f300f300f400f100dd00dd00b4008300b400c400cf00c800cb00d900d3",
            INIT_0D => X"00cc00c300c000bf00a300a600cd00e100e300d500b100a90091009200b200da",
            INIT_0E => X"00f400f200f200f700e600ca00d900c0008600c200e000e800ea00d700ce00d1",
            INIT_0F => X"00cf00d000ca00cf00e000b4009a00cc00dc00c900c400bc00ab0092009a00c7",
            INIT_10 => X"00f500f300f300f500e300d100df00ae008700ba00c100c100dd00cc00c100c9",
            INIT_11 => X"00ca00cd00cd00c600dc00d000a300bc00cb00d100df00cb00a1008b009400b2",
            INIT_12 => X"00f200f100f300f200e500cd00c200a4008c00c100bd00b800ca00c400c000c4",
            INIT_13 => X"00c700ca00d000c600d700e000bc00c800e600ee00ed00e300bc00ba00ca00d3",
            INIT_14 => X"00ea00ee00f300f400df00a000a9009c008600b100b300ac00ae00ae00b400b7",
            INIT_15 => X"00bb00be00bc00be00cd00dc00d000c400d900e600f600f400f400f400f400f4",
            INIT_16 => X"00d300e600f200f200d800b600be0097006a006e009300a0009e009f00a600aa",
            INIT_17 => X"00a900a3009e00a600ad00bd00c600af00b700e000f800f300f400f400f400f4",
            INIT_18 => X"00c400da00e900e100bd00b400c3009f005d005c008d00a000ba00a8008f008c",
            INIT_19 => X"008b0089009200a700980083008f009600bc00e300f300f400f400f400f400f4",
            INIT_1A => X"00c300c700d300c100a4009500a20089009600aa00b200a600bd00cd00a60092",
            INIT_1B => X"009900ac00c000d300af00800080008a00a000b100bf00d300ef00f500f300f3",
            INIT_1C => X"00c200cf00c800a2009c0088008e008900a200b200b1009f009600a30095008b",
            INIT_1D => X"008d0092009200930086007c007f0085009500a300ad00a600cc00f500f300f4",
            INIT_1E => X"00c300d000ad006e0071008b00b400b90085009a007f00570049004c0059005f",
            INIT_1F => X"005c0060005e00580056005600630067006d0074008f009b00af00e800f500f5",
            INIT_20 => X"00b700aa00a100650060008800b500a10080008400810087008c007d007d006a",
            INIT_21 => X"0035002b002c0027004d004700230028002000500091009700a700db00f600f3",
            INIT_22 => X"00ca00c100c2007c0078009200990049006900870083009400b8009f00a90083",
            INIT_23 => X"006600760084007a00af00aa006f0073006f009100b200b500bb00c500f200f4",
            INIT_24 => X"00d800c800b800720073009d00820024004f009500810063006f0081009d0084",
            INIT_25 => X"00b100c100b700b900c800c100ba00bd00b500c700b60097009400a200e800f6",
            INIT_26 => X"00d900cc00bb00710060008b0071003d004e00700073005d00550053005e007d",
            INIT_27 => X"00bf009f007f008a00a00095008c008f008a00bd009f00630073009a00e200f7",
            INIT_28 => X"00d500d000c700750049005c00630054004b004100610069005f00570067005f",
            INIT_29 => X"008600a200990097009600900089008f00930099008f006f0073009200de00f7",
            INIT_2A => X"00cc00ce00cc008300650051005c005a0046002d003900450062006f007d0057",
            INIT_2B => X"004a00660070006700620065005e007d0073005200710095009a008900d400f8",
            INIT_2C => X"00d100d000ce00750069007a0056005e005600360033002f0066008300ad0063",
            INIT_2D => X"002d0064009e00820079008a007c00ab00bb004b005f00ab0098007500cf00fa",
            INIT_2E => X"00dd00d600cc0068003b007400720080007c00410034003000380046006c004b",
            INIT_2F => X"0030005f00a6008f009100a7008f00af00af004a004800620054006800d600fb",
            INIT_30 => X"00d700d400c90063002f0044008000b0008700500038002d00280027002b002f",
            INIT_31 => X"0037003c0050006e007d00930090008b005c0043004600430045006d00d900fb",
            INIT_32 => X"00cf00cf00cb009d00730075008500aa007e006500480030002800290029002d",
            INIT_33 => X"00320027005300c000da00dc00c700c9006b00340038003f005a007e00d200f7",
            INIT_34 => X"00bc00c000ce00d800bf009a008600a1007900730068003e0021002200230029",
            INIT_35 => X"00330031005500b300c700c000be00bb0060002700260042006f008500d100f5",
            INIT_36 => X"00bf00c600cd00c600b5009e008400a000720076006f004600270026002c0031",
            INIT_37 => X"0044005d0069007e0087009600ad00a600480028002a00470071008200cf00f2",
            INIT_38 => X"00ce00d100c600b800ab00a300820085006b006f0068004d0032002f00350039",
            INIT_39 => X"003f0048005700680078009100a800b000450028003000470066007e00d400ee",
            INIT_3A => X"00c700c200c200bd00b200a600860065006300690060004f003e0036003b003e",
            INIT_3B => X"00410045004e0057006400740081008f00570027002c00470059008500df00e8",
            INIT_3C => X"00c100bc00be00bc00bd00bc00900050005a00630058004600490045004a004e",
            INIT_3D => X"004e004e0056005d00610066006d0072005e00300030004a006400ad00e800e7",
            INIT_3E => X"00c400c700d000cd00c800bb00a50055004c004c004e00540054005900620063",
            INIT_3F => X"005e00630072007c007d00810080007f0070005b00540060009400cc00e100df",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY29;


    MEM_GOLD_LAYER0_ENTITY0 : if BRAM_NAME = "gold_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00a0001200400104005100bc01010000000000470000001c0000000000ba0000",
            INIT_01 => X"0000000000000031000000000092000000000000000000000000000000000000",
            INIT_02 => X"000000000000000001040000000000020000000000000000000000a800000038",
            INIT_03 => X"0000000000000000000000020000000000000000000000000000005300370000",
            INIT_04 => X"0000000000000000000000000000000000000000000f00000000000000000000",
            INIT_05 => X"000000a8017a013400370113008200b7003500000000002d00790000014d0062",
            INIT_06 => X"00000000000000000000007e001000350000006a000000d10000000000000000",
            INIT_07 => X"00b000b0000000a00033007700d2008100c600000000000800a9005700000065",
            INIT_08 => X"00c8000000a1003c00000058007a00000000000000060000005c000000000000",
            INIT_09 => X"0000002c00e6000000770048000000ff00240000000000190000003600000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000005d004d00b5006c00aa00000000000000000000003f0000001b0030",
            INIT_0C => X"0015000000000000011900b300000012000000aa000000bd00b6002600000000",
            INIT_0D => X"0028000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000c001240144014f00d00068001700000040000000000009005700160000",
            INIT_0F => X"00cf005d00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000a8000100b8001e0028009600900015006300000000",
            INIT_11 => X"00000000000000000000000000000000000000000000000000000000011b009e",
            INIT_12 => X"00000000006c0000000000000000007900f80043000400ff0067001200110000",
            INIT_13 => X"0000001c00000069004100000086004e0031000000000091006c005100170026",
            INIT_14 => X"0046000000b000fd00e0000000780000001000000000000000000000005900ab",
            INIT_15 => X"00c100fb00ef006a008f00db003b00530014001000000000007b004600ab0062",
            INIT_16 => X"005a013c00a2006d008c007a01230051009700a10000000000000000003c0000",
            INIT_17 => X"000700000000000000000000000001040000000000000000001e004f00a2012f",
            INIT_18 => X"008c00000000015b013a0161008300a1007201380012000000000088007000dc",
            INIT_19 => X"00e000ad013e00cd00ae00000000000000000000000000000000000000c8001f",
            INIT_1A => X"00bf0046004b004e001b00260000001e0073013b009f0036001e000600aa00a5",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000006a0043007601010066007c000000000000000000000000",
            INIT_1E => X"000000000000000000000000000000590069000000310000000000000000003d",
            INIT_1F => X"0000000000100031007200ed000000000000000000000000000000000070012c",
            INIT_20 => X"017f00d0000000000000000000320000006700080039002100de006d00440076",
            INIT_21 => X"0084014100eb00000000000000000000000000000000000000b20078006e003f",
            INIT_22 => X"007f009200000000000000000000001c01910000001e00340087014800000000",
            INIT_23 => X"0000000000000000000000000058004a0046000000000000000000f300d700c5",
            INIT_24 => X"0000000000000000000000000118006b000000000031000000fe003a007101a4",
            INIT_25 => X"013000b600000000000000000000000000e3000000f300000000000000000000",
            INIT_26 => X"00000000000000000000000000000000000000000000000000000169004d00c7",
            INIT_27 => X"00f500aa002a00000100007800520000000000000000007601c0000000000000",
            INIT_28 => X"00000000000000000000000000000000000000000000000000000000007d0000",
            INIT_29 => X"00000000001100000000000000000074000000c80139000600b9000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000005c00000000000000000000000000000000",
            INIT_2C => X"000000000000000000450000000000c300eb016c01a101d500d401b401db0149",
            INIT_2D => X"000000000000007c0083005c0000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000079017600d100a000d4004d02030255",
            INIT_2F => X"0218022a027001b6012900000063000000000000000000590000000000000000",
            INIT_30 => X"00000000003d00da000000000000000000a8004a00dd005f014801d600220000",
            INIT_31 => X"0000000000af00000000000e0090018a00000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000000f900d4009000420137013d",
            INIT_33 => X"013800b700160000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000145019b00b80115014f01060000002c000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000b9016d019d0000029f",
            INIT_36 => X"00000000000000000000000000fb012100fa0000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000d30000000000d00083009f00000000",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000000000003d",
            INIT_39 => X"000f00000000000000000000000000000000000000000000006f003800000000",
            INIT_3A => X"0034003400000000008b00000079007a018e014300a000540000000000000000",
            INIT_3B => X"0000009000e40124009a00a400c20000002800a6000000080000000000000000",
            INIT_3C => X"006f000b000000e400db00ec016e009d005f01d9000000000000000000000000",
            INIT_3D => X"00000000000000000000000000000000000000000000000000000000008b001f",
            INIT_3E => X"001c000000000000003300000000000000000000000000000000000e00000000",
            INIT_3F => X"000000000000000000000000011b0000000000000000000000000000000000c1",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY0;


    MEM_GOLD_LAYER0_ENTITY1 : if BRAM_NAME = "gold_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009f009300000000000000000000000000f5000000dc00000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000000000000000000c500f5006f",
            INIT_02 => X"009e003c00d60000000000210000000000000000000000480260016100d3018f",
            INIT_03 => X"000200c101a300d10079008f01a4002f00000000000000000052005b007100b2",
            INIT_04 => X"0000002d006200b7009600e900dc0000010500080047006f00b001c501ed01db",
            INIT_05 => X"01b602dc01dc00000000000000000000000000fd00c000530000000000000000",
            INIT_06 => X"0000000000000000003700000000000000000000000000000000000001a700c7",
            INIT_07 => X"00c000b3006101040000000000700000004500c7016701c101ac011100e300d2",
            INIT_08 => X"00000031000000000000000000000000000000fe009f004a00000000000000ec",
            INIT_09 => X"00b3002500000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000000000000000000000000000000000000000000000000000840000002b",
            INIT_0B => X"00c20104008b00c2009d0074013100e100b900000000000000f100f7010c0000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000089000000270061",
            INIT_0E => X"0000000700000000000000000072006b00900000000000000000000000000007",
            INIT_0F => X"0000000000000000001f00000000003000000000000000000000000000000000",
            INIT_10 => X"0003004300000000000000000000018b00de0179003800a000530113010d009d",
            INIT_11 => X"000000000000004e001700d70025000000dc0000000000000000000000000000",
            INIT_12 => X"000000000014002a000d000000000000000000000000009900e5007c00a000df",
            INIT_13 => X"00a600c6007300a000230015000000230000000000000018001a000000000000",
            INIT_14 => X"00000000000000360000008200730057015800180045001e0066009c008c0000",
            INIT_15 => X"00000000000000670000001c0051000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000009000000000000018100cf00d0000000c500d5",
            INIT_17 => X"00b100cf00620000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000a200b40029009f005800530094006c006a00000000",
            INIT_19 => X"000000000000000000000000000000000050002c007e000000000063000000c0",
            INIT_1A => X"000000000000008500000000000000000022000000000000006700b000180012",
            INIT_1B => X"004900300000000000000000000000000000001d005900380028000000000000",
            INIT_1C => X"001c000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00d6007700710000000b0010000000110000000900000000000000000008001f",
            INIT_1E => X"00000092005300a200830000009000eb005400cc0000000b0000000000000000",
            INIT_1F => X"0000009300db009000b700b700a90032004d0020000c001b0000000000000000",
            INIT_20 => X"00100084000901500123011e000000000030006c00bb00890000000000000018",
            INIT_21 => X"0000004a00000000000000000000000000000000000000000000000000a000a7",
            INIT_22 => X"0051001200670000002800a9009c00000000000000000000000000000000002e",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000005000000000000000000480000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000007100bc0000",
            INIT_26 => X"00a500c90000005d0025000000000000002f0000000000000075003100490197",
            INIT_27 => X"0091013c005b0047007f001f0042000000410000004e013c000e000000ae006d",
            INIT_28 => X"007d00b40000011600a100010000003e0000000e00fc007d00d900fa00bb0182",
            INIT_29 => X"01020105014d000000000000000000000000003e004f000a0000000000000000",
            INIT_2A => X"000000000000000000000000000000000000001a005c000000000000019f00fc",
            INIT_2B => X"00c200e100940080010600b2007a00eb0107001100a5008e000000f5008e0074",
            INIT_2C => X"00370026000000000000000000a8014c0088000000000000000003050212002c",
            INIT_2D => X"0000006d0000000000750000010100a900000000000000000000000000000000",
            INIT_2E => X"0000000000000000001200c90054000000000000000000000000006a00000000",
            INIT_2F => X"00a001aa016a00000054006100000000000200000000000000a8000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000e10026001b00000000009700b400440000002c000000000083",
            INIT_32 => X"0000000000000056004a00240000000000000000000000000000000000000000",
            INIT_33 => X"00000000005f001300000000000a000000440091000a0000004800a300000000",
            INIT_34 => X"000700000000000000000000000000000000000000a9016700ac00bd015501ba",
            INIT_35 => X"000c009a0079008300140002000000a200170000000000000000000000000000",
            INIT_36 => X"00000000000000000000000e0080000a00270000006e0045010700ca000900f9",
            INIT_37 => X"00cd026602bc035e0077004d000000b5005f0119000000000000000000250000",
            INIT_38 => X"0000000000000006011700c50000000000000088005f0000008f013c01250000",
            INIT_39 => X"0000000000420000001f00ff008a00b800000000000000000000000000000000",
            INIT_3A => X"0000000000a4006b000000000000000000000000009f0060009a00d900340028",
            INIT_3B => X"0168016401780000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000c9011b0115004000770173007e000c002300000000",
            INIT_3D => X"0000000000000000000000000000000000be00a20000000000000137021c028e",
            INIT_3E => X"0000003e004900000000000000000073008a0093005a005300ff000000000000",
            INIT_3F => X"00000000000000000000000000000000000000000000008100a701810043005b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY1;


    MEM_GOLD_LAYER0_ENTITY2 : if BRAM_NAME = "gold_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009c0000000000000000000000000000000000000000000000000000000f0071",
            INIT_01 => X"00000000000000000000002d00000000000a002b000000000072004f003200c7",
            INIT_02 => X"003a000000530000000001db01760128008300cc009e002c003f0104008c0000",
            INIT_03 => X"0000012900640000007b0000008a007e005c000a000000000000004300000051",
            INIT_04 => X"0000000000000021002b00000000017800f100010024008d0079004200580060",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000030044",
            INIT_06 => X"000e00000096002b000000100008000000000000001f00000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000000000000000000000000003b",
            INIT_08 => X"00000000000000000050005a00f800620000000000e200000000000000000000",
            INIT_09 => X"00000000000000000000000000000000000000000000000000000051008700ae",
            INIT_0A => X"0000009000cf011a00e3010d00000000000000000091000000000052013800ae",
            INIT_0B => X"0047005000000197007c006a007f00f9002b00bc010100ef0000000000000098",
            INIT_0C => X"00e30000003d00210000017b010a003301c30162013b00890059013b00e70030",
            INIT_0D => X"01150113017f0000000000000000000000000063009b01320000000000000000",
            INIT_0E => X"00a50000000f0027000801aa00ca000001620000000000000000000001380164",
            INIT_0F => X"01580000009501920032002d015400420114007c0049015e00da012e0212026d",
            INIT_10 => X"003f000000000014000000000000007600000000000000000000000000000000",
            INIT_11 => X"0000000b00000009005500000036004900000000009c00000000000000000000",
            INIT_12 => X"00000000000000000000000000000000002b001c00000000000000aa010d0000",
            INIT_13 => X"00e000cf0074010e00b1004e0000000000000000000000000000000000710000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000034006100590000006e017c00320000010000c500a001d300ee009c00e8",
            INIT_16 => X"0190014e007500ed006900ff00fc00e6002e005500de000000d4006501260084",
            INIT_17 => X"0094007b00520000000000000000000000000000000000000000000000540000",
            INIT_18 => X"000000000000003e0000000000080083004f000300000000004c007300000000",
            INIT_19 => X"0000001600000000008300800032000000000069000000f5007700bf00ad0078",
            INIT_1A => X"005a0079000000fb0011000000a900760037000000000000001a000000000000",
            INIT_1B => X"00000008000000000000000000000000000000000000005a002a000800070000",
            INIT_1C => X"001a00000000001b000000000044008d0000003e000000000000006000000000",
            INIT_1D => X"001000000000001f001b00660010004800000000000000000000000000000000",
            INIT_1E => X"000000970037003d0059014a00be0086007300e100000000000000000000001c",
            INIT_1F => X"00000000002e0000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000002c002a00890048003700810039000100f800000000",
            INIT_21 => X"00000000000000000000000000000000003700000000003e0000003000000000",
            INIT_22 => X"00000000000000000000000000000000000000ee00d100b2015200d900ec001b",
            INIT_23 => X"008e009b00a600de006f0068000000420000000000000000000000000000000d",
            INIT_24 => X"00be0000003b00d300000000000000000000000000000000000000dd0151015c",
            INIT_25 => X"015600e600a90115009c0000000000000000000000000042000000000012010e",
            INIT_26 => X"00520078010f0000000000af0008002b00070000000000000000001700000055",
            INIT_27 => X"00b800000037000000000047000000390054000000000000000e003f00000000",
            INIT_28 => X"0000000000190000000000000000000000000000000000390047000000ad0075",
            INIT_29 => X"0000000c003f00f0000000000000000000000000000000000000000000f4010e",
            INIT_2A => X"019101530000000001a20166000000d100000017003b00000000000400150039",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000290000000000000000000000000000",
            INIT_2D => X"00000000000000000066000000000085003f0000000500a30000000000450000",
            INIT_2E => X"000000000060003c0000000000280005000000000000009200000000006d0000",
            INIT_2F => X"000000220095003e0000004a00a2000000000000000000000000000000000000",
            INIT_30 => X"0000000001110000003c00ab001600ce0000000000c7007f002b009600a50043",
            INIT_31 => X"00ba00dd001e0026015b00ab00d7003f000000f400da00000161015a013900f2",
            INIT_32 => X"00b2011b0190007b011400000000000000980000000000000044000000000000",
            INIT_33 => X"0000000000370000002300a60000000000000000000000000000000000000000",
            INIT_34 => X"007000a5010e00c6000000e000de0089008300190086007800a0005100540000",
            INIT_35 => X"0000000000000000000000000000003100000000000000000000000000000000",
            INIT_36 => X"000000000000000000e4011800cd002d00c40000003b00910096007d00000000",
            INIT_37 => X"0076002600000000000000000000000000560000000000d4003d0000002c0000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000048008a00be005d009700000056004e004d0003005c0000000100dd",
            INIT_3A => X"001a0000002a0020000000000055000000000000000000000000000000410000",
            INIT_3B => X"0000000000be002f002b000000000000001c0000000000000000000000000000",
            INIT_3C => X"00000026000000550000004900b00000000000000000001e0022003e00930025",
            INIT_3D => X"00340054003d004c00be0000000000290000006d000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000000000000000002b0000000000df",
            INIT_3F => X"00000000005a000000cf00860000006d001e0000000000320000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY3 : if BRAM_NAME = "gold_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000022004100000082002d004400ea010e0000",
            INIT_01 => X"000000000027002f000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000cf008700a400de00c200bf00c300cc00e4000000000000000000030000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000820070000000e4009d000000ae0073001000000000",
            INIT_05 => X"000000000000000000000000000000000000000000000000001b000000540000",
            INIT_06 => X"00000000000000000000000000000031007d00ed007e007201090000000000d3",
            INIT_07 => X"0023000000000000000000000000000000000000000000ca00b8009e00a60000",
            INIT_08 => X"003a00660000004e0092008f0083004e0006007c00db00b50136000000000000",
            INIT_09 => X"00000000000000000000004d0000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000040000000bc00f8001500e40031000000000000",
            INIT_0B => X"00000000000000000000000000000000000000000000000000000000004900a5",
            INIT_0C => X"006500000000000000000000005c003400c4000000000000002d006900700000",
            INIT_0D => X"0000006400b50084006f00000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000003b0000005c00c3000000bc00ae002a0078",
            INIT_0F => X"00000000000000000000000000000000004b0000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000094006e00ae00b90077012c006e00bc0077000000000000",
            INIT_12 => X"00000000000000470000000000190000005d0082007e0070008200aa00e30000",
            INIT_13 => X"0000000000000000000000000000007000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000011500ae00e000fe01450116",
            INIT_15 => X"0059011c00f5000000000000000000000000000000000000005a0057003400bc",
            INIT_16 => X"00ac0096006400660034003200000000000000000000004e008000a7005e000b",
            INIT_17 => X"0000000000000000000000000000000000250000000000c10000000000400060",
            INIT_18 => X"004b004001080120000900e200d300570169016d0215000401b9000000000000",
            INIT_19 => X"01b701da000000000000007300410000008f00af000000000000000000000000",
            INIT_1A => X"0000000000000000037c02790120014900000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000016000000000004b000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000000008009e013b01bf00eb003b000000be000000000000000000000134",
            INIT_1E => X"001e014200000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000e3000000000000006900d100fe00eb000e00000000000000000000",
            INIT_20 => X"00000000016300cc016c00d000ca00b400730000000000000065002600940156",
            INIT_21 => X"00000000006c0000000000860000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000001ec022f004200db0262",
            INIT_23 => X"005f009e008c000000c6017a00310027000d00000000006a0000001101b70000",
            INIT_24 => X"0170012000000000000000000051008c0148008200c400a400a1009701390000",
            INIT_25 => X"0000000000000000010000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000062002900e6011c0109009f0000000000000000000000000000",
            INIT_27 => X"0000000002360000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000008400aa00330040000000000000004600f500000000",
            INIT_29 => X"0000000000000000000000000000000000c80000019401f9008a000000000000",
            INIT_2A => X"028f026b016a01d2035600000127000000260000000000000000000000000000",
            INIT_2B => X"00000000000000000000000000000000008e020000d80135002a000000000000",
            INIT_2C => X"00000008000000000000000000fb000000000000000000000000000000000000",
            INIT_2D => X"0000008701cf003f0124000000110000000000f401120000012d000000590000",
            INIT_2E => X"004f00880084000000bc0000000000c7011501c9008201bf009a000000000046",
            INIT_2F => X"0000000000000000000000000089000001790000000000000000000000000028",
            INIT_30 => X"00d701ba019b00a602a201a8037400b301c70026027b02310064005e007a0053",
            INIT_31 => X"005a00d700ca0000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000001a009c00000000002b00780051000000b1009d",
            INIT_33 => X"00bb000000000000000000000000000000000000000000000000000000000078",
            INIT_34 => X"0000005000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000ce005901270017000000b3000000000037000000000000",
            INIT_36 => X"0000000000000000000000000224007f004000f3007200000175016801980000",
            INIT_37 => X"001100000000011e0000004501030000000000000000000000b5000000000078",
            INIT_38 => X"000000000000000000000000000000000000000002c801de0134012c02670182",
            INIT_39 => X"0154013801650000000000000000000000000000000000ad0000000000000010",
            INIT_3A => X"0000000000590000000000c3000000000000000000c1000000000010001a0153",
            INIT_3B => X"000000200000000000000000000001a501d1008901a00096000400af01340000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000033007500000000006f00000000002e000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000001e00000029002a017e01b50155",
            INIT_3F => X"00bd016801ea0081018f01e80000006f000000000016009100f100d3003d0000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY3;


    MEM_GOLD_LAYER0_ENTITY4 : if BRAM_NAME = "gold_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000e700000000010c0114000000e300b9000000fe00f2009200f601820143",
            INIT_02 => X"00810104013a0000000100cb00000000005c000000000021001a003600690064",
            INIT_03 => X"00930000012e00b3003600000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000500000000000000000000000000000000000000000000",
            INIT_05 => X"006600000038016600b50000011900000000004f00be0072001c013400900000",
            INIT_06 => X"0089004e002400110000000000010000000c0094002e0000000f008a00000000",
            INIT_07 => X"000000a400000000005e00600000009f000000810000000000ae000000000000",
            INIT_08 => X"000000000000000000000000000000000000000000000000002b000000000010",
            INIT_09 => X"000000cd013d0029000000600000000000000000000000000000000000000000",
            INIT_0A => X"000000000000000000b100000000001f0000000000000000002e000000000000",
            INIT_0B => X"0016000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000a3005e0000009600980000006300c3000000000000",
            INIT_0D => X"0000000000000000000000000000000000000018000000000000008700000000",
            INIT_0E => X"00000000000000000000000000000000000000cd00db014600d60089010b0000",
            INIT_0F => X"0072010400410000000000000071000000a700d2001b00a20075000900500130",
            INIT_10 => X"00c5000001150094000000000000000000000000000000000000008200000045",
            INIT_11 => X"00fd00460000000d0000000000000000003c0000000000190000000000000145",
            INIT_12 => X"0088002001e60066000e017200390000002100e6006900000024014c00000000",
            INIT_13 => X"012200000000000000000000006200000000008b000000000000000000000000",
            INIT_14 => X"0000000000050031000000000000000700000000000000000000005000b50055",
            INIT_15 => X"000000d100000000000b00000000000000000000000000000000000000000117",
            INIT_16 => X"0105000000ad00e800000000000d0070000000000000000e0000007b002f0000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000007c00bc0000001400a100000000000000000000000000000000",
            INIT_19 => X"0000000000000000007b0000000000140021000000160000000c000000760081",
            INIT_1A => X"00000000000d000000000000000000000000000000000000006a004400000062",
            INIT_1B => X"007d00000000003d005b00000084006100000000000000000000000000000000",
            INIT_1C => X"000000a700d1002d00000124001b0012011200250057005d008f006b004b007d",
            INIT_1D => X"01ad005700840000019c01b1000000b901f5009100eb01d200ae00b60079007f",
            INIT_1E => X"01390058009500fd009300000000003f004b00000010000000000000001600dd",
            INIT_1F => X"006a0000000000a900000000003e000000000000000000000000000000000000",
            INIT_20 => X"014000a9003500a20047004500af004900920000000000000000000000330000",
            INIT_21 => X"006200000000000000aa00000000001d00000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000000000000000000000000002e0050000000000000",
            INIT_23 => X"0000000000250034001c00000000003300000000000000120049001600b90000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000cf009d00f500bc001b00780000003c0064017700b1010c010100db00ec",
            INIT_26 => X"00aa00b800560137007a013100e800a0000000fd000e0072002000a70000000f",
            INIT_27 => X"005c0000000000150088000000000000000000000000000000000000014b001a",
            INIT_28 => X"004500000000000000000000004d001800000000000000120086003300410009",
            INIT_29 => X"0000000000050000000000000000003e00000022001800f10039001c00000000",
            INIT_2A => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000450030000000000065000000000023000000000000000000000000",
            INIT_2C => X"0000000000000000000000000032004600000000001700240000000000000060",
            INIT_2D => X"00000000000000000000002300aa000800000000000000000000000000000000",
            INIT_2E => X"0000014e011a0173010d00bb00010069007b011e000000000048004b000b0049",
            INIT_2F => X"0126015000a40000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000012000b002100dd00a4006d003500ab00a900000000",
            INIT_31 => X"00000000000000000000000000000000001c0000000000000000000000000000",
            INIT_32 => X"0000000000650000000000000000000000070010002f006400e900ca00000108",
            INIT_33 => X"00c0008a000000000000000000000000000000000000004e008200ab00cc0081",
            INIT_34 => X"0053006d00b8008100000000000000000000000000000000000001d1003a00e6",
            INIT_35 => X"008a005000710000000000000000000000000041000000000016000000000000",
            INIT_36 => X"0000000000000084000000000045000000000000008900920068008700ce0033",
            INIT_37 => X"0000002100b30000005600460036006700140000000000000000000000000000",
            INIT_38 => X"00000000000000470000000000000000000200000000000000f6010b0113010e",
            INIT_39 => X"004c0000009f0006004800000000000000000000000000000000000000c60000",
            INIT_3A => X"002600a20000002700770000000000dc00b5019f0000001800000049000f0069",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000540019000000000055003c000000380003000000000000",
            INIT_3E => X"00950062000200000010000000000000000000000000003500000000004c0098",
            INIT_3F => X"000b00190000000000b50000001b000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY4;


    MEM_GOLD_LAYER0_ENTITY5 : if BRAM_NAME = "gold_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000001200000000001d0090008800f200000080006f",
            INIT_01 => X"00aa00ef00f50000000000000000000000220000000000010000000e000000a9",
            INIT_02 => X"004b0097008a00a200d6000000b8000000000043000000000000000000000000",
            INIT_03 => X"0058000000000053004800000000000000000000000000000000000000000000",
            INIT_04 => X"014100000000019b000e0000004e010a00750032004d0000013a015601220000",
            INIT_05 => X"017201d40000000000000000000000000000000600ce00000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000aa00c8",
            INIT_07 => X"000000bb0000000000000000016000440000011c000000000000002c00620000",
            INIT_08 => X"000000000000000000000000000000000000000000000000000000000000002c",
            INIT_09 => X"000000b30000000000e5000000000060005800ec00000000017400000000002e",
            INIT_0A => X"0000000000000000000000000000000000000057000000000000000000000000",
            INIT_0B => X"00000000002e000000000000000c000000120000006b00000009000000000000",
            INIT_0C => X"0000006c00210029006e00820000005f008a009201790174019100bb00530000",
            INIT_0D => X"004b004100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000000000000000000003f00580048000000000000000001730000000001f8",
            INIT_0F => X"01ce0000009a00830000003c00690000006200000000000000000000002c0000",
            INIT_10 => X"000000150089000000b800ac0054006f000000de015a01d900c6012200810019",
            INIT_11 => X"0000000000000022009f00000000014400000000000000000000000000000000",
            INIT_12 => X"000000000000000000920000000000fb000000000169005600cb018c00070000",
            INIT_13 => X"00d90044003c0000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000000000000000000011000f90077016a0043000000d70000000000000000",
            INIT_15 => X"00000000000000000000000000000000009f0000000000420134000000fb00a9",
            INIT_16 => X"0000005400000000004b0019004c000000580000006500290000000000000063",
            INIT_17 => X"00000000000000000000003c00000000002b000400810064007700f200380000",
            INIT_18 => X"000000d70000000000000000000000000000000000000000000000000053007c",
            INIT_19 => X"00000000007b001a005400000161004000000174004200000000008500000017",
            INIT_1A => X"0018004a002e0000004d00ea00000000000f0000001a00000098000000000000",
            INIT_1B => X"0000008e0000000b00000035015200000000012400b90000000000d200000000",
            INIT_1C => X"0098000000740052000b005c01d1009e013100400111010b0027000000000000",
            INIT_1D => X"0000001501570000000000000000000000000000000000000000000000000000",
            INIT_1E => X"000000550000000000000000000000000000010d00000000000000c7005d004a",
            INIT_1F => X"0000000000000000000000000000000000080000000000000000002100c20000",
            INIT_20 => X"004f0043000000000000000000b9004e00000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000017000000000000000000000000000000690000",
            INIT_22 => X"000000db010a0000000000000000004d000000be002200480000006901440000",
            INIT_23 => X"000000c40000002600ef0000011e005500000127000000000087004e0058007f",
            INIT_24 => X"001f000000cf000000aa00d3002200000056000000e401a800ca0129017c0141",
            INIT_25 => X"00c001690184000000000000000000000000000000000000000000000000006f",
            INIT_26 => X"000000000000000000000000000000370000000000000102005e000000000082",
            INIT_27 => X"0064000000dc0000000000000000000000f90000000001ba0184000000ac00a4",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY5;



end a1;