-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_18k_layer1_entity1 is
    generic (
        DEVICE: string := "7SERIES"
        );
  
    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(10-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
  end ifmap_18k_layer1_entity1;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"001c00000000001a000400000000000000000003002f00000000000900040011",
       INIT_01 => X"00000000004a000c000000000000001b001f00000000000000000046009c0085",
       INIT_02 => X"002800000000000000200041001b0000000000000000000f0046000000000000",
       INIT_03 => X"0000000000000000000000000000000000020000000000000000000000000000",
       INIT_04 => X"0000000400070012000000000011000000000000000000000000000800000000",
       INIT_05 => X"0000000000000000001300000000000000000000000000000000000000140013",
       INIT_06 => X"00040000002800220000009d00a300a200a500a4009d00ac00b700ad0094007c",
       INIT_07 => X"007c00840092009200a200ad00a800ac00a0008c00a900a0007a003a002e003e",
       INIT_08 => X"004e006e008b0089006a00ac00b000af008e00730048002d0007001e000a0027",
       INIT_09 => X"003a0067004d002b00a400aa00a20059004d00270015000c0033002d001b0025",
       INIT_0A => X"003a0017001f00940060004e00470043002f001f0000003100390017001c002f",
       INIT_0B => X"00160012008e00990025003b00450031002d0000003e002a001000120017000e",
       INIT_0C => X"002a0062009f002f0032003e002d002f0000003200280010000e0026001c000a",
       INIT_0D => X"002c006200370026002e00270029001e002f002d00090022004100140000002b",
       INIT_0E => X"000e0055002200360030000d005400420026000f002d00790010000500240000",
       INIT_0F => X"0035002000080028002d0034001d000600090062008a00000015002300000017",
       INIT_10 => X"001a0000000000060000000000000000000000000000000000000006003a0000",
       INIT_11 => X"0000000000000000000000000000000000000000000000000034000000000000",
       INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_14 => X"0000000000000000000000000022002300250020001e002700260024001d0017",
       INIT_15 => X"001a00260024001e00180023002c002a001f00280020000f001d000e001d0000",
       INIT_16 => X"00090020002b001c00060039002800210027001a000000060021002e00000000",
       INIT_17 => X"00000025002c0000004c00210029000f00240004000000000048000000090000",
       INIT_18 => X"0000004a00000026000200560009000b00000000000000590000000000060000",
       INIT_19 => X"002b0000000a0000001a003e0013000000000000008e00000000001400000000",
       INIT_1A => X"0000000000200000003f0036000000000000006600000000000a001500000000",
       INIT_1B => X"00000000000000380042000000000000004200000000001d000f000800000002",
       INIT_1C => X"0000002100040011000000000024000000250000001e00210023000000000000",
       INIT_1D => X"002c0000000f00270000000200050000000c003000340014002a000400000078",
       INIT_1E => X"0000000000220000000000000008000900010000000000200014000000400000",
       INIT_1F => X"0000000000000000000000000000000000000000000000210043000000000000",
       INIT_20 => X"00000000000000000000000000000000000000000000005d0000000000000000",
       INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_22 => X"0000000000000000000400000000002b0030002d002c002f00290030003a0037",
       INIT_23 => X"002a002500260027002a0031002c00350030002e002d0000001f0029003b000c",
       INIT_24 => X"00000000000e001f0025001c0029002e00350032003b002d0023000000000000",
       INIT_25 => X"000000000004001a000000000023003200250019000000000000000000000000",
       INIT_26 => X"0006000000110000000000120018000000000000000000000000000000000000",
       INIT_27 => X"0000000500000000000b00380003000300000000000000000000000000000000",
       INIT_28 => X"0000000000000007003a00070000000000000000000000000000000000000000",
       INIT_29 => X"00000000000000000002000000000000000000000000000000000000000d0000",
       INIT_2A => X"0000000000000000001a000500000000000f0003001800040000000800000000",
       INIT_2B => X"000000000000000000000000000000080011000a00000000001f000000000000",
       INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_30 => X"00000000000000000000000000000000000a0011000800080004000c000c000b",
       INIT_31 => X"000b0021002d00230011000800060000000a000a000c00080000000500230042",
       INIT_32 => X"000000000000000a0017000a0035003300050008000500370016000900000000",
       INIT_33 => X"000000000000000e000c000000000005000800080000000000020000001a0004",
       INIT_34 => X"001000060000000e000100000002000e00000000000900000007000000000000",
       INIT_35 => X"000000000000000f000000060003003e00280000000000000000001400150007",
       INIT_36 => X"0000000000000000001c00180012000000310000001100000011000000000000",
       INIT_37 => X"000000000000000000000002003500350021000e0000000900000005000e0000",
       INIT_38 => X"000000010000000000000026000000000000000000260030000000000000000c",
       INIT_39 => X"00000004000000230009000000000000004e0036001100000000001800030000",
       INIT_3A => X"0007000000000000001e0051003700000000000000000005000a00350021000c",
       INIT_3B => X"0000005600280004000500030000000000000000000000000000001600000018",
       INIT_3C => X"003f0000000000000000000000000000000000000000000000000018004f000b",
       INIT_3D => X"0000000000000000000000000000000000000014000000000000002200000003",
       INIT_3E => X"001200000000000000000000000000000000000d0013000a000e000900150008",
       INIT_3F => X"0006000c001c0022001b0013000600020008000b0009000d000f0036000f001a",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
