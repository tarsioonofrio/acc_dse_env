library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    4309, -4548, 1922, -1687, 1872, -2230, -4892, -4908, 8348, -4973, -5603, 15533, 2609, 7923, 8185, -989, 951, -10732, -2628, -784, -8448, -3995, -1956, 6940, 1563, 12563, 5468, -3873, -5359, 9306, -3817, -11036,

    -- weights
    -- filter=0 channel=0
    -9, 3, 6, -40, -35, -2, -36, -20, 2,
    -- filter=0 channel=1
    -20, -7, -19, -18, 2, -20, 17, 20, -8,
    -- filter=0 channel=2
    23, 23, 5, -14, 19, -5, 10, -9, -15,
    -- filter=0 channel=3
    7, -17, 13, -18, -17, 31, -5, 7, 20,
    -- filter=0 channel=4
    11, -3, 14, 0, 5, -10, 14, -5, 9,
    -- filter=0 channel=5
    18, 24, 17, 13, -1, 8, 6, -7, -10,
    -- filter=0 channel=6
    34, 15, 29, 6, -3, 20, -5, 26, -5,
    -- filter=0 channel=7
    10, -5, 2, -18, -22, -15, 12, -3, -11,
    -- filter=0 channel=8
    23, 5, 27, 0, 0, 24, -6, 0, 24,
    -- filter=0 channel=9
    11, -5, 7, 23, 16, 13, 10, -4, 11,
    -- filter=0 channel=10
    6, 2, 27, 31, 29, -10, 6, 21, 13,
    -- filter=0 channel=11
    -16, 6, -13, 3, 18, -9, -3, 20, -9,
    -- filter=0 channel=12
    17, -1, 14, 0, 1, 16, -4, 6, 30,
    -- filter=0 channel=13
    0, 14, 8, -22, -13, -12, 0, 3, 6,
    -- filter=0 channel=14
    -4, -2, -14, 6, 9, -5, -14, -1, 18,
    -- filter=0 channel=15
    -6, 2, -15, -14, -11, -3, 7, 1, 10,
    -- filter=1 channel=0
    13, 2, 31, -6, 3, 23, 15, 9, 12,
    -- filter=1 channel=1
    3, -3, 18, -3, -16, -6, -11, 0, 4,
    -- filter=1 channel=2
    -10, 9, 4, -26, -21, -12, -9, -26, -17,
    -- filter=1 channel=3
    12, 13, 11, 0, -19, -16, -5, 8, 20,
    -- filter=1 channel=4
    -29, -22, -29, 4, -13, -30, -24, -6, -5,
    -- filter=1 channel=5
    -16, 23, -13, 9, -8, 0, -8, 0, -12,
    -- filter=1 channel=6
    -28, -6, 3, -5, -21, 18, -1, -6, -11,
    -- filter=1 channel=7
    0, 9, 5, -4, -3, 7, -5, 11, -6,
    -- filter=1 channel=8
    -5, -31, -8, -19, -6, -14, -10, -3, 0,
    -- filter=1 channel=9
    -2, -12, -2, 24, 24, 22, -10, 17, 24,
    -- filter=1 channel=10
    -4, 11, -25, 0, -11, -16, 11, -13, -21,
    -- filter=1 channel=11
    20, -12, -13, 13, 16, 14, 12, 19, 17,
    -- filter=1 channel=12
    -7, 11, 27, 4, -9, 24, -2, 5, 17,
    -- filter=1 channel=13
    -17, -16, 0, -12, -19, 21, 14, 19, 2,
    -- filter=1 channel=14
    -8, -14, -1, -14, 10, -8, -7, 15, 10,
    -- filter=1 channel=15
    -16, 16, 37, -6, 21, 12, 10, 5, -6,
    -- filter=2 channel=0
    3, 7, -11, -18, 8, 19, 15, -10, 0,
    -- filter=2 channel=1
    10, -16, -6, -13, -10, -9, -15, 14, -8,
    -- filter=2 channel=2
    -20, 14, -10, -14, -14, 18, 7, -19, 20,
    -- filter=2 channel=3
    3, -20, -8, 15, 10, 0, -5, -1, -21,
    -- filter=2 channel=4
    4, 8, -1, 6, -7, -10, 12, 17, 9,
    -- filter=2 channel=5
    17, 0, 0, 0, -3, -12, -20, 15, 9,
    -- filter=2 channel=6
    3, -11, -2, -6, -11, 6, 15, 0, -20,
    -- filter=2 channel=7
    11, -17, -12, 3, -7, 7, -4, 20, -20,
    -- filter=2 channel=8
    -15, -11, -20, 4, 19, 2, 9, 4, -4,
    -- filter=2 channel=9
    7, -7, 6, -14, -7, 2, -5, 14, -8,
    -- filter=2 channel=10
    -6, -4, 7, -5, -14, 1, -1, 0, -16,
    -- filter=2 channel=11
    9, -21, 6, -4, -15, -3, 4, 3, 17,
    -- filter=2 channel=12
    -6, -11, -15, -8, -5, 12, 1, 18, 3,
    -- filter=2 channel=13
    -14, -17, -5, -13, -1, 18, -16, -11, -13,
    -- filter=2 channel=14
    -14, -1, -1, -8, -16, -17, 8, -14, 10,
    -- filter=2 channel=15
    3, -15, 14, 6, -19, -15, -12, -7, 0,
    -- filter=3 channel=0
    12, 1, -14, 0, 3, 3, 7, 18, 10,
    -- filter=3 channel=1
    -16, -7, -1, 7, 14, 9, 5, -7, -21,
    -- filter=3 channel=2
    16, 20, -8, -15, -11, -5, 10, 17, 13,
    -- filter=3 channel=3
    -20, -15, 6, -1, -10, 10, -14, 0, 15,
    -- filter=3 channel=4
    -16, -16, -16, 20, -11, 16, -17, 0, 13,
    -- filter=3 channel=5
    0, 10, -12, -13, 15, 0, 5, -6, 3,
    -- filter=3 channel=6
    -1, 20, 5, -20, -20, 0, 20, -1, 18,
    -- filter=3 channel=7
    13, -3, -20, -3, -5, 7, 2, -14, 4,
    -- filter=3 channel=8
    -1, 12, 15, -12, -15, -3, 14, -15, -11,
    -- filter=3 channel=9
    15, 14, -7, 13, -13, 13, -19, 11, -18,
    -- filter=3 channel=10
    20, -20, 2, 13, -3, -20, -19, -6, -2,
    -- filter=3 channel=11
    -17, 10, 0, -8, 5, 0, -19, 9, 9,
    -- filter=3 channel=12
    19, -16, -11, 7, -8, 0, 2, -19, 14,
    -- filter=3 channel=13
    -5, -1, -6, 6, -16, -15, -12, -12, 13,
    -- filter=3 channel=14
    -1, 16, -3, 20, 0, -11, 16, -6, 13,
    -- filter=3 channel=15
    -7, 9, -9, -17, -16, -17, 15, 19, -13,
    -- filter=4 channel=0
    16, 17, 3, 26, -2, 24, 5, 27, 0,
    -- filter=4 channel=1
    0, 0, 5, -9, 14, 0, -6, -9, -14,
    -- filter=4 channel=2
    2, -14, 10, 8, 1, 8, 6, 1, 0,
    -- filter=4 channel=3
    10, -18, -25, -13, 6, 3, 4, -6, -17,
    -- filter=4 channel=4
    -12, -15, 10, -1, -1, 14, 10, 0, 16,
    -- filter=4 channel=5
    1, -4, 4, 10, 12, 20, 5, 11, -2,
    -- filter=4 channel=6
    -14, 24, 12, -14, 19, 17, -13, 24, -1,
    -- filter=4 channel=7
    16, -13, -12, 11, 16, 0, -9, 2, -7,
    -- filter=4 channel=8
    -9, -28, -2, -4, -15, -24, -20, -3, 2,
    -- filter=4 channel=9
    -15, -11, 11, 11, -6, 15, 10, -19, -16,
    -- filter=4 channel=10
    -1, -18, -12, -3, 12, -18, 4, 7, -8,
    -- filter=4 channel=11
    8, 2, -8, 20, -2, 17, 17, -20, 0,
    -- filter=4 channel=12
    5, 6, -22, 12, 9, -13, 12, -6, -6,
    -- filter=4 channel=13
    0, -2, 0, -9, -4, -3, -6, 2, 5,
    -- filter=4 channel=14
    5, 17, 6, -21, 7, -19, -20, 15, -13,
    -- filter=4 channel=15
    34, 28, 36, 15, 19, 27, 17, 0, 35,
    -- filter=5 channel=0
    6, 13, -8, -5, 22, 1, 26, -8, -6,
    -- filter=5 channel=1
    -19, 17, 4, 8, -8, -4, -10, 16, -16,
    -- filter=5 channel=2
    6, 20, 0, -17, -17, 16, 20, 19, -10,
    -- filter=5 channel=3
    -11, -15, 0, -1, 9, 7, 0, -4, -22,
    -- filter=5 channel=4
    -6, -9, -18, 14, -14, -2, -6, 15, 6,
    -- filter=5 channel=5
    -9, 9, 18, -16, -2, 11, -4, -17, -4,
    -- filter=5 channel=6
    -7, -19, 9, -13, 0, 19, -21, -12, 6,
    -- filter=5 channel=7
    -6, 10, -8, -18, -4, -13, 9, 5, -15,
    -- filter=5 channel=8
    -12, 12, 14, 9, 5, 13, 21, 5, -3,
    -- filter=5 channel=9
    14, 10, 4, -2, 19, 0, -16, 12, 6,
    -- filter=5 channel=10
    -21, -6, -17, 8, -16, -4, -6, -15, 2,
    -- filter=5 channel=11
    19, 16, -18, 5, 16, -16, -18, 16, 6,
    -- filter=5 channel=12
    22, 0, -9, 9, 0, 6, 22, -15, -9,
    -- filter=5 channel=13
    12, 7, -10, 13, 26, -17, 4, 25, 11,
    -- filter=5 channel=14
    9, -17, -6, 11, -11, 1, 9, 7, 13,
    -- filter=5 channel=15
    -8, 3, -19, 14, 0, -5, 21, -4, 7,
    -- filter=6 channel=0
    17, 18, -12, -13, -4, -2, -10, 8, -9,
    -- filter=6 channel=1
    -4, 19, -1, 5, 4, 15, -19, 12, 14,
    -- filter=6 channel=2
    -5, -15, 6, 6, 13, 14, 12, -16, 3,
    -- filter=6 channel=3
    10, -20, -12, 19, -16, -12, -14, 3, -14,
    -- filter=6 channel=4
    3, -19, -9, 17, -3, 4, 12, -17, -10,
    -- filter=6 channel=5
    12, -16, 18, -18, -17, 16, -2, 2, 7,
    -- filter=6 channel=6
    -14, -20, -18, 2, 0, -18, 1, -13, -6,
    -- filter=6 channel=7
    -4, 0, -14, -6, -6, -19, 14, -19, 9,
    -- filter=6 channel=8
    2, -2, 7, 5, -9, -4, -18, 7, -12,
    -- filter=6 channel=9
    3, -15, -19, 17, 1, 4, -6, -9, 0,
    -- filter=6 channel=10
    -8, -16, -4, 11, -20, -20, 17, 15, 0,
    -- filter=6 channel=11
    -16, 8, 12, -9, -11, 2, 16, 6, -17,
    -- filter=6 channel=12
    -12, 8, 17, -5, -18, 11, -14, -18, 20,
    -- filter=6 channel=13
    6, 19, -14, -8, -14, 16, -4, 13, 18,
    -- filter=6 channel=14
    4, -7, 11, -8, -18, -12, -19, -10, 0,
    -- filter=6 channel=15
    -3, 0, -3, -9, -8, -7, 10, -7, -13,
    -- filter=7 channel=0
    7, 15, 31, -9, -9, 32, -19, 25, 19,
    -- filter=7 channel=1
    -2, -3, -6, 20, -8, 0, 19, 8, -5,
    -- filter=7 channel=2
    12, 0, 2, -22, -23, -6, 6, -15, -25,
    -- filter=7 channel=3
    19, 29, 9, 15, 17, 32, -7, 20, 19,
    -- filter=7 channel=4
    -6, -19, 4, 9, -24, -16, -13, 9, 18,
    -- filter=7 channel=5
    -17, -18, -11, 0, 5, -4, 0, 17, 7,
    -- filter=7 channel=6
    -15, -13, -10, 13, 4, -19, 1, 20, 9,
    -- filter=7 channel=7
    -14, 11, -7, 5, 0, -11, -10, 18, 9,
    -- filter=7 channel=8
    11, 11, -9, 12, 2, -9, 2, 2, -22,
    -- filter=7 channel=9
    -12, -1, -22, 0, -4, -12, -15, -16, 18,
    -- filter=7 channel=10
    6, 4, 7, 16, -1, 1, 3, -5, -10,
    -- filter=7 channel=11
    -6, 12, 18, -17, -18, -12, -3, 2, 18,
    -- filter=7 channel=12
    24, 12, -7, 30, 11, 29, 0, -7, 19,
    -- filter=7 channel=13
    13, 6, -10, 12, 14, 33, 13, 18, 16,
    -- filter=7 channel=14
    10, 13, 20, -8, 9, -11, 10, 15, 17,
    -- filter=7 channel=15
    1, 22, 20, -6, -18, 15, -6, 16, -1,
    -- filter=8 channel=0
    1, 10, -26, -7, -17, 13, -13, 1, 14,
    -- filter=8 channel=1
    -10, 2, -9, 5, -9, 4, 19, 14, -14,
    -- filter=8 channel=2
    -19, -10, -1, 10, -14, -16, 7, 16, -1,
    -- filter=8 channel=3
    -11, 17, -23, 11, 6, -22, 22, -14, -11,
    -- filter=8 channel=4
    -16, 3, -8, -3, 15, -14, -3, -18, -7,
    -- filter=8 channel=5
    -13, 6, 5, 5, 4, 20, 18, 6, 23,
    -- filter=8 channel=6
    7, -9, 13, 16, -14, 13, 8, 20, 22,
    -- filter=8 channel=7
    -12, -8, -6, 5, 21, 6, -20, 20, -7,
    -- filter=8 channel=8
    21, -12, 19, 13, 19, 14, 10, 23, -4,
    -- filter=8 channel=9
    20, -12, 6, 14, -4, 0, -18, -2, 14,
    -- filter=8 channel=10
    -4, 22, 22, 8, -14, 9, -17, -15, 25,
    -- filter=8 channel=11
    -4, 18, -1, -1, 0, -13, -2, -9, 0,
    -- filter=8 channel=12
    -10, -12, -20, 17, -7, -18, 18, -21, -23,
    -- filter=8 channel=13
    0, 3, 5, 24, -17, -7, 0, -9, 8,
    -- filter=8 channel=14
    0, 4, 18, -1, -2, -5, 9, 11, 2,
    -- filter=8 channel=15
    9, 0, -19, -13, 19, -21, 8, -1, -22,
    -- filter=9 channel=0
    -1, 16, 20, -10, -7, -16, -9, -21, -18,
    -- filter=9 channel=1
    -7, 16, 6, 6, 10, 17, -9, 8, -5,
    -- filter=9 channel=2
    12, -13, 9, -18, 0, -3, 3, 2, -13,
    -- filter=9 channel=3
    9, 2, 7, 16, 9, 4, -21, 8, -10,
    -- filter=9 channel=4
    12, 26, 27, 24, 0, -9, 14, 29, 28,
    -- filter=9 channel=5
    -13, -6, -18, 19, 19, 15, 21, 5, 7,
    -- filter=9 channel=6
    -4, -12, 9, -3, 5, 15, 27, 25, -3,
    -- filter=9 channel=7
    12, -20, -2, -2, -9, -9, 0, -8, -20,
    -- filter=9 channel=8
    -8, 16, 15, 9, 21, -9, -3, -12, 20,
    -- filter=9 channel=9
    -19, 13, -14, -15, 5, 18, 10, -5, 21,
    -- filter=9 channel=10
    5, -4, -9, 11, -6, -3, 19, 1, 4,
    -- filter=9 channel=11
    -12, 19, -19, -17, -16, -9, 6, 4, 12,
    -- filter=9 channel=12
    -9, 18, 3, 12, -8, 2, -16, 15, -8,
    -- filter=9 channel=13
    2, -8, 1, 19, -8, -15, -15, 14, -9,
    -- filter=9 channel=14
    10, 11, -3, 20, 17, -16, 14, 14, 13,
    -- filter=9 channel=15
    -6, 11, -13, 9, 17, 5, 3, 12, -4,
    -- filter=10 channel=0
    23, -4, 10, 30, 20, -4, 16, 0, -16,
    -- filter=10 channel=1
    -2, 9, -16, 1, -11, -20, -12, -12, 17,
    -- filter=10 channel=2
    15, 19, -12, -14, -19, -10, -16, 18, 17,
    -- filter=10 channel=3
    0, -18, -24, -18, 1, -18, 13, -2, -4,
    -- filter=10 channel=4
    4, 1, -13, 23, -8, 19, 0, 16, 11,
    -- filter=10 channel=5
    -1, -15, 9, 20, -14, -7, -15, 18, -3,
    -- filter=10 channel=6
    20, -4, -4, 3, 2, 17, -16, 21, 19,
    -- filter=10 channel=7
    -15, -7, -7, 13, 11, -5, -19, 9, -4,
    -- filter=10 channel=8
    -12, -15, -2, -13, -18, 19, -9, 13, -13,
    -- filter=10 channel=9
    -21, -17, -14, 16, 0, 11, -23, -3, -16,
    -- filter=10 channel=10
    -13, -2, 18, 12, 10, 8, -1, -15, -11,
    -- filter=10 channel=11
    -1, 4, -2, -17, -20, -7, 7, -12, -16,
    -- filter=10 channel=12
    8, -12, -15, 17, -17, 7, 14, 2, -23,
    -- filter=10 channel=13
    6, 21, 8, 15, -13, 18, 14, -19, -14,
    -- filter=10 channel=14
    -8, -19, -9, 12, 2, 14, 4, -9, -3,
    -- filter=10 channel=15
    25, -9, 4, -2, 26, 6, 28, -12, 0,
    -- filter=11 channel=0
    11, 6, -14, -13, -6, -14, -6, -25, 13,
    -- filter=11 channel=1
    -6, -3, -10, -15, -21, 0, 18, 10, -16,
    -- filter=11 channel=2
    -9, 11, -15, 16, -9, -4, -10, 0, -6,
    -- filter=11 channel=3
    6, 0, 19, 16, -7, 17, -5, -13, -5,
    -- filter=11 channel=4
    5, 5, -13, 15, 9, -6, -20, 3, 2,
    -- filter=11 channel=5
    -12, 7, 16, 14, 3, -13, -10, -3, -16,
    -- filter=11 channel=6
    -13, 11, 20, -10, 21, 12, 5, 11, -7,
    -- filter=11 channel=7
    4, 21, 29, 24, 28, 25, 11, 30, 5,
    -- filter=11 channel=8
    22, 19, 6, 13, -6, 6, -6, -1, 28,
    -- filter=11 channel=9
    1, 31, 0, 11, 15, 28, -2, 14, 29,
    -- filter=11 channel=10
    10, 10, 30, 12, -4, 29, -1, -2, 29,
    -- filter=11 channel=11
    12, 15, -5, 10, 5, 1, 4, 17, 17,
    -- filter=11 channel=12
    24, -2, 28, 22, 20, 8, -4, -1, 17,
    -- filter=11 channel=13
    13, -28, -17, -23, -23, -4, -12, -18, -1,
    -- filter=11 channel=14
    15, 3, -13, 13, 1, 12, 0, 9, 17,
    -- filter=11 channel=15
    5, -35, -32, -30, 3, 7, -30, -28, 1,
    -- filter=12 channel=0
    14, -9, -11, -8, 5, -13, -5, 3, 10,
    -- filter=12 channel=1
    10, -2, 15, -10, -2, -9, 19, 16, 14,
    -- filter=12 channel=2
    -7, 12, -18, 13, -8, -6, 11, 11, 5,
    -- filter=12 channel=3
    6, 5, 11, -17, 27, 11, -16, -9, 13,
    -- filter=12 channel=4
    14, -12, 7, 25, -4, 12, 17, 18, 14,
    -- filter=12 channel=5
    17, 17, -8, 5, -1, -6, 14, -2, 0,
    -- filter=12 channel=6
    -18, 0, 11, 23, 2, 2, 24, -2, 11,
    -- filter=12 channel=7
    -16, 19, 2, 16, -14, -23, -22, -1, 11,
    -- filter=12 channel=8
    11, 8, -14, -19, 6, 7, 0, 7, 10,
    -- filter=12 channel=9
    13, -24, -22, -13, -7, -18, -9, -11, 15,
    -- filter=12 channel=10
    -7, -8, 16, 24, 20, 17, 8, 5, -14,
    -- filter=12 channel=11
    20, -5, -17, -10, -2, -18, -19, -16, 8,
    -- filter=12 channel=12
    4, 17, 24, 24, 25, 29, 6, -5, 1,
    -- filter=12 channel=13
    5, 22, 22, 8, 3, 24, -4, 17, -5,
    -- filter=12 channel=14
    -10, -20, -6, 3, -10, -2, 20, -13, -3,
    -- filter=12 channel=15
    8, -7, 18, -2, -27, -21, -7, -25, -24,
    -- filter=13 channel=0
    -3, -6, -17, -7, -25, -21, -25, -31, 0,
    -- filter=13 channel=1
    -20, -9, 16, 0, 12, 15, -19, 19, -7,
    -- filter=13 channel=2
    6, 9, 18, 22, 8, -11, 4, 10, -3,
    -- filter=13 channel=3
    1, -4, 8, 18, -5, 14, 6, 28, 15,
    -- filter=13 channel=4
    3, -28, -28, -19, -18, -8, -31, -8, -28,
    -- filter=13 channel=5
    -17, -2, -5, 11, 10, 7, 11, 4, -23,
    -- filter=13 channel=6
    -32, -23, -36, -31, -27, -38, -14, -11, -8,
    -- filter=13 channel=7
    12, 2, 9, -24, 10, 0, -23, -22, -1,
    -- filter=13 channel=8
    38, 6, 36, 36, 22, 17, 29, 30, 19,
    -- filter=13 channel=9
    -20, -22, 11, -4, -1, -5, -8, -6, -12,
    -- filter=13 channel=10
    10, 23, 0, 5, -2, 23, 4, 22, -1,
    -- filter=13 channel=11
    -13, 0, -16, 9, 20, 16, 0, 9, -18,
    -- filter=13 channel=12
    -7, 16, 21, 9, 24, 36, 24, 27, 32,
    -- filter=13 channel=13
    21, 25, 35, 15, 21, 27, -7, -1, 27,
    -- filter=13 channel=14
    -18, -13, 7, 6, -20, 20, -10, 14, -4,
    -- filter=13 channel=15
    -35, -21, -17, -23, -23, -10, -44, -46, -21,
    -- filter=14 channel=0
    -22, 22, -10, 0, -7, 22, -25, 0, 15,
    -- filter=14 channel=1
    -16, 11, -11, -11, 5, -1, -18, -17, 17,
    -- filter=14 channel=2
    -21, 0, -14, 10, -16, -18, -15, -24, 0,
    -- filter=14 channel=3
    12, 0, -9, 1, -15, -10, -4, 10, 20,
    -- filter=14 channel=4
    -1, -8, 3, -34, -20, -23, -1, 1, -21,
    -- filter=14 channel=5
    15, -1, 6, 3, 24, 12, -12, 8, -1,
    -- filter=14 channel=6
    3, 11, 21, -9, -11, 8, -1, -14, -9,
    -- filter=14 channel=7
    21, 10, 2, 2, 30, 0, 26, -4, 17,
    -- filter=14 channel=8
    -29, -20, -25, -19, -4, -5, -10, -31, -1,
    -- filter=14 channel=9
    17, -2, -12, 28, 27, 16, 8, 15, 3,
    -- filter=14 channel=10
    4, -12, 10, 2, -19, -16, 8, -21, -1,
    -- filter=14 channel=11
    19, 9, -18, 6, -12, 11, 12, -4, 13,
    -- filter=14 channel=12
    21, -5, 32, 1, 7, 25, 21, 2, 22,
    -- filter=14 channel=13
    -26, 11, 19, -25, -21, -8, -30, -3, -1,
    -- filter=14 channel=14
    1, 9, 13, 6, 9, -13, -16, -21, -10,
    -- filter=14 channel=15
    -4, 1, 12, 10, -21, 24, -2, 15, 4,
    -- filter=15 channel=0
    13, 4, -10, 11, 0, 8, -8, -12, -4,
    -- filter=15 channel=1
    15, -18, 17, 16, 1, -15, -20, -3, 3,
    -- filter=15 channel=2
    0, 17, 0, 11, 0, -12, -3, -6, 3,
    -- filter=15 channel=3
    6, 4, 6, 10, 30, -3, 10, -9, -7,
    -- filter=15 channel=4
    15, 19, 15, -11, 8, 8, -8, 14, -6,
    -- filter=15 channel=5
    -6, -22, 3, -17, 1, -2, -23, -22, 2,
    -- filter=15 channel=6
    -18, -24, -17, -7, 0, -14, -23, -5, -25,
    -- filter=15 channel=7
    -15, -22, -26, -3, -8, -4, 0, 11, -11,
    -- filter=15 channel=8
    -5, 13, -7, 19, 31, 2, 22, 20, 22,
    -- filter=15 channel=9
    0, -2, -20, 12, -23, -21, -15, -24, 15,
    -- filter=15 channel=10
    -14, -8, 15, 5, -11, 18, 12, -13, 21,
    -- filter=15 channel=11
    -20, -15, 16, -11, 15, -20, 17, -20, -16,
    -- filter=15 channel=12
    -7, -3, -5, 20, 10, -4, 23, -7, 19,
    -- filter=15 channel=13
    31, 0, 8, 23, 24, -4, 7, -6, -8,
    -- filter=15 channel=14
    15, 8, -11, -8, 0, 4, -21, -14, -12,
    -- filter=15 channel=15
    5, -4, -9, -27, -28, -22, 6, -25, 1,
    -- filter=16 channel=0
    28, 15, 2, 8, 28, 22, 24, 25, -9,
    -- filter=16 channel=1
    15, 0, 12, 7, 12, 19, -14, 18, 15,
    -- filter=16 channel=2
    -16, -1, 1, -5, 13, -14, 0, -24, -18,
    -- filter=16 channel=3
    -16, 7, 0, -11, -19, -3, 0, -4, 9,
    -- filter=16 channel=4
    -31, -1, -12, -3, 6, 9, -26, -3, -23,
    -- filter=16 channel=5
    -2, -1, -10, 0, 14, 13, -12, -3, -12,
    -- filter=16 channel=6
    2, 7, -18, 9, -17, -23, 6, -20, -21,
    -- filter=16 channel=7
    -12, 20, 1, 17, 5, 29, 10, 11, 11,
    -- filter=16 channel=8
    -13, -6, -11, 8, -20, -16, -3, -6, -10,
    -- filter=16 channel=9
    -5, 3, 13, 23, 0, -11, -1, 4, 25,
    -- filter=16 channel=10
    -17, -12, 10, 5, -12, 10, -22, 12, -4,
    -- filter=16 channel=11
    1, -2, 15, 16, 11, -14, -16, 0, 14,
    -- filter=16 channel=12
    -6, -16, 9, -12, 7, 2, 22, 19, 3,
    -- filter=16 channel=13
    -8, -4, 6, -14, 6, -26, -23, 0, -7,
    -- filter=16 channel=14
    9, 5, 21, 18, 4, 3, -16, -14, -13,
    -- filter=16 channel=15
    5, 9, 0, -16, -2, -7, -5, -22, -12,
    -- filter=17 channel=0
    -5, 16, 14, 30, 18, 22, 22, 31, 23,
    -- filter=17 channel=1
    20, -9, 14, -3, 12, -11, -4, 14, -12,
    -- filter=17 channel=2
    -17, 17, -9, -4, -15, -21, 14, 9, -21,
    -- filter=17 channel=3
    35, 28, -20, 22, 22, -5, 36, 25, -21,
    -- filter=17 channel=4
    -15, -30, -21, -21, -1, -12, -21, 11, -9,
    -- filter=17 channel=5
    -31, -23, 10, -21, -18, 9, -7, 18, 17,
    -- filter=17 channel=6
    -21, -13, -15, -22, -22, -7, -18, -11, -17,
    -- filter=17 channel=7
    -8, 2, -10, -1, 0, 11, -14, -17, -3,
    -- filter=17 channel=8
    11, 4, 12, 21, 4, -9, 27, 14, 6,
    -- filter=17 channel=9
    -14, -13, -25, 3, -18, 3, 11, 13, 8,
    -- filter=17 channel=10
    -14, 5, -14, 8, -17, 2, -3, -12, -16,
    -- filter=17 channel=11
    -16, -2, -10, -3, -2, 4, -1, 16, 16,
    -- filter=17 channel=12
    0, 1, -25, 25, 1, 0, 12, 23, -2,
    -- filter=17 channel=13
    39, 34, 21, 27, 0, -1, 27, 32, 8,
    -- filter=17 channel=14
    -3, 3, 11, 16, 3, 2, 10, -7, -17,
    -- filter=17 channel=15
    -16, 2, 34, -9, 9, 24, 6, -16, 1,
    -- filter=18 channel=0
    8, 26, 26, 17, 15, -13, 7, 29, 23,
    -- filter=18 channel=1
    -11, 0, 3, 3, 5, 15, -4, -12, 17,
    -- filter=18 channel=2
    7, 13, -6, -1, -12, 14, 11, -13, -12,
    -- filter=18 channel=3
    6, -23, -10, -18, -16, -14, 3, -24, -26,
    -- filter=18 channel=4
    8, -19, -12, -17, 5, -8, -10, -21, -25,
    -- filter=18 channel=5
    -11, 13, -17, -14, -18, 7, -10, 8, -6,
    -- filter=18 channel=6
    5, -10, 6, 12, -10, -10, -5, 11, -16,
    -- filter=18 channel=7
    14, 23, 13, 19, -4, -3, 4, -8, 14,
    -- filter=18 channel=8
    -23, -8, -18, -27, -3, -21, -12, -5, -30,
    -- filter=18 channel=9
    8, 0, -13, 24, 13, -3, -6, -7, 19,
    -- filter=18 channel=10
    0, -18, 1, -4, 8, -24, -2, 10, 4,
    -- filter=18 channel=11
    -1, -3, 12, 16, -6, 20, -9, -19, -11,
    -- filter=18 channel=12
    22, 18, -8, -3, -14, 10, 3, 17, -2,
    -- filter=18 channel=13
    7, -23, -8, -8, -13, -19, -13, -24, -25,
    -- filter=18 channel=14
    20, -2, -1, 20, 11, 20, -4, 7, -11,
    -- filter=18 channel=15
    26, 9, 19, 6, -1, 23, 20, 21, 15,
    -- filter=19 channel=0
    -10, -12, -1, 0, -8, 11, 20, 13, 10,
    -- filter=19 channel=1
    -4, 0, 0, 16, 17, 3, 6, 19, -12,
    -- filter=19 channel=2
    7, 9, 1, -10, 2, -18, 16, -7, 11,
    -- filter=19 channel=3
    -20, -15, -16, 20, 0, -20, -1, 5, 6,
    -- filter=19 channel=4
    0, 14, -8, -14, -11, -4, -9, 18, -19,
    -- filter=19 channel=5
    17, 6, -19, 4, 12, -18, 13, -7, -9,
    -- filter=19 channel=6
    8, -18, 18, 20, -11, -5, 0, -4, -20,
    -- filter=19 channel=7
    15, 15, 16, -3, -13, -21, -2, 8, -5,
    -- filter=19 channel=8
    0, -21, -2, 10, -15, 19, -10, 13, -2,
    -- filter=19 channel=9
    19, -19, 0, 2, 0, -6, 5, 19, -14,
    -- filter=19 channel=10
    11, -18, 3, 16, 20, 7, -6, -8, -18,
    -- filter=19 channel=11
    -16, -15, 3, -10, -8, -16, 4, -17, -4,
    -- filter=19 channel=12
    17, -11, -12, -12, 8, -19, -21, -20, -3,
    -- filter=19 channel=13
    -1, -5, -16, -13, -5, -14, 6, 21, -21,
    -- filter=19 channel=14
    2, 2, -6, 20, 20, 13, 13, -2, 14,
    -- filter=19 channel=15
    -12, 0, -9, -18, -11, 5, 12, -2, -6,
    -- filter=20 channel=0
    28, 31, 21, 30, 33, 33, -11, 24, 11,
    -- filter=20 channel=1
    20, -3, 9, -1, -3, -17, -1, 5, 3,
    -- filter=20 channel=2
    5, 1, -2, -32, -32, -2, -26, 0, -27,
    -- filter=20 channel=3
    37, 36, 32, 17, 20, -2, -8, -7, -3,
    -- filter=20 channel=4
    -25, -47, -25, -12, -33, -13, -13, -37, -8,
    -- filter=20 channel=5
    8, 2, -6, 12, 6, 18, 2, 10, 27,
    -- filter=20 channel=6
    -12, -23, 8, -30, -14, 13, 6, -20, -14,
    -- filter=20 channel=7
    -5, 17, -4, 18, 21, 22, 25, 32, 22,
    -- filter=20 channel=8
    -12, -2, -46, -31, -22, -10, -24, -25, -10,
    -- filter=20 channel=9
    19, 13, 20, -13, -5, 18, 5, 27, -10,
    -- filter=20 channel=10
    -3, -30, -18, -27, -10, -16, -16, 4, -28,
    -- filter=20 channel=11
    -15, -1, 14, -6, -5, -1, -5, 19, -16,
    -- filter=20 channel=12
    38, 1, 37, 24, 23, 24, 22, 22, 22,
    -- filter=20 channel=13
    -3, 16, -10, -10, -6, 19, -2, 5, -9,
    -- filter=20 channel=14
    4, 7, -8, -12, 3, 18, -9, 20, 18,
    -- filter=20 channel=15
    9, -10, -4, -34, -25, 18, -8, -2, -1,
    -- filter=21 channel=0
    17, 9, 5, 19, 30, 4, 31, -3, 26,
    -- filter=21 channel=1
    -6, 3, -18, -15, -9, 8, -16, 0, 12,
    -- filter=21 channel=2
    20, -5, 16, -20, 6, 7, 0, 19, -6,
    -- filter=21 channel=3
    0, 1, -13, 37, 15, -3, 27, 28, 20,
    -- filter=21 channel=4
    -20, -11, 4, 17, 3, -11, 20, -12, 21,
    -- filter=21 channel=5
    -13, -27, 8, 0, -22, 14, -7, -8, 14,
    -- filter=21 channel=6
    -11, -2, 15, -16, -17, -7, -4, 3, 10,
    -- filter=21 channel=7
    -12, -18, -21, 7, -28, 5, -30, -31, -11,
    -- filter=21 channel=8
    -2, -15, 10, 19, -2, -8, -12, 5, -19,
    -- filter=21 channel=9
    3, -19, -28, -30, -31, -32, -33, -6, -29,
    -- filter=21 channel=10
    8, -20, -22, 0, -12, -6, 1, -13, 6,
    -- filter=21 channel=11
    -2, -17, 19, 2, 11, 8, -7, 5, 5,
    -- filter=21 channel=12
    6, -19, -23, 10, 1, -13, 31, -12, -13,
    -- filter=21 channel=13
    13, 31, 10, 7, 43, 36, 50, 21, 36,
    -- filter=21 channel=14
    -8, 13, 19, 5, -11, 9, -17, 6, -13,
    -- filter=21 channel=15
    8, 14, 10, 0, 23, 36, 21, 32, 36,
    -- filter=22 channel=0
    24, 28, 7, 28, 4, -16, 18, -9, -32,
    -- filter=22 channel=1
    2, 2, -20, -1, 4, -14, 10, -19, 21,
    -- filter=22 channel=2
    8, -3, 2, 23, 17, 18, 28, 24, 7,
    -- filter=22 channel=3
    44, 44, 12, -3, -14, -30, -22, -44, -54,
    -- filter=22 channel=4
    51, 25, 47, 23, 51, 38, 42, 48, 42,
    -- filter=22 channel=5
    24, -8, 0, 20, 8, 21, 2, -7, 16,
    -- filter=22 channel=6
    9, 12, 16, 40, 25, 51, 38, 43, 24,
    -- filter=22 channel=7
    -18, 4, -5, -30, -30, -26, -12, -11, -9,
    -- filter=22 channel=8
    5, -18, -16, -10, -13, -8, -2, 9, 1,
    -- filter=22 channel=9
    -8, -8, 22, 27, 3, 19, 4, 21, 18,
    -- filter=22 channel=10
    12, 20, 8, 21, 17, 27, 5, 7, 14,
    -- filter=22 channel=11
    19, 8, -9, 18, -8, -5, -9, -17, -8,
    -- filter=22 channel=12
    45, 23, 5, 30, 11, 24, -4, -16, -13,
    -- filter=22 channel=13
    7, 43, 38, 23, -2, -11, -6, -29, -36,
    -- filter=22 channel=14
    -9, 2, 0, 6, -15, -5, -19, 17, 19,
    -- filter=22 channel=15
    -4, -2, -9, -15, -20, -27, 5, -15, -31,
    -- filter=23 channel=0
    11, 13, -20, -4, 2, 0, -14, 18, 0,
    -- filter=23 channel=1
    -2, -18, 10, -6, 8, 5, -16, 2, -8,
    -- filter=23 channel=2
    16, -3, -5, -15, 23, -14, 15, 3, 3,
    -- filter=23 channel=3
    9, 0, 15, 1, -19, -13, 0, -11, -17,
    -- filter=23 channel=4
    22, 9, 24, 28, 19, 30, 27, 16, -8,
    -- filter=23 channel=5
    19, 11, -7, -11, 23, 21, -4, -16, 6,
    -- filter=23 channel=6
    -4, -3, 11, 12, 18, -4, 22, -3, 25,
    -- filter=23 channel=7
    8, 9, -14, -18, 18, -13, -20, 12, 19,
    -- filter=23 channel=8
    -6, 14, -21, -23, 4, -10, -24, 17, -18,
    -- filter=23 channel=9
    -13, 6, 5, -4, 6, 16, -5, -12, 0,
    -- filter=23 channel=10
    16, -15, 19, 11, 16, 24, -6, -22, 6,
    -- filter=23 channel=11
    -8, 16, 2, 0, -9, -3, 18, 19, 13,
    -- filter=23 channel=12
    12, 6, -7, -7, -2, 17, 2, -21, -13,
    -- filter=23 channel=13
    15, 22, 23, -7, 15, 9, 17, -16, -9,
    -- filter=23 channel=14
    -5, -20, -20, 12, -20, -2, 16, -15, 17,
    -- filter=23 channel=15
    12, 16, 7, 0, -6, 0, 29, -6, 9,
    -- filter=24 channel=0
    11, 3, 0, 16, -15, 25, -8, 7, -6,
    -- filter=24 channel=1
    15, 14, 15, 11, 3, -6, 12, -15, 8,
    -- filter=24 channel=2
    -12, 0, -7, -5, -30, 0, -5, 11, -10,
    -- filter=24 channel=3
    0, 14, 3, 10, -7, 12, -11, 11, 15,
    -- filter=24 channel=4
    -26, -12, -36, -3, -19, -2, -30, -20, -15,
    -- filter=24 channel=5
    18, -17, 12, 8, 18, 22, 1, 18, -14,
    -- filter=24 channel=6
    5, 5, -19, -3, -7, 4, -14, -23, 0,
    -- filter=24 channel=7
    31, 35, 13, 33, 11, 11, 30, 14, 14,
    -- filter=24 channel=8
    -22, -22, 1, -14, -28, 5, 0, -31, 0,
    -- filter=24 channel=9
    12, 8, 21, 25, 24, 26, 26, 0, 18,
    -- filter=24 channel=10
    1, -12, -3, -15, -7, -15, -24, 3, -18,
    -- filter=24 channel=11
    15, -14, 13, 15, -17, 13, 16, 11, 13,
    -- filter=24 channel=12
    16, -6, 30, -10, 19, 0, -1, 7, -4,
    -- filter=24 channel=13
    -20, -29, -8, 5, 5, -12, -8, -13, -8,
    -- filter=24 channel=14
    10, 0, -21, -19, 19, 18, -13, 13, -1,
    -- filter=24 channel=15
    -8, 11, 12, -6, -2, 11, -19, -9, 18,
    -- filter=25 channel=0
    -8, -5, -5, 5, 0, -11, 9, -6, 16,
    -- filter=25 channel=1
    -10, -11, 1, -6, 6, 5, -6, -4, 6,
    -- filter=25 channel=2
    -10, 1, 24, 12, 26, -6, 23, 25, -6,
    -- filter=25 channel=3
    -8, 3, 0, -8, 5, 6, -1, -10, -10,
    -- filter=25 channel=4
    27, 33, 23, 1, 9, 9, 1, -4, 14,
    -- filter=25 channel=5
    33, 22, 5, 0, 26, 14, 20, 0, 18,
    -- filter=25 channel=6
    20, 33, 24, 3, 30, 32, 33, 26, 1,
    -- filter=25 channel=7
    -31, -25, -31, -10, -15, -13, -9, -1, 1,
    -- filter=25 channel=8
    -11, -19, -21, -17, -19, -14, 8, 10, 1,
    -- filter=25 channel=9
    -6, 0, 3, 12, -3, -13, -28, -28, 9,
    -- filter=25 channel=10
    21, -11, 10, 15, -1, -12, -14, -5, -25,
    -- filter=25 channel=11
    15, -16, -3, -8, 14, 0, 2, -13, 8,
    -- filter=25 channel=12
    -14, -11, 10, -27, -24, 3, 14, -15, -19,
    -- filter=25 channel=13
    13, 32, 0, 27, 11, 25, -3, 25, -2,
    -- filter=25 channel=14
    -6, -10, -2, 3, 2, -1, 0, 10, 10,
    -- filter=25 channel=15
    48, 30, 12, 58, 44, 23, 60, 40, 49,
    -- filter=26 channel=0
    8, -20, -21, 12, 13, 0, 7, -1, -22,
    -- filter=26 channel=1
    2, 7, -19, -9, -11, -4, 7, -13, 1,
    -- filter=26 channel=2
    -3, -15, -19, 9, -17, 13, 11, -5, 15,
    -- filter=26 channel=3
    7, -12, 8, 27, 29, -10, 27, -8, -25,
    -- filter=26 channel=4
    11, 12, 0, 1, 0, -9, 17, -16, -12,
    -- filter=26 channel=5
    -6, -16, 6, -17, -4, -24, -20, 7, -6,
    -- filter=26 channel=6
    -5, 0, -28, -24, -12, -22, -15, 10, -29,
    -- filter=26 channel=7
    -3, 0, 24, -6, -9, -14, 10, -22, -3,
    -- filter=26 channel=8
    36, 30, 30, 44, 37, 51, 41, 49, 31,
    -- filter=26 channel=9
    -25, -19, 20, -6, -4, -10, 16, -13, -7,
    -- filter=26 channel=10
    0, 19, 20, 18, -3, 27, -7, -12, 11,
    -- filter=26 channel=11
    1, 19, 11, 20, 20, -14, 16, 17, -15,
    -- filter=26 channel=12
    -11, -12, -3, 29, -1, -24, 27, -1, -27,
    -- filter=26 channel=13
    0, 24, 12, 2, 25, 17, 16, 21, 13,
    -- filter=26 channel=14
    13, 14, -18, 12, -18, -3, -3, 16, -5,
    -- filter=26 channel=15
    -28, -30, 5, -3, -13, -23, -26, -10, -5,
    -- filter=27 channel=0
    -14, 21, -21, 7, -15, 0, 9, 6, 16,
    -- filter=27 channel=1
    12, -19, -7, -19, -14, -12, -4, 12, 13,
    -- filter=27 channel=2
    8, 3, -5, 12, -12, 8, -16, -12, 4,
    -- filter=27 channel=3
    -14, -4, -19, -5, 18, -14, -15, 18, 7,
    -- filter=27 channel=4
    -20, 12, -9, 12, -21, -8, 17, 9, 14,
    -- filter=27 channel=5
    6, 13, -8, 11, 16, -14, 3, 14, -18,
    -- filter=27 channel=6
    19, 0, 19, 17, -11, -7, -9, 17, -5,
    -- filter=27 channel=7
    2, -10, -7, 6, -20, -13, -10, 8, -5,
    -- filter=27 channel=8
    -19, 3, -19, 13, 11, -10, -5, -21, -3,
    -- filter=27 channel=9
    -21, -12, -3, 15, -3, 6, -11, -4, 3,
    -- filter=27 channel=10
    1, 0, -15, 1, 12, -10, -12, 17, 17,
    -- filter=27 channel=11
    11, -15, -4, 5, 14, 9, -17, 14, -8,
    -- filter=27 channel=12
    -18, -11, -18, 17, 4, 2, -9, 19, 17,
    -- filter=27 channel=13
    0, -20, -1, -18, -19, 1, -21, -2, -17,
    -- filter=27 channel=14
    0, -12, 6, 13, 11, -20, 15, 19, 17,
    -- filter=27 channel=15
    -21, -11, -14, 5, -6, -20, 16, 0, -9,
    -- filter=28 channel=0
    4, -11, 5, 4, 19, -7, -16, 2, 11,
    -- filter=28 channel=1
    -20, -11, -21, 4, -16, -7, 18, -6, 17,
    -- filter=28 channel=2
    -8, -16, -7, 12, 4, 11, 3, -15, -23,
    -- filter=28 channel=3
    8, -7, -6, 20, 6, 16, 7, 19, -12,
    -- filter=28 channel=4
    9, 10, -22, -22, -2, 10, 12, 7, 7,
    -- filter=28 channel=5
    0, 6, -4, -21, 6, 12, -14, 14, 15,
    -- filter=28 channel=6
    3, 3, -5, -6, -17, -1, 13, 17, 5,
    -- filter=28 channel=7
    20, 0, 19, 16, 20, 27, 11, -9, 8,
    -- filter=28 channel=8
    -13, 11, -21, 3, 4, -13, 3, -26, 7,
    -- filter=28 channel=9
    12, 0, 16, -15, -17, 0, -12, -2, -16,
    -- filter=28 channel=10
    0, -22, 3, 7, -19, 11, -14, -12, 2,
    -- filter=28 channel=11
    -6, -11, -10, 20, -15, 3, 8, 9, -1,
    -- filter=28 channel=12
    20, -9, 10, 9, -6, -7, 21, -7, 4,
    -- filter=28 channel=13
    -11, 16, -14, 16, -18, -20, -17, 17, 1,
    -- filter=28 channel=14
    -8, -9, 3, -16, 5, -21, -15, -14, -2,
    -- filter=28 channel=15
    14, 9, 0, -16, 12, -11, -14, -18, 15,
    -- filter=29 channel=0
    16, 17, -17, 4, 11, -22, 10, 18, -10,
    -- filter=29 channel=1
    -4, -5, 7, 5, -14, -16, -4, 13, -7,
    -- filter=29 channel=2
    7, 17, 5, 13, 14, 0, -25, -24, -19,
    -- filter=29 channel=3
    24, 12, -19, 18, -8, -27, 11, 13, -12,
    -- filter=29 channel=4
    6, -16, -11, -3, -11, -20, 0, 1, 12,
    -- filter=29 channel=5
    -6, -14, 12, 4, 0, 5, 18, 15, 18,
    -- filter=29 channel=6
    1, -19, 17, 9, 8, -2, -17, -22, -17,
    -- filter=29 channel=7
    37, 34, 25, 17, 36, 21, 37, 35, 35,
    -- filter=29 channel=8
    3, 19, 24, -1, 29, -4, -4, 16, 0,
    -- filter=29 channel=9
    17, 0, -2, 21, 26, 10, -5, 15, 16,
    -- filter=29 channel=10
    21, -6, 1, -8, 5, 9, -15, 23, 20,
    -- filter=29 channel=11
    -1, 7, -14, 0, 0, 6, 13, 16, 5,
    -- filter=29 channel=12
    -12, 12, 2, -3, 3, 7, 2, 7, 5,
    -- filter=29 channel=13
    -12, -33, 2, -24, 2, -29, -2, -30, -10,
    -- filter=29 channel=14
    2, -13, 13, -16, -17, -18, 3, 6, -9,
    -- filter=29 channel=15
    -11, -11, -33, -13, -30, -3, -14, -10, 6,
    -- filter=30 channel=0
    -20, 16, -19, 17, 12, -10, -12, 7, -5,
    -- filter=30 channel=1
    -2, -21, -9, 6, 9, 3, -15, -13, 16,
    -- filter=30 channel=2
    -13, 7, -1, -14, 10, 0, 18, -16, 4,
    -- filter=30 channel=3
    -2, 0, 5, -13, -13, 13, 17, -1, -8,
    -- filter=30 channel=4
    -20, -9, -20, -5, 17, -12, -9, 15, 19,
    -- filter=30 channel=5
    -20, -10, 17, 17, 1, -7, -3, 14, -1,
    -- filter=30 channel=6
    8, -1, -5, 11, -4, 19, -7, 3, 5,
    -- filter=30 channel=7
    3, -12, 12, 14, -5, -11, 13, -7, 15,
    -- filter=30 channel=8
    -1, 4, 5, 19, 2, -18, -3, 13, -8,
    -- filter=30 channel=9
    14, 4, 2, -15, -16, 16, 4, 5, 2,
    -- filter=30 channel=10
    -16, -4, 10, 8, -15, 18, -19, -10, -20,
    -- filter=30 channel=11
    13, 13, -20, -10, 14, 12, 13, 5, -9,
    -- filter=30 channel=12
    -11, -2, -9, 6, -19, 2, -13, 9, -20,
    -- filter=30 channel=13
    6, 0, 20, -5, -3, 10, 3, -4, -8,
    -- filter=30 channel=14
    14, -8, -11, 3, 12, -20, 1, -12, 18,
    -- filter=30 channel=15
    -10, 13, 0, 2, -12, 6, 8, -2, -16,
    -- filter=31 channel=0
    3, -18, 16, -5, 10, -17, 0, -6, -3,
    -- filter=31 channel=1
    -1, -9, -11, 2, 16, -14, 20, -18, -17,
    -- filter=31 channel=2
    -18, -8, 1, -2, 10, 11, 19, 1, 5,
    -- filter=31 channel=3
    5, 24, -8, 25, 22, -6, 19, 21, 21,
    -- filter=31 channel=4
    9, 7, 12, -20, 8, 15, -22, -16, -12,
    -- filter=31 channel=5
    -25, -26, -24, -25, 8, 2, -12, 13, -11,
    -- filter=31 channel=6
    2, -9, -8, -21, -19, -3, 2, 14, -6,
    -- filter=31 channel=7
    -27, 5, -17, -17, -20, -16, -15, 0, 1,
    -- filter=31 channel=8
    10, 14, -6, 23, 23, 1, 12, 9, 24,
    -- filter=31 channel=9
    -18, 5, -27, -32, -22, -18, -10, -22, 9,
    -- filter=31 channel=10
    -15, 3, -9, 10, 18, -15, -1, -20, 3,
    -- filter=31 channel=11
    9, -1, 14, -20, 5, -18, 4, 12, -7,
    -- filter=31 channel=12
    -8, 9, 7, 12, -2, 8, -10, 0, 3,
    -- filter=31 channel=13
    30, -6, 25, 13, 0, 31, 17, 0, 21,
    -- filter=31 channel=14
    -7, -16, 14, 6, -4, 6, -13, 0, -11,
    -- filter=31 channel=15
    -6, -5, 1, 0, -21, -16, -32, 2, 5,

    others => 0);
end iwght_package;
