library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    16, 16, 10, 9, 6, 8, 12, 13, 5, 11, 20, 15, 7, 2, 1, 
    0, 3, 9, 11, 10, 0, 3, 5, 41, 0, 0, 0, 0, 5, 0, 
    15, 31, 8, 10, 12, 76, 44, 19, 0, 0, 33, 18, 0, 0, 0, 
    0, 0, 1, 3, 0, 3, 0, 8, 1, 41, 45, 36, 28, 0, 0, 
    39, 0, 17, 14, 0, 10, 51, 19, 13, 0, 17, 11, 0, 0, 0, 
    105, 43, 39, 58, 127, 124, 37, 20, 0, 0, 83, 60, 14, 3, 0, 
    94, 42, 46, 19, 30, 26, 79, 44, 23, 0, 86, 19, 1, 0, 2, 
    88, 59, 7, 0, 11, 59, 128, 80, 44, 30, 77, 35, 15, 37, 32, 
    95, 79, 65, 14, 19, 105, 50, 0, 1, 18, 53, 72, 21, 3, 0, 
    113, 94, 64, 12, 46, 36, 27, 0, 23, 75, 53, 0, 0, 0, 15, 
    53, 84, 80, 0, 0, 0, 34, 114, 60, 0, 0, 0, 0, 0, 1, 
    86, 103, 76, 33, 196, 135, 71, 72, 39, 17, 12, 21, 20, 23, 30, 
    16, 68, 81, 109, 163, 21, 22, 19, 15, 7, 6, 7, 31, 42, 14, 
    35, 10, 77, 144, 57, 21, 15, 16, 22, 20, 31, 44, 36, 11, 74, 
    41, 24, 28, 80, 36, 38, 49, 28, 12, 11, 27, 26, 3, 27, 31, 
    
    -- channel=1
    122, 124, 128, 128, 128, 124, 129, 139, 135, 113, 97, 100, 105, 113, 112, 
    129, 131, 135, 130, 131, 123, 114, 116, 78, 60, 37, 45, 70, 93, 107, 
    96, 103, 130, 133, 135, 113, 62, 53, 49, 47, 23, 25, 23, 62, 89, 
    20, 92, 114, 136, 114, 89, 53, 37, 27, 59, 20, 35, 14, 31, 85, 
    0, 61, 89, 135, 67, 61, 26, 25, 22, 62, 36, 24, 34, 20, 66, 
    4, 34, 77, 95, 54, 40, 24, 32, 13, 92, 20, 12, 38, 22, 27, 
    9, 3, 68, 80, 85, 67, 32, 23, 11, 70, 1, 17, 30, 31, 32, 
    12, 0, 44, 53, 82, 69, 10, 26, 22, 75, 17, 13, 36, 36, 61, 
    1, 5, 0, 35, 49, 32, 28, 32, 51, 39, 49, 13, 36, 60, 102, 
    13, 13, 0, 25, 16, 51, 48, 15, 44, 40, 10, 20, 52, 98, 104, 
    15, 15, 0, 71, 0, 22, 31, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 2, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 13, 0, 8, 0, 0, 0, 7, 0, 0, 0, 0, 
    22, 23, 0, 0, 37, 11, 15, 0, 0, 0, 16, 0, 0, 0, 0, 
    18, 33, 0, 0, 0, 0, 42, 0, 0, 0, 23, 0, 0, 0, 0, 
    29, 50, 0, 0, 0, 35, 11, 0, 0, 0, 7, 0, 0, 0, 0, 
    50, 60, 7, 5, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    46, 47, 32, 11, 28, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 
    53, 44, 34, 23, 44, 22, 24, 54, 14, 0, 0, 0, 6, 27, 27, 
    65, 54, 40, 50, 98, 48, 37, 41, 32, 24, 27, 30, 37, 37, 41, 
    38, 41, 32, 87, 56, 26, 25, 20, 20, 22, 32, 39, 42, 45, 50, 
    53, 35, 42, 88, 27, 26, 26, 24, 25, 32, 38, 49, 44, 55, 57, 
    48, 42, 30, 60, 19, 25, 30, 23, 26, 35, 38, 32, 45, 66, 46, 
    
    -- channel=3
    17, 26, 21, 21, 16, 25, 15, 10, 10, 11, 17, 21, 24, 10, 6, 
    11, 14, 17, 19, 25, 80, 14, 16, 17, 56, 55, 28, 20, 15, 11, 
    17, 22, 15, 16, 13, 65, 53, 25, 28, 107, 112, 102, 48, 5, 29, 
    43, 29, 12, 17, 27, 51, 77, 61, 65, 94, 121, 70, 72, 15, 18, 
    132, 106, 34, 61, 158, 118, 126, 83, 56, 84, 121, 70, 70, 42, 0, 
    152, 176, 61, 44, 193, 161, 161, 91, 56, 120, 155, 93, 76, 73, 34, 
    163, 163, 54, 28, 89, 151, 172, 135, 81, 143, 149, 83, 71, 88, 64, 
    184, 201, 68, 54, 59, 175, 175, 120, 91, 127, 148, 85, 77, 88, 67, 
    220, 215, 130, 128, 75, 110, 97, 90, 85, 64, 77, 74, 54, 67, 33, 
    232, 216, 159, 143, 103, 78, 125, 144, 79, 90, 64, 26, 38, 41, 30, 
    208, 201, 159, 212, 225, 110, 165, 200, 125, 67, 56, 76, 90, 95, 83, 
    166, 226, 186, 247, 229, 162, 133, 132, 122, 114, 125, 137, 153, 154, 153, 
    148, 151, 215, 249, 187, 137, 127, 124, 123, 128, 144, 154, 157, 164, 186, 
    168, 138, 166, 250, 145, 142, 136, 123, 133, 145, 155, 162, 162, 178, 175, 
    172, 159, 137, 147, 115, 127, 141, 142, 145, 159, 146, 151, 186, 200, 150, 
    
    -- channel=4
    113, 109, 108, 111, 113, 98, 113, 124, 119, 110, 104, 98, 95, 98, 106, 
    109, 104, 108, 115, 108, 60, 97, 103, 117, 58, 29, 42, 70, 92, 98, 
    109, 118, 114, 118, 119, 143, 127, 88, 38, 13, 41, 40, 44, 58, 81, 
    56, 3, 104, 110, 103, 76, 38, 40, 44, 34, 79, 61, 72, 47, 55, 
    48, 0, 101, 57, 0, 3, 61, 54, 62, 12, 35, 47, 36, 40, 38, 
    67, 42, 106, 118, 101, 88, 62, 48, 47, 0, 81, 87, 40, 43, 18, 
    49, 58, 98, 123, 55, 37, 73, 64, 62, 0, 92, 54, 39, 27, 41, 
    43, 47, 28, 73, 37, 25, 120, 92, 77, 36, 93, 71, 35, 56, 82, 
    52, 34, 70, 32, 59, 102, 81, 48, 26, 85, 76, 112, 56, 53, 64, 
    82, 49, 76, 4, 45, 51, 36, 19, 36, 96, 101, 43, 2, 54, 109, 
    37, 48, 88, 0, 3, 0, 0, 75, 63, 43, 0, 0, 0, 28, 40, 
    30, 55, 40, 0, 157, 116, 56, 55, 31, 12, 2, 2, 0, 0, 4, 
    0, 22, 24, 78, 136, 4, 4, 7, 8, 0, 0, 0, 0, 5, 0, 
    4, 0, 0, 139, 50, 0, 3, 0, 0, 0, 2, 9, 7, 0, 28, 
    5, 0, 5, 67, 35, 20, 25, 9, 0, 0, 0, 0, 0, 0, 10, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 5, 13, 0, 
    18, 50, 0, 0, 0, 62, 5, 10, 0, 0, 0, 0, 0, 10, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 28, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 12, 22, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 34, 38, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 42, 15, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 46, 7, 0, 0, 0, 0, 7, 4, 
    72, 29, 0, 0, 46, 49, 28, 25, 7, 0, 0, 0, 0, 0, 0, 
    0, 38, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 79, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 20, 
    0, 0, 0, 73, 3, 12, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    1, 0, 6, 0, 0, 2, 0, 0, 0, 0, 0, 9, 3, 0, 0, 
    1, 1, 6, 0, 13, 29, 0, 0, 0, 27, 0, 0, 4, 18, 0, 
    0, 57, 3, 0, 9, 7, 0, 0, 11, 81, 0, 0, 0, 10, 31, 
    0, 101, 0, 12, 0, 32, 0, 0, 0, 104, 0, 0, 0, 0, 85, 
    0, 29, 0, 102, 0, 0, 0, 0, 0, 148, 0, 0, 0, 0, 30, 
    0, 8, 0, 30, 104, 0, 0, 0, 0, 257, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 97, 86, 0, 0, 0, 203, 0, 0, 4, 21, 0, 
    0, 0, 0, 0, 67, 95, 0, 0, 0, 128, 0, 0, 33, 0, 0, 
    0, 0, 0, 47, 0, 9, 0, 0, 31, 0, 14, 0, 31, 32, 14, 
    0, 0, 0, 85, 0, 8, 57, 0, 0, 0, 0, 0, 45, 46, 0, 
    94, 0, 0, 220, 0, 0, 75, 0, 0, 0, 0, 20, 13, 10, 0, 
    78, 65, 0, 150, 0, 0, 0, 0, 0, 0, 2, 6, 5, 0, 0, 
    0, 82, 133, 0, 0, 0, 0, 0, 0, 3, 8, 5, 0, 4, 14, 
    0, 0, 172, 0, 0, 4, 0, 0, 6, 4, 0, 0, 0, 35, 0, 
    0, 0, 11, 0, 0, 22, 8, 0, 12, 0, 0, 4, 58, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 27, 40, 24, 0, 0, 
    27, 7, 0, 0, 0, 0, 5, 21, 23, 0, 6, 0, 13, 13, 0, 
    52, 41, 0, 0, 39, 21, 5, 22, 15, 17, 23, 21, 32, 38, 0, 
    26, 16, 0, 0, 0, 0, 10, 22, 42, 36, 1, 7, 20, 38, 46, 
    43, 14, 0, 0, 0, 0, 0, 15, 24, 21, 3, 28, 28, 33, 23, 
    33, 50, 23, 0, 0, 0, 0, 0, 1, 0, 0, 15, 21, 0, 0, 
    42, 42, 34, 14, 0, 0, 0, 18, 22, 0, 0, 0, 2, 0, 0, 
    9, 25, 40, 47, 16, 14, 25, 46, 17, 0, 0, 30, 28, 0, 0, 
    28, 22, 28, 78, 102, 89, 47, 23, 44, 65, 98, 114, 104, 66, 59, 
    62, 39, 45, 31, 0, 32, 59, 65, 91, 108, 121, 124, 135, 129, 131, 
    149, 64, 47, 0, 50, 118, 115, 113, 117, 129, 143, 150, 132, 133, 167, 
    157, 140, 57, 27, 88, 124, 126, 118, 121, 134, 136, 131, 142, 167, 116, 
    154, 149, 110, 72, 96, 101, 103, 120, 130, 142, 133, 137, 162, 166, 151, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 63, 5, 0, 0, 29, 54, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 31, 72, 34, 34, 26, 0, 1, 
    20, 67, 1, 2, 0, 30, 55, 33, 28, 33, 11, 7, 3, 4, 8, 
    62, 104, 3, 61, 125, 87, 16, 14, 0, 71, 59, 31, 34, 25, 0, 
    28, 45, 0, 0, 0, 7, 46, 35, 19, 127, 13, 0, 25, 30, 41, 
    51, 28, 0, 0, 19, 76, 27, 37, 9, 96, 9, 23, 33, 56, 29, 
    61, 52, 48, 27, 62, 60, 0, 0, 1, 44, 15, 3, 29, 9, 0, 
    60, 65, 18, 54, 33, 0, 7, 39, 50, 13, 0, 0, 0, 24, 29, 
    36, 56, 20, 83, 21, 11, 56, 86, 21, 0, 0, 9, 52, 36, 0, 
    68, 57, 7, 155, 151, 119, 81, 4, 7, 29, 69, 96, 72, 48, 44, 
    14, 40, 67, 142, 0, 0, 1, 4, 30, 52, 60, 61, 74, 71, 64, 
    70, 24, 81, 36, 0, 58, 53, 52, 57, 70, 81, 86, 65, 66, 101, 
    65, 68, 51, 0, 36, 64, 66, 57, 59, 67, 64, 55, 64, 98, 29, 
    61, 68, 58, 0, 30, 35, 35, 55, 81, 84, 65, 69, 125, 96, 55, 
    
    -- channel=10
    125, 123, 128, 131, 131, 121, 137, 145, 133, 108, 87, 90, 100, 113, 108, 
    130, 136, 135, 136, 130, 117, 139, 114, 77, 35, 31, 41, 54, 81, 105, 
    86, 86, 134, 138, 139, 118, 73, 47, 20, 18, 29, 16, 24, 41, 76, 
    48, 51, 133, 134, 119, 74, 60, 25, 13, 24, 44, 31, 9, 9, 50, 
    30, 58, 130, 96, 87, 88, 61, 28, 12, 8, 55, 41, 17, 9, 33, 
    34, 41, 126, 99, 28, 56, 60, 47, 26, 7, 65, 28, 16, 12, 11, 
    34, 44, 85, 105, 47, 51, 65, 48, 32, 21, 50, 27, 14, 12, 33, 
    41, 36, 55, 86, 54, 51, 57, 33, 29, 46, 40, 30, 6, 33, 59, 
    38, 33, 32, 19, 67, 38, 43, 32, 26, 83, 33, 17, 8, 38, 97, 
    36, 37, 30, 11, 40, 31, 28, 46, 49, 25, 10, 0, 9, 91, 114, 
    9, 46, 37, 12, 48, 37, 11, 14, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 63, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 27, 10, 0, 
    20, 47, 0, 0, 0, 86, 2, 22, 0, 0, 0, 0, 0, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 20, 0, 0, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 26, 107, 13, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 6, 33, 0, 58, 0, 3, 0, 0, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 18, 40, 0, 33, 0, 0, 8, 23, 0, 
    0, 0, 0, 0, 0, 92, 3, 0, 0, 19, 49, 36, 35, 0, 0, 
    0, 1, 0, 5, 0, 0, 0, 0, 6, 33, 31, 6, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 21, 3, 
    136, 37, 0, 0, 88, 74, 77, 65, 14, 1, 0, 6, 0, 0, 0, 
    0, 108, 8, 28, 31, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 
    0, 7, 112, 46, 0, 0, 0, 0, 0, 0, 8, 22, 3, 0, 63, 
    0, 1, 31, 90, 28, 36, 29, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    3, 0, 0, 3, 5, 0, 5, 2, 5, 11, 9, 0, 0, 10, 11, 
    0, 0, 0, 7, 0, 0, 46, 20, 25, 0, 10, 21, 0, 0, 6, 
    46, 0, 3, 3, 1, 0, 52, 5, 0, 0, 28, 0, 48, 0, 0, 
    92, 0, 11, 0, 31, 0, 9, 36, 14, 0, 57, 18, 33, 44, 0, 
    62, 0, 65, 0, 0, 38, 56, 58, 36, 0, 0, 77, 0, 39, 0, 
    91, 0, 80, 80, 0, 18, 42, 27, 70, 0, 92, 74, 0, 17, 30, 
    77, 45, 7, 66, 0, 0, 1, 48, 59, 0, 81, 56, 0, 0, 38, 
    77, 0, 48, 17, 0, 0, 103, 16, 30, 0, 44, 60, 0, 3, 4, 
    65, 0, 152, 0, 81, 0, 11, 15, 0, 43, 0, 68, 0, 0, 0, 
    0, 0, 117, 0, 56, 34, 0, 3, 55, 22, 56, 0, 0, 0, 17, 
    0, 2, 97, 0, 95, 51, 0, 15, 76, 36, 0, 0, 0, 0, 12, 
    0, 0, 3, 0, 163, 63, 0, 0, 6, 0, 0, 0, 0, 0, 5, 
    31, 0, 0, 48, 117, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 62, 31, 0, 13, 2, 0, 0, 0, 0, 0, 0, 40, 
    43, 0, 12, 0, 17, 0, 0, 0, 0, 0, 15, 0, 0, 18, 49, 
    
    -- channel=13
    101, 112, 111, 111, 107, 107, 116, 121, 107, 81, 70, 79, 93, 100, 95, 
    110, 119, 115, 113, 108, 123, 106, 94, 58, 42, 36, 40, 50, 71, 90, 
    68, 70, 111, 117, 110, 84, 65, 37, 30, 38, 37, 37, 32, 32, 80, 
    45, 56, 104, 110, 99, 62, 62, 32, 25, 25, 56, 34, 28, 24, 55, 
    35, 62, 100, 74, 102, 79, 65, 46, 27, 29, 58, 46, 35, 31, 31, 
    15, 51, 106, 72, 51, 65, 83, 54, 43, 33, 54, 35, 28, 28, 34, 
    28, 48, 70, 97, 53, 64, 57, 53, 43, 32, 45, 36, 26, 28, 43, 
    39, 53, 38, 74, 38, 49, 49, 38, 44, 52, 49, 36, 21, 39, 72, 
    40, 39, 28, 43, 47, 33, 48, 41, 35, 58, 28, 28, 25, 62, 94, 
    42, 37, 40, 26, 38, 35, 42, 58, 37, 31, 20, 8, 34, 83, 87, 
    21, 40, 38, 40, 72, 32, 15, 20, 15, 9, 0, 0, 0, 0, 0, 
    0, 4, 36, 55, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 9, 1, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 24, 3, 0, 0, 49, 37, 34, 3, 0, 0, 
    0, 3, 0, 0, 0, 6, 11, 10, 20, 59, 35, 26, 21, 0, 12, 
    33, 35, 0, 21, 34, 24, 32, 14, 14, 50, 37, 6, 20, 0, 0, 
    55, 75, 0, 5, 107, 68, 47, 21, 0, 75, 50, 24, 31, 19, 0, 
    56, 61, 14, 0, 49, 63, 71, 41, 14, 90, 49, 17, 25, 35, 11, 
    66, 77, 10, 0, 27, 88, 62, 56, 26, 71, 57, 20, 35, 36, 16, 
    83, 99, 30, 57, 13, 60, 33, 25, 34, 16, 34, 21, 24, 22, 0, 
    105, 101, 45, 74, 28, 23, 54, 45, 19, 38, 20, 7, 14, 9, 0, 
    111, 88, 51, 112, 60, 22, 81, 95, 39, 17, 16, 28, 34, 43, 29, 
    116, 122, 76, 130, 103, 80, 75, 74, 60, 60, 67, 74, 82, 83, 80, 
    77, 102, 118, 113, 76, 68, 65, 65, 64, 69, 78, 80, 85, 92, 96, 
    88, 75, 115, 117, 70, 75, 66, 63, 71, 77, 85, 93, 90, 97, 101, 
    86, 86, 79, 90, 63, 77, 83, 75, 76, 80, 76, 84, 102, 98, 73, 
    
    -- channel=15
    56, 56, 58, 57, 56, 53, 66, 73, 59, 38, 32, 39, 43, 49, 44, 
    58, 67, 61, 60, 56, 23, 49, 45, 30, 0, 0, 0, 8, 33, 40, 
    17, 50, 65, 66, 64, 35, 16, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 59, 63, 36, 19, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 39, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    130, 128, 128, 128, 129, 130, 130, 129, 130, 128, 129, 128, 128, 128, 128, 
    133, 130, 130, 130, 130, 130, 130, 129, 128, 147, 139, 126, 130, 129, 129, 
    138, 135, 131, 130, 129, 131, 134, 139, 161, 131, 116, 136, 131, 131, 131, 
    115, 122, 127, 131, 133, 134, 129, 124, 77, 56, 31, 63, 127, 127, 129, 
    180, 180, 129, 138, 135, 120, 95, 120, 110, 128, 161, 181, 186, 167, 129, 
    13, 11, 84, 156, 150, 209, 212, 203, 181, 124, 62, 28, 17, 26, 125, 
    177, 187, 152, 94, 82, 76, 15, 0, 27, 138, 180, 198, 184, 176, 171, 
    42, 0, 76, 97, 110, 18, 0, 96, 154, 124, 68, 24, 12, 9, 42, 
    0, 60, 15, 44, 105, 142, 152, 138, 78, 111, 110, 124, 144, 158, 134, 
    78, 178, 171, 172, 163, 143, 118, 91, 91, 84, 86, 80, 47, 52, 59, 
    61, 59, 84, 109, 128, 147, 149, 144, 125, 110, 83, 58, 34, 17, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 59, 27, 
    0, 0, 7, 0, 0, 0, 47, 145, 110, 109, 122, 91, 14, 20, 34, 
    0, 0, 0, 0, 0, 0, 0, 59, 98, 35, 0, 0, 30, 38, 62, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 30, 40, 60, 
    
    -- channel=17
    13, 14, 14, 14, 14, 14, 14, 14, 16, 14, 11, 13, 14, 14, 14, 
    12, 13, 13, 13, 13, 13, 14, 14, 12, 0, 5, 14, 13, 13, 13, 
    13, 14, 14, 13, 14, 13, 13, 1, 0, 0, 14, 15, 12, 14, 13, 
    7, 7, 12, 15, 14, 0, 20, 0, 0, 0, 0, 27, 7, 10, 12, 
    0, 0, 14, 14, 14, 3, 23, 8, 12, 1, 0, 0, 0, 14, 9, 
    10, 17, 15, 12, 12, 0, 1, 3, 3, 0, 0, 5, 0, 33, 10, 
    0, 0, 0, 14, 0, 0, 0, 4, 33, 8, 1, 0, 3, 0, 8, 
    6, 19, 5, 27, 1, 5, 29, 0, 0, 0, 0, 0, 4, 6, 18, 
    80, 4, 19, 23, 12, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    12, 44, 11, 15, 19, 23, 8, 0, 0, 0, 1, 20, 15, 16, 32, 
    20, 31, 26, 20, 24, 26, 77, 35, 54, 52, 35, 28, 40, 36, 35, 
    0, 30, 32, 26, 29, 30, 82, 90, 82, 56, 60, 54, 34, 34, 29, 
    4, 36, 35, 31, 32, 31, 54, 50, 61, 69, 48, 34, 35, 33, 27, 
    
    -- channel=18
    84, 84, 84, 84, 84, 84, 84, 83, 82, 84, 86, 84, 84, 84, 84, 
    86, 85, 85, 85, 85, 85, 85, 84, 86, 86, 79, 86, 85, 85, 85, 
    83, 84, 85, 85, 85, 87, 85, 87, 85, 77, 62, 75, 86, 85, 86, 
    91, 89, 86, 85, 86, 86, 77, 82, 67, 67, 59, 74, 91, 88, 87, 
    70, 73, 82, 82, 87, 87, 75, 87, 81, 89, 84, 74, 73, 76, 88, 
    44, 43, 71, 73, 77, 79, 71, 74, 79, 88, 72, 59, 50, 54, 89, 
    56, 61, 78, 59, 76, 26, 18, 31, 63, 85, 80, 70, 69, 62, 74, 
    0, 13, 13, 43, 74, 52, 42, 57, 63, 65, 51, 41, 36, 49, 51, 
    0, 70, 47, 57, 77, 87, 91, 78, 53, 61, 63, 61, 55, 55, 57, 
    26, 71, 78, 87, 84, 88, 82, 68, 69, 51, 51, 41, 31, 24, 27, 
    0, 0, 0, 0, 0, 9, 32, 35, 31, 26, 19, 13, 12, 15, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 39, 
    
    -- channel=19
    285, 284, 284, 284, 284, 285, 285, 284, 283, 284, 287, 284, 284, 284, 285, 
    286, 285, 285, 285, 284, 284, 285, 284, 279, 260, 269, 281, 285, 285, 286, 
    285, 285, 287, 286, 286, 285, 285, 271, 254, 239, 225, 283, 286, 286, 288, 
    279, 283, 284, 287, 288, 275, 276, 275, 256, 245, 232, 251, 287, 287, 289, 
    207, 225, 285, 283, 286, 280, 265, 282, 282, 285, 266, 251, 233, 267, 292, 
    227, 238, 251, 241, 270, 225, 248, 261, 283, 290, 255, 237, 217, 230, 286, 
    186, 202, 231, 256, 241, 148, 127, 170, 218, 271, 264, 249, 247, 241, 257, 
    110, 163, 154, 203, 262, 234, 231, 222, 222, 210, 178, 164, 169, 196, 206, 
    127, 240, 220, 231, 266, 273, 272, 255, 235, 222, 243, 222, 215, 214, 211, 
    166, 221, 226, 231, 234, 234, 225, 199, 195, 180, 172, 161, 146, 146, 167, 
    39, 74, 71, 77, 86, 111, 137, 142, 143, 129, 117, 116, 137, 135, 147, 
    0, 17, 48, 2, 0, 0, 103, 72, 74, 81, 101, 117, 125, 144, 149, 
    0, 0, 0, 0, 0, 0, 59, 171, 147, 126, 102, 106, 98, 128, 176, 
    4, 0, 0, 0, 0, 0, 0, 14, 4, 26, 41, 78, 121, 146, 197, 
    23, 0, 0, 0, 0, 0, 0, 0, 10, 55, 102, 117, 132, 163, 207, 
    
    -- channel=20
    61, 60, 60, 60, 60, 61, 61, 61, 62, 62, 59, 61, 61, 60, 60, 
    63, 61, 61, 62, 62, 62, 62, 63, 66, 94, 78, 56, 61, 61, 61, 
    67, 64, 62, 62, 59, 63, 64, 82, 101, 85, 54, 64, 63, 63, 62, 
    50, 57, 61, 63, 61, 83, 63, 72, 25, 12, 0, 3, 63, 63, 63, 
    133, 117, 71, 68, 65, 68, 37, 58, 41, 57, 90, 121, 128, 90, 65, 
    0, 0, 29, 91, 92, 133, 137, 124, 98, 73, 22, 0, 0, 0, 57, 
    127, 119, 88, 42, 52, 75, 16, 0, 0, 63, 101, 124, 112, 113, 94, 
    12, 0, 61, 50, 63, 0, 0, 49, 109, 92, 55, 18, 1, 0, 0, 
    0, 10, 0, 0, 31, 78, 86, 79, 22, 40, 44, 61, 81, 106, 92, 
    14, 98, 88, 84, 77, 67, 54, 38, 37, 38, 39, 44, 17, 23, 28, 
    78, 68, 72, 88, 101, 103, 88, 81, 75, 66, 51, 32, 5, 0, 19, 
    49, 13, 17, 14, 21, 15, 0, 0, 0, 0, 0, 0, 8, 46, 19, 
    29, 33, 54, 55, 33, 25, 0, 38, 11, 38, 86, 88, 28, 25, 23, 
    62, 23, 25, 28, 24, 24, 0, 19, 75, 55, 0, 3, 49, 40, 42, 
    84, 24, 22, 22, 17, 16, 10, 25, 0, 0, 42, 61, 45, 40, 39, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 15, 13, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 70, 9, 0, 0, 0, 0, 0, 0, 0, 15, 51, 66, 46, 0, 
    0, 0, 0, 10, 12, 85, 113, 93, 50, 0, 0, 0, 0, 0, 0, 
    96, 97, 49, 0, 0, 0, 0, 0, 0, 0, 41, 69, 77, 63, 48, 
    29, 0, 0, 0, 0, 0, 0, 0, 30, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 24, 0, 15, 19, 31, 60, 63, 37, 
    44, 90, 82, 78, 60, 44, 25, 0, 7, 0, 20, 20, 0, 0, 0, 
    39, 40, 52, 82, 104, 116, 114, 106, 89, 74, 50, 25, 0, 0, 0, 
    14, 22, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 46, 28, 8, 1, 65, 60, 17, 25, 53, 31, 0, 0, 0, 
    0, 0, 4, 5, 2, 2, 2, 45, 54, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 66, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 57, 0, 0, 0, 
    4, 47, 78, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 93, 5, 
    0, 20, 0, 0, 8, 0, 30, 32, 47, 0, 0, 0, 0, 98, 8, 
    6, 66, 26, 44, 0, 0, 22, 57, 88, 0, 0, 0, 9, 0, 65, 
    101, 60, 0, 98, 0, 0, 27, 0, 0, 0, 0, 0, 7, 5, 24, 
    282, 0, 0, 19, 16, 0, 0, 0, 0, 0, 11, 0, 8, 3, 0, 
    104, 7, 16, 7, 9, 0, 0, 0, 0, 0, 0, 0, 2, 10, 30, 
    0, 39, 0, 8, 25, 43, 24, 20, 5, 0, 0, 15, 32, 3, 32, 
    0, 78, 0, 0, 0, 27, 125, 0, 0, 0, 19, 11, 9, 3, 45, 
    0, 28, 16, 0, 0, 6, 222, 1, 0, 0, 0, 8, 18, 35, 59, 
    0, 0, 7, 0, 0, 2, 103, 20, 0, 10, 28, 38, 8, 41, 53, 
    0, 0, 0, 0, 0, 1, 34, 27, 23, 61, 9, 2, 24, 34, 47, 
    
    -- channel=23
    15, 15, 15, 15, 15, 15, 15, 13, 13, 16, 20, 15, 15, 15, 15, 
    14, 15, 15, 14, 14, 14, 14, 13, 14, 0, 2, 13, 15, 15, 15, 
    9, 10, 14, 14, 14, 14, 15, 7, 1, 32, 17, 11, 14, 13, 15, 
    30, 28, 17, 12, 13, 4, 7, 32, 65, 86, 92, 56, 22, 21, 18, 
    0, 0, 4, 5, 11, 27, 27, 26, 36, 36, 9, 0, 0, 0, 18, 
    114, 104, 36, 0, 0, 0, 0, 0, 0, 39, 80, 97, 98, 64, 22, 
    0, 0, 0, 45, 47, 65, 71, 94, 64, 12, 0, 0, 0, 0, 0, 
    59, 95, 28, 0, 35, 104, 114, 32, 0, 17, 50, 72, 80, 92, 67, 
    122, 75, 93, 70, 40, 16, 7, 38, 75, 51, 59, 42, 18, 4, 18, 
    32, 8, 16, 20, 30, 43, 59, 67, 61, 72, 60, 66, 78, 63, 54, 
    11, 23, 16, 3, 0, 0, 15, 24, 32, 40, 54, 65, 82, 75, 47, 
    32, 41, 59, 61, 48, 48, 129, 152, 133, 130, 123, 102, 35, 33, 41, 
    46, 18, 0, 13, 33, 35, 0, 0, 0, 0, 0, 0, 27, 35, 39, 
    39, 37, 33, 35, 37, 38, 0, 0, 0, 0, 38, 31, 21, 26, 29, 
    30, 44, 45, 46, 46, 50, 24, 0, 38, 29, 8, 15, 24, 32, 35, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    73, 73, 73, 73, 73, 73, 73, 72, 73, 72, 73, 74, 73, 73, 74, 
    71, 73, 73, 72, 72, 72, 72, 73, 69, 26, 47, 73, 73, 73, 74, 
    65, 68, 72, 73, 75, 69, 71, 46, 16, 20, 42, 62, 72, 73, 74, 
    86, 81, 76, 72, 72, 47, 69, 61, 108, 117, 134, 123, 77, 78, 77, 
    0, 0, 58, 65, 69, 70, 97, 79, 94, 69, 24, 0, 0, 31, 76, 
    148, 161, 85, 21, 23, 0, 0, 0, 26, 72, 117, 141, 128, 148, 80, 
    0, 0, 2, 83, 72, 21, 73, 125, 140, 48, 0, 0, 0, 0, 15, 
    44, 132, 24, 48, 64, 149, 183, 60, 0, 14, 48, 85, 106, 125, 110, 
    179, 92, 136, 121, 82, 45, 30, 32, 74, 47, 47, 19, 0, 0, 0, 
    35, 0, 0, 0, 0, 4, 19, 33, 32, 28, 16, 12, 39, 40, 46, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 47, 63, 57, 
    0, 18, 25, 16, 1, 3, 136, 135, 103, 105, 119, 103, 40, 23, 79, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 71, 92, 
    0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 66, 79, 47, 66, 79, 
    0, 27, 25, 20, 21, 25, 18, 0, 61, 84, 48, 41, 61, 75, 88, 
    
    -- channel=26
    68, 67, 67, 67, 67, 67, 67, 68, 68, 66, 62, 67, 67, 67, 67, 
    68, 67, 67, 67, 67, 67, 67, 68, 67, 57, 36, 57, 68, 67, 67, 
    65, 66, 68, 68, 68, 67, 63, 63, 39, 21, 27, 38, 68, 68, 68, 
    54, 61, 67, 69, 68, 69, 51, 60, 35, 35, 36, 55, 62, 64, 66, 
    8, 9, 32, 67, 67, 64, 68, 63, 58, 51, 36, 24, 23, 19, 60, 
    26, 33, 68, 58, 45, 37, 11, 16, 25, 43, 38, 40, 40, 40, 59, 
    0, 0, 10, 20, 49, 12, 0, 11, 38, 55, 41, 29, 16, 27, 18, 
    0, 6, 31, 31, 34, 31, 42, 58, 28, 19, 16, 12, 20, 22, 33, 
    0, 41, 30, 47, 44, 47, 35, 12, 9, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 23, 
    4, 0, 0, 0, 0, 0, 5, 36, 50, 48, 35, 20, 22, 27, 31, 
    10, 0, 0, 0, 0, 0, 10, 77, 65, 22, 22, 34, 32, 29, 33, 
    14, 0, 0, 0, 0, 0, 0, 19, 14, 37, 43, 32, 30, 34, 37, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 44, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 58, 23, 56, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    155, 139, 32, 3, 0, 0, 0, 0, 0, 0, 48, 100, 124, 85, 0, 
    0, 0, 2, 54, 38, 124, 138, 113, 71, 0, 0, 0, 0, 0, 4, 
    164, 171, 82, 0, 0, 0, 7, 0, 0, 21, 69, 101, 84, 103, 91, 
    35, 0, 34, 61, 0, 0, 0, 6, 91, 52, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 49, 0, 0, 14, 4, 35, 79, 110, 72, 
    98, 127, 134, 126, 110, 83, 61, 38, 46, 17, 60, 36, 12, 17, 17, 
    100, 92, 112, 143, 164, 170, 158, 145, 121, 104, 75, 50, 11, 0, 0, 
    0, 26, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 30, 61, 22, 0, 0, 155, 34, 5, 22, 84, 55, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 64, 41, 56, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 54, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 37, 15, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41, 0, 26, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 38, 24, 15, 0, 0, 
    0, 0, 0, 17, 0, 54, 0, 0, 0, 0, 0, 0, 35, 0, 0, 
    11, 0, 0, 0, 35, 127, 0, 0, 0, 7, 28, 34, 0, 14, 0, 
    0, 0, 17, 0, 0, 3, 0, 66, 8, 1, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 28, 0, 17, 0, 34, 10, 2, 0, 
    0, 4, 0, 0, 0, 0, 4, 3, 0, 30, 2, 9, 0, 0, 0, 
    31, 0, 25, 9, 0, 0, 0, 0, 6, 14, 0, 0, 0, 0, 0, 
    36, 0, 22, 43, 23, 0, 0, 37, 0, 0, 0, 0, 13, 0, 0, 
    74, 4, 0, 21, 12, 6, 0, 22, 28, 49, 46, 0, 0, 0, 0, 
    128, 6, 1, 7, 4, 1, 0, 21, 54, 0, 0, 0, 0, 0, 0, 
    88, 15, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    51, 51, 51, 51, 51, 51, 51, 53, 53, 49, 48, 51, 51, 51, 51, 
    51, 51, 51, 51, 51, 51, 50, 52, 48, 36, 27, 46, 51, 51, 51, 
    50, 51, 52, 51, 52, 52, 45, 40, 14, 14, 11, 32, 50, 51, 50, 
    35, 41, 46, 52, 54, 53, 40, 47, 34, 33, 35, 31, 40, 42, 46, 
    0, 0, 29, 50, 51, 51, 47, 48, 45, 37, 14, 0, 0, 4, 40, 
    39, 47, 46, 33, 34, 0, 0, 2, 11, 32, 33, 41, 48, 35, 37, 
    0, 0, 8, 30, 34, 6, 0, 21, 35, 37, 22, 14, 13, 13, 6, 
    0, 33, 22, 29, 35, 50, 51, 33, 12, 14, 16, 19, 21, 29, 21, 
    20, 40, 42, 45, 33, 25, 12, 10, 15, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 26, 
    10, 0, 30, 26, 14, 7, 26, 31, 19, 25, 39, 49, 43, 41, 34, 
    22, 4, 21, 21, 12, 12, 32, 143, 152, 128, 84, 59, 47, 32, 25, 
    23, 13, 14, 16, 13, 13, 58, 207, 163, 93, 63, 45, 31, 22, 19, 
    19, 20, 14, 12, 17, 13, 23, 77, 67, 58, 45, 24, 24, 23, 21, 
    
    -- channel=30
    129, 130, 130, 130, 130, 130, 131, 129, 130, 130, 132, 130, 130, 130, 131, 
    130, 131, 131, 130, 131, 130, 131, 130, 127, 118, 140, 134, 130, 130, 131, 
    132, 131, 132, 131, 131, 129, 134, 123, 127, 111, 120, 148, 131, 132, 133, 
    132, 131, 132, 131, 131, 121, 137, 118, 112, 102, 97, 122, 135, 134, 134, 
    123, 135, 150, 132, 132, 124, 123, 128, 129, 129, 133, 135, 128, 155, 140, 
    88, 95, 117, 118, 132, 122, 145, 147, 156, 135, 107, 93, 76, 110, 139, 
    112, 132, 125, 121, 104, 44, 64, 76, 102, 129, 133, 131, 134, 129, 146, 
    72, 66, 72, 114, 125, 85, 92, 100, 118, 104, 77, 68, 73, 81, 93, 
    71, 108, 85, 100, 126, 132, 138, 117, 105, 110, 122, 110, 118, 122, 111, 
    106, 123, 127, 127, 127, 122, 109, 95, 99, 81, 87, 77, 71, 73, 83, 
    27, 52, 45, 56, 66, 83, 91, 92, 86, 73, 67, 64, 67, 57, 72, 
    0, 17, 6, 0, 0, 0, 45, 0, 16, 20, 27, 33, 56, 64, 70, 
    0, 0, 0, 0, 0, 0, 61, 47, 33, 31, 41, 49, 36, 59, 86, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 52, 71, 101, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 39, 52, 62, 78, 103, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 21, 14, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 53, 133, 101, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    93, 92, 102, 124, 124, 132, 131, 128, 124, 137, 154, 136, 136, 128, 135, 
    102, 100, 115, 129, 125, 133, 134, 133, 130, 146, 146, 134, 144, 138, 139, 
    110, 110, 116, 124, 119, 125, 120, 148, 150, 141, 100, 161, 150, 140, 139, 
    127, 108, 130, 145, 139, 128, 126, 91, 137, 120, 66, 136, 158, 146, 169, 
    126, 107, 109, 121, 140, 145, 140, 121, 72, 44, 45, 8, 40, 64, 95, 
    0, 9, 21, 14, 0, 12, 35, 58, 39, 22, 1, 0, 19, 46, 57, 
    20, 38, 44, 23, 53, 44, 28, 13, 0, 0, 25, 102, 94, 87, 101, 
    16, 0, 0, 5, 45, 64, 73, 86, 103, 105, 98, 88, 86, 41, 0, 
    72, 102, 85, 91, 108, 122, 109, 78, 59, 38, 7, 59, 79, 72, 98, 
    32, 2, 50, 90, 78, 52, 64, 98, 114, 80, 76, 92, 110, 101, 71, 
    63, 61, 71, 92, 107, 103, 81, 75, 39, 87, 115, 97, 57, 34, 21, 
    43, 77, 66, 48, 17, 39, 102, 56, 40, 49, 50, 37, 10, 6, 0, 
    54, 97, 100, 66, 70, 66, 39, 22, 42, 39, 13, 7, 15, 0, 0, 
    34, 36, 18, 10, 13, 21, 20, 12, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 9, 17, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 3, 0, 10, 7, 7, 13, 7, 5, 13, 
    0, 1, 1, 0, 4, 7, 8, 5, 12, 0, 22, 17, 10, 9, 19, 
    0, 15, 17, 12, 18, 15, 5, 15, 23, 0, 37, 18, 9, 17, 25, 
    0, 28, 25, 28, 26, 29, 17, 11, 0, 0, 0, 0, 25, 22, 39, 
    0, 3, 4, 17, 14, 17, 7, 0, 0, 0, 0, 20, 36, 10, 29, 
    1, 10, 0, 7, 0, 1, 0, 0, 0, 0, 23, 26, 8, 27, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 23, 7, 41, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 19, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 27, 17, 7, 13, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 6, 6, 
    0, 0, 0, 5, 4, 2, 0, 0, 14, 0, 2, 4, 4, 8, 10, 
    11, 13, 10, 9, 9, 8, 5, 3, 23, 0, 6, 6, 9, 10, 2, 
    
    -- channel=34
    85, 63, 90, 94, 95, 88, 91, 92, 87, 95, 86, 90, 89, 93, 89, 
    80, 56, 81, 82, 85, 77, 85, 89, 85, 89, 67, 89, 87, 93, 82, 
    73, 45, 67, 69, 74, 70, 76, 70, 72, 69, 50, 76, 77, 78, 78, 
    58, 26, 52, 53, 60, 55, 65, 50, 44, 51, 19, 32, 61, 57, 45, 
    29, 15, 29, 29, 35, 38, 45, 57, 30, 22, 12, 2, 0, 22, 17, 
    1, 4, 9, 1, 24, 27, 38, 40, 18, 15, 2, 25, 7, 35, 3, 
    16, 9, 15, 14, 47, 49, 53, 42, 36, 35, 26, 42, 49, 13, 0, 
    32, 28, 38, 45, 63, 70, 73, 63, 61, 44, 23, 36, 38, 9, 0, 
    51, 42, 50, 74, 79, 73, 64, 54, 45, 37, 19, 34, 40, 29, 27, 
    38, 43, 51, 58, 58, 56, 51, 48, 38, 47, 45, 47, 29, 16, 0, 
    47, 57, 56, 49, 44, 50, 51, 22, 9, 40, 33, 24, 3, 0, 0, 
    32, 49, 46, 24, 21, 33, 40, 5, 0, 13, 4, 0, 0, 0, 0, 
    17, 27, 26, 5, 2, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    261, 239, 289, 291, 301, 291, 297, 295, 290, 302, 291, 300, 293, 300, 294, 
    256, 230, 279, 277, 289, 273, 282, 293, 284, 265, 252, 294, 290, 298, 293, 
    249, 213, 261, 264, 268, 261, 257, 245, 262, 234, 205, 278, 279, 277, 281, 
    228, 195, 229, 248, 244, 245, 239, 213, 177, 160, 127, 125, 208, 235, 231, 
    148, 129, 139, 142, 160, 167, 184, 183, 158, 138, 131, 129, 135, 170, 126, 
    110, 107, 126, 121, 141, 134, 165, 159, 139, 138, 147, 190, 146, 167, 103, 
    129, 121, 121, 136, 180, 192, 190, 180, 168, 169, 179, 210, 199, 122, 111, 
    160, 164, 176, 198, 225, 237, 241, 227, 227, 186, 169, 182, 189, 136, 106, 
    174, 178, 200, 238, 238, 235, 225, 208, 190, 187, 161, 181, 187, 168, 163, 
    165, 167, 201, 208, 218, 207, 207, 195, 191, 205, 198, 188, 159, 129, 105, 
    205, 202, 199, 185, 183, 215, 186, 131, 124, 169, 165, 142, 100, 79, 56, 
    164, 193, 175, 133, 131, 154, 169, 129, 117, 119, 97, 89, 64, 49, 31, 
    134, 154, 148, 122, 116, 111, 101, 92, 86, 88, 67, 60, 52, 34, 26, 
    59, 60, 58, 59, 63, 64, 69, 62, 73, 57, 50, 37, 33, 29, 29, 
    23, 22, 30, 35, 42, 46, 49, 41, 62, 57, 30, 29, 26, 31, 5, 
    
    -- channel=36
    31, 13, 21, 35, 38, 46, 52, 61, 49, 57, 72, 61, 59, 56, 51, 
    49, 30, 39, 55, 58, 63, 66, 67, 56, 101, 72, 57, 69, 68, 59, 
    61, 42, 50, 65, 68, 70, 77, 86, 79, 125, 38, 81, 89, 83, 65, 
    81, 46, 69, 83, 89, 75, 84, 69, 116, 113, 63, 113, 101, 99, 102, 
    106, 91, 100, 99, 117, 115, 105, 99, 52, 32, 29, 0, 19, 81, 89, 
    1, 1, 28, 15, 0, 3, 10, 32, 29, 26, 0, 0, 39, 47, 54, 
    6, 33, 40, 6, 18, 15, 0, 0, 0, 0, 0, 61, 77, 62, 113, 
    0, 0, 0, 0, 0, 3, 14, 29, 44, 80, 75, 62, 59, 58, 0, 
    19, 58, 29, 21, 33, 57, 63, 51, 23, 28, 0, 35, 51, 49, 78, 
    8, 0, 0, 35, 34, 11, 22, 57, 71, 49, 40, 60, 89, 101, 79, 
    18, 13, 23, 47, 56, 58, 67, 71, 25, 61, 94, 95, 73, 61, 52, 
    9, 35, 51, 39, 12, 5, 71, 48, 44, 57, 65, 65, 41, 42, 43, 
    24, 61, 74, 52, 68, 73, 48, 35, 56, 63, 44, 34, 50, 30, 24, 
    56, 58, 49, 36, 41, 51, 51, 47, 14, 28, 39, 31, 32, 21, 22, 
    32, 25, 26, 24, 21, 19, 30, 43, 29, 55, 25, 27, 24, 20, 46, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 0, 7, 3, 18, 0, 0, 0, 
    7, 0, 7, 11, 3, 0, 0, 0, 29, 54, 0, 49, 96, 39, 32, 
    70, 38, 50, 62, 69, 67, 52, 52, 7, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 23, 0, 0, 0, 0, 
    0, 33, 0, 0, 0, 12, 2, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 9, 28, 0, 0, 0, 32, 42, 28, 
    0, 0, 0, 15, 38, 22, 0, 3, 0, 27, 42, 37, 23, 18, 21, 
    0, 0, 0, 0, 0, 0, 46, 9, 0, 7, 20, 18, 0, 6, 9, 
    22, 43, 62, 31, 28, 27, 7, 0, 23, 22, 3, 3, 15, 2, 0, 
    22, 28, 15, 9, 13, 20, 11, 5, 0, 0, 9, 1, 1, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 12, 7, 3, 2, 0, 0, 0, 15, 
    
    -- channel=38
    0, 34, 25, 0, 0, 0, 0, 0, 14, 0, 0, 4, 0, 0, 3, 
    0, 31, 31, 0, 1, 0, 0, 0, 6, 0, 60, 22, 0, 0, 13, 
    0, 22, 36, 0, 0, 0, 0, 4, 31, 0, 127, 47, 0, 0, 22, 
    0, 28, 18, 21, 0, 6, 0, 0, 0, 0, 18, 17, 112, 8, 33, 
    0, 15, 0, 34, 9, 21, 12, 0, 0, 0, 5, 16, 43, 0, 15, 
    32, 19, 0, 26, 3, 0, 7, 0, 0, 0, 64, 34, 0, 34, 0, 
    15, 0, 0, 61, 24, 0, 0, 0, 0, 0, 60, 10, 0, 0, 0, 
    0, 0, 14, 20, 8, 0, 0, 0, 0, 0, 43, 28, 0, 0, 0, 
    0, 0, 53, 25, 0, 0, 0, 0, 4, 0, 30, 0, 0, 0, 0, 
    0, 38, 16, 0, 1, 0, 0, 0, 17, 5, 0, 0, 0, 0, 0, 
    45, 0, 0, 0, 15, 42, 0, 0, 61, 13, 0, 0, 0, 0, 0, 
    78, 0, 0, 0, 2, 53, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    50, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 2, 0, 13, 4, 4, 4, 0, 36, 0, 0, 0, 0, 1, 0, 
    0, 8, 4, 6, 3, 2, 0, 0, 74, 0, 0, 0, 0, 8, 0, 
    
    -- channel=39
    89, 79, 75, 61, 55, 42, 30, 31, 27, 22, 8, 17, 24, 24, 21, 
    65, 52, 45, 33, 27, 18, 12, 16, 19, 0, 1, 11, 12, 11, 12, 
    41, 31, 20, 15, 5, 8, 6, 0, 0, 7, 7, 0, 0, 0, 0, 
    9, 15, 0, 0, 0, 0, 0, 10, 0, 17, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 58, 70, 62, 80, 30, 4, 0, 
    86, 75, 67, 73, 84, 83, 83, 80, 73, 80, 94, 77, 37, 4, 30, 
    80, 60, 65, 72, 75, 94, 110, 120, 122, 104, 58, 1, 14, 0, 5, 
    112, 116, 128, 129, 110, 101, 97, 79, 57, 26, 0, 0, 14, 48, 92, 
    78, 52, 73, 81, 76, 61, 57, 64, 63, 76, 64, 37, 29, 25, 0, 
    117, 119, 98, 72, 86, 91, 74, 38, 25, 44, 41, 25, 1, 0, 7, 
    98, 99, 85, 62, 41, 52, 48, 45, 51, 20, 8, 19, 25, 39, 24, 
    77, 77, 74, 74, 89, 64, 39, 53, 47, 42, 34, 43, 49, 43, 45, 
    60, 41, 42, 48, 36, 32, 52, 56, 38, 41, 51, 49, 46, 56, 60, 
    33, 36, 47, 53, 48, 41, 47, 49, 72, 63, 50, 49, 55, 61, 56, 
    49, 54, 58, 59, 65, 66, 59, 43, 40, 53, 50, 54, 58, 59, 32, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    76, 92, 99, 85, 84, 77, 79, 72, 83, 75, 61, 80, 78, 80, 83, 
    64, 81, 83, 70, 72, 63, 58, 64, 76, 25, 44, 78, 67, 66, 75, 
    53, 64, 72, 64, 64, 59, 45, 24, 41, 0, 57, 43, 43, 49, 66, 
    19, 41, 22, 21, 25, 43, 33, 47, 0, 0, 14, 0, 0, 3, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 38, 41, 69, 61, 10, 0, 
    67, 71, 44, 62, 96, 79, 71, 37, 47, 60, 107, 139, 64, 52, 24, 
    57, 38, 20, 70, 64, 85, 96, 109, 127, 111, 105, 43, 25, 0, 0, 
    89, 102, 131, 133, 109, 99, 91, 66, 48, 3, 10, 36, 40, 48, 123, 
    39, 10, 45, 69, 52, 36, 39, 58, 75, 73, 104, 62, 45, 38, 1, 
    66, 114, 87, 47, 63, 90, 73, 26, 22, 51, 54, 26, 0, 0, 0, 
    65, 72, 56, 25, 9, 36, 27, 3, 50, 21, 0, 0, 0, 2, 0, 
    64, 50, 32, 32, 65, 62, 0, 21, 31, 16, 5, 6, 14, 9, 0, 
    30, 0, 0, 3, 0, 0, 16, 28, 4, 0, 15, 17, 0, 13, 20, 
    0, 0, 3, 15, 12, 7, 10, 11, 53, 26, 9, 13, 13, 23, 18, 
    12, 23, 27, 31, 36, 38, 26, 2, 30, 0, 15, 12, 18, 23, 0, 
    
    -- channel=42
    3, 1, 13, 27, 33, 44, 53, 57, 55, 60, 64, 64, 65, 63, 63, 
    21, 17, 33, 46, 51, 56, 56, 53, 60, 62, 37, 65, 71, 67, 66, 
    34, 29, 46, 61, 67, 61, 61, 52, 50, 47, 14, 46, 67, 68, 66, 
    38, 31, 52, 57, 75, 64, 66, 47, 26, 0, 0, 16, 6, 55, 65, 
    0, 0, 10, 17, 25, 26, 17, 10, 0, 0, 0, 0, 33, 47, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 61, 33, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 23, 55, 48, 60, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 38, 43, 28, 22, 
    0, 0, 0, 0, 0, 0, 0, 1, 13, 17, 29, 37, 29, 27, 40, 
    0, 0, 0, 0, 0, 0, 4, 7, 0, 12, 22, 23, 15, 7, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 2, 6, 0, 0, 2, 7, 2, 0, 31, 48, 1, 0, 0, 0, 
    0, 16, 12, 0, 1, 0, 4, 59, 37, 18, 55, 52, 10, 16, 11, 
    19, 14, 39, 33, 25, 11, 8, 0, 95, 79, 84, 163, 125, 61, 75, 
    102, 86, 96, 119, 112, 112, 85, 63, 3, 0, 17, 0, 10, 9, 74, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 
    7, 4, 15, 10, 10, 0, 0, 0, 0, 0, 0, 25, 0, 55, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 39, 67, 22, 0, 0, 0, 
    21, 66, 38, 9, 20, 44, 40, 2, 0, 0, 0, 0, 2, 0, 50, 
    0, 0, 0, 30, 0, 0, 0, 31, 50, 6, 1, 11, 58, 65, 57, 
    5, 0, 5, 28, 72, 44, 21, 38, 22, 50, 71, 58, 32, 22, 31, 
    36, 17, 14, 18, 0, 24, 39, 7, 23, 26, 32, 34, 8, 18, 7, 
    47, 63, 62, 43, 64, 64, 15, 7, 40, 39, 4, 17, 15, 3, 0, 
    57, 50, 28, 17, 20, 32, 29, 19, 0, 0, 13, 8, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 17, 27, 0, 8, 0, 0, 0, 19, 
    
    -- channel=44
    20, 0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 0, 5, 0, 0, 
    22, 0, 0, 7, 0, 5, 0, 0, 0, 69, 0, 0, 14, 0, 0, 
    25, 0, 0, 5, 0, 1, 15, 0, 0, 115, 0, 0, 21, 0, 0, 
    29, 0, 0, 0, 1, 0, 2, 42, 66, 11, 0, 7, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 18, 13, 16, 0, 0, 0, 34, 13, 
    0, 0, 26, 0, 0, 0, 0, 17, 0, 0, 0, 0, 114, 0, 74, 
    0, 21, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 38, 111, 
    0, 0, 0, 0, 0, 0, 0, 25, 0, 65, 0, 0, 3, 83, 0, 
    14, 1, 0, 0, 8, 6, 0, 0, 0, 14, 0, 1, 1, 26, 0, 
    4, 0, 0, 7, 0, 0, 0, 29, 0, 0, 0, 28, 35, 41, 6, 
    0, 0, 5, 23, 0, 0, 50, 30, 0, 0, 23, 22, 26, 9, 28, 
    0, 0, 40, 3, 0, 0, 30, 23, 0, 0, 23, 3, 17, 15, 16, 
    0, 13, 12, 14, 7, 0, 0, 4, 15, 0, 10, 0, 26, 1, 4, 
    9, 0, 0, 0, 0, 0, 0, 5, 0, 45, 1, 11, 5, 0, 7, 
    2, 0, 0, 0, 0, 0, 2, 18, 0, 55, 3, 5, 0, 0, 45, 
    
    -- channel=45
    9, 1, 15, 20, 32, 36, 41, 46, 41, 46, 44, 47, 46, 49, 48, 
    18, 10, 26, 34, 42, 42, 46, 46, 43, 37, 23, 49, 50, 53, 51, 
    29, 18, 35, 48, 50, 47, 49, 34, 32, 34, 8, 30, 48, 53, 51, 
    38, 32, 51, 59, 64, 57, 53, 39, 2, 0, 0, 0, 8, 45, 47, 
    4, 1, 10, 10, 21, 16, 11, 3, 0, 0, 0, 23, 30, 53, 19, 
    0, 0, 9, 6, 15, 3, 0, 0, 0, 0, 11, 51, 58, 51, 22, 
    0, 0, 0, 0, 0, 1, 1, 4, 7, 11, 27, 45, 57, 38, 17, 
    0, 11, 14, 10, 8, 3, 0, 1, 3, 14, 18, 39, 42, 41, 54, 
    0, 0, 0, 0, 0, 0, 0, 1, 13, 32, 35, 35, 30, 33, 34, 
    0, 0, 0, 0, 0, 0, 6, 2, 0, 16, 24, 27, 11, 8, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 8, 
    
    -- channel=46
    121, 121, 145, 142, 144, 138, 140, 134, 139, 142, 138, 141, 133, 138, 137, 
    118, 116, 140, 131, 139, 127, 132, 139, 135, 120, 132, 141, 131, 138, 137, 
    113, 106, 130, 120, 127, 119, 116, 124, 134, 93, 120, 147, 128, 131, 135, 
    104, 90, 110, 117, 112, 112, 108, 91, 89, 78, 71, 79, 130, 117, 120, 
    81, 72, 75, 83, 87, 93, 98, 89, 71, 65, 67, 50, 65, 67, 62, 
    50, 49, 50, 56, 57, 55, 77, 73, 69, 64, 69, 79, 37, 83, 30, 
    65, 57, 54, 73, 91, 87, 86, 77, 68, 70, 85, 100, 76, 51, 34, 
    71, 67, 72, 87, 105, 112, 115, 108, 114, 86, 93, 88, 81, 35, 22, 
    86, 99, 108, 122, 120, 123, 118, 103, 92, 72, 67, 78, 84, 69, 82, 
    71, 78, 101, 105, 109, 100, 99, 95, 104, 100, 91, 84, 79, 61, 52, 
    110, 101, 99, 93, 103, 119, 86, 61, 67, 91, 88, 70, 48, 37, 25, 
    99, 100, 83, 66, 64, 84, 81, 62, 61, 59, 49, 48, 25, 21, 8, 
    78, 85, 80, 66, 68, 64, 50, 45, 47, 47, 29, 29, 20, 12, 7, 
    34, 35, 32, 33, 34, 36, 38, 30, 35, 18, 22, 13, 11, 9, 7, 
    6, 8, 12, 14, 17, 19, 24, 16, 41, 16, 11, 8, 8, 12, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    69, 91, 84, 81, 87, 83, 81, 80, 76, 80, 81, 84, 79, 86, 106, 
    79, 105, 100, 116, 126, 166, 167, 158, 167, 164, 165, 159, 115, 121, 120, 
    81, 102, 116, 134, 72, 52, 73, 67, 62, 58, 67, 82, 131, 114, 120, 
    75, 99, 87, 64, 75, 80, 62, 72, 88, 89, 82, 72, 93, 117, 121, 
    77, 96, 96, 93, 92, 97, 93, 90, 104, 97, 89, 88, 102, 109, 119, 
    89, 109, 143, 96, 64, 65, 69, 77, 77, 72, 72, 92, 113, 110, 111, 
    92, 81, 43, 138, 181, 132, 113, 115, 114, 112, 115, 117, 117, 121, 126, 
    95, 111, 78, 0, 37, 137, 164, 130, 121, 119, 110, 112, 108, 108, 112, 
    98, 119, 120, 109, 60, 17, 81, 172, 195, 161, 129, 111, 114, 117, 118, 
    97, 120, 122, 128, 126, 22, 15, 13, 32, 94, 162, 206, 192, 149, 121, 
    100, 119, 122, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 101, 
    168, 196, 202, 204, 209, 186, 129, 137, 169, 137, 131, 122, 125, 148, 151, 
    44, 47, 40, 39, 36, 39, 41, 66, 94, 99, 105, 113, 124, 127, 127, 
    59, 60, 56, 41, 30, 25, 22, 21, 12, 4, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 
    
    -- channel=49
    16, 0, 0, 0, 6, 0, 0, 2, 0, 0, 0, 0, 6, 6, 4, 
    6, 0, 0, 0, 32, 29, 23, 28, 24, 26, 22, 26, 10, 0, 0, 
    7, 0, 0, 8, 29, 46, 35, 49, 33, 31, 35, 31, 19, 0, 0, 
    4, 0, 0, 23, 29, 24, 25, 28, 24, 17, 32, 19, 32, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 15, 25, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 2, 0, 0, 0, 25, 29, 23, 12, 0, 0, 0, 0, 0, 0, 
    21, 4, 1, 0, 0, 24, 31, 29, 24, 7, 16, 12, 12, 1, 0, 
    20, 0, 0, 0, 10, 0, 16, 52, 18, 19, 19, 17, 44, 15, 3, 
    20, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 
    22, 2, 4, 7, 12, 12, 11, 9, 0, 2, 0, 0, 0, 0, 0, 
    27, 14, 15, 22, 24, 25, 24, 27, 29, 28, 32, 29, 29, 30, 41, 
    35, 26, 26, 31, 29, 32, 29, 35, 31, 32, 33, 37, 36, 40, 6, 
    
    -- channel=50
    57, 86, 69, 53, 64, 69, 66, 65, 62, 65, 68, 68, 69, 77, 78, 
    62, 83, 79, 27, 27, 31, 35, 31, 35, 38, 43, 42, 76, 81, 84, 
    58, 79, 72, 46, 33, 28, 16, 33, 41, 41, 37, 41, 63, 83, 81, 
    59, 78, 66, 28, 39, 40, 36, 30, 42, 41, 38, 41, 56, 79, 86, 
    63, 76, 82, 73, 61, 62, 61, 64, 68, 64, 59, 71, 76, 82, 84, 
    69, 77, 69, 74, 72, 68, 71, 75, 73, 70, 69, 72, 82, 80, 82, 
    71, 67, 39, 40, 59, 71, 82, 87, 84, 80, 79, 81, 81, 82, 85, 
    74, 84, 80, 25, 0, 33, 63, 77, 83, 82, 78, 79, 81, 81, 84, 
    72, 82, 83, 81, 19, 0, 0, 38, 53, 60, 73, 84, 84, 81, 83, 
    69, 79, 83, 80, 22, 0, 0, 0, 0, 0, 22, 45, 48, 61, 78, 
    69, 84, 84, 76, 35, 0, 0, 4, 13, 0, 0, 0, 19, 43, 74, 
    51, 63, 59, 58, 56, 55, 31, 40, 71, 64, 60, 64, 62, 78, 79, 
    2, 15, 12, 5, 0, 0, 0, 2, 9, 5, 4, 7, 9, 8, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    222, 256, 232, 211, 224, 231, 225, 222, 223, 226, 228, 227, 235, 250, 260, 
    231, 264, 257, 183, 190, 219, 214, 219, 221, 224, 228, 227, 266, 264, 269, 
    227, 260, 256, 195, 177, 161, 156, 171, 178, 179, 185, 196, 253, 266, 273, 
    226, 258, 221, 156, 176, 185, 166, 169, 186, 180, 178, 187, 209, 265, 270, 
    239, 254, 254, 228, 212, 210, 217, 219, 223, 217, 211, 235, 253, 264, 270, 
    252, 247, 240, 267, 242, 241, 247, 252, 248, 245, 243, 253, 264, 263, 268, 
    256, 246, 167, 144, 231, 274, 270, 273, 272, 265, 265, 265, 265, 266, 270, 
    262, 278, 257, 180, 84, 169, 255, 279, 268, 262, 259, 262, 263, 262, 265, 
    264, 278, 275, 264, 129, 71, 100, 163, 225, 255, 269, 268, 265, 263, 269, 
    260, 268, 274, 256, 139, 35, 59, 72, 75, 88, 124, 184, 233, 261, 271, 
    258, 270, 272, 252, 176, 98, 67, 112, 151, 106, 105, 86, 139, 206, 240, 
    212, 227, 221, 217, 215, 205, 182, 205, 223, 211, 213, 216, 218, 227, 230, 
    125, 138, 130, 121, 115, 114, 113, 126, 135, 130, 131, 133, 140, 138, 130, 
    67, 72, 71, 62, 51, 49, 47, 48, 46, 36, 34, 35, 36, 37, 69, 
    42, 39, 39, 35, 35, 45, 41, 41, 44, 39, 32, 29, 48, 75, 80, 
    
    -- channel=52
    19, 17, 31, 26, 27, 30, 34, 29, 28, 30, 30, 32, 19, 19, 35, 
    19, 28, 29, 52, 42, 63, 76, 57, 62, 64, 64, 55, 33, 42, 40, 
    23, 31, 35, 33, 12, 0, 2, 0, 0, 0, 0, 0, 33, 41, 40, 
    16, 25, 40, 18, 25, 22, 26, 17, 32, 44, 37, 29, 17, 45, 42, 
    21, 25, 26, 34, 35, 39, 36, 27, 36, 44, 37, 18, 19, 32, 36, 
    32, 36, 64, 26, 0, 0, 0, 3, 4, 7, 8, 16, 37, 36, 31, 
    36, 37, 44, 86, 90, 49, 29, 29, 31, 33, 34, 38, 39, 42, 43, 
    34, 34, 24, 1, 28, 71, 74, 49, 41, 43, 37, 37, 33, 34, 32, 
    35, 44, 46, 45, 73, 39, 76, 115, 112, 79, 42, 29, 35, 40, 37, 
    39, 47, 48, 64, 135, 48, 40, 36, 57, 103, 117, 138, 113, 68, 37, 
    40, 41, 45, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    98, 112, 126, 130, 133, 122, 71, 65, 87, 61, 55, 45, 45, 58, 60, 
    34, 21, 18, 24, 29, 31, 25, 35, 63, 66, 73, 76, 83, 88, 92, 
    83, 78, 77, 71, 73, 65, 59, 61, 61, 59, 52, 48, 46, 45, 13, 
    55, 42, 38, 39, 45, 26, 25, 27, 31, 26, 33, 46, 37, 6, 89, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 28, 29, 32, 28, 35, 24, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 93, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 74, 62, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 102, 105, 43, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 21, 12, 0, 0, 40, 101, 134, 103, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    90, 95, 105, 112, 116, 113, 74, 58, 72, 48, 48, 39, 30, 45, 46, 
    0, 0, 0, 0, 0, 2, 4, 18, 35, 45, 50, 55, 61, 62, 60, 
    13, 25, 24, 14, 13, 12, 7, 5, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    
    -- channel=54
    53, 6, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    47, 17, 0, 0, 16, 9, 0, 18, 0, 4, 1, 29, 21, 0, 0, 
    43, 13, 0, 0, 0, 1, 0, 22, 0, 0, 4, 25, 34, 0, 0, 
    27, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 
    1, 12, 0, 0, 0, 0, 0, 0, 0, 0, 1, 31, 0, 0, 0, 
    4, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    19, 0, 0, 7, 85, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 100, 88, 9, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 22, 58, 65, 62, 29, 27, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 26, 14, 11, 0, 73, 58, 68, 39, 9, 
    42, 0, 0, 0, 0, 0, 0, 80, 0, 0, 0, 0, 95, 18, 8, 
    46, 4, 2, 7, 16, 0, 16, 60, 0, 0, 10, 1, 10, 1, 7, 
    2, 0, 0, 0, 0, 0, 4, 21, 0, 5, 2, 13, 12, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 53, 
    0, 0, 0, 1, 0, 10, 0, 5, 0, 0, 0, 0, 32, 30, 0, 
    
    -- channel=55
    52, 70, 68, 38, 42, 48, 43, 45, 48, 45, 43, 43, 50, 44, 43, 
    59, 66, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 37, 38, 
    57, 67, 47, 0, 15, 19, 3, 12, 28, 26, 30, 19, 21, 42, 41, 
    63, 70, 37, 10, 12, 26, 20, 13, 10, 0, 0, 8, 23, 40, 43, 
    67, 68, 70, 55, 45, 38, 46, 46, 40, 44, 40, 49, 56, 50, 52, 
    55, 51, 30, 70, 85, 82, 79, 77, 78, 76, 72, 60, 51, 51, 53, 
    46, 75, 51, 0, 0, 40, 54, 54, 54, 51, 48, 49, 47, 42, 43, 
    42, 56, 72, 95, 26, 0, 0, 37, 42, 42, 46, 49, 53, 54, 56, 
    37, 38, 38, 46, 45, 16, 0, 0, 0, 4, 38, 52, 49, 47, 52, 
    29, 29, 34, 18, 8, 7, 14, 18, 2, 0, 0, 0, 0, 15, 46, 
    30, 37, 35, 48, 115, 126, 98, 104, 110, 117, 116, 103, 83, 63, 41, 
    0, 0, 0, 0, 0, 0, 8, 3, 3, 22, 28, 37, 35, 25, 23, 
    32, 50, 54, 47, 41, 43, 44, 33, 20, 13, 9, 5, 2, 0, 0, 
    0, 0, 0, 1, 0, 6, 9, 8, 12, 16, 18, 19, 21, 29, 79, 
    16, 26, 27, 23, 22, 39, 36, 32, 34, 36, 27, 23, 48, 74, 4, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    81, 84, 69, 59, 64, 73, 71, 73, 76, 74, 74, 70, 83, 86, 80, 
    80, 77, 68, 0, 0, 0, 0, 0, 0, 0, 0, 5, 62, 63, 72, 
    75, 77, 46, 5, 27, 52, 27, 46, 61, 59, 58, 59, 52, 70, 73, 
    79, 78, 34, 42, 37, 42, 45, 42, 36, 16, 26, 45, 65, 65, 68, 
    80, 79, 74, 52, 52, 49, 53, 54, 47, 42, 54, 70, 81, 72, 74, 
    80, 59, 25, 75, 102, 103, 101, 95, 95, 95, 94, 89, 70, 74, 81, 
    81, 80, 62, 0, 0, 49, 74, 75, 75, 70, 68, 66, 65, 61, 64, 
    83, 80, 89, 122, 30, 0, 14, 58, 63, 61, 69, 70, 73, 72, 76, 
    80, 74, 72, 66, 9, 18, 0, 0, 0, 7, 54, 73, 69, 67, 71, 
    77, 68, 68, 32, 0, 0, 6, 20, 10, 0, 0, 0, 0, 28, 65, 
    73, 68, 68, 61, 141, 150, 124, 160, 164, 124, 168, 131, 153, 104, 71, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 15, 14, 0, 0, 
    37, 34, 34, 30, 30, 24, 24, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 9, 12, 12, 28, 95, 
    9, 15, 17, 19, 17, 36, 37, 40, 39, 40, 29, 18, 60, 95, 5, 
    
    -- channel=58
    9, 12, 27, 28, 23, 30, 35, 33, 36, 37, 36, 36, 34, 40, 39, 
    4, 8, 20, 69, 59, 51, 57, 48, 54, 51, 47, 41, 32, 38, 39, 
    5, 6, 26, 41, 45, 42, 50, 46, 40, 42, 44, 46, 23, 37, 36, 
    8, 6, 33, 74, 55, 54, 60, 58, 62, 67, 60, 55, 52, 33, 31, 
    14, 8, 12, 23, 12, 14, 12, 19, 15, 20, 23, 17, 29, 27, 26, 
    22, 20, 10, 1, 22, 19, 22, 24, 23, 23, 26, 27, 25, 31, 29, 
    29, 27, 41, 29, 0, 8, 27, 29, 31, 31, 28, 27, 27, 29, 27, 
    31, 30, 34, 43, 41, 0, 0, 28, 36, 33, 32, 29, 28, 28, 23, 
    36, 40, 44, 46, 43, 8, 18, 8, 0, 10, 17, 31, 30, 28, 24, 
    39, 47, 44, 48, 27, 0, 0, 8, 19, 14, 0, 0, 0, 10, 23, 
    33, 40, 42, 44, 36, 45, 23, 22, 43, 44, 26, 41, 24, 43, 35, 
    9, 8, 8, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 5, 2, 4, 11, 5, 3, 5, 7, 7, 4, 3, 2, 1, 1, 
    12, 3, 1, 4, 6, 3, 10, 12, 15, 13, 11, 9, 2, 4, 17, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 6, 0, 18, 44, 75, 65, 58, 65, 63, 58, 44, 0, 1, 0, 
    7, 1, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 
    0, 0, 0, 0, 6, 15, 6, 5, 11, 7, 6, 4, 0, 0, 0, 
    0, 5, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 135, 113, 21, 0, 0, 0, 0, 0, 0, 1, 8, 7, 
    0, 0, 0, 0, 17, 131, 78, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 105, 165, 122, 55, 16, 0, 0, 0, 0, 
    2, 0, 0, 10, 6, 44, 19, 0, 37, 121, 191, 176, 114, 43, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    117, 123, 134, 141, 150, 97, 65, 89, 104, 49, 69, 36, 67, 87, 77, 
    0, 0, 0, 0, 0, 0, 0, 35, 48, 61, 70, 80, 86, 91, 92, 
    53, 65, 55, 42, 36, 34, 29, 26, 13, 8, 6, 3, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    
    -- channel=60
    0, 0, 34, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 87, 0, 0, 19, 3, 14, 5, 6, 0, 0, 0, 0, 
    0, 0, 9, 54, 8, 0, 18, 0, 0, 2, 0, 5, 0, 0, 0, 
    0, 0, 30, 46, 0, 0, 23, 0, 10, 29, 0, 0, 0, 0, 0, 
    0, 0, 0, 31, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 80, 1, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 91, 80, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 208, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 181, 0, 0, 0, 6, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 5, 107, 0, 0, 7, 31, 0, 15, 0, 0, 0, 
    0, 15, 15, 14, 8, 16, 2, 0, 2, 14, 0, 0, 3, 0, 0, 
    0, 3, 11, 8, 10, 9, 6, 0, 19, 7, 11, 5, 4, 15, 10, 
    20, 3, 4, 0, 8, 0, 0, 0, 0, 8, 0, 1, 0, 0, 0, 
    26, 5, 0, 0, 2, 0, 4, 0, 0, 0, 8, 3, 0, 0, 32, 
    
    -- channel=61
    16, 22, 32, 40, 36, 37, 40, 38, 40, 40, 40, 38, 39, 44, 39, 
    12, 13, 30, 97, 101, 98, 95, 98, 101, 93, 92, 75, 51, 40, 40, 
    13, 9, 32, 99, 103, 99, 109, 108, 94, 95, 94, 89, 51, 37, 38, 
    17, 12, 49, 124, 88, 89, 92, 97, 94, 103, 97, 90, 71, 32, 30, 
    26, 15, 20, 36, 28, 25, 25, 35, 30, 32, 33, 29, 42, 29, 28, 
    29, 20, 8, 29, 33, 32, 37, 41, 39, 34, 35, 33, 31, 34, 31, 
    30, 37, 37, 11, 6, 29, 37, 39, 39, 38, 35, 33, 31, 31, 30, 
    30, 34, 43, 67, 28, 7, 20, 40, 41, 38, 37, 34, 33, 32, 26, 
    36, 39, 40, 48, 51, 29, 16, 7, 15, 29, 34, 40, 36, 31, 28, 
    41, 42, 41, 44, 39, 18, 26, 36, 27, 10, 0, 2, 11, 26, 35, 
    34, 43, 40, 54, 71, 69, 47, 52, 66, 55, 55, 50, 41, 46, 38, 
    6, 14, 7, 6, 3, 7, 8, 10, 8, 8, 10, 12, 11, 8, 11, 
    22, 30, 28, 25, 23, 24, 22, 20, 18, 16, 14, 12, 13, 17, 13, 
    18, 22, 21, 21, 21, 19, 20, 21, 21, 19, 18, 18, 19, 13, 3, 
    26, 22, 23, 22, 22, 28, 31, 29, 29, 28, 24, 21, 9, 0, 0, 
    
    -- channel=62
    106, 120, 96, 87, 103, 101, 97, 97, 94, 97, 98, 97, 101, 108, 117, 
    113, 131, 117, 63, 77, 94, 89, 88, 90, 96, 94, 101, 124, 123, 124, 
    113, 127, 117, 67, 54, 43, 37, 50, 54, 51, 62, 74, 120, 125, 126, 
    107, 125, 95, 50, 64, 69, 59, 65, 73, 65, 67, 71, 91, 124, 128, 
    108, 123, 117, 96, 96, 97, 98, 97, 100, 97, 97, 109, 113, 122, 128, 
    117, 115, 121, 124, 104, 103, 106, 108, 105, 105, 107, 115, 125, 122, 125, 
    121, 100, 60, 84, 138, 137, 126, 125, 124, 120, 123, 123, 124, 125, 129, 
    126, 126, 106, 43, 25, 106, 144, 132, 122, 120, 120, 120, 122, 121, 125, 
    126, 129, 127, 115, 13, 32, 62, 105, 132, 131, 130, 120, 121, 123, 127, 
    124, 124, 127, 111, 32, 15, 23, 25, 35, 51, 91, 121, 137, 134, 127, 
    124, 124, 126, 104, 41, 0, 4, 35, 35, 10, 17, 8, 58, 88, 112, 
    120, 125, 123, 122, 125, 107, 95, 112, 115, 102, 107, 103, 108, 113, 116, 
    51, 56, 49, 48, 46, 46, 48, 62, 67, 70, 72, 76, 81, 79, 78, 
    28, 39, 35, 31, 22, 21, 22, 23, 19, 13, 12, 11, 10, 13, 30, 
    4, 11, 9, 8, 8, 10, 6, 9, 7, 4, 3, 7, 23, 28, 47, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 31, 0, 7, 0, 0, 0, 0, 10, 13, 0, 0, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 52, 12, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 34, 27, 30, 
    23, 0, 31, 0, 0, 15, 26, 0, 2, 17, 24, 0, 43, 38, 9, 
    0, 0, 44, 30, 40, 30, 15, 16, 45, 39, 28, 19, 52, 11, 15, 
    14, 0, 8, 36, 5, 39, 27, 35, 28, 0, 23, 59, 28, 36, 46, 
    0, 0, 55, 47, 61, 21, 34, 54, 34, 59, 62, 52, 94, 80, 0, 
    15, 60, 27, 11, 28, 80, 48, 35, 66, 55, 56, 50, 40, 0, 0, 
    46, 0, 0, 0, 0, 0, 30, 69, 64, 79, 63, 52, 37, 11, 0, 
    0, 0, 0, 0, 25, 6, 37, 78, 82, 62, 28, 52, 52, 34, 30, 
    75, 119, 42, 0, 0, 21, 54, 106, 107, 60, 65, 56, 31, 50, 17, 
    0, 50, 89, 40, 0, 0, 12, 0, 0, 65, 62, 70, 72, 0, 0, 
    4, 0, 0, 73, 57, 0, 0, 0, 44, 68, 99, 64, 0, 0, 0, 
    
    -- channel=65
    32, 33, 44, 29, 4, 62, 38, 49, 47, 46, 23, 73, 6, 49, 40, 
    31, 44, 32, 26, 8, 49, 28, 57, 35, 49, 23, 80, 7, 62, 29, 
    28, 32, 32, 23, 12, 58, 57, 41, 34, 18, 42, 82, 20, 41, 37, 
    16, 56, 33, 19, 46, 66, 44, 19, 66, 20, 66, 78, 24, 36, 0, 
    24, 61, 4, 38, 67, 48, 13, 72, 50, 70, 58, 70, 41, 32, 0, 
    19, 61, 31, 12, 60, 52, 56, 56, 50, 48, 41, 89, 39, 29, 0, 
    23, 53, 44, 31, 50, 65, 60, 60, 53, 57, 58, 63, 36, 49, 0, 
    24, 45, 41, 39, 33, 60, 59, 69, 58, 65, 66, 56, 33, 44, 0, 
    42, 48, 33, 33, 60, 31, 65, 54, 57, 54, 59, 59, 46, 40, 11, 
    40, 25, 22, 43, 26, 62, 50, 50, 57, 47, 51, 50, 21, 34, 58, 
    6, 49, 34, 43, 56, 28, 69, 47, 39, 44, 50, 48, 43, 49, 36, 
    51, 65, 44, 61, 17, 59, 52, 52, 49, 38, 55, 56, 55, 59, 32, 
    49, 65, 48, 63, 47, 54, 51, 43, 57, 45, 52, 45, 43, 62, 37, 
    17, 66, 70, 59, 60, 59, 61, 39, 72, 50, 50, 50, 18, 62, 40, 
    24, 36, 89, 84, 58, 57, 57, 55, 55, 56, 47, 37, 38, 44, 87, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 3, 11, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 12, 17, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 15, 6, 0, 0, 0, 0, 0, 
    0, 9, 2, 0, 0, 0, 0, 0, 0, 4, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=67
    48, 13, 26, 47, 11, 5, 35, 35, 52, 67, 60, 68, 61, 23, 45, 
    77, 39, 51, 59, 6, 0, 30, 31, 61, 51, 57, 72, 96, 40, 70, 
    62, 67, 67, 51, 5, 12, 33, 37, 72, 27, 65, 82, 137, 90, 100, 
    32, 52, 54, 52, 12, 42, 54, 23, 38, 59, 56, 88, 154, 121, 94, 
    43, 108, 107, 22, 60, 91, 51, 26, 63, 68, 87, 93, 135, 134, 71, 
    45, 99, 151, 83, 56, 89, 84, 108, 102, 98, 93, 85, 127, 137, 59, 
    49, 77, 124, 139, 101, 92, 86, 91, 98, 102, 107, 114, 119, 119, 79, 
    71, 87, 112, 135, 132, 51, 104, 111, 117, 103, 101, 138, 132, 123, 50, 
    88, 99, 107, 117, 119, 150, 101, 129, 124, 132, 122, 126, 132, 105, 67, 
    104, 104, 68, 91, 100, 98, 152, 147, 146, 150, 126, 122, 97, 56, 84, 
    89, 79, 70, 85, 83, 100, 131, 172, 160, 135, 132, 120, 101, 96, 104, 
    120, 127, 88, 82, 105, 103, 142, 162, 163, 136, 138, 115, 90, 99, 118, 
    107, 166, 168, 110, 93, 109, 131, 106, 133, 154, 137, 123, 77, 65, 96, 
    56, 26, 139, 166, 122, 87, 87, 94, 72, 137, 145, 110, 57, 50, 118, 
    51, 10, 15, 138, 180, 147, 106, 101, 76, 113, 109, 108, 55, 58, 86, 
    
    -- channel=68
    48, 48, 36, 61, 78, 26, 64, 57, 88, 102, 99, 40, 122, 63, 55, 
    54, 51, 75, 57, 79, 48, 80, 45, 78, 60, 100, 26, 107, 4, 68, 
    103, 108, 72, 68, 78, 24, 37, 76, 83, 94, 76, 27, 97, 69, 70, 
    83, 18, 58, 70, 41, 49, 123, 125, 38, 69, 32, 74, 119, 72, 111, 
    71, 38, 83, 62, 45, 76, 107, 13, 70, 62, 103, 117, 108, 82, 126, 
    93, 52, 90, 62, 37, 70, 55, 32, 77, 87, 96, 47, 128, 88, 116, 
    64, 39, 79, 85, 80, 72, 57, 59, 75, 61, 46, 52, 106, 76, 106, 
    91, 61, 64, 91, 45, 58, 60, 55, 56, 32, 47, 52, 63, 91, 128, 
    51, 53, 97, 101, 77, 54, 34, 58, 54, 73, 75, 63, 100, 111, 96, 
    67, 115, 105, 84, 100, 71, 60, 38, 57, 65, 63, 73, 88, 57, 49, 
    117, 62, 87, 55, 62, 77, 32, 65, 62, 78, 74, 72, 75, 58, 61, 
    28, 5, 92, 69, 95, 58, 57, 77, 73, 66, 44, 67, 101, 84, 115, 
    122, 146, 125, 110, 114, 69, 82, 124, 97, 62, 56, 74, 81, 99, 119, 
    92, 116, 154, 118, 115, 118, 120, 86, 19, 69, 67, 85, 132, 65, 95, 
    106, 73, 72, 146, 125, 101, 112, 116, 110, 94, 107, 110, 52, 42, 39, 
    
    -- channel=69
    0, 0, 0, 0, 5, 0, 0, 0, 0, 14, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 7, 21, 0, 0, 0, 2, 0, 0, 0, 0, 
    13, 20, 0, 0, 0, 0, 0, 0, 18, 3, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 13, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 21, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 8, 11, 14, 0, 0, 0, 0, 0, 0, 0, 31, 23, 0, 
    0, 18, 0, 0, 8, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 74, 0, 0, 0, 0, 5, 45, 52, 0, 0, 0, 0, 0, 0, 
    0, 48, 78, 0, 0, 0, 0, 0, 0, 1, 0, 0, 33, 0, 0, 
    9, 0, 23, 52, 0, 0, 0, 0, 0, 33, 58, 13, 0, 0, 0, 
    
    -- channel=70
    0, 0, 29, 9, 0, 95, 0, 38, 7, 28, 0, 123, 0, 65, 10, 
    0, 0, 0, 8, 0, 62, 6, 59, 0, 24, 0, 155, 0, 58, 0, 
    0, 23, 1, 0, 0, 70, 24, 0, 45, 0, 50, 136, 0, 2, 0, 
    0, 99, 0, 0, 2, 65, 0, 0, 99, 0, 52, 94, 0, 0, 0, 
    0, 138, 0, 0, 100, 2, 0, 83, 0, 36, 0, 57, 0, 0, 0, 
    0, 141, 3, 0, 46, 15, 0, 58, 0, 0, 0, 101, 0, 15, 0, 
    0, 77, 57, 0, 0, 8, 0, 0, 0, 15, 8, 15, 0, 26, 0, 
    0, 64, 37, 0, 5, 0, 45, 0, 0, 0, 0, 44, 0, 8, 0, 
    12, 18, 0, 0, 44, 0, 18, 0, 0, 0, 0, 17, 0, 0, 0, 
    1, 0, 0, 50, 11, 41, 17, 13, 0, 0, 0, 0, 0, 0, 50, 
    0, 68, 0, 42, 8, 0, 99, 0, 0, 0, 0, 0, 0, 1, 18, 
    14, 14, 0, 31, 0, 34, 52, 4, 0, 0, 12, 0, 0, 46, 0, 
    31, 100, 0, 0, 0, 49, 14, 0, 74, 0, 0, 0, 0, 41, 0, 
    0, 69, 147, 13, 0, 0, 0, 0, 53, 18, 6, 0, 0, 89, 43, 
    0, 0, 117, 139, 7, 0, 0, 0, 0, 24, 6, 0, 0, 0, 133, 
    
    -- channel=71
    36, 41, 42, 43, 34, 36, 25, 23, 0, 0, 10, 17, 2, 3, 32, 
    38, 36, 29, 39, 32, 10, 11, 29, 22, 22, 14, 17, 27, 53, 31, 
    0, 0, 26, 25, 27, 54, 51, 17, 12, 0, 18, 18, 15, 28, 30, 
    26, 50, 29, 26, 42, 25, 0, 0, 25, 35, 28, 0, 0, 20, 2, 
    32, 27, 39, 17, 27, 10, 7, 52, 27, 26, 0, 0, 0, 19, 16, 
    13, 8, 29, 68, 21, 0, 8, 23, 3, 0, 0, 0, 0, 14, 21, 
    37, 27, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 
    16, 21, 22, 2, 4, 0, 0, 0, 0, 2, 0, 0, 3, 0, 0, 
    37, 31, 1, 2, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 46, 
    0, 6, 25, 35, 33, 13, 0, 0, 0, 0, 0, 0, 0, 34, 26, 
    63, 48, 22, 22, 8, 23, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 24, 22, 0, 0, 0, 0, 7, 33, 
    7, 27, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 46, 53, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    51, 40, 72, 53, 0, 58, 38, 43, 28, 24, 18, 78, 0, 26, 51, 
    59, 65, 44, 54, 0, 24, 12, 57, 49, 58, 16, 92, 35, 106, 58, 
    0, 6, 41, 22, 0, 80, 100, 38, 36, 0, 41, 102, 53, 73, 53, 
    22, 109, 45, 26, 51, 103, 26, 0, 63, 43, 97, 99, 38, 68, 0, 
    34, 94, 65, 12, 80, 68, 7, 101, 80, 96, 53, 43, 51, 57, 0, 
    0, 62, 62, 86, 104, 35, 24, 91, 67, 45, 28, 104, 35, 57, 0, 
    50, 75, 59, 57, 14, 20, 48, 36, 10, 21, 42, 57, 35, 75, 5, 
    26, 68, 75, 39, 77, 10, 33, 31, 47, 71, 39, 46, 47, 48, 0, 
    76, 80, 26, 30, 12, 58, 41, 33, 44, 26, 21, 37, 0, 0, 32, 
    55, 9, 19, 34, 38, 0, 39, 63, 33, 33, 32, 21, 12, 46, 71, 
    0, 66, 38, 71, 58, 59, 64, 39, 42, 3, 17, 22, 24, 58, 94, 
    110, 160, 93, 85, 47, 48, 52, 21, 25, 20, 45, 18, 0, 56, 55, 
    0, 3, 77, 88, 60, 66, 21, 0, 0, 35, 28, 14, 5, 25, 45, 
    15, 0, 4, 82, 84, 80, 49, 65, 81, 19, 35, 0, 0, 52, 75, 
    1, 39, 14, 24, 73, 108, 95, 72, 8, 0, 0, 2, 72, 93, 130, 
    
    -- channel=74
    14, 13, 10, 2, 2, 0, 15, 9, 34, 25, 25, 16, 54, 7, 13, 
    25, 32, 22, 5, 7, 0, 1, 13, 24, 25, 25, 20, 55, 22, 30, 
    22, 5, 10, 10, 1, 2, 25, 27, 3, 28, 6, 35, 63, 37, 34, 
    12, 11, 37, 11, 7, 37, 47, 15, 14, 10, 44, 53, 51, 41, 38, 
    18, 14, 34, 32, 12, 49, 47, 11, 46, 47, 57, 57, 63, 38, 29, 
    24, 11, 31, 40, 49, 53, 43, 38, 61, 60, 61, 48, 67, 27, 35, 
    23, 23, 34, 50, 68, 69, 61, 74, 58, 54, 53, 74, 59, 43, 34, 
    24, 20, 36, 42, 48, 78, 56, 71, 71, 80, 78, 48, 73, 40, 35, 
    26, 43, 36, 34, 60, 36, 70, 67, 79, 76, 74, 70, 60, 39, 15, 
    36, 33, 25, 18, 23, 52, 53, 64, 78, 73, 68, 71, 48, 21, 22, 
    36, 18, 35, 21, 49, 27, 52, 77, 65, 74, 64, 68, 61, 28, 37, 
    38, 81, 85, 47, 29, 46, 60, 77, 68, 65, 66, 75, 73, 37, 37, 
    45, 46, 85, 94, 63, 28, 65, 69, 34, 60, 76, 73, 62, 34, 39, 
    29, 34, 37, 76, 102, 76, 66, 40, 55, 63, 60, 75, 42, 7, 25, 
    32, 8, 41, 54, 77, 99, 90, 78, 64, 46, 46, 40, 42, 41, 70, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 0, 0, 0, 32, 0, 
    0, 0, 0, 0, 0, 27, 18, 0, 0, 0, 0, 1, 0, 0, 0, 
    37, 19, 0, 10, 0, 0, 0, 0, 21, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 33, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 
    0, 38, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 3, 0, 
    0, 0, 27, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 30, 25, 55, 0, 1, 0, 0, 5, 0, 0, 31, 35, 0, 
    0, 32, 5, 9, 13, 94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 13, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 2, 7, 1, 0, 0, 0, 0, 0, 0, 
    88, 91, 0, 0, 0, 0, 24, 67, 73, 0, 11, 0, 0, 26, 5, 
    0, 127, 99, 0, 0, 0, 0, 0, 0, 18, 0, 3, 31, 0, 0, 
    0, 0, 93, 77, 0, 0, 0, 0, 24, 37, 75, 0, 0, 0, 0, 
    
    -- channel=76
    0, 18, 0, 0, 69, 0, 9, 0, 0, 0, 40, 0, 127, 0, 0, 
    0, 23, 0, 0, 81, 0, 0, 0, 0, 0, 30, 0, 73, 0, 19, 
    42, 0, 0, 13, 68, 0, 0, 30, 0, 71, 0, 0, 41, 0, 0, 
    22, 0, 37, 33, 0, 0, 37, 33, 0, 18, 0, 0, 0, 0, 88, 
    45, 0, 59, 37, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 131, 
    78, 0, 0, 74, 0, 0, 16, 0, 11, 0, 0, 0, 36, 0, 147, 
    56, 0, 0, 7, 29, 0, 0, 2, 3, 0, 0, 0, 4, 0, 100, 
    34, 0, 0, 0, 0, 52, 0, 0, 0, 0, 21, 0, 70, 0, 120, 
    0, 0, 1, 0, 0, 47, 0, 0, 11, 0, 0, 15, 20, 13, 67, 
    9, 13, 47, 0, 0, 0, 5, 0, 0, 20, 6, 19, 51, 7, 0, 
    71, 0, 40, 0, 0, 32, 0, 5, 16, 17, 4, 3, 26, 0, 0, 
    0, 0, 59, 0, 6, 0, 0, 0, 0, 35, 0, 19, 29, 0, 0, 
    1, 0, 0, 37, 37, 0, 0, 62, 0, 0, 0, 34, 53, 0, 11, 
    49, 0, 0, 0, 38, 14, 0, 0, 0, 0, 0, 54, 89, 0, 0, 
    58, 15, 0, 0, 0, 20, 18, 0, 35, 0, 6, 0, 31, 0, 0, 
    
    -- channel=77
    10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 1, 
    3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 7, 1, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 30, 0, 3, 
    0, 0, 5, 10, 4, 0, 0, 0, 0, 12, 14, 0, 12, 1, 9, 
    0, 0, 7, 7, 3, 0, 9, 4, 0, 0, 0, 0, 7, 0, 9, 
    1, 0, 0, 16, 1, 28, 50, 26, 15, 12, 22, 1, 1, 0, 20, 
    6, 0, 0, 7, 47, 66, 69, 61, 55, 60, 65, 55, 17, 0, 13, 
    0, 0, 0, 2, 66, 53, 63, 73, 81, 84, 72, 56, 70, 2, 0, 
    4, 0, 0, 0, 25, 74, 67, 73, 78, 72, 70, 62, 59, 13, 4, 
    0, 0, 0, 0, 0, 24, 70, 74, 76, 77, 67, 67, 55, 10, 0, 
    0, 3, 0, 0, 0, 12, 47, 73, 72, 70, 72, 72, 58, 13, 0, 
    25, 50, 21, 0, 0, 9, 52, 78, 67, 69, 81, 77, 58, 6, 0, 
    0, 0, 24, 8, 0, 0, 38, 54, 37, 76, 73, 80, 60, 0, 0, 
    5, 0, 0, 14, 15, 0, 0, 19, 28, 67, 70, 70, 35, 0, 0, 
    3, 1, 0, 0, 15, 14, 0, 0, 13, 46, 41, 39, 28, 9, 1, 
    
    -- channel=78
    17, 0, 15, 27, 0, 13, 13, 23, 32, 44, 21, 48, 3, 23, 15, 
    33, 10, 25, 31, 0, 7, 19, 19, 29, 27, 22, 53, 19, 18, 31, 
    34, 41, 30, 25, 0, 9, 16, 19, 48, 8, 40, 58, 49, 44, 41, 
    10, 35, 15, 15, 0, 35, 30, 9, 27, 14, 35, 58, 76, 57, 31, 
    11, 75, 36, 1, 36, 42, 3, 9, 36, 35, 45, 66, 66, 66, 10, 
    9, 75, 79, 13, 32, 38, 16, 51, 41, 43, 35, 48, 59, 77, 0, 
    7, 49, 77, 65, 32, 30, 23, 29, 32, 36, 35, 36, 53, 66, 10, 
    28, 56, 59, 66, 45, 2, 41, 33, 36, 24, 24, 64, 32, 64, 9, 
    41, 47, 59, 66, 65, 37, 37, 46, 40, 48, 41, 47, 48, 51, 18, 
    50, 56, 35, 53, 56, 62, 53, 53, 53, 51, 42, 40, 26, 18, 43, 
    35, 48, 23, 52, 37, 40, 71, 66, 58, 50, 49, 40, 30, 42, 60, 
    44, 45, 26, 45, 54, 52, 64, 66, 65, 41, 46, 36, 30, 54, 70, 
    68, 115, 75, 44, 43, 63, 65, 42, 74, 56, 54, 34, 14, 44, 59, 
    17, 34, 108, 83, 45, 49, 51, 33, 31, 57, 55, 30, 12, 33, 65, 
    15, 0, 33, 104, 91, 57, 46, 54, 35, 53, 55, 46, 3, 24, 65, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=80
    22, 0, 25, 17, 20, 18, 24, 16, 21, 3, 0, 0, 0, 0, 15, 
    41, 39, 29, 22, 22, 15, 17, 14, 9, 0, 0, 17, 10, 12, 10, 
    45, 23, 25, 36, 31, 36, 21, 24, 26, 0, 0, 0, 14, 25, 7, 
    63, 30, 40, 37, 46, 48, 47, 35, 37, 39, 24, 15, 10, 0, 16, 
    59, 26, 34, 38, 37, 40, 28, 0, 23, 40, 46, 36, 4, 20, 16, 
    25, 31, 12, 39, 54, 22, 30, 82, 60, 11, 38, 42, 0, 8, 10, 
    0, 70, 61, 47, 26, 52, 92, 0, 0, 0, 38, 11, 0, 0, 7, 
    14, 22, 67, 68, 37, 55, 42, 59, 70, 56, 25, 17, 0, 0, 2, 
    26, 18, 50, 69, 58, 91, 77, 108, 104, 124, 119, 13, 0, 5, 17, 
    37, 31, 65, 60, 73, 69, 91, 0, 26, 33, 0, 0, 0, 6, 11, 
    43, 59, 85, 69, 0, 64, 60, 63, 93, 11, 8, 0, 0, 44, 57, 
    69, 31, 60, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 42, 65, 
    33, 52, 41, 78, 26, 31, 10, 1, 0, 0, 0, 0, 0, 0, 11, 
    39, 58, 64, 43, 56, 0, 25, 39, 4, 0, 0, 0, 0, 0, 20, 
    34, 10, 43, 23, 17, 20, 42, 54, 37, 30, 14, 21, 23, 16, 2, 
    
    -- channel=81
    74, 104, 95, 97, 96, 99, 91, 90, 63, 65, 59, 56, 62, 70, 52, 
    92, 89, 98, 100, 102, 107, 105, 101, 77, 68, 61, 66, 69, 63, 67, 
    71, 88, 101, 104, 106, 104, 102, 118, 99, 72, 85, 74, 73, 71, 69, 
    72, 89, 96, 106, 106, 107, 105, 104, 102, 96, 96, 73, 64, 75, 71, 
    67, 89, 98, 104, 107, 104, 83, 85, 81, 99, 97, 56, 71, 69, 67, 
    94, 77, 100, 98, 96, 100, 51, 69, 56, 82, 66, 43, 63, 66, 70, 
    104, 89, 80, 75, 92, 78, 61, 52, 70, 73, 42, 37, 56, 65, 66, 
    66, 100, 70, 81, 86, 75, 89, 80, 62, 55, 39, 40, 59, 67, 57, 
    76, 96, 73, 69, 64, 79, 63, 76, 66, 58, 21, 35, 72, 77, 27, 
    66, 99, 62, 13, 80, 77, 48, 83, 60, 45, 45, 46, 74, 90, 7, 
    72, 90, 57, 4, 56, 48, 44, 80, 43, 47, 45, 47, 73, 91, 14, 
    74, 79, 65, 62, 67, 70, 81, 47, 36, 35, 31, 46, 61, 77, 51, 
    88, 78, 77, 79, 80, 68, 74, 61, 53, 44, 36, 45, 59, 54, 73, 
    72, 83, 67, 77, 48, 73, 85, 63, 72, 62, 66, 75, 70, 79, 54, 
    74, 86, 74, 85, 77, 80, 87, 76, 76, 77, 84, 86, 79, 71, 82, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    60, 33, 44, 46, 47, 33, 32, 36, 34, 12, 24, 19, 21, 29, 35, 
    82, 73, 51, 55, 51, 45, 31, 33, 24, 0, 19, 27, 44, 37, 30, 
    71, 76, 58, 60, 63, 54, 45, 28, 50, 43, 29, 24, 29, 37, 37, 
    93, 72, 67, 68, 71, 64, 56, 43, 47, 63, 45, 23, 20, 23, 39, 
    68, 78, 74, 70, 68, 62, 67, 71, 37, 50, 63, 40, 25, 32, 40, 
    57, 78, 77, 77, 62, 106, 105, 84, 77, 56, 52, 28, 10, 21, 33, 
    20, 111, 115, 101, 89, 115, 121, 99, 77, 89, 62, 18, 6, 18, 23, 
    44, 81, 118, 100, 131, 131, 98, 142, 145, 141, 82, 24, 20, 49, 14, 
    57, 95, 123, 78, 134, 128, 96, 99, 109, 87, 58, 5, 7, 81, 46, 
    59, 89, 149, 64, 71, 110, 92, 91, 46, 19, 5, 0, 9, 101, 83, 
    70, 90, 131, 58, 0, 18, 33, 45, 34, 0, 0, 10, 7, 85, 122, 
    73, 78, 100, 78, 26, 30, 26, 17, 0, 0, 0, 0, 12, 27, 112, 
    60, 82, 75, 94, 58, 50, 56, 36, 17, 0, 0, 0, 0, 11, 37, 
    60, 73, 78, 61, 63, 53, 62, 63, 46, 39, 34, 35, 30, 24, 41, 
    70, 66, 72, 67, 70, 66, 56, 57, 49, 45, 46, 58, 56, 43, 40, 
    
    -- channel=84
    68, 13, 62, 50, 65, 61, 65, 51, 70, 46, 36, 35, 27, 21, 46, 
    71, 89, 66, 60, 61, 57, 61, 53, 69, 46, 36, 37, 29, 42, 37, 
    86, 71, 64, 71, 67, 73, 68, 61, 64, 34, 0, 29, 35, 46, 33, 
    92, 66, 76, 67, 75, 78, 73, 72, 64, 65, 59, 65, 47, 28, 38, 
    78, 58, 69, 76, 73, 79, 61, 38, 59, 59, 65, 95, 42, 48, 43, 
    41, 65, 50, 73, 94, 54, 53, 80, 99, 39, 62, 91, 36, 47, 39, 
    0, 74, 76, 78, 51, 67, 102, 37, 0, 19, 69, 54, 27, 37, 41, 
    43, 18, 78, 76, 49, 64, 55, 56, 64, 63, 64, 59, 32, 12, 41, 
    36, 14, 57, 84, 89, 87, 86, 114, 109, 126, 150, 70, 11, 27, 73, 
    52, 19, 61, 116, 65, 71, 102, 1, 54, 68, 19, 13, 11, 14, 76, 
    47, 41, 88, 119, 17, 92, 87, 71, 121, 64, 59, 42, 11, 28, 100, 
    60, 30, 67, 27, 27, 0, 0, 54, 54, 39, 37, 39, 35, 48, 82, 
    33, 47, 50, 75, 57, 57, 21, 26, 15, 8, 8, 2, 12, 42, 40, 
    48, 40, 63, 53, 77, 26, 23, 50, 23, 12, 10, 0, 8, 7, 48, 
    37, 10, 41, 20, 28, 26, 51, 58, 50, 40, 29, 32, 35, 45, 20, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 5, 6, 0, 
    12, 0, 0, 0, 0, 0, 0, 44, 27, 0, 0, 19, 12, 0, 0, 
    0, 12, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 20, 1, 0, 52, 53, 71, 99, 23, 0, 0, 0, 
    0, 0, 0, 0, 119, 5, 33, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 10, 31, 0, 62, 61, 45, 70, 4, 30, 30, 0, 17, 7, 
    11, 0, 5, 0, 0, 0, 0, 0, 0, 10, 12, 13, 19, 11, 45, 
    0, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 5, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 15, 0, 3, 0, 0, 0, 10, 0, 2, 4, 0, 1, 25, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 4, 17, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 1, 1, 1, 
    0, 1, 0, 11, 0, 0, 0, 0, 12, 0, 0, 0, 0, 17, 3, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 34, 3, 0, 26, 2, 6, 
    160, 0, 8, 0, 0, 58, 0, 0, 0, 35, 0, 0, 30, 4, 18, 
    129, 71, 0, 0, 17, 9, 0, 0, 10, 0, 0, 0, 15, 12, 3, 
    0, 134, 0, 0, 51, 0, 0, 20, 0, 0, 0, 0, 38, 35, 0, 
    0, 105, 0, 0, 52, 32, 0, 9, 13, 0, 0, 0, 85, 84, 0, 
    0, 112, 0, 0, 130, 47, 0, 53, 0, 0, 0, 0, 71, 133, 0, 
    0, 73, 0, 0, 43, 17, 6, 54, 0, 0, 0, 17, 35, 150, 0, 
    0, 16, 7, 0, 0, 0, 2, 0, 0, 0, 0, 30, 68, 56, 15, 
    10, 0, 0, 24, 0, 0, 16, 0, 0, 0, 0, 9, 40, 10, 45, 
    0, 50, 0, 22, 0, 7, 31, 0, 0, 0, 0, 9, 0, 11, 0, 
    0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 18, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 21, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 9, 0, 0, 0, 10, 19, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 34, 39, 38, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    12, 59, 0, 1, 0, 0, 0, 0, 0, 0, 0, 5, 7, 10, 0, 
    10, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 6, 0, 3, 0, 0, 0, 1, 34, 42, 2, 0, 0, 3, 
    0, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 3, 1, 0, 0, 4, 32, 0, 0, 0, 0, 0, 0, 0, 
    15, 15, 27, 7, 0, 56, 33, 0, 0, 14, 0, 0, 0, 0, 0, 
    44, 1, 4, 8, 38, 24, 0, 58, 90, 54, 0, 0, 6, 0, 0, 
    0, 36, 1, 0, 53, 27, 24, 30, 21, 30, 6, 0, 6, 48, 0, 
    0, 47, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 34, 0, 
    0, 39, 25, 0, 0, 0, 0, 53, 0, 0, 9, 10, 14, 58, 0, 
    0, 4, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 16, 26, 0, 
    0, 7, 6, 44, 13, 44, 29, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 7, 11, 24, 34, 28, 35, 16, 0, 0, 
    0, 0, 0, 0, 0, 8, 2, 0, 14, 20, 25, 47, 35, 28, 0, 
    0, 21, 0, 11, 18, 2, 0, 0, 0, 0, 0, 3, 0, 0, 17, 
    
    -- channel=90
    94, 94, 96, 93, 100, 101, 88, 79, 60, 35, 36, 41, 39, 44, 37, 
    95, 104, 101, 105, 108, 110, 110, 99, 84, 44, 31, 42, 47, 55, 45, 
    100, 89, 108, 111, 113, 118, 114, 112, 101, 72, 65, 62, 57, 51, 52, 
    84, 99, 106, 109, 117, 120, 116, 103, 100, 101, 102, 78, 49, 52, 55, 
    72, 90, 108, 114, 118, 112, 90, 90, 96, 87, 89, 72, 39, 50, 51, 
    30, 105, 108, 114, 117, 86, 85, 66, 58, 67, 75, 46, 33, 43, 48, 
    52, 73, 105, 96, 91, 104, 82, 64, 70, 77, 65, 27, 24, 42, 46, 
    66, 64, 95, 90, 88, 106, 113, 86, 84, 79, 70, 26, 17, 47, 59, 
    74, 69, 93, 88, 70, 83, 101, 79, 64, 66, 36, 5, 16, 51, 51, 
    81, 70, 77, 71, 25, 76, 78, 63, 94, 25, 15, 21, 22, 53, 60, 
    84, 71, 73, 54, 24, 24, 24, 59, 39, 17, 5, 9, 32, 52, 58, 
    77, 77, 64, 76, 74, 43, 57, 49, 8, 0, 0, 0, 10, 51, 42, 
    81, 84, 82, 70, 81, 64, 60, 64, 34, 17, 7, 1, 23, 22, 50, 
    74, 65, 80, 68, 57, 65, 75, 76, 57, 52, 49, 54, 57, 57, 46, 
    71, 81, 78, 79, 75, 88, 84, 73, 72, 67, 73, 79, 79, 74, 58, 
    
    -- channel=91
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 6, 0, 
    31, 0, 0, 0, 6, 0, 0, 56, 3, 0, 1, 9, 17, 0, 4, 
    22, 12, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 1, 0, 7, 
    0, 22, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 1, 35, 30, 3, 75, 60, 99, 90, 14, 10, 0, 0, 
    0, 8, 0, 0, 125, 27, 11, 0, 0, 17, 0, 0, 13, 0, 0, 
    0, 22, 30, 0, 6, 118, 71, 92, 45, 7, 41, 9, 0, 54, 0, 
    6, 0, 10, 0, 0, 0, 0, 0, 7, 10, 4, 41, 24, 65, 12, 
    0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 42, 
    0, 24, 0, 7, 11, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    32, 6, 15, 3, 11, 14, 18, 2, 47, 8, 0, 18, 0, 0, 34, 
    19, 25, 12, 1, 0, 9, 30, 8, 44, 37, 0, 0, 0, 23, 0, 
    52, 0, 13, 1, 0, 14, 26, 0, 5, 50, 0, 38, 8, 0, 8, 
    29, 0, 7, 0, 12, 18, 20, 25, 0, 0, 19, 64, 6, 0, 1, 
    3, 0, 6, 5, 2, 20, 9, 0, 54, 0, 7, 90, 0, 2, 0, 
    0, 16, 0, 12, 21, 0, 63, 15, 35, 0, 39, 59, 0, 5, 0, 
    0, 0, 13, 21, 0, 10, 20, 22, 0, 1, 76, 51, 0, 0, 4, 
    37, 0, 24, 0, 0, 8, 37, 0, 1, 0, 100, 65, 0, 0, 66, 
    24, 0, 6, 74, 0, 0, 88, 3, 3, 39, 72, 21, 0, 0, 131, 
    34, 0, 0, 192, 0, 0, 66, 0, 100, 28, 6, 26, 0, 0, 141, 
    43, 0, 10, 114, 11, 0, 0, 0, 52, 43, 9, 0, 0, 0, 78, 
    12, 9, 0, 39, 42, 0, 10, 51, 37, 3, 10, 0, 0, 0, 0, 
    12, 0, 32, 0, 75, 38, 0, 44, 39, 20, 22, 0, 0, 0, 0, 
    35, 0, 39, 23, 27, 0, 0, 47, 0, 25, 7, 0, 17, 11, 0, 
    0, 6, 17, 1, 16, 8, 21, 7, 21, 13, 0, 0, 19, 30, 0, 
    
    -- channel=93
    112, 110, 121, 129, 131, 128, 124, 108, 89, 67, 81, 80, 81, 85, 82, 
    108, 113, 121, 130, 134, 139, 141, 139, 119, 66, 73, 87, 100, 99, 88, 
    97, 104, 123, 129, 132, 136, 142, 134, 135, 112, 111, 106, 105, 98, 97, 
    91, 104, 119, 127, 131, 145, 143, 129, 125, 135, 126, 105, 95, 97, 98, 
    81, 108, 124, 125, 134, 127, 114, 121, 113, 124, 116, 89, 80, 89, 94, 
    65, 114, 122, 120, 117, 91, 85, 75, 88, 98, 99, 67, 66, 81, 91, 
    73, 95, 109, 107, 100, 92, 95, 100, 94, 91, 84, 60, 58, 80, 85, 
    104, 92, 108, 94, 95, 111, 123, 102, 90, 91, 91, 56, 52, 89, 81, 
    128, 104, 107, 85, 82, 90, 114, 93, 86, 70, 55, 45, 51, 83, 79, 
    131, 97, 90, 82, 43, 86, 107, 125, 116, 58, 61, 71, 63, 83, 83, 
    133, 104, 83, 81, 53, 34, 67, 96, 76, 49, 37, 60, 74, 72, 83, 
    126, 125, 85, 115, 106, 110, 113, 89, 35, 24, 22, 22, 55, 70, 83, 
    134, 132, 106, 88, 102, 107, 124, 116, 83, 60, 48, 43, 52, 64, 74, 
    121, 114, 123, 99, 90, 113, 124, 133, 108, 103, 104, 107, 104, 100, 89, 
    130, 136, 135, 131, 123, 138, 128, 123, 118, 121, 126, 127, 125, 117, 104, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 14, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 11, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 8, 7, 7, 3, 31, 17, 26, 12, 6, 0, 0, 0, 0, 0, 
    3, 41, 27, 19, 16, 38, 36, 7, 7, 13, 0, 0, 0, 0, 0, 
    0, 36, 28, 28, 45, 33, 11, 46, 49, 45, 0, 0, 0, 2, 0, 
    0, 33, 30, 9, 57, 46, 9, 36, 42, 36, 12, 0, 0, 29, 0, 
    0, 34, 49, 0, 57, 42, 7, 15, 0, 0, 0, 0, 0, 45, 0, 
    0, 29, 46, 0, 0, 9, 5, 12, 0, 0, 0, 0, 0, 50, 22, 
    1, 5, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 43, 
    0, 8, 5, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 14, 2, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    26, 24, 50, 47, 51, 55, 49, 39, 13, 15, 16, 13, 13, 15, 7, 
    27, 36, 53, 49, 53, 57, 63, 62, 37, 13, 17, 21, 24, 22, 18, 
    19, 28, 49, 55, 51, 62, 62, 68, 49, 18, 19, 30, 32, 29, 24, 
    19, 28, 46, 49, 53, 69, 64, 59, 56, 57, 49, 33, 30, 29, 26, 
    24, 28, 43, 50, 58, 50, 40, 28, 43, 58, 43, 16, 23, 24, 26, 
    32, 34, 32, 40, 49, 6, 0, 1, 25, 29, 25, 10, 13, 22, 26, 
    10, 30, 17, 21, 20, 2, 15, 0, 0, 0, 4, 0, 2, 17, 23, 
    23, 20, 15, 17, 3, 10, 29, 0, 0, 0, 0, 0, 4, 5, 10, 
    35, 19, 6, 14, 0, 27, 22, 28, 19, 18, 9, 0, 5, 6, 0, 
    42, 17, 0, 0, 3, 17, 28, 15, 23, 7, 1, 0, 12, 0, 0, 
    37, 26, 0, 0, 1, 10, 34, 45, 27, 7, 0, 7, 14, 9, 0, 
    48, 29, 7, 5, 19, 11, 21, 11, 0, 0, 0, 0, 16, 26, 0, 
    53, 39, 23, 20, 22, 38, 38, 18, 0, 0, 0, 0, 0, 20, 7, 
    35, 46, 30, 34, 18, 29, 40, 39, 20, 12, 14, 9, 11, 17, 9, 
    39, 37, 43, 36, 31, 40, 47, 44, 43, 44, 43, 42, 38, 33, 28, 
    
    -- channel=96
    14, 36, 39, 47, 47, 39, 34, 32, 32, 54, 27, 6, 3, 0, 0, 
    39, 27, 35, 36, 34, 26, 19, 18, 11, 8, 0, 0, 0, 0, 0, 
    46, 54, 30, 24, 16, 9, 8, 4, 1, 0, 0, 17, 0, 0, 0, 
    7, 6, 6, 5, 2, 6, 0, 0, 0, 2, 42, 0, 0, 12, 9, 
    0, 7, 11, 13, 8, 4, 7, 9, 0, 0, 0, 0, 0, 0, 0, 
    6, 9, 9, 11, 5, 0, 0, 27, 114, 165, 0, 0, 7, 0, 0, 
    9, 13, 13, 3, 0, 88, 109, 97, 46, 0, 40, 14, 0, 0, 0, 
    15, 14, 0, 0, 13, 0, 5, 0, 0, 0, 96, 154, 14, 0, 0, 
    16, 4, 8, 41, 34, 9, 8, 0, 132, 152, 127, 98, 0, 0, 0, 
    8, 0, 18, 0, 15, 0, 12, 92, 115, 182, 199, 12, 0, 52, 91, 
    30, 168, 73, 0, 0, 0, 0, 91, 127, 141, 60, 148, 134, 116, 132, 
    34, 16, 0, 0, 0, 0, 27, 94, 99, 0, 0, 33, 77, 73, 0, 
    10, 6, 3, 0, 0, 0, 3, 101, 67, 0, 0, 0, 58, 69, 0, 
    0, 20, 62, 78, 104, 185, 209, 221, 148, 0, 37, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 
    
    -- channel=97
    201, 200, 200, 202, 187, 176, 170, 157, 141, 126, 109, 99, 55, 54, 83, 
    188, 174, 163, 160, 148, 138, 136, 130, 122, 115, 113, 70, 32, 74, 94, 
    134, 121, 126, 124, 122, 118, 119, 120, 119, 116, 94, 26, 53, 94, 97, 
    107, 114, 116, 116, 119, 121, 121, 123, 120, 110, 32, 42, 80, 105, 100, 
    108, 116, 117, 116, 119, 122, 113, 105, 101, 67, 27, 57, 81, 95, 101, 
    116, 115, 116, 114, 112, 103, 91, 64, 46, 6, 10, 0, 58, 57, 90, 
    118, 115, 110, 107, 99, 38, 0, 0, 7, 57, 26, 0, 24, 35, 59, 
    115, 112, 110, 74, 36, 44, 14, 21, 56, 55, 0, 0, 0, 37, 49, 
    112, 103, 56, 20, 0, 23, 55, 44, 5, 0, 0, 0, 42, 54, 33, 
    111, 102, 0, 15, 0, 39, 55, 0, 0, 0, 5, 0, 19, 0, 0, 
    118, 22, 0, 0, 13, 32, 57, 0, 0, 0, 16, 25, 0, 0, 0, 
    76, 23, 0, 0, 27, 26, 37, 0, 0, 12, 13, 52, 0, 0, 24, 
    62, 23, 0, 0, 31, 6, 21, 0, 0, 25, 2, 24, 21, 0, 38, 
    58, 35, 6, 0, 9, 0, 0, 0, 0, 22, 0, 3, 21, 12, 33, 
    54, 27, 10, 9, 15, 14, 15, 16, 20, 42, 4, 9, 29, 30, 35, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 15, 39, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 76, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 83, 77, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 51, 80, 95, 82, 9, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 78, 82, 81, 70, 35, 27, 42, 32, 
    0, 35, 21, 0, 0, 0, 0, 73, 71, 0, 0, 54, 65, 42, 0, 
    0, 0, 14, 0, 0, 0, 20, 75, 49, 0, 0, 0, 37, 11, 0, 
    0, 0, 11, 0, 0, 12, 43, 76, 39, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 16, 25, 29, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 13, 33, 41, 37, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 82, 110, 143, 183, 213, 23, 1, 1, 0, 
    0, 0, 0, 0, 18, 70, 103, 49, 39, 93, 236, 164, 0, 3, 0, 
    0, 0, 0, 16, 50, 42, 62, 76, 92, 168, 277, 179, 63, 0, 45, 
    0, 0, 8, 66, 45, 26, 82, 227, 275, 301, 261, 99, 54, 78, 153, 
    0, 109, 77, 45, 9, 8, 115, 251, 266, 216, 257, 213, 157, 185, 158, 
    25, 143, 151, 30, 0, 29, 113, 245, 203, 107, 47, 200, 227, 174, 77, 
    8, 63, 122, 21, 4, 68, 193, 252, 147, 30, 14, 53, 193, 86, 0, 
    0, 62, 120, 46, 73, 140, 189, 248, 132, 58, 50, 5, 112, 46, 0, 
    0, 47, 82, 63, 81, 126, 142, 148, 105, 67, 65, 0, 0, 0, 0, 
    5, 21, 24, 3, 0, 1, 0, 0, 0, 8, 38, 0, 0, 0, 0, 
    
    -- channel=100
    46, 78, 84, 95, 96, 84, 78, 80, 66, 83, 68, 50, 57, 38, 29, 
    79, 66, 68, 63, 59, 52, 47, 53, 44, 41, 27, 42, 44, 0, 23, 
    70, 73, 51, 42, 37, 28, 27, 33, 30, 26, 27, 54, 14, 0, 32, 
    30, 20, 20, 21, 19, 20, 17, 19, 22, 31, 86, 30, 21, 43, 41, 
    10, 15, 18, 22, 16, 21, 35, 31, 1, 0, 6, 0, 28, 33, 31, 
    14, 15, 20, 25, 18, 0, 0, 2, 68, 109, 0, 39, 41, 22, 27, 
    16, 16, 25, 19, 4, 73, 115, 121, 91, 0, 0, 61, 6, 43, 30, 
    17, 21, 7, 0, 49, 21, 41, 0, 0, 0, 27, 120, 53, 8, 0, 
    17, 12, 36, 50, 68, 52, 0, 0, 55, 72, 85, 107, 0, 0, 0, 
    5, 0, 50, 16, 62, 21, 0, 35, 47, 102, 111, 1, 0, 19, 70, 
    0, 100, 101, 33, 49, 0, 0, 37, 106, 151, 76, 71, 81, 92, 151, 
    31, 30, 23, 46, 1, 0, 0, 31, 127, 18, 25, 14, 53, 97, 35, 
    20, 20, 18, 26, 0, 0, 0, 46, 100, 0, 6, 20, 55, 107, 27, 
    11, 24, 65, 86, 92, 150, 168, 176, 159, 22, 61, 45, 59, 59, 20, 
    11, 26, 8, 0, 0, 0, 5, 13, 21, 22, 59, 60, 21, 20, 15, 
    
    -- channel=101
    0, 0, 13, 19, 27, 21, 23, 17, 13, 47, 14, 3, 10, 36, 1, 
    9, 2, 19, 23, 24, 18, 18, 12, 7, 2, 0, 0, 9, 0, 0, 
    39, 43, 24, 16, 11, 2, 1, 0, 0, 0, 0, 16, 0, 0, 0, 
    12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 23, 9, 0, 4, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 72, 125, 0, 0, 49, 0, 3, 
    0, 0, 1, 0, 0, 49, 61, 63, 48, 0, 0, 0, 0, 62, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 0, 0, 
    1, 0, 0, 37, 37, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 11, 0, 0, 0, 61, 127, 0, 0, 0, 2, 
    0, 127, 22, 0, 5, 0, 0, 0, 21, 71, 25, 124, 18, 36, 98, 
    9, 0, 8, 0, 0, 0, 0, 0, 26, 0, 0, 14, 18, 28, 1, 
    6, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 43, 12, 
    0, 13, 64, 63, 97, 158, 169, 174, 139, 5, 27, 0, 50, 24, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 42, 13, 0, 0, 0, 
    
    -- channel=102
    2, 0, 1, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 42, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 25, 0, 0, 22, 0, 
    0, 0, 0, 0, 1, 0, 2, 0, 0, 10, 0, 40, 7, 0, 0, 
    1, 0, 0, 0, 9, 8, 8, 8, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 48, 33, 7, 28, 0, 23, 0, 50, 0, 0, 
    0, 0, 0, 16, 44, 22, 0, 0, 0, 189, 98, 0, 0, 13, 0, 
    0, 0, 30, 0, 0, 32, 0, 25, 48, 116, 0, 0, 0, 26, 54, 
    0, 32, 0, 21, 0, 38, 131, 140, 8, 0, 0, 0, 32, 64, 25, 
    38, 143, 0, 31, 0, 66, 230, 39, 0, 0, 53, 0, 6, 0, 0, 
    137, 28, 0, 0, 0, 89, 200, 11, 0, 0, 54, 209, 0, 0, 0, 
    61, 15, 0, 0, 38, 98, 187, 0, 0, 17, 0, 162, 42, 0, 0, 
    44, 30, 28, 0, 102, 18, 95, 0, 0, 66, 0, 8, 108, 0, 24, 
    22, 33, 8, 0, 73, 42, 37, 20, 0, 99, 0, 0, 26, 0, 15, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 0, 0, 4, 22, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 69, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 35, 17, 0, 0, 108, 53, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 59, 92, 40, 0, 0, 
    0, 0, 0, 0, 24, 21, 39, 131, 175, 117, 63, 2, 38, 42, 79, 
    0, 0, 0, 18, 17, 13, 62, 68, 23, 28, 11, 14, 66, 112, 64, 
    0, 60, 68, 46, 28, 33, 52, 46, 51, 0, 0, 111, 101, 61, 9, 
    0, 0, 47, 42, 35, 90, 88, 55, 0, 0, 0, 0, 29, 13, 0, 
    0, 41, 69, 52, 68, 64, 76, 62, 38, 46, 52, 15, 45, 23, 26, 
    0, 43, 64, 85, 118, 134, 78, 53, 57, 67, 81, 34, 4, 20, 13, 
    0, 15, 10, 8, 0, 0, 0, 0, 0, 33, 28, 31, 6, 24, 34, 
    0, 36, 82, 91, 78, 80, 70, 60, 51, 28, 12, 33, 43, 43, 45, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 52, 73, 54, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 42, 97, 50, 0, 0, 141, 7, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 88, 120, 48, 27, 0, 0, 
    0, 0, 0, 23, 0, 26, 26, 156, 249, 252, 93, 0, 0, 32, 106, 
    0, 0, 0, 0, 0, 0, 74, 158, 66, 54, 36, 0, 65, 156, 94, 
    0, 148, 16, 22, 0, 9, 104, 71, 65, 0, 0, 112, 145, 70, 0, 
    0, 0, 0, 4, 0, 89, 150, 76, 0, 0, 0, 0, 11, 0, 0, 
    0, 23, 42, 0, 50, 77, 117, 83, 0, 33, 10, 21, 30, 0, 0, 
    0, 24, 47, 39, 145, 158, 143, 72, 0, 62, 43, 12, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 3, 
    0, 16, 49, 66, 47, 50, 39, 25, 13, 0, 0, 0, 10, 12, 23, 
    
    -- channel=106
    198, 200, 203, 204, 192, 171, 163, 150, 130, 102, 95, 75, 27, 10, 62, 
    187, 170, 166, 149, 134, 120, 118, 111, 100, 90, 83, 62, 0, 28, 76, 
    115, 111, 107, 104, 98, 94, 98, 98, 95, 91, 42, 7, 36, 63, 76, 
    81, 87, 90, 91, 95, 97, 103, 107, 103, 88, 21, 0, 58, 85, 80, 
    81, 90, 92, 91, 93, 94, 88, 96, 100, 92, 13, 21, 72, 74, 74, 
    89, 90, 90, 90, 81, 69, 52, 42, 29, 2, 0, 59, 0, 51, 65, 
    93, 91, 88, 73, 54, 26, 4, 0, 0, 0, 33, 30, 12, 0, 31, 
    90, 89, 65, 56, 23, 7, 4, 0, 39, 48, 42, 39, 0, 0, 6, 
    87, 67, 40, 0, 0, 0, 0, 24, 49, 40, 53, 39, 13, 13, 32, 
    69, 44, 31, 0, 0, 0, 0, 25, 21, 33, 0, 14, 28, 23, 27, 
    46, 16, 0, 0, 0, 0, 0, 20, 29, 0, 0, 0, 9, 9, 3, 
    37, 0, 0, 0, 0, 0, 0, 28, 33, 0, 0, 0, 0, 13, 0, 
    17, 0, 0, 0, 0, 5, 25, 23, 23, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    0, 0, 7, 14, 12, 12, 15, 2, 15, 60, 5, 0, 11, 42, 0, 
    2, 0, 14, 13, 11, 8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 42, 17, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 44, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 66, 83, 0, 0, 53, 0, 0, 
    0, 0, 0, 0, 0, 93, 104, 121, 69, 0, 10, 0, 0, 61, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 
    0, 0, 4, 34, 42, 50, 0, 0, 22, 17, 17, 0, 0, 0, 0, 
    0, 0, 0, 15, 12, 19, 13, 29, 2, 110, 103, 0, 0, 0, 35, 
    0, 176, 0, 5, 0, 0, 0, 5, 64, 89, 128, 154, 35, 60, 115, 
    8, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 99, 14, 39, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 9, 100, 26, 21, 
    0, 14, 83, 67, 158, 221, 233, 235, 103, 30, 32, 2, 89, 10, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 35, 0, 0, 0, 0, 
    
    -- channel=108
    24, 37, 19, 29, 36, 32, 18, 38, 26, 0, 22, 14, 54, 0, 26, 
    15, 33, 43, 34, 27, 27, 19, 25, 22, 22, 0, 56, 24, 0, 25, 
    28, 33, 25, 26, 16, 18, 18, 15, 16, 6, 0, 25, 16, 0, 35, 
    14, 14, 16, 20, 15, 15, 5, 14, 12, 21, 51, 0, 20, 23, 22, 
    14, 19, 19, 22, 8, 7, 0, 0, 0, 46, 42, 12, 26, 25, 16, 
    16, 20, 23, 21, 0, 0, 0, 13, 19, 0, 0, 243, 0, 42, 23, 
    17, 23, 33, 0, 0, 4, 25, 56, 0, 0, 0, 214, 84, 0, 14, 
    19, 26, 0, 30, 15, 0, 6, 0, 0, 0, 0, 170, 100, 0, 0, 
    26, 0, 41, 0, 53, 0, 0, 0, 0, 0, 80, 171, 0, 0, 0, 
    0, 0, 183, 0, 79, 0, 0, 0, 0, 88, 0, 49, 0, 5, 73, 
    0, 0, 88, 50, 36, 0, 0, 0, 138, 82, 12, 0, 50, 65, 109, 
    0, 12, 0, 85, 0, 0, 0, 0, 197, 0, 19, 0, 0, 145, 11, 
    0, 0, 0, 67, 0, 0, 0, 0, 205, 0, 57, 42, 0, 126, 0, 
    0, 0, 0, 43, 0, 0, 0, 12, 62, 0, 19, 64, 0, 24, 0, 
    0, 10, 0, 28, 0, 0, 6, 10, 11, 0, 35, 43, 0, 0, 0, 
    
    -- channel=109
    288, 274, 275, 269, 258, 240, 234, 219, 199, 163, 162, 141, 65, 61, 139, 
    259, 243, 242, 237, 224, 207, 205, 191, 181, 173, 154, 104, 49, 95, 159, 
    186, 192, 199, 199, 190, 189, 193, 184, 182, 173, 93, 44, 81, 134, 155, 
    172, 184, 186, 187, 191, 196, 199, 193, 181, 155, 45, 37, 137, 160, 162, 
    181, 192, 192, 192, 193, 183, 156, 166, 159, 134, 45, 51, 132, 151, 152, 
    192, 194, 190, 187, 173, 140, 92, 63, 34, 19, 46, 52, 24, 119, 140, 
    194, 194, 189, 167, 119, 49, 18, 4, 20, 6, 28, 69, 16, 31, 95, 
    192, 191, 149, 110, 55, 43, 32, 48, 69, 43, 30, 32, 48, 23, 65, 
    192, 162, 62, 14, 10, 0, 0, 36, 27, 31, 45, 62, 80, 57, 47, 
    173, 117, 36, 8, 13, 1, 0, 18, 17, 6, 2, 63, 42, 28, 29, 
    132, 7, 13, 13, 10, 9, 0, 15, 17, 1, 0, 0, 12, 10, 12, 
    113, 14, 13, 17, 8, 0, 0, 19, 32, 15, 17, 0, 10, 18, 29, 
    87, 17, 4, 13, 8, 27, 16, 16, 32, 11, 32, 10, 0, 11, 30, 
    88, 32, 0, 0, 0, 0, 0, 0, 0, 7, 14, 13, 0, 6, 17, 
    83, 39, 8, 12, 0, 4, 8, 12, 14, 3, 9, 12, 12, 12, 11, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 28, 68, 98, 82, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 31, 51, 25, 22, 62, 124, 13, 0, 0, 0, 
    0, 0, 0, 0, 1, 10, 16, 8, 5, 65, 128, 61, 0, 0, 0, 
    0, 0, 0, 32, 13, 19, 50, 116, 136, 147, 114, 0, 1, 7, 63, 
    0, 20, 0, 21, 0, 6, 83, 130, 127, 109, 149, 62, 55, 81, 64, 
    0, 96, 50, 4, 0, 10, 69, 122, 87, 46, 39, 149, 107, 79, 31, 
    0, 18, 56, 0, 0, 41, 112, 120, 34, 7, 0, 52, 99, 19, 0, 
    0, 26, 63, 0, 31, 49, 98, 118, 18, 28, 0, 0, 79, 1, 0, 
    0, 17, 50, 36, 69, 97, 106, 107, 52, 41, 24, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 15, 0, 0, 0, 0, 
    
    -- channel=111
    196, 203, 214, 217, 207, 191, 182, 169, 149, 116, 107, 80, 6, 36, 75, 
    202, 184, 189, 186, 169, 152, 148, 136, 125, 110, 92, 31, 0, 44, 88, 
    143, 146, 147, 140, 131, 124, 124, 117, 111, 111, 5, 0, 16, 64, 86, 
    116, 119, 120, 118, 123, 126, 120, 112, 104, 82, 0, 3, 74, 94, 98, 
    113, 123, 125, 121, 124, 102, 89, 95, 73, 12, 0, 10, 71, 94, 94, 
    122, 123, 122, 117, 109, 46, 0, 0, 0, 0, 0, 0, 0, 51, 85, 
    123, 123, 115, 106, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 
    123, 120, 73, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    121, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    9, 9, 11, 27, 18, 5, 7, 9, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 4, 20, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 7, 15, 8, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 16, 17, 9, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 61, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 19, 17, 
    73, 74, 51, 0, 0, 19, 5, 0, 0, 0, 0, 0, 0, 26, 35, 
    42, 38, 47, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 29, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 
    7, 60, 158, 125, 81, 58, 21, 7, 0, 0, 0, 0, 0, 0, 0, 
    138, 151, 164, 94, 59, 67, 14, 21, 0, 0, 0, 0, 0, 0, 0, 
    219, 188, 81, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 63, 46, 24, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    20, 13, 35, 54, 38, 0, 0, 0, 0, 6, 35, 0, 0, 1, 7, 
    34, 44, 17, 0, 0, 3, 0, 2, 0, 0, 0, 8, 0, 0, 0, 
    
    -- channel=113
    26, 26, 30, 26, 44, 49, 40, 31, 27, 29, 28, 25, 27, 30, 28, 
    25, 24, 29, 40, 54, 75, 64, 60, 42, 34, 39, 41, 43, 42, 38, 
    26, 25, 28, 44, 63, 83, 90, 95, 78, 53, 46, 47, 44, 36, 34, 
    30, 30, 20, 59, 75, 86, 95, 103, 98, 76, 61, 51, 41, 37, 46, 
    42, 46, 25, 48, 81, 84, 83, 90, 106, 103, 101, 79, 61, 57, 63, 
    37, 31, 0, 44, 62, 89, 78, 80, 96, 102, 105, 96, 81, 66, 58, 
    25, 23, 22, 11, 65, 75, 70, 89, 90, 85, 93, 108, 82, 61, 39, 
    31, 36, 35, 41, 23, 77, 72, 96, 91, 75, 90, 98, 81, 61, 49, 
    39, 38, 36, 55, 41, 42, 62, 85, 89, 74, 86, 91, 91, 72, 51, 
    45, 39, 26, 0, 55, 28, 77, 75, 88, 79, 85, 88, 88, 60, 59, 
    17, 8, 0, 35, 61, 63, 80, 76, 88, 85, 79, 84, 85, 67, 63, 
    0, 0, 12, 29, 48, 77, 76, 52, 73, 83, 82, 75, 78, 82, 58, 
    21, 23, 28, 40, 40, 58, 73, 61, 80, 89, 69, 76, 74, 82, 71, 
    36, 45, 47, 45, 53, 60, 65, 67, 77, 77, 65, 70, 77, 76, 80, 
    43, 45, 56, 65, 75, 69, 67, 68, 74, 72, 75, 70, 69, 78, 72, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 20, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 18, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 20, 35, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 64, 76, 51, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    93, 92, 25, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 50, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=115
    77, 70, 77, 77, 65, 64, 57, 61, 50, 42, 36, 25, 14, 11, 6, 
    75, 68, 66, 50, 39, 34, 45, 32, 38, 39, 30, 29, 28, 34, 34, 
    67, 66, 44, 32, 11, 0, 0, 3, 37, 64, 61, 63, 57, 55, 43, 
    58, 61, 47, 0, 0, 0, 0, 0, 7, 48, 66, 57, 63, 50, 34, 
    92, 112, 99, 10, 0, 26, 30, 0, 0, 0, 15, 38, 58, 55, 44, 
    155, 165, 141, 10, 15, 25, 36, 17, 6, 0, 0, 10, 42, 66, 58, 
    157, 157, 152, 65, 12, 42, 38, 18, 28, 11, 0, 0, 30, 57, 53, 
    144, 151, 146, 127, 71, 20, 30, 15, 44, 35, 0, 0, 19, 33, 46, 
    157, 183, 198, 130, 156, 99, 80, 23, 41, 42, 14, 0, 10, 24, 29, 
    228, 259, 253, 225, 141, 126, 68, 40, 36, 44, 33, 5, 2, 9, 1, 
    301, 284, 165, 112, 68, 62, 32, 29, 36, 38, 32, 9, 0, 25, 0, 
    240, 207, 139, 94, 28, 0, 35, 14, 8, 20, 35, 26, 0, 27, 22, 
    117, 108, 102, 88, 71, 31, 29, 31, 9, 36, 65, 35, 13, 7, 34, 
    75, 73, 66, 51, 40, 38, 18, 18, 11, 23, 55, 34, 6, 4, 13, 
    51, 37, 22, 1, 3, 34, 24, 10, 0, 0, 4, 15, 9, 0, 0, 
    
    -- channel=116
    53, 55, 48, 57, 79, 87, 72, 62, 50, 52, 54, 51, 45, 32, 28, 
    54, 54, 52, 67, 88, 111, 117, 95, 66, 47, 37, 23, 13, 8, 18, 
    59, 57, 65, 78, 111, 116, 129, 126, 75, 34, 42, 46, 47, 53, 59, 
    54, 47, 39, 53, 117, 108, 104, 113, 128, 114, 92, 88, 51, 44, 44, 
    0, 0, 38, 85, 99, 90, 91, 117, 131, 135, 134, 113, 55, 41, 38, 
    39, 60, 93, 62, 78, 69, 124, 135, 115, 123, 135, 128, 77, 59, 55, 
    73, 73, 64, 54, 58, 110, 138, 127, 108, 113, 131, 123, 107, 76, 75, 
    59, 47, 60, 65, 45, 12, 81, 106, 114, 122, 132, 131, 118, 80, 46, 
    44, 30, 4, 23, 67, 63, 70, 110, 126, 128, 125, 133, 113, 84, 83, 
    0, 8, 85, 141, 116, 127, 90, 134, 123, 123, 122, 139, 122, 90, 45, 
    67, 92, 169, 157, 149, 175, 137, 127, 126, 129, 134, 136, 104, 56, 39, 
    170, 167, 95, 77, 101, 121, 82, 82, 114, 117, 97, 110, 95, 59, 61, 
    97, 88, 75, 56, 59, 50, 91, 106, 94, 94, 98, 122, 104, 64, 63, 
    62, 53, 80, 100, 85, 60, 63, 82, 98, 109, 136, 128, 111, 75, 62, 
    75, 90, 76, 57, 44, 56, 70, 73, 63, 66, 75, 89, 86, 58, 58, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 34, 6, 0, 0, 0, 0, 0, 0, 13, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    0, 0, 2, 10, 20, 21, 0, 0, 0, 0, 0, 0, 0, 2, 2, 
    0, 0, 1, 48, 27, 51, 10, 28, 0, 0, 0, 0, 0, 0, 0, 
    88, 80, 8, 2, 0, 5, 0, 0, 4, 0, 0, 0, 0, 5, 0, 
    24, 18, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 10, 35, 22, 0, 0, 5, 1, 16, 43, 0, 6, 10, 5, 
    20, 35, 18, 0, 0, 0, 0, 5, 0, 0, 3, 23, 17, 4, 5, 
    
    -- channel=118
    0, 0, 18, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 8, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 6, 9, 15, 30, 4, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 7, 9, 11, 13, 17, 25, 8, 0, 0, 0, 0, 
    17, 14, 0, 0, 11, 55, 5, 0, 3, 10, 23, 5, 7, 0, 0, 
    12, 0, 0, 0, 1, 60, 0, 0, 7, 0, 0, 30, 27, 0, 0, 
    0, 0, 0, 0, 8, 54, 0, 4, 17, 0, 0, 37, 8, 14, 0, 
    7, 6, 0, 0, 0, 25, 0, 19, 25, 0, 0, 7, 11, 9, 0, 
    18, 28, 0, 0, 0, 0, 4, 0, 23, 0, 0, 0, 26, 1, 0, 
    19, 14, 0, 0, 0, 0, 16, 0, 19, 1, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 3, 15, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 43, 0, 27, 26, 9, 0, 0, 35, 0, 
    0, 0, 0, 0, 0, 0, 28, 0, 16, 57, 0, 0, 0, 8, 6, 
    0, 3, 0, 0, 0, 0, 0, 0, 7, 36, 20, 0, 0, 0, 19, 
    0, 0, 0, 0, 26, 15, 0, 0, 0, 0, 18, 7, 0, 3, 0, 
    
    -- channel=119
    28, 25, 23, 14, 0, 0, 5, 18, 25, 21, 22, 25, 28, 33, 40, 
    28, 27, 17, 12, 0, 0, 0, 0, 7, 23, 28, 38, 42, 42, 37, 
    21, 22, 6, 0, 0, 0, 0, 0, 0, 27, 17, 11, 7, 5, 0, 
    22, 28, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 4, 
    63, 67, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 10, 17, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 20, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 20, 5, 9, 42, 23, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    18, 31, 63, 41, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 3, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    32, 26, 31, 18, 16, 31, 23, 19, 23, 18, 11, 8, 10, 19, 24, 
    31, 28, 27, 10, 18, 7, 15, 23, 16, 27, 38, 50, 56, 55, 42, 
    23, 23, 0, 9, 7, 20, 13, 18, 47, 59, 47, 36, 20, 7, 0, 
    29, 38, 39, 28, 22, 36, 39, 26, 14, 9, 23, 8, 19, 16, 16, 
    105, 118, 59, 11, 26, 48, 61, 32, 23, 20, 15, 22, 29, 27, 28, 
    70, 51, 17, 20, 49, 72, 27, 24, 37, 28, 23, 26, 19, 11, 8, 
    30, 29, 39, 44, 11, 6, 14, 29, 47, 35, 22, 30, 11, 0, 0, 
    53, 63, 43, 36, 72, 82, 40, 38, 51, 37, 26, 28, 21, 18, 21, 
    74, 101, 139, 97, 75, 48, 42, 33, 40, 36, 40, 32, 36, 11, 0, 
    160, 129, 32, 8, 12, 3, 24, 20, 46, 43, 42, 30, 27, 0, 0, 
    77, 40, 0, 0, 0, 0, 1, 0, 30, 26, 17, 25, 22, 22, 0, 
    0, 0, 5, 27, 8, 15, 47, 20, 17, 34, 50, 37, 6, 6, 0, 
    0, 2, 10, 27, 25, 34, 13, 17, 41, 62, 58, 25, 17, 0, 1, 
    20, 26, 0, 0, 0, 10, 24, 9, 7, 1, 0, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    11, 12, 11, 15, 32, 37, 31, 11, 8, 8, 2, 0, 0, 0, 0, 
    10, 11, 12, 21, 42, 53, 50, 46, 18, 13, 18, 17, 16, 16, 16, 
    10, 8, 15, 12, 49, 62, 74, 76, 44, 31, 35, 35, 28, 22, 20, 
    11, 13, 18, 38, 52, 66, 75, 89, 85, 53, 45, 48, 24, 24, 28, 
    30, 39, 51, 41, 53, 50, 72, 91, 93, 90, 80, 63, 46, 49, 51, 
    46, 48, 44, 42, 44, 64, 79, 75, 81, 95, 94, 77, 63, 58, 52, 
    38, 39, 38, 44, 40, 46, 69, 78, 74, 81, 89, 81, 68, 43, 32, 
    39, 45, 54, 44, 57, 55, 77, 83, 75, 78, 87, 84, 62, 47, 33, 
    51, 58, 70, 95, 65, 70, 57, 93, 74, 74, 83, 85, 68, 55, 43, 
    75, 81, 81, 62, 76, 68, 71, 86, 75, 74, 82, 88, 71, 51, 32, 
    77, 78, 77, 59, 59, 66, 63, 64, 77, 77, 80, 82, 70, 48, 49, 
    47, 35, 23, 40, 58, 58, 47, 52, 54, 64, 67, 79, 72, 54, 52, 
    22, 22, 26, 33, 34, 44, 55, 49, 56, 61, 67, 78, 72, 61, 48, 
    25, 31, 41, 40, 36, 40, 50, 56, 56, 55, 48, 63, 71, 57, 53, 
    32, 34, 37, 42, 43, 46, 52, 55, 53, 49, 51, 54, 53, 53, 46, 
    
    -- channel=123
    0, 0, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 9, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 21, 12, 2, 0, 8, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    17, 11, 0, 0, 18, 40, 0, 0, 0, 0, 0, 0, 0, 13, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 33, 
    0, 0, 38, 0, 47, 0, 13, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 12, 58, 82, 56, 55, 24, 25, 0, 0, 0, 0, 0, 0, 0, 
    134, 122, 0, 0, 0, 15, 0, 0, 21, 0, 0, 0, 0, 4, 0, 
    39, 39, 15, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 51, 33, 0, 0, 5, 5, 40, 48, 0, 7, 3, 14, 
    32, 49, 21, 0, 1, 0, 0, 1, 0, 0, 19, 32, 11, 3, 2, 
    
    -- channel=124
    0, 7, 0, 3, 0, 0, 18, 0, 9, 6, 8, 13, 8, 0, 5, 
    0, 8, 0, 0, 4, 0, 0, 8, 7, 0, 0, 0, 0, 0, 9, 
    0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 2, 5, 10, 15, 19, 
    0, 0, 26, 6, 0, 0, 0, 0, 0, 0, 0, 19, 1, 12, 8, 
    0, 0, 64, 55, 0, 0, 0, 22, 0, 0, 0, 0, 0, 7, 7, 
    0, 0, 49, 62, 0, 0, 5, 12, 0, 0, 1, 0, 0, 1, 16, 
    0, 0, 0, 125, 0, 0, 11, 0, 0, 9, 3, 0, 7, 0, 27, 
    0, 0, 16, 0, 78, 0, 15, 0, 0, 14, 8, 0, 0, 0, 3, 
    0, 0, 0, 76, 1, 79, 0, 26, 0, 0, 3, 6, 0, 13, 38, 
    0, 0, 33, 89, 0, 37, 0, 38, 0, 0, 0, 17, 0, 38, 11, 
    0, 37, 155, 0, 10, 0, 3, 0, 0, 0, 2, 6, 3, 0, 32, 
    53, 22, 42, 14, 53, 0, 0, 58, 0, 0, 0, 8, 27, 0, 50, 
    11, 4, 0, 0, 15, 29, 0, 9, 0, 0, 0, 8, 36, 7, 0, 
    0, 0, 18, 27, 0, 0, 4, 0, 0, 0, 0, 1, 17, 10, 0, 
    25, 18, 3, 14, 0, 0, 20, 21, 10, 2, 0, 0, 15, 9, 8, 
    
    -- channel=125
    11, 11, 16, 19, 19, 19, 20, 17, 15, 14, 13, 13, 13, 18, 21, 
    10, 12, 16, 15, 20, 11, 18, 19, 20, 23, 29, 35, 36, 40, 40, 
    8, 10, 16, 11, 11, 12, 13, 21, 26, 38, 36, 42, 39, 37, 38, 
    12, 15, 37, 20, 0, 9, 17, 27, 30, 20, 28, 36, 43, 43, 50, 
    36, 42, 50, 24, 0, 7, 19, 24, 26, 24, 22, 27, 53, 71, 71, 
    39, 34, 38, 22, 16, 14, 7, 9, 19, 25, 23, 12, 47, 76, 69, 
    26, 30, 36, 51, 21, 4, 10, 13, 15, 19, 21, 10, 33, 49, 44, 
    30, 40, 44, 44, 62, 38, 38, 24, 10, 12, 16, 10, 15, 32, 52, 
    39, 51, 68, 58, 56, 62, 51, 33, 1, 4, 12, 8, 6, 29, 61, 
    66, 65, 43, 47, 26, 46, 36, 31, 1, 2, 12, 7, 2, 40, 73, 
    53, 52, 31, 14, 0, 10, 8, 14, 11, 7, 17, 11, 18, 62, 77, 
    10, 9, 25, 25, 19, 0, 10, 27, 2, 1, 15, 21, 40, 65, 80, 
    13, 15, 27, 37, 39, 35, 24, 22, 7, 0, 11, 12, 45, 69, 71, 
    28, 36, 37, 43, 53, 59, 42, 36, 24, 7, 0, 5, 27, 69, 71, 
    38, 47, 58, 68, 71, 67, 58, 69, 71, 58, 43, 43, 57, 76, 79, 
    
    -- channel=126
    33, 28, 35, 33, 31, 29, 21, 25, 15, 13, 10, 5, 0, 0, 0, 
    32, 26, 29, 20, 17, 23, 22, 14, 11, 10, 1, 0, 0, 0, 0, 
    30, 28, 14, 18, 7, 0, 1, 2, 12, 17, 17, 16, 14, 15, 8, 
    24, 24, 0, 0, 1, 0, 0, 0, 3, 29, 31, 19, 15, 8, 0, 
    28, 36, 20, 0, 0, 17, 8, 0, 0, 0, 13, 17, 14, 4, 0, 
    67, 74, 48, 0, 0, 17, 17, 5, 0, 0, 0, 10, 12, 12, 6, 
    74, 72, 62, 0, 0, 31, 18, 9, 12, 0, 0, 2, 8, 18, 11, 
    66, 64, 59, 51, 0, 0, 0, 4, 23, 12, 0, 0, 9, 11, 3, 
    69, 78, 69, 27, 59, 16, 26, 1, 26, 20, 2, 0, 8, 2, 0, 
    87, 108, 118, 91, 76, 48, 34, 9, 21, 23, 13, 0, 3, 0, 0, 
    139, 127, 65, 63, 45, 41, 22, 15, 20, 20, 14, 0, 0, 0, 0, 
    132, 111, 54, 35, 0, 0, 14, 0, 11, 14, 13, 4, 0, 1, 0, 
    57, 54, 45, 33, 15, 0, 16, 7, 8, 24, 26, 16, 0, 0, 0, 
    29, 25, 26, 17, 9, 3, 0, 0, 0, 14, 38, 15, 0, 0, 0, 
    15, 9, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 12, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 20, 8, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 27, 20, 
    0, 0, 10, 16, 20, 1, 0, 21, 19, 6, 0, 4, 17, 33, 26, 
    
    -- channel=128
    0, 0, 40, 55, 37, 47, 42, 37, 14, 6, 15, 31, 51, 54, 57, 
    0, 0, 36, 76, 33, 43, 67, 61, 74, 57, 0, 62, 65, 66, 70, 
    0, 0, 0, 45, 73, 70, 69, 88, 107, 49, 17, 91, 82, 70, 65, 
    0, 0, 0, 76, 93, 76, 8, 17, 21, 46, 86, 77, 102, 117, 114, 
    33, 3, 60, 73, 49, 101, 88, 72, 37, 57, 81, 78, 113, 106, 87, 
    80, 81, 88, 64, 61, 103, 98, 60, 10, 36, 76, 93, 114, 82, 63, 
    82, 83, 107, 60, 65, 71, 63, 60, 51, 54, 70, 89, 121, 90, 60, 
    88, 90, 75, 57, 80, 83, 84, 50, 88, 79, 92, 162, 148, 132, 108, 
    77, 72, 54, 65, 90, 52, 57, 59, 64, 83, 54, 35, 101, 149, 114, 
    75, 57, 76, 91, 102, 135, 123, 69, 13, 43, 84, 56, 29, 48, 86, 
    91, 84, 83, 82, 82, 92, 92, 116, 98, 80, 68, 36, 58, 73, 57, 
    98, 85, 75, 107, 110, 117, 63, 89, 90, 81, 28, 71, 64, 63, 49, 
    92, 87, 84, 104, 109, 119, 87, 106, 104, 72, 49, 70, 83, 80, 45, 
    94, 76, 77, 94, 84, 30, 90, 88, 81, 65, 39, 52, 53, 41, 46, 
    105, 60, 73, 98, 97, 86, 99, 70, 59, 25, 46, 41, 36, 29, 63, 
    
    -- channel=129
    25, 87, 73, 66, 60, 74, 74, 77, 44, 30, 75, 69, 78, 81, 80, 
    26, 64, 70, 63, 34, 46, 55, 60, 50, 16, 93, 55, 63, 69, 71, 
    26, 40, 80, 66, 38, 0, 31, 50, 34, 39, 58, 47, 45, 51, 52, 
    32, 70, 85, 43, 42, 9, 27, 26, 38, 62, 31, 55, 34, 27, 46, 
    45, 67, 50, 25, 54, 22, 18, 11, 34, 47, 47, 56, 36, 35, 65, 
    47, 52, 44, 42, 47, 24, 10, 23, 30, 42, 41, 56, 37, 34, 61, 
    53, 54, 42, 47, 27, 29, 14, 35, 23, 29, 44, 56, 44, 37, 48, 
    50, 54, 27, 67, 29, 22, 15, 28, 31, 50, 34, 63, 53, 35, 49, 
    35, 52, 37, 62, 24, 24, 20, 2, 66, 40, 40, 39, 72, 39, 70, 
    42, 54, 43, 31, 35, 25, 17, 19, 30, 53, 36, 53, 60, 48, 58, 
    43, 34, 44, 38, 37, 18, 42, 34, 21, 33, 50, 56, 46, 36, 49, 
    47, 29, 56, 30, 26, 26, 50, 39, 33, 27, 65, 44, 44, 41, 40, 
    45, 46, 59, 28, 5, 46, 49, 42, 33, 37, 56, 43, 43, 41, 43, 
    45, 50, 66, 34, 22, 54, 44, 44, 42, 47, 52, 45, 39, 56, 49, 
    45, 50, 64, 35, 26, 33, 36, 48, 36, 59, 49, 49, 44, 55, 47, 
    
    -- channel=130
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 25, 7, 7, 4, 14, 0, 0, 25, 18, 12, 9, 
    0, 0, 0, 0, 43, 31, 0, 7, 11, 3, 18, 38, 43, 41, 33, 
    0, 0, 0, 4, 33, 49, 4, 0, 0, 1, 41, 42, 62, 54, 41, 
    14, 0, 23, 4, 19, 50, 41, 11, 0, 3, 36, 43, 63, 35, 16, 
    28, 24, 28, 6, 25, 42, 31, 8, 5, 6, 28, 54, 64, 38, 10, 
    23, 18, 13, 18, 21, 34, 35, 14, 27, 18, 28, 46, 63, 59, 26, 
    26, 16, 6, 30, 42, 30, 43, 9, 21, 14, 19, 32, 44, 62, 40, 
    25, 11, 29, 26, 51, 48, 40, 34, 0, 1, 19, 0, 10, 35, 27, 
    35, 15, 34, 38, 43, 59, 58, 42, 1, 13, 10, 0, 0, 5, 0, 
    42, 28, 37, 41, 46, 31, 33, 44, 45, 13, 0, 2, 10, 9, 0, 
    39, 31, 30, 58, 52, 36, 25, 32, 31, 6, 0, 7, 17, 5, 0, 
    34, 23, 19, 52, 44, 5, 34, 24, 21, 0, 0, 1, 7, 1, 0, 
    29, 10, 6, 51, 45, 3, 14, 6, 2, 0, 0, 0, 0, 0, 1, 
    16, 5, 0, 45, 45, 30, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=131
    0, 20, 127, 123, 111, 110, 113, 121, 126, 54, 103, 147, 144, 141, 137, 
    0, 2, 108, 137, 173, 125, 144, 160, 165, 113, 129, 187, 171, 163, 158, 
    0, 0, 80, 122, 216, 169, 105, 122, 139, 142, 167, 205, 208, 203, 194, 
    29, 41, 108, 134, 210, 211, 142, 103, 99, 141, 211, 229, 251, 229, 225, 
    165, 152, 186, 131, 172, 214, 192, 132, 114, 141, 198, 239, 253, 199, 181, 
    194, 190, 192, 155, 182, 202, 182, 130, 133, 148, 183, 243, 259, 207, 159, 
    187, 183, 154, 184, 169, 179, 165, 152, 169, 167, 183, 241, 263, 253, 188, 
    183, 181, 147, 186, 198, 197, 188, 152, 183, 156, 184, 175, 265, 250, 233, 
    181, 156, 176, 179, 234, 225, 198, 164, 118, 153, 164, 111, 130, 194, 210, 
    202, 171, 202, 205, 208, 228, 245, 211, 138, 152, 141, 131, 129, 135, 141, 
    219, 185, 213, 214, 218, 189, 192, 214, 207, 143, 132, 134, 154, 138, 117, 
    213, 191, 202, 237, 227, 192, 192, 200, 189, 133, 120, 144, 165, 141, 120, 
    202, 178, 192, 234, 196, 139, 190, 182, 165, 119, 125, 131, 133, 137, 120, 
    193, 158, 165, 231, 199, 152, 158, 145, 124, 98, 110, 117, 104, 107, 132, 
    168, 152, 134, 230, 213, 177, 129, 119, 93, 86, 104, 115, 107, 101, 124, 
    
    -- channel=132
    21, 0, 64, 71, 60, 70, 69, 62, 47, 46, 8, 39, 60, 68, 72, 
    21, 9, 63, 63, 23, 46, 64, 61, 70, 81, 0, 64, 69, 71, 74, 
    21, 19, 26, 46, 25, 67, 70, 85, 108, 49, 17, 81, 72, 61, 62, 
    0, 0, 0, 87, 45, 50, 15, 36, 32, 15, 70, 46, 53, 92, 93, 
    61, 16, 70, 98, 20, 58, 63, 76, 40, 31, 56, 61, 86, 123, 100, 
    87, 77, 98, 78, 33, 60, 84, 58, 19, 17, 52, 71, 97, 117, 107, 
    101, 86, 109, 71, 63, 47, 56, 25, 43, 40, 44, 64, 96, 89, 85, 
    110, 88, 83, 26, 55, 60, 56, 34, 71, 53, 83, 117, 121, 118, 104, 
    118, 83, 40, 21, 58, 24, 28, 61, 41, 80, 59, 72, 87, 146, 100, 
    103, 65, 56, 66, 73, 88, 74, 44, 30, 39, 85, 67, 34, 57, 88, 
    99, 98, 63, 56, 57, 84, 64, 72, 77, 82, 76, 39, 51, 75, 63, 
    102, 114, 53, 63, 72, 77, 46, 59, 72, 94, 36, 67, 56, 65, 66, 
    105, 122, 79, 71, 97, 67, 65, 85, 97, 83, 57, 70, 76, 81, 59, 
    111, 125, 92, 67, 73, 9, 78, 89, 90, 79, 54, 63, 70, 50, 53, 
    127, 115, 94, 67, 75, 79, 100, 79, 85, 50, 62, 56, 56, 42, 69, 
    
    -- channel=133
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 2, 34, 47, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 75, 26, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 56, 13, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 14, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 17, 14, 3, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    0, 177, 52, 0, 0, 13, 0, 5, 0, 0, 148, 4, 0, 0, 0, 
    0, 104, 105, 33, 0, 0, 16, 20, 0, 0, 181, 0, 0, 0, 0, 
    0, 33, 163, 33, 54, 0, 0, 31, 0, 23, 62, 19, 0, 0, 0, 
    0, 67, 98, 0, 93, 0, 0, 0, 4, 105, 0, 73, 0, 0, 27, 
    0, 51, 0, 0, 98, 0, 0, 0, 16, 70, 35, 69, 0, 0, 38, 
    0, 4, 0, 0, 49, 0, 0, 0, 3, 54, 31, 86, 0, 0, 0, 
    0, 0, 0, 31, 0, 10, 0, 35, 0, 28, 27, 80, 0, 0, 0, 
    0, 8, 0, 116, 0, 0, 0, 0, 30, 4, 0, 58, 76, 0, 8, 
    0, 8, 0, 48, 0, 0, 0, 0, 59, 0, 0, 0, 86, 0, 92, 
    0, 0, 5, 0, 6, 0, 0, 0, 0, 29, 0, 4, 15, 0, 38, 
    0, 0, 42, 0, 0, 0, 44, 8, 0, 0, 4, 14, 4, 0, 0, 
    0, 0, 74, 0, 0, 0, 17, 0, 0, 0, 56, 0, 12, 0, 0, 
    0, 0, 62, 0, 0, 6, 27, 0, 0, 0, 37, 0, 0, 0, 0, 
    0, 0, 67, 15, 0, 4, 0, 0, 0, 0, 19, 0, 0, 40, 4, 
    0, 0, 39, 53, 0, 0, 0, 0, 0, 39, 4, 3, 0, 14, 6, 
    
    -- channel=135
    41, 0, 0, 0, 0, 0, 0, 0, 6, 10, 6, 0, 0, 0, 0, 
    40, 7, 0, 0, 33, 0, 0, 0, 0, 6, 24, 0, 0, 0, 0, 
    37, 22, 0, 0, 20, 18, 0, 0, 0, 11, 13, 0, 0, 0, 0, 
    91, 94, 33, 0, 0, 32, 49, 19, 12, 6, 0, 2, 9, 0, 0, 
    17, 18, 0, 0, 9, 5, 4, 0, 9, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 15, 35, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 15, 15, 17, 29, 15, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 6, 20, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 4, 17, 39, 37, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 38, 24, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=137
    5, 37, 26, 25, 25, 27, 31, 43, 61, 19, 67, 62, 45, 42, 33, 
    7, 20, 10, 29, 73, 39, 27, 48, 30, 3, 127, 65, 53, 44, 35, 
    7, 8, 46, 53, 70, 27, 0, 0, 0, 52, 101, 55, 62, 72, 72, 
    109, 140, 148, 16, 48, 56, 80, 43, 38, 66, 47, 90, 77, 40, 52, 
    73, 120, 62, 18, 70, 43, 33, 7, 32, 51, 57, 95, 70, 31, 50, 
    56, 57, 40, 40, 68, 36, 7, 24, 64, 70, 56, 82, 71, 57, 58, 
    51, 51, 0, 49, 47, 54, 31, 61, 49, 65, 62, 83, 70, 81, 83, 
    39, 38, 0, 71, 54, 48, 41, 39, 33, 41, 19, 0, 33, 40, 69, 
    43, 42, 52, 70, 69, 103, 82, 29, 35, 23, 39, 35, 0, 0, 46, 
    61, 74, 57, 60, 46, 19, 42, 70, 77, 58, 0, 21, 60, 35, 12, 
    63, 45, 63, 67, 73, 28, 42, 36, 30, 3, 15, 51, 42, 14, 16, 
    56, 40, 74, 57, 41, 20, 63, 51, 30, 0, 55, 24, 38, 25, 21, 
    52, 32, 65, 55, 3, 0, 33, 18, 0, 2, 29, 18, 0, 5, 29, 
    42, 28, 57, 63, 37, 82, 10, 4, 0, 0, 28, 22, 5, 29, 35, 
    14, 38, 42, 52, 47, 22, 0, 0, 0, 27, 17, 25, 27, 35, 14, 
    
    -- channel=138
    0, 11, 75, 78, 77, 83, 93, 86, 72, 57, 22, 97, 108, 109, 109, 
    0, 0, 57, 58, 47, 74, 61, 75, 81, 53, 45, 95, 105, 106, 107, 
    0, 0, 40, 71, 37, 57, 49, 49, 48, 31, 70, 78, 85, 89, 93, 
    55, 21, 72, 77, 31, 50, 57, 51, 36, 39, 62, 67, 84, 86, 75, 
    77, 73, 84, 76, 41, 52, 57, 47, 27, 34, 60, 84, 94, 103, 88, 
    84, 81, 85, 72, 51, 53, 55, 37, 34, 36, 59, 78, 98, 105, 99, 
    97, 87, 94, 58, 64, 46, 53, 27, 52, 39, 56, 82, 97, 97, 105, 
    96, 78, 79, 53, 68, 51, 39, 51, 36, 64, 60, 72, 69, 99, 84, 
    95, 73, 65, 76, 54, 64, 63, 57, 62, 61, 61, 70, 72, 69, 75, 
    94, 80, 71, 66, 71, 61, 45, 58, 76, 56, 75, 62, 62, 74, 75, 
    90, 84, 59, 80, 74, 76, 58, 60, 62, 78, 49, 64, 62, 65, 59, 
    91, 84, 63, 69, 76, 66, 70, 69, 72, 68, 56, 62, 56, 65, 57, 
    92, 92, 70, 67, 75, 57, 65, 74, 70, 57, 53, 55, 58, 49, 58, 
    91, 93, 71, 63, 74, 67, 80, 67, 62, 50, 53, 53, 51, 48, 55, 
    79, 81, 72, 50, 69, 76, 64, 53, 53, 38, 51, 51, 51, 54, 53, 
    
    -- channel=139
    0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 46, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 38, 0, 0, 0, 44, 71, 58, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 33, 0, 0, 0, 0, 8, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 12, 5, 0, 0, 0, 14, 6, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 11, 10, 0, 0, 0, 
    0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 6, 0, 3, 0, 0, 0, 0, 7, 7, 15, 126, 37, 12, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 113, 79, 42, 
    0, 0, 0, 0, 19, 43, 0, 0, 0, 0, 25, 0, 0, 0, 56, 
    0, 0, 0, 0, 0, 0, 30, 15, 0, 15, 0, 0, 0, 0, 3, 
    0, 0, 6, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 9, 0, 19, 46, 12, 18, 20, 0, 9, 5, 41, 16, 0, 
    0, 0, 17, 0, 0, 0, 20, 21, 17, 12, 6, 0, 0, 8, 0, 
    24, 0, 22, 20, 0, 0, 28, 20, 9, 0, 7, 0, 0, 0, 17, 
    
    -- channel=140
    1, 0, 0, 8, 9, 0, 3, 0, 14, 115, 0, 0, 0, 0, 7, 
    2, 0, 0, 0, 0, 35, 0, 0, 14, 90, 0, 0, 5, 3, 8, 
    5, 0, 0, 0, 0, 101, 21, 0, 8, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 61, 0, 17, 52, 40, 0, 0, 0, 0, 4, 42, 0, 
    14, 0, 0, 80, 0, 0, 31, 74, 0, 0, 0, 0, 0, 62, 0, 
    1, 0, 5, 45, 0, 6, 48, 20, 0, 0, 0, 0, 0, 57, 3, 
    7, 0, 57, 0, 13, 0, 45, 0, 12, 0, 0, 0, 0, 2, 29, 
    27, 0, 98, 0, 27, 13, 0, 63, 0, 0, 20, 0, 0, 20, 0, 
    53, 0, 0, 0, 0, 0, 34, 54, 0, 32, 0, 67, 0, 0, 0, 
    13, 7, 0, 0, 0, 0, 0, 7, 83, 0, 32, 0, 0, 12, 0, 
    0, 53, 0, 0, 0, 60, 0, 0, 13, 61, 0, 0, 0, 24, 12, 
    0, 44, 0, 0, 21, 23, 0, 0, 26, 61, 0, 5, 0, 33, 20, 
    8, 20, 0, 0, 72, 7, 0, 10, 31, 41, 0, 7, 5, 0, 11, 
    18, 30, 0, 0, 32, 27, 19, 14, 31, 8, 0, 6, 27, 0, 0, 
    15, 1, 0, 0, 17, 40, 49, 0, 44, 0, 0, 0, 8, 0, 0, 
    
    -- channel=141
    17, 28, 93, 79, 74, 80, 89, 80, 82, 58, 47, 95, 107, 102, 106, 
    18, 19, 75, 65, 63, 59, 62, 72, 77, 73, 57, 79, 89, 93, 98, 
    22, 19, 59, 68, 57, 61, 47, 48, 51, 51, 52, 50, 62, 68, 73, 
    71, 52, 64, 56, 47, 65, 72, 62, 52, 45, 55, 52, 69, 58, 47, 
    64, 56, 57, 57, 48, 54, 63, 55, 45, 41, 52, 53, 63, 56, 39, 
    55, 51, 53, 61, 52, 51, 59, 50, 54, 45, 48, 44, 52, 53, 37, 
    52, 55, 62, 69, 53, 47, 57, 45, 56, 42, 48, 53, 51, 58, 46, 
    46, 52, 92, 70, 57, 49, 49, 60, 52, 47, 53, 31, 45, 52, 41, 
    47, 43, 90, 72, 56, 65, 59, 67, 50, 60, 69, 69, 37, 40, 36, 
    47, 45, 63, 62, 47, 45, 51, 65, 73, 65, 68, 74, 72, 70, 51, 
    44, 43, 49, 64, 62, 61, 50, 54, 65, 69, 60, 68, 68, 67, 61, 
    42, 46, 42, 59, 65, 68, 68, 66, 67, 69, 61, 61, 67, 68, 66, 
    42, 41, 35, 55, 67, 72, 71, 65, 66, 62, 58, 57, 57, 59, 65, 
    44, 41, 23, 48, 69, 92, 73, 66, 64, 54, 58, 59, 60, 57, 65, 
    35, 42, 18, 43, 56, 65, 60, 63, 61, 52, 56, 61, 63, 60, 58, 
    
    -- channel=142
    0, 25, 49, 36, 33, 37, 31, 37, 28, 0, 54, 51, 43, 44, 40, 
    0, 4, 58, 53, 62, 39, 58, 64, 62, 17, 66, 73, 61, 56, 52, 
    0, 0, 56, 43, 97, 49, 42, 58, 60, 57, 76, 96, 85, 82, 74, 
    0, 0, 45, 47, 108, 78, 33, 25, 35, 70, 95, 109, 105, 98, 110, 
    53, 62, 77, 39, 85, 96, 73, 41, 46, 68, 95, 118, 113, 79, 92, 
    82, 84, 85, 50, 83, 89, 69, 44, 48, 64, 86, 126, 119, 79, 73, 
    81, 79, 57, 77, 68, 77, 57, 66, 65, 78, 83, 123, 123, 105, 73, 
    78, 80, 31, 93, 76, 85, 77, 50, 88, 68, 79, 104, 139, 115, 110, 
    72, 70, 58, 77, 100, 91, 72, 52, 58, 57, 64, 27, 77, 98, 115, 
    84, 70, 86, 88, 97, 108, 112, 79, 31, 59, 52, 49, 41, 46, 67, 
    98, 75, 101, 88, 91, 71, 96, 97, 83, 50, 52, 49, 59, 48, 42, 
    99, 79, 101, 103, 95, 75, 80, 82, 75, 38, 49, 57, 68, 46, 37, 
    92, 78, 99, 104, 75, 52, 85, 78, 64, 38, 53, 50, 55, 57, 41, 
    85, 66, 89, 107, 73, 44, 61, 58, 43, 35, 44, 42, 32, 45, 49, 
    78, 66, 70, 113, 88, 67, 47, 47, 25, 30, 39, 41, 32, 36, 51, 
    
    -- channel=143
    0, 2, 1, 0, 0, 4, 3, 0, 0, 0, 0, 0, 2, 2, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=144
    90, 80, 92, 109, 78, 65, 50, 29, 71, 114, 113, 117, 79, 64, 71, 
    122, 119, 124, 145, 113, 120, 147, 180, 176, 161, 130, 106, 128, 120, 92, 
    139, 139, 142, 93, 32, 21, 26, 18, 34, 57, 87, 97, 118, 115, 103, 
    138, 137, 141, 122, 50, 112, 113, 112, 88, 72, 67, 128, 116, 65, 84, 
    142, 135, 170, 136, 60, 111, 138, 100, 104, 116, 90, 76, 108, 85, 16, 
    148, 151, 112, 80, 87, 79, 80, 104, 110, 98, 135, 120, 111, 140, 138, 
    123, 160, 129, 83, 3, 75, 85, 61, 58, 82, 82, 86, 149, 191, 144, 
    127, 147, 69, 69, 98, 66, 51, 62, 98, 94, 68, 97, 106, 99, 117, 
    83, 79, 37, 158, 34, 69, 63, 4, 0, 0, 0, 0, 0, 59, 122, 
    112, 95, 72, 39, 51, 49, 60, 93, 119, 110, 129, 115, 110, 111, 79, 
    117, 93, 0, 19, 15, 36, 0, 28, 64, 48, 40, 9, 75, 17, 71, 
    123, 119, 40, 0, 0, 3, 86, 84, 30, 97, 39, 81, 112, 74, 77, 
    120, 12, 0, 49, 19, 0, 0, 0, 0, 0, 34, 32, 33, 0, 21, 
    91, 123, 79, 58, 39, 7, 0, 0, 0, 79, 128, 86, 12, 0, 54, 
    117, 92, 61, 68, 33, 15, 0, 0, 0, 24, 68, 73, 0, 0, 20, 
    
    -- channel=145
    25, 26, 17, 18, 24, 25, 31, 41, 35, 26, 29, 30, 22, 44, 31, 
    16, 17, 10, 0, 0, 0, 0, 0, 0, 15, 30, 33, 27, 27, 50, 
    12, 13, 0, 0, 0, 0, 0, 0, 0, 0, 25, 31, 23, 25, 60, 
    12, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 27, 20, 30, 43, 
    15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 22, 4, 34, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 13, 13, 
    22, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 13, 12, 
    13, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    15, 0, 34, 0, 2, 8, 0, 0, 17, 29, 0, 16, 21, 0, 34, 
    1, 0, 7, 0, 2, 0, 0, 9, 0, 0, 0, 0, 0, 0, 39, 
    6, 0, 13, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 0, 10, 2, 0, 10, 15, 0, 49, 0, 0, 10, 0, 0, 42, 
    0, 0, 10, 0, 0, 1, 15, 14, 22, 49, 7, 0, 0, 15, 37, 
    0, 0, 0, 0, 0, 0, 19, 22, 20, 9, 0, 0, 0, 24, 20, 
    0, 0, 0, 0, 0, 0, 11, 9, 8, 3, 0, 0, 2, 17, 30, 
    
    -- channel=146
    64, 59, 69, 45, 39, 39, 39, 39, 53, 68, 59, 64, 57, 42, 31, 
    87, 85, 86, 52, 56, 64, 61, 72, 79, 63, 48, 62, 68, 50, 42, 
    92, 92, 89, 42, 49, 63, 66, 63, 65, 55, 60, 65, 63, 37, 32, 
    91, 91, 78, 74, 54, 73, 72, 92, 86, 79, 48, 69, 64, 44, 9, 
    90, 91, 75, 66, 62, 68, 89, 80, 81, 77, 86, 71, 73, 76, 51, 
    83, 89, 53, 38, 27, 56, 65, 58, 59, 62, 75, 57, 86, 91, 91, 
    64, 69, 42, 34, 35, 60, 65, 44, 49, 55, 22, 27, 59, 82, 86, 
    52, 28, 23, 39, 36, 22, 22, 15, 0, 0, 4, 0, 15, 55, 93, 
    57, 14, 8, 26, 11, 21, 18, 11, 0, 0, 9, 0, 10, 42, 53, 
    68, 21, 16, 0, 0, 9, 7, 31, 47, 61, 62, 55, 71, 32, 34, 
    70, 31, 0, 0, 0, 0, 2, 3, 7, 26, 20, 23, 27, 21, 21, 
    82, 26, 2, 6, 0, 0, 0, 0, 0, 17, 24, 37, 0, 5, 11, 
    79, 44, 5, 37, 3, 0, 0, 0, 0, 17, 36, 37, 0, 0, 9, 
    74, 73, 44, 36, 9, 0, 0, 0, 0, 14, 60, 54, 0, 0, 20, 
    76, 69, 54, 17, 1, 0, 0, 0, 0, 0, 14, 31, 0, 0, 22, 
    
    -- channel=147
    252, 245, 251, 196, 200, 205, 215, 229, 255, 263, 250, 262, 246, 213, 212, 
    291, 289, 277, 188, 186, 197, 192, 211, 235, 239, 231, 255, 261, 220, 230, 
    298, 298, 277, 175, 180, 197, 197, 189, 179, 171, 210, 259, 240, 201, 196, 
    297, 292, 266, 198, 207, 258, 246, 250, 244, 235, 202, 244, 256, 202, 167, 
    297, 290, 224, 196, 201, 216, 237, 229, 236, 244, 247, 226, 276, 262, 220, 
    284, 276, 234, 156, 146, 193, 185, 192, 194, 206, 214, 225, 276, 300, 298, 
    245, 225, 187, 183, 155, 186, 201, 162, 172, 187, 151, 157, 216, 260, 308, 
    217, 146, 173, 163, 169, 145, 116, 106, 99, 105, 92, 99, 152, 185, 278, 
    212, 132, 150, 116, 146, 140, 178, 136, 110, 127, 138, 98, 140, 175, 242, 
    242, 123, 121, 75, 96, 106, 99, 143, 199, 176, 185, 177, 186, 150, 197, 
    244, 141, 89, 82, 43, 76, 125, 73, 145, 130, 133, 161, 99, 163, 173, 
    248, 117, 99, 129, 53, 29, 77, 87, 74, 165, 158, 155, 114, 94, 166, 
    247, 185, 97, 161, 100, 22, 13, 24, 46, 171, 208, 164, 45, 66, 149, 
    229, 230, 178, 142, 116, 57, 14, 28, 60, 135, 197, 163, 32, 62, 171, 
    233, 217, 180, 106, 101, 66, 38, 47, 60, 89, 127, 138, 28, 62, 182, 
    
    -- channel=148
    53, 50, 53, 79, 53, 22, 14, 0, 34, 73, 81, 75, 56, 54, 74, 
    54, 54, 68, 92, 61, 50, 65, 96, 100, 112, 110, 66, 83, 114, 83, 
    65, 64, 75, 74, 0, 0, 0, 0, 0, 0, 42, 52, 80, 120, 98, 
    65, 71, 67, 72, 0, 0, 6, 0, 0, 0, 4, 73, 74, 60, 83, 
    66, 71, 90, 64, 0, 0, 25, 0, 0, 0, 0, 0, 43, 53, 0, 
    64, 85, 46, 24, 7, 0, 0, 0, 10, 0, 23, 33, 29, 66, 63, 
    47, 97, 67, 28, 0, 0, 0, 0, 0, 0, 25, 25, 74, 93, 72, 
    62, 107, 16, 37, 13, 15, 0, 22, 50, 49, 34, 54, 37, 6, 22, 
    28, 43, 8, 116, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    52, 74, 49, 40, 8, 27, 24, 8, 58, 32, 56, 47, 37, 55, 0, 
    45, 67, 0, 20, 18, 14, 0, 8, 18, 10, 7, 0, 19, 0, 0, 
    34, 100, 18, 0, 11, 19, 54, 88, 0, 56, 0, 23, 97, 49, 0, 
    17, 0, 0, 15, 13, 9, 17, 10, 0, 0, 0, 26, 36, 0, 0, 
    0, 35, 25, 28, 9, 27, 2, 0, 0, 32, 52, 74, 36, 0, 0, 
    19, 5, 10, 34, 16, 21, 0, 0, 0, 3, 16, 46, 17, 0, 0, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 50, 55, 60, 93, 93, 52, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 
    0, 0, 17, 29, 3, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 16, 22, 0, 33, 0, 0, 0, 0, 
    0, 22, 9, 0, 0, 0, 11, 0, 1, 30, 10, 24, 63, 68, 0, 
    4, 18, 2, 0, 13, 0, 0, 1, 56, 53, 27, 65, 60, 9, 16, 
    0, 0, 0, 60, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 64, 0, 36, 3, 16, 30, 29, 21, 40, 34, 50, 14, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 45, 0, 0, 0, 57, 58, 27, 39, 0, 23, 21, 59, 0, 
    0, 0, 0, 6, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 21, 0, 0, 0, 0, 0, 43, 47, 28, 0, 0, 0, 
    0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 13, 42, 0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 1, 3, 25, 26, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 21, 8, 35, 36, 2, 28, 0, 0, 40, 
    0, 0, 0, 0, 40, 0, 0, 0, 0, 12, 109, 12, 0, 0, 68, 
    0, 0, 0, 0, 122, 30, 0, 0, 0, 0, 0, 85, 0, 0, 0, 
    0, 0, 0, 0, 74, 24, 0, 4, 7, 15, 0, 85, 31, 0, 0, 
    39, 0, 0, 0, 61, 16, 0, 0, 0, 21, 9, 56, 104, 0, 0, 
    23, 0, 0, 0, 11, 0, 0, 0, 24, 0, 0, 69, 79, 55, 33, 
    0, 0, 94, 0, 0, 0, 0, 0, 0, 10, 0, 27, 95, 63, 148, 
    0, 0, 83, 0, 54, 14, 7, 0, 0, 26, 0, 0, 53, 0, 158, 
    0, 0, 43, 0, 43, 0, 31, 97, 0, 16, 0, 0, 8, 0, 208, 
    0, 0, 0, 0, 0, 40, 51, 0, 98, 0, 0, 51, 0, 43, 145, 
    0, 0, 66, 0, 0, 17, 73, 0, 147, 1, 2, 22, 0, 23, 216, 
    0, 0, 0, 0, 0, 0, 1, 18, 46, 185, 0, 0, 0, 53, 202, 
    4, 0, 0, 0, 0, 0, 0, 21, 53, 86, 43, 0, 0, 92, 170, 
    0, 0, 0, 0, 0, 0, 0, 3, 16, 26, 44, 0, 0, 70, 204, 
    
    -- channel=151
    23, 19, 19, 0, 15, 42, 48, 57, 28, 6, 0, 0, 30, 13, 18, 
    21, 20, 16, 5, 15, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 12, 13, 57, 116, 141, 141, 144, 121, 69, 4, 11, 0, 0, 0, 
    12, 8, 17, 54, 102, 88, 97, 111, 123, 135, 60, 0, 12, 14, 0, 
    9, 14, 0, 63, 97, 79, 84, 111, 103, 100, 102, 46, 20, 36, 63, 
    0, 0, 50, 85, 66, 97, 103, 88, 81, 86, 61, 40, 18, 13, 13, 
    2, 0, 0, 83, 128, 112, 109, 112, 109, 87, 63, 28, 0, 0, 9, 
    0, 0, 24, 29, 71, 82, 79, 59, 29, 36, 45, 19, 35, 45, 17, 
    32, 42, 19, 0, 81, 57, 93, 118, 154, 156, 147, 154, 137, 83, 25, 
    24, 26, 1, 46, 46, 56, 37, 32, 41, 37, 31, 34, 26, 48, 39, 
    22, 49, 64, 57, 47, 52, 106, 57, 51, 68, 72, 90, 51, 94, 55, 
    39, 20, 34, 106, 73, 33, 0, 26, 24, 37, 68, 21, 25, 15, 40, 
    60, 128, 96, 60, 76, 63, 46, 50, 60, 89, 88, 73, 45, 65, 73, 
    66, 55, 69, 48, 66, 64, 59, 63, 55, 15, 20, 43, 44, 60, 74, 
    69, 79, 82, 52, 58, 59, 64, 65, 60, 56, 39, 54, 58, 57, 92, 
    
    -- channel=152
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=153
    90, 98, 78, 30, 52, 73, 101, 133, 109, 75, 67, 69, 91, 91, 77, 
    86, 87, 57, 0, 0, 0, 0, 0, 0, 5, 35, 68, 59, 38, 78, 
    74, 72, 49, 8, 71, 97, 105, 100, 70, 40, 74, 82, 46, 14, 49, 
    74, 64, 50, 0, 81, 70, 50, 45, 70, 86, 58, 41, 59, 65, 38, 
    70, 59, 0, 0, 61, 31, 10, 45, 43, 50, 57, 87, 91, 92, 140, 
    53, 28, 50, 1, 7, 41, 30, 13, 7, 28, 8, 34, 87, 73, 75, 
    42, 0, 0, 25, 100, 41, 26, 32, 44, 25, 6, 18, 0, 0, 62, 
    16, 0, 49, 32, 7, 15, 17, 0, 0, 0, 0, 0, 0, 23, 76, 
    56, 13, 46, 0, 41, 25, 48, 84, 167, 174, 152, 172, 162, 61, 65, 
    48, 0, 0, 2, 4, 0, 0, 14, 0, 0, 0, 0, 2, 0, 85, 
    48, 0, 28, 14, 3, 10, 92, 11, 25, 31, 29, 92, 5, 65, 89, 
    37, 0, 22, 77, 18, 6, 0, 0, 20, 0, 51, 6, 0, 0, 71, 
    43, 87, 105, 23, 26, 14, 5, 12, 27, 142, 106, 38, 0, 32, 111, 
    61, 19, 18, 11, 19, 1, 27, 32, 45, 0, 0, 0, 0, 45, 86, 
    31, 45, 33, 0, 12, 9, 31, 33, 30, 22, 9, 0, 9, 41, 117, 
    
    -- channel=154
    74, 76, 70, 69, 39, 44, 50, 59, 73, 77, 81, 71, 74, 88, 72, 
    72, 73, 74, 38, 0, 0, 0, 3, 9, 40, 67, 70, 76, 92, 72, 
    71, 71, 66, 28, 0, 0, 0, 0, 0, 0, 27, 72, 85, 78, 76, 
    71, 70, 59, 12, 0, 0, 0, 0, 0, 0, 24, 42, 68, 83, 75, 
    69, 70, 42, 0, 0, 0, 0, 0, 0, 0, 0, 28, 60, 74, 74, 
    56, 66, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 71, 71, 
    55, 54, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 30, 54, 
    55, 43, 4, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    56, 26, 23, 11, 0, 0, 0, 0, 0, 6, 8, 11, 2, 0, 18, 
    51, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 22, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 11, 0, 2, 
    23, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 24, 14, 0, 0, 0, 
    4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 75, 86, 112, 143, 127, 85, 29, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 32, 0, 0, 11, 43, 
    0, 0, 0, 0, 5, 0, 0, 19, 0, 0, 30, 57, 0, 0, 17, 
    0, 0, 63, 11, 28, 55, 34, 24, 27, 23, 0, 19, 0, 0, 0, 
    25, 16, 0, 0, 80, 18, 20, 47, 59, 41, 71, 63, 18, 0, 0, 
    28, 48, 47, 0, 0, 13, 5, 3, 1, 29, 30, 74, 133, 107, 8, 
    30, 61, 0, 0, 43, 19, 30, 39, 90, 83, 55, 98, 101, 72, 55, 
    0, 0, 17, 83, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 82, 
    0, 0, 77, 0, 68, 19, 77, 63, 69, 81, 88, 82, 76, 49, 57, 
    0, 0, 0, 0, 14, 32, 0, 4, 50, 0, 3, 0, 32, 0, 41, 
    14, 11, 30, 0, 0, 26, 125, 32, 75, 20, 0, 63, 16, 112, 47, 
    13, 0, 0, 8, 0, 0, 2, 5, 3, 0, 0, 0, 9, 0, 17, 
    0, 24, 0, 19, 0, 0, 0, 0, 0, 121, 83, 17, 0, 6, 28, 
    24, 0, 0, 29, 12, 0, 0, 0, 0, 19, 57, 19, 0, 6, 0, 
    
    -- channel=156
    0, 0, 8, 57, 0, 0, 0, 0, 0, 0, 13, 0, 13, 1, 15, 
    0, 0, 26, 125, 10, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 
    0, 0, 24, 195, 0, 0, 0, 22, 1, 0, 0, 0, 35, 46, 0, 
    0, 13, 16, 158, 0, 0, 73, 0, 0, 0, 26, 0, 0, 40, 21, 
    0, 16, 92, 97, 0, 2, 20, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 41, 58, 141, 0, 0, 24, 7, 2, 0, 0, 0, 0, 0, 0, 
    0, 56, 27, 35, 1, 13, 19, 16, 0, 0, 33, 0, 0, 0, 0, 
    22, 109, 0, 101, 11, 20, 1, 45, 12, 0, 29, 6, 0, 0, 0, 
    34, 116, 0, 95, 0, 0, 0, 12, 0, 0, 30, 0, 0, 19, 0, 
    29, 184, 0, 91, 0, 32, 0, 0, 25, 0, 19, 0, 0, 59, 0, 
    4, 164, 15, 27, 38, 0, 0, 120, 0, 41, 1, 0, 70, 0, 0, 
    18, 214, 0, 0, 96, 23, 0, 48, 0, 0, 0, 6, 126, 0, 0, 
    0, 82, 24, 0, 50, 64, 4, 0, 0, 0, 14, 112, 79, 0, 0, 
    0, 25, 66, 11, 8, 74, 0, 0, 0, 0, 0, 100, 52, 0, 0, 
    8, 9, 48, 49, 3, 28, 7, 0, 0, 0, 0, 10, 65, 0, 0, 
    
    -- channel=157
    53, 51, 60, 50, 44, 55, 51, 53, 48, 46, 47, 48, 57, 47, 44, 
    53, 53, 56, 28, 14, 11, 3, 3, 10, 23, 28, 51, 51, 46, 38, 
    52, 52, 54, 44, 16, 28, 26, 24, 17, 13, 18, 57, 60, 46, 25, 
    52, 52, 49, 39, 22, 35, 25, 7, 18, 21, 32, 29, 59, 64, 40, 
    53, 55, 26, 18, 13, 6, 6, 10, 13, 8, 21, 35, 50, 65, 71, 
    53, 55, 50, 40, 3, 13, 14, 6, 6, 11, 5, 18, 41, 53, 53, 
    61, 56, 50, 40, 26, 16, 17, 15, 12, 15, 17, 9, 14, 19, 47, 
    73, 48, 52, 55, 13, 32, 25, 22, 10, 7, 14, 5, 2, 12, 37, 
    73, 52, 54, 20, 33, 25, 31, 49, 62, 57, 66, 62, 50, 40, 32, 
    66, 43, 30, 27, 8, 19, 8, 4, 26, 10, 12, 12, 16, 17, 19, 
    59, 47, 43, 28, 21, 12, 32, 33, 20, 37, 33, 42, 30, 36, 24, 
    46, 35, 21, 48, 34, 14, 1, 17, 8, 25, 36, 28, 18, 12, 8, 
    40, 63, 41, 38, 34, 27, 17, 16, 17, 40, 53, 57, 24, 18, 12, 
    41, 39, 41, 34, 25, 33, 22, 21, 19, 10, 15, 45, 20, 13, 11, 
    29, 31, 41, 23, 23, 27, 24, 24, 22, 23, 21, 37, 26, 17, 17, 
    
    -- channel=158
    109, 107, 105, 77, 86, 85, 89, 93, 115, 122, 114, 122, 97, 91, 85, 
    130, 129, 117, 68, 89, 100, 99, 114, 129, 132, 116, 119, 122, 99, 112, 
    137, 137, 120, 40, 80, 77, 78, 67, 68, 74, 118, 120, 102, 85, 108, 
    136, 132, 117, 56, 110, 130, 103, 118, 111, 104, 91, 131, 111, 73, 76, 
    138, 128, 98, 67, 105, 104, 108, 110, 114, 117, 106, 117, 129, 103, 75, 
    138, 121, 87, 38, 85, 92, 80, 92, 96, 100, 112, 120, 144, 137, 137, 
    112, 94, 82, 56, 55, 82, 85, 67, 76, 87, 69, 87, 127, 143, 149, 
    94, 50, 82, 56, 72, 63, 51, 45, 59, 61, 42, 59, 92, 93, 156, 
    75, 27, 69, 47, 65, 63, 75, 39, 12, 26, 23, 5, 41, 73, 144, 
    96, 18, 68, 9, 49, 40, 52, 79, 91, 87, 88, 86, 94, 59, 118, 
    104, 23, 24, 20, 12, 42, 50, 13, 84, 48, 54, 72, 34, 66, 96, 
    106, 18, 57, 34, 0, 10, 55, 31, 52, 76, 65, 75, 33, 57, 103, 
    111, 38, 22, 66, 23, 0, 0, 5, 18, 89, 80, 43, 5, 29, 87, 
    101, 100, 62, 62, 44, 2, 0, 2, 24, 81, 101, 49, 0, 32, 98, 
    105, 93, 63, 39, 41, 16, 3, 9, 20, 39, 65, 52, 0, 30, 101, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
