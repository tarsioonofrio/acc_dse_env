library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 44, 
    32, 0, 0, 1, 27, 0, 0, 
    20, 0, 7, 87, 75, 80, 105, 
    0, 0, 157, 60, 58, 66, 62, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    14, 0, 0, 21, 32, 13, 65, 
    0, 64, 1, 0, 86, 0, 0, 
    0, 0, 55, 0, 0, 0, 0, 
    0, 56, 69, 59, 5, 0, 32, 
    0, 29, 0, 0, 45, 10, 75, 
    162, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 15, 0, 24, 
    196, 0, 0, 0, 62, 64, 0, 
    158, 173, 26, 0, 100, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 169, 204, 191, 165, 
    212, 0, 60, 0, 0, 0, 49, 
    73, 0, 39, 0, 0, 24, 0, 
    0, 131, 0, 71, 0, 0, 0, 
    0, 0, 96, 0, 112, 110, 130, 
    164, 0, 351, 275, 53, 78, 0, 
    0, 172, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 35, 0, 0, 0, 
    117, 0, 0, 77, 0, 0, 8, 
    30, 167, 0, 0, 0, 0, 0, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 164, 144, 0, 
    148, 0, 288, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 45, 
    49, 34, 0, 40, 0, 0, 0, 
    0, 0, 220, 0, 0, 242, 0, 
    0, 0, 0, 190, 0, 0, 0, 
    0, 186, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 7, 0, 0, 
    50, 0, 16, 20, 175, 0, 14, 
    129, 0, 115, 30, 316, 0, 43, 
    205, 115, 117, 32, 110, 0, 29, 
    117, 237, 60, 85, 0, 39, 57, 
    92, 267, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    47, 9, 115, 0, 89, 36, 71, 
    13, 114, 24, 0, 44, 0, 0, 
    0, 0, 48, 0, 78, 0, 0, 
    0, 0, 6, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 72, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    128, 186, 0, 68, 0, 0, 100, 
    0, 357, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 129, 0, 
    50, 0, 0, 33, 0, 160, 144, 
    249, 0, 0, 292, 0, 203, 87, 
    184, 0, 0, 155, 0, 149, 0, 
    159, 20, 0, 0, 58, 0, 0, 
    0, 0, 292, 44, 104, 0, 25, 
    26, 0, 84, 54, 0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 0, 13, 0, 0, 
    0, 39, 46, 12, 0, 15, 0, 
    29, 0, 5, 53, 0, 37, 0, 
    32, 36, 0, 35, 42, 13, 0, 
    0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 114, 0, 0, 
    0, 64, 68, 0, 0, 0, 0, 
    0, 0, 47, 0, 0, 21, 0, 
    0, 0, 0, 87, 0, 0, 0, 
    0, 7, 153, 0, 78, 33, 0, 
    0, 0, 136, 27, 0, 0, 0, 
    0, 125, 0, 0, 0, 0, 0, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 
    0, 0, 13, 14, 24, 81, 25, 
    0, 0, 0, 0, 2, 0, 1, 
    
    -- channel=26
    0, 0, 161, 55, 214, 0, 28, 
    650, 175, 101, 0, 441, 0, 0, 
    461, 0, 0, 0, 1068, 0, 0, 
    256, 0, 240, 132, 445, 0, 6, 
    290, 1046, 25, 0, 0, 0, 0, 
    29, 760, 0, 0, 0, 0, 0, 
    0, 0, 215, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    82, 1, 96, 118, 49, 19, 78, 
    35, 16, 0, 30, 13, 0, 11, 
    9, 0, 0, 0, 53, 0, 0, 
    34, 88, 97, 22, 0, 51, 0, 
    0, 0, 0, 62, 60, 23, 7, 
    58, 8, 0, 5, 0, 0, 0, 
    0, 102, 23, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 16, 0, 131, 0, 
    0, 0, 0, 168, 0, 127, 29, 
    0, 0, 0, 304, 0, 211, 44, 
    77, 0, 0, 0, 0, 135, 0, 
    0, 0, 18, 0, 11, 0, 0, 
    0, 0, 283, 0, 89, 0, 0, 
    0, 0, 169, 93, 27, 0, 0, 
    
    -- channel=32
    0, 0, 55, 0, 0, 0, 0, 
    0, 0, 0, 31, 0, 33, 0, 
    7, 0, 30, 93, 119, 0, 20, 
    0, 0, 2, 0, 30, 32, 37, 
    51, 50, 0, 171, 0, 0, 47, 
    0, 387, 30, 0, 57, 66, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 9, 0, 
    43, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 73, 20, 0, 0, 28, 0, 
    0, 0, 13, 14, 0, 47, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 32, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 78, 126, 
    0, 0, 11, 150, 194, 197, 155, 
    
    -- channel=36
    2, 12, 0, 24, 0, 0, 19, 
    0, 86, 0, 0, 35, 28, 31, 
    128, 79, 51, 27, 0, 18, 3, 
    84, 16, 26, 83, 73, 20, 71, 
    126, 123, 7, 15, 9, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 43, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 71, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 59, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    78, 82, 53, 121, 68, 22, 82, 
    0, 125, 60, 14, 46, 69, 20, 
    89, 0, 46, 0, 0, 77, 0, 
    0, 37, 63, 139, 125, 57, 67, 
    0, 22, 87, 0, 3, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 0, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 76, 32, 9, 30, 51, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    33, 19, 25, 35, 0, 6, 27, 
    8, 84, 44, 44, 27, 36, 0, 
    0, 0, 33, 63, 0, 65, 6, 
    0, 52, 0, 35, 0, 37, 8, 
    0, 43, 23, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 83, 
    5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 71, 95, 46, 
    0, 0, 0, 10, 35, 9, 0, 
    
    -- channel=44
    355, 378, 260, 185, 98, 23, 194, 
    59, 260, 139, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 83, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    83, 66, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 0, 71, 
    0, 0, 0, 65, 63, 252, 140, 
    92, 0, 0, 92, 112, 152, 14, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 74, 0, 
    143, 0, 270, 205, 325, 319, 312, 
    335, 266, 398, 225, 269, 348, 248, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 
    76, 0, 0, 179, 54, 0, 90, 
    221, 0, 0, 0, 0, 49, 0, 
    269, 174, 0, 147, 0, 0, 0, 
    20, 176, 0, 0, 43, 38, 71, 
    0, 223, 121, 102, 122, 87, 196, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    0, 0, 186, 0, 253, 9, 0, 
    46, 42, 198, 0, 54, 0, 0, 
    0, 33, 0, 0, 426, 0, 0, 
    0, 0, 19, 0, 23, 0, 0, 
    0, 0, 0, 224, 0, 0, 139, 
    0, 490, 0, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 0, 66, 
    
    -- channel=54
    0, 0, 0, 0, 63, 0, 0, 
    180, 0, 0, 0, 46, 0, 41, 
    0, 146, 0, 0, 394, 0, 0, 
    0, 97, 0, 0, 80, 0, 0, 
    0, 44, 46, 0, 0, 99, 32, 
    0, 0, 0, 0, 108, 4, 0, 
    17, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    124, 127, 98, 149, 136, 81, 99, 
    97, 141, 137, 82, 19, 60, 32, 
    41, 20, 0, 45, 0, 41, 44, 
    17, 19, 0, 62, 0, 48, 58, 
    2, 49, 92, 10, 93, 87, 72, 
    0, 0, 139, 35, 57, 49, 33, 
    0, 24, 104, 31, 24, 21, 14, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 77, 
    218, 0, 0, 62, 87, 193, 0, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 183, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 10, 7, 59, 0, 
    36, 0, 23, 102, 106, 154, 162, 
    249, 92, 172, 161, 149, 156, 160, 
    
    -- channel=61
    19, 8, 0, 68, 24, 85, 61, 
    141, 116, 86, 151, 111, 119, 169, 
    222, 295, 14, 203, 250, 220, 81, 
    252, 235, 4, 122, 175, 147, 40, 
    106, 255, 210, 75, 111, 34, 12, 
    30, 219, 144, 0, 30, 0, 0, 
    94, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 50, 0, 0, 0, 
    100, 0, 0, 101, 65, 17, 78, 
    15, 122, 99, 42, 14, 61, 2, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    142, 198, 109, 116, 3, 0, 129, 
    0, 135, 0, 0, 49, 16, 41, 
    73, 0, 0, 5, 40, 32, 0, 
    123, 163, 64, 21, 173, 46, 0, 
    100, 0, 0, 0, 8, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 0, 
    16, 0, 0, 107, 0, 46, 0, 
    50, 0, 0, 83, 0, 15, 0, 
    116, 0, 0, 0, 0, 0, 0, 
    0, 0, 65, 87, 0, 0, 0, 
    0, 300, 97, 4, 14, 0, 63, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=67
    0, 0, 0, 0, 0, 3, 36, 
    0, 0, 0, 0, 38, 0, 75, 
    67, 0, 0, 6, 101, 0, 73, 
    36, 0, 0, 0, 131, 28, 0, 
    185, 5, 0, 0, 0, 0, 61, 
    132, 245, 0, 146, 335, 353, 332, 
    404, 126, 317, 315, 378, 395, 427, 
    
    -- channel=68
    61, 95, 93, 28, 44, 23, 30, 
    0, 101, 23, 0, 53, 0, 37, 
    0, 32, 60, 0, 49, 0, 5, 
    0, 15, 0, 0, 32, 0, 9, 
    0, 0, 0, 6, 0, 0, 42, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=69
    224, 96, 52, 85, 0, 0, 200, 
    0, 0, 0, 0, 0, 0, 0, 
    171, 91, 134, 0, 0, 0, 0, 
    0, 0, 59, 0, 73, 0, 27, 
    0, 0, 0, 0, 0, 0, 89, 
    199, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 28, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 
    111, 0, 0, 15, 26, 36, 30, 
    
    -- channel=71
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=72
    35, 75, 25, 48, 64, 88, 44, 
    0, 0, 60, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 27, 23, 59, 75, 
    0, 0, 32, 65, 59, 39, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    0, 0, 0, 0, 85, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 6, 0, 
    65, 53, 124, 19, 167, 231, 90, 
    10, 0, 151, 22, 97, 24, 103, 
    
    -- channel=76
    0, 17, 93, 0, 0, 0, 0, 
    0, 0, 63, 0, 0, 0, 0, 
    0, 0, 83, 66, 0, 0, 84, 
    179, 0, 175, 0, 0, 0, 28, 
    256, 0, 0, 176, 54, 0, 15, 
    126, 55, 0, 91, 0, 1, 55, 
    0, 563, 0, 0, 31, 45, 101, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=78
    62, 55, 0, 0, 49, 0, 120, 
    88, 112, 0, 0, 260, 0, 0, 
    247, 0, 28, 0, 345, 0, 34, 
    318, 228, 157, 0, 107, 0, 42, 
    108, 182, 0, 0, 0, 0, 125, 
    253, 0, 0, 0, 0, 39, 62, 
    40, 160, 0, 21, 44, 69, 0, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 78, 85, 0, 
    84, 10, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 76, 0, 0, 12, 
    0, 0, 0, 0, 0, 20, 146, 
    0, 0, 0, 139, 147, 124, 182, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 
    37, 0, 7, 45, 82, 55, 22, 
    34, 66, 0, 89, 153, 56, 8, 
    35, 23, 32, 18, 48, 23, 44, 
    0, 191, 25, 17, 41, 0, 0, 
    0, 97, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 53, 0, 0, 
    0, 0, 216, 0, 0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    0, 0, 0, 52, 182, 3, 0, 
    66, 358, 147, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 0, 0, 0, 0, 
    0, 163, 118, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    112, 72, 50, 0, 101, 0, 92, 
    320, 214, 37, 0, 97, 0, 69, 
    0, 0, 0, 0, 283, 0, 0, 
    0, 144, 0, 0, 0, 0, 0, 
    0, 197, 113, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=96
    0, 0, 85, 290, 265, 150, 99, 
    0, 4, 0, 4, 0, 0, 0, 
    15, 0, 13, 0, 0, 24, 0, 
    0, 34, 0, 91, 0, 30, 0, 
    0, 0, 0, 0, 83, 32, 93, 
    131, 0, 364, 188, 83, 15, 72, 
    0, 249, 144, 40, 0, 20, 0, 
    
    -- channel=97
    144, 99, 4, 7, 0, 0, 94, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    208, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 45, 
    0, 0, 0, 107, 81, 27, 1, 
    
    -- channel=98
    232, 146, 63, 117, 44, 160, 231, 
    314, 182, 0, 0, 51, 0, 15, 
    36, 0, 0, 0, 151, 0, 0, 
    0, 95, 0, 0, 0, 0, 35, 
    0, 0, 0, 37, 0, 0, 328, 
    23, 0, 0, 0, 21, 118, 167, 
    111, 0, 5, 199, 171, 194, 185, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 0, 
    0, 2, 43, 0, 193, 0, 0, 
    0, 2, 0, 0, 34, 0, 0, 
    0, 0, 74, 94, 0, 41, 23, 
    0, 255, 85, 15, 28, 27, 0, 
    11, 0, 0, 0, 0, 0, 32, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 137, 14, 0, 0, 18, 
    0, 0, 0, 62, 30, 13, 33, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 38, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 3, 0, 0, 0, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 0, 0, 52, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 83, 0, 
    0, 0, 265, 182, 280, 116, 109, 
    82, 0, 214, 20, 12, 36, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    0, 0, 64, 0, 151, 0, 94, 
    0, 8, 0, 0, 15, 0, 0, 
    188, 0, 450, 49, 7, 60, 273, 
    125, 141, 59, 57, 0, 0, 0, 
    0, 0, 0, 57, 49, 0, 2, 
    245, 0, 438, 0, 87, 65, 0, 
    0, 124, 158, 0, 0, 0, 0, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 46, 0, 0, 90, 
    0, 2, 0, 0, 0, 178, 23, 
    65, 222, 0, 0, 0, 178, 0, 
    0, 0, 51, 34, 0, 55, 0, 
    0, 0, 0, 0, 0, 0, 37, 
    0, 47, 0, 62, 11, 11, 0, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 20, 48, 0, 0, 0, 0, 
    22, 0, 128, 82, 87, 126, 77, 
    8, 0, 16, 13, 59, 68, 88, 
    
    -- channel=113
    0, 0, 0, 121, 135, 249, 112, 
    0, 0, 125, 80, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 60, 132, 
    0, 0, 0, 173, 177, 155, 144, 
    36, 0, 182, 66, 100, 49, 36, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 51, 0, 0, 0, 0, 
    0, 0, 253, 6, 44, 112, 54, 
    0, 0, 98, 15, 26, 46, 30, 
    
    -- channel=115
    40, 23, 20, 36, 11, 0, 29, 
    0, 45, 0, 0, 74, 8, 15, 
    39, 52, 52, 0, 56, 35, 16, 
    0, 25, 35, 22, 86, 32, 60, 
    0, 6, 0, 0, 0, 0, 1, 
    0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 246, 0, 0, 
    0, 0, 0, 0, 105, 0, 0, 
    0, 0, 108, 0, 14, 0, 0, 
    85, 220, 0, 0, 0, 0, 0, 
    242, 0, 0, 17, 0, 0, 67, 
    0, 57, 0, 64, 62, 81, 128, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 55, 0, 
    0, 0, 77, 60, 0, 21, 49, 
    20, 0, 0, 21, 4, 0, 11, 
    20, 76, 191, 84, 0, 62, 0, 
    21, 6, 21, 13, 83, 66, 12, 
    0, 37, 0, 0, 4, 0, 0, 
    
    -- channel=121
    2, 135, 0, 126, 0, 0, 17, 
    0, 0, 0, 0, 0, 110, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 130, 0, 0, 0, 
    67, 0, 0, 0, 56, 0, 0, 
    0, 0, 0, 85, 0, 0, 17, 
    0, 2, 91, 70, 66, 21, 8, 
    
    -- channel=122
    0, 0, 0, 116, 33, 17, 43, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    75, 0, 88, 166, 8, 13, 44, 
    2, 32, 6, 0, 0, 0, 0, 
    
    -- channel=123
    61, 91, 17, 33, 50, 60, 45, 
    0, 0, 76, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 88, 0, 19, 16, 
    0, 0, 0, 5, 0, 0, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=125
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    20, 0, 43, 16, 89, 0, 32, 
    0, 48, 59, 0, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 
    0, 11, 58, 0, 73, 4, 32, 
    0, 0, 6, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=130
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=132
    0, 0, 0, 150, 118, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 0, 0, 
    0, 0, 0, 0, 87, 0, 0, 
    0, 0, 278, 253, 0, 3, 0, 
    0, 273, 0, 0, 0, 0, 0, 
    
    -- channel=133
    49, 0, 0, 302, 0, 41, 34, 
    0, 133, 0, 20, 93, 0, 0, 
    46, 102, 0, 0, 0, 93, 0, 
    12, 0, 219, 13, 0, 79, 36, 
    0, 0, 0, 0, 328, 0, 0, 
    0, 0, 242, 0, 0, 0, 9, 
    0, 273, 0, 0, 0, 53, 0, 
    
    -- channel=134
    0, 0, 0, 0, 143, 0, 42, 
    0, 122, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 160, 0, 
    0, 0, 0, 92, 0, 0, 0, 
    0, 0, 60, 0, 0, 224, 0, 
    0, 0, 239, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 195, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 163, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    0, 0, 0, 0, 0, 0, 0, 
    104, 0, 0, 83, 0, 50, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 188, 53, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=137
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 243, 0, 0, 0, 0, 0, 
    0, 0, 81, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=140
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=141
    0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 48, 0, 88, 
    46, 0, 0, 0, 198, 33, 106, 
    59, 72, 0, 0, 0, 0, 0, 
    0, 47, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=142
    0, 0, 0, 0, 291, 0, 0, 
    0, 107, 98, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 81, 0, 0, 358, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    110, 0, 0, 6, 44, 0, 0, 
    
    -- channel=143
    0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 
    0, 0, 0, 95, 72, 0, 0, 
    0, 0, 211, 4, 0, 0, 0, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 33, 0, 0, 
    105, 0, 0, 0, 169, 0, 0, 
    88, 0, 0, 0, 0, 0, 0, 
    60, 122, 0, 4, 0, 0, 0, 
    143, 196, 0, 0, 0, 0, 0, 
    0, 95, 0, 0, 0, 5, 17, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=146
    230, 158, 89, 299, 165, 78, 190, 
    181, 360, 20, 0, 0, 0, 0, 
    0, 113, 0, 0, 79, 0, 0, 
    0, 145, 0, 0, 0, 0, 0, 
    0, 167, 0, 0, 43, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=147
    0, 0, 0, 146, 0, 4, 0, 
    0, 36, 0, 17, 67, 0, 0, 
    0, 0, 0, 0, 33, 0, 0, 
    0, 0, 19, 53, 0, 0, 20, 
    0, 68, 0, 0, 103, 0, 12, 
    0, 0, 162, 0, 0, 0, 0, 
    0, 0, 21, 18, 0, 30, 0, 
    
    -- channel=148
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=152
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=153
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 5, 25, 0, 
    
    -- channel=155
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=156
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=157
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=160
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=161
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    172, 0, 24, 0, 0, 0, 0, 
    0, 0, 126, 0, 31, 0, 58, 
    201, 0, 0, 0, 0, 0, 1, 
    60, 251, 0, 124, 0, 55, 47, 
    0, 473, 0, 23, 7, 14, 27, 
    
    -- channel=162
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 83, 0, 
    0, 0, 0, 29, 0, 59, 0, 
    0, 0, 0, 0, 0, 98, 0, 
    0, 0, 0, 0, 188, 0, 0, 
    0, 0, 359, 13, 0, 0, 0, 
    
    -- channel=163
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=165
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 12, 22, 0, 
    0, 0, 51, 8, 131, 61, 0, 
    22, 0, 0, 56, 0, 0, 0, 
    88, 188, 57, 70, 46, 90, 38, 
    226, 162, 186, 159, 189, 133, 154, 
    0, 216, 145, 64, 84, 81, 129, 
    
    -- channel=166
    136, 251, 25, 0, 0, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 35, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    84, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=167
    54, 70, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 59, 0, 54, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 267, 0, 0, 0, 0, 
    0, 0, 69, 0, 0, 0, 0, 
    
    -- channel=168
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 80, 
    0, 0, 0, 0, 0, 87, 0, 
    0, 11, 0, 0, 0, 49, 0, 
    0, 0, 218, 0, 0, 55, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    76, 51, 0, 0, 0, 0, 0, 
    
    -- channel=169
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=170
    0, 0, 0, 16, 0, 0, 0, 
    0, 0, 0, 0, 37, 9, 28, 
    69, 32, 47, 0, 31, 0, 0, 
    0, 0, 50, 64, 72, 0, 20, 
    0, 16, 0, 0, 41, 10, 0, 
    0, 103, 69, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=171
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=172
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 77, 0, 19, 0, 0, 
    
    -- channel=173
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 41, 33, 169, 
    0, 0, 203, 282, 236, 172, 76, 
    
    -- channel=174
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    3, 0, 0, 5, 0, 0, 65, 
    105, 35, 33, 0, 98, 22, 65, 
    57, 75, 89, 5, 158, 75, 0, 
    0, 88, 23, 18, 88, 21, 14, 
    0, 18, 102, 0, 16, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=177
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=178
    0, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 127, 0, 115, 0, 
    0, 0, 0, 297, 0, 101, 0, 
    0, 0, 0, 0, 0, 75, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=179
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=180
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=181
    0, 0, 0, 0, 0, 0, 0, 
    46, 0, 0, 0, 0, 0, 202, 
    0, 211, 0, 0, 156, 172, 0, 
    0, 115, 0, 0, 0, 197, 0, 
    0, 0, 68, 0, 0, 102, 0, 
    0, 0, 154, 0, 0, 0, 0, 
    101, 0, 11, 0, 0, 0, 0, 
    
    -- channel=182
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=183
    122, 317, 0, 0, 0, 24, 101, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 108, 
    0, 0, 0, 0, 0, 221, 181, 
    0, 0, 0, 164, 208, 139, 0, 
    
    -- channel=184
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=185
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=186
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=187
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 15, 27, 6, 
    
    -- channel=188
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=189
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=190
    0, 0, 0, 0, 0, 0, 0, 
    0, 117, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 46, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 56, 87, 87, 5, 
    
    -- channel=191
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=192
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 
    90, 0, 14, 0, 157, 86, 0, 
    17, 11, 0, 2, 0, 19, 0, 
    0, 60, 0, 0, 0, 0, 0, 
    128, 118, 461, 72, 113, 71, 44, 
    189, 222, 249, 98, 91, 79, 118, 
    
    -- channel=193
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=194
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=195
    0, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 142, 
    37, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 28, 
    27, 0, 0, 0, 8, 0, 16, 
    174, 0, 12, 98, 0, 92, 143, 
    340, 106, 0, 89, 54, 145, 81, 
    
    -- channel=196
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=197
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 
    0, 0, 0, 0, 0, 0, 41, 
    0, 0, 0, 0, 0, 26, 0, 
    0, 0, 0, 38, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=198
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=199
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 37, 210, 236, 
    88, 0, 8, 240, 283, 338, 232, 
    
    -- channel=200
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=201
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=202
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=203
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=204
    0, 82, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 
    0, 0, 15, 58, 65, 13, 0, 
    
    -- channel=205
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=206
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=207
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=208
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=209
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=211
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=212
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=213
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=214
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=215
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 200, 0, 0, 
    0, 0, 0, 0, 206, 0, 0, 
    0, 0, 193, 0, 20, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 
    194, 281, 0, 42, 0, 131, 96, 
    251, 17, 0, 59, 122, 136, 175, 
    
    -- channel=216
    0, 0, 0, 89, 43, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 
    0, 12, 0, 0, 21, 12, 0, 
    0, 0, 135, 62, 3, 84, 0, 
    0, 0, 14, 0, 150, 85, 0, 
    62, 0, 80, 25, 0, 0, 0, 
    0, 296, 0, 0, 0, 0, 0, 
    
    -- channel=217
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=218
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 79, 0, 
    0, 0, 0, 48, 0, 28, 0, 
    0, 0, 0, 160, 0, 0, 51, 
    0, 0, 0, 0, 10, 0, 0, 
    0, 0, 137, 61, 0, 0, 0, 
    0, 0, 124, 56, 0, 12, 0, 
    
    -- channel=219
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=220
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=221
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=222
    139, 57, 142, 149, 169, 64, 142, 
    31, 127, 67, 0, 0, 0, 0, 
    0, 0, 86, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 56, 0, 38, 26, 
    103, 0, 68, 96, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 
    
    -- channel=223
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=224
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=225
    0, 0, 0, 253, 179, 105, 121, 
    0, 57, 4, 0, 0, 0, 0, 
    0, 57, 46, 0, 0, 21, 0, 
    0, 64, 0, 56, 0, 0, 0, 
    0, 0, 0, 0, 157, 0, 0, 
    45, 0, 370, 173, 43, 38, 0, 
    0, 79, 0, 0, 0, 9, 0, 
    
    -- channel=226
    0, 64, 0, 0, 18, 57, 0, 
    12, 72, 65, 82, 7, 117, 33, 
    75, 0, 0, 164, 0, 94, 123, 
    149, 150, 0, 42, 35, 0, 22, 
    107, 139, 96, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=227
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=228
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=229
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=230
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=231
    84, 74, 0, 2, 0, 0, 188, 
    0, 0, 0, 0, 21, 0, 156, 
    0, 538, 0, 0, 99, 0, 0, 
    0, 0, 257, 3, 321, 0, 0, 
    0, 0, 74, 0, 0, 0, 25, 
    438, 0, 0, 140, 0, 0, 0, 
    386, 0, 0, 0, 0, 0, 0, 
    
    -- channel=232
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=233
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=234
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=235
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=236
    0, 0, 0, 25, 0, 0, 0, 
    0, 0, 0, 18, 7, 14, 0, 
    0, 75, 0, 0, 0, 0, 0, 
    0, 0, 95, 14, 0, 21, 0, 
    0, 0, 0, 1, 100, 0, 0, 
    0, 60, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=237
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 72, 
    0, 0, 0, 58, 0, 200, 0, 
    
    -- channel=238
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=239
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 187, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=240
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 96, 0, 0, 0, 
    0, 38, 0, 0, 0, 0, 0, 
    
    -- channel=241
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=242
    11, 12, 17, 27, 0, 7, 0, 
    0, 40, 0, 7, 0, 51, 0, 
    0, 0, 0, 70, 0, 0, 45, 
    0, 0, 0, 18, 0, 0, 52, 
    68, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=243
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 
    194, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 160, 
    0, 0, 0, 192, 236, 272, 289, 
    
    -- channel=244
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=246
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=248
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=249
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=250
    0, 0, 0, 20, 0, 136, 91, 
    269, 3, 5, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 
    0, 40, 180, 0, 94, 0, 35, 
    45, 0, 0, 83, 0, 0, 45, 
    129, 0, 0, 67, 51, 70, 126, 
    
    -- channel=251
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    319, 322, 130, 170, 0, 0, 124, 
    0, 141, 0, 0, 0, 0, 0, 
    0, 82, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=253
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 
    113, 104, 0, 63, 72, 127, 0, 
    17, 88, 0, 19, 80, 63, 0, 
    29, 0, 0, 0, 0, 0, 0, 
    0, 20, 124, 0, 0, 0, 0, 
    95, 0, 0, 0, 0, 0, 0, 
    
    -- channel=254
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=255
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
