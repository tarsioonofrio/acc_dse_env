library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_36k_layer0_entity5 is
    generic (
        BRAM_SIZE: string := 36Kb;
        BRAM_SIZE_ADD: integer := 8;
        DEVICE: string := 7SERIES;
        INPUT_SIZE : integer := 8;
        READ_WIDTH : integer := 0
        );
  
    port (reset   : in std_logic;
          clock   : in std_logic;
          chip_en : in std_logic;
          wr_en   : in std_logic;
          data_in : in std_logic_vector(INPUT_SIZE-1 downto 0);
          address : in std_logic_vector(BRAM_SIZE_ADD-1 downto 0);
  
          data_av  : out std_logic;
          data_out : out std_logic_vector(INPUT_SIZE-1 downto 0);
  
          n_read  : out std_logic_vector(31 downto 0);
          n_write : out std_logic_vector(31 downto 0)
          );
  end ifmap_36k_layer0_entity5;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => "7SERIES",             -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"009c00b000b300c000b900ab00ad00ad00af00b300b600b800b900b800b600b5",
       INIT_01 => X"00b300b300b700b900ba00ba00bb00bd00bb00bb00bc00c300c500c400ca00b7",
       INIT_02 => X"009b00b300b800c300be00a2009f00a400a300a500a900b000ab00ae00a400a7",
       INIT_03 => X"00ac00a600a800a600a900af00ab00a900aa00ae00bf00cc00ce00d000d700be",
       INIT_04 => X"009a00b200b900c400cb00c100b200a800a000af00be00c400c300c500be00bc",
       INIT_05 => X"00c400c300c200c300c400c600c100bf00c000c400cd00cd00ce00d000d700bf",
       INIT_06 => X"009a00b200bc00c300ca00c500bc0080006c0098009a009b009e009500950094",
       INIT_07 => X"00a700a100a300ad00a800a300ae009f00bc00d000cc00ce00cc00cd00d400bc",
       INIT_08 => X"009a00b100bb00bf00c600c400bd007e0080008b006a006b0073007800760071",
       INIT_09 => X"007700720072007e007600700088007000a000cb00c900ce00ce00cd00d600be",
       INIT_0A => X"009700ae00bb00bd00c500c800b7009300a900a8009100a500aa00920095009d",
       INIT_0B => X"00b400b200b000bd00b000b300bc00b100c400d000cf00d000d000d100d800be",
       INIT_0C => X"009800ac00b900bd00c200c6009300600095009700900098009800790080008b",
       INIT_0D => X"009c009700aa00a2009600ad009600a4009c00a600cc00d200d300cf00d400bc",
       INIT_0E => X"009b00ac00b600bb00c200b500770065007b008300830078009200870087007f",
       INIT_0F => X"007b007b0083007b006d0084007b009f007b008400bf00c700c900c900d000ba",
       INIT_10 => X"00a100af00b400b900c000ba00ab00af00a200a500ac00a600af00ac00ad00aa",
       INIT_11 => X"00ac00b200b200af00a300ac00b200be00ac00b000c800cd00c800c900d100b9",
       INIT_12 => X"00ac00b700b400ba00be00c000c200b700a000a500a200a3009f009e00a400a2",
       INIT_13 => X"00a700ae00ac00a200a000a300a500b600c800c600ca00cd00ca00ca00d000b8",
       INIT_14 => X"00b100c400ba00be00c000c100c100b700a300a700a5009f00a400a600aa00ac",
       INIT_15 => X"00a800a600a600ab00a800ad00ab00b200c700c600c700c700c800c800d000b8",
       INIT_16 => X"00b700cc00c300c800c900bb00be00c600c200c100c100c100c100c200c600c6",
       INIT_17 => X"00c600c300c300c600c500c400c400c500c900cb00c900c900ca00c800d100bb",
       INIT_18 => X"00b900cd00c600b200a6008d009a00c400ca00ca00c700c500c500c700c900ca",
       INIT_19 => X"00c900c700c600c400c400c600c700c600c700ca00cb00ce00cf00ce00d400bd",
       INIT_1A => X"00ba00d000c800a50090007c005f006b008f00b300c700c700c500c600c900cc",
       INIT_1B => X"00cc00cd00ce00cc00c900c900cd00cd00cc00cb00cb00cb00ca00ca00cf00b7",
       INIT_1C => X"00ba00d400d000cc00ce00c1008f005b00510065008e00b500c600cc00cf00cf",
       INIT_1D => X"00cf00cf00cf00ca00c500c500c600c500c500c500c500c500c400c500cc00b5",
       INIT_1E => X"00b800d600d200ce00d100d400cf00b300740053005d008000ae00cb00d200ce",
       INIT_1F => X"00cc00ca00ca00c900c600c700c900c900c800ca00c900c700c600c600cb00b4",
       INIT_20 => X"00ba00d700d600d500d600d600d400d900af005b004900560065008a00b500cc",
       INIT_21 => X"00d000cb00c700c600c700c900c900c800c800ca00c900c900ca00c800cc00b6",
       INIT_22 => X"00bb00d800d800d900db00d900d600d300cc007b00440052004f005100610082",
       INIT_23 => X"00a500bc00c900ca00c400c100c700c600c600c700c800c800c900c700cc00b6",
       INIT_24 => X"00bc00d900d500d600d800d800d600d200d4008800460053004e00500050004d",
       INIT_25 => X"00530066007e0097009f00b200c900cc00cb00c900c800c600c700c500c900b4",
       INIT_26 => X"00bb00da00d600d500d700d800d700d800cc0070002d0037003a0045004d0051",
       INIT_27 => X"0050004d0046003e003b004f007c00a000b500c400cd00cd00cb00c800ca00b4",
       INIT_28 => X"00bc00d800d200d100d300d600d400d4009a005f003a00210030003e0041004d",
       INIT_29 => X"00520054005400480038002f003f0048004e006b0084009e00b500c100ca00b6",
       INIT_2A => X"00b800d200ce00cf00d100d300d400c800910085008f0061002d0032002e005a",
       INIT_2B => X"0096009e007f004700610070005800410043008200a500a200a800b500c500b0",
       INIT_2C => X"00b700d200cd00d000d300d400d500d200d100d100d400bf00940093009300a6",
       INIT_2D => X"00c800d000c3009d00a600b500b400a2009f00b400c100c500c300c100c700b1",
       INIT_2E => X"00ae00c400c300c200c200be00bb00b900b800b500b700b500b200b000ae00ad",
       INIT_2F => X"00aa00a400a600ac00aa00a600aa00b000af00a5009d009b009d00a300af009e",
       INIT_30 => X"0070006c007000690067006400610060005c005a005e00570054005300570067",
       INIT_31 => X"00730070006f00700071007300740076007a007b007c007b0079007a0084007c",
       INIT_32 => X"00750073007100700071006f00710071006f0070006f006e006e006d006e006b",
       INIT_33 => X"00730073006c006e006f006d0068006b006d006e007000700064005f00620065",
       INIT_34 => X"007100660069006a006a00660061005d005f005e005900550052004e004f004e",
       INIT_35 => X"0050004f0047004400430041004100410041004200420041003c003700470064",
       INIT_36 => X"0054003c0041004000400040003e003c00420040003d00380039003c003d003f",
       INIT_37 => X"004000430041003b0038003a003b003c003a0039003800380038004800750080",
       INIT_38 => X"0053003b003f003e003f0041003d003f0043003e003c0039003a003a003c003d",
       INIT_39 => X"004100440040003e003d003c003e003d003a003a003d0041005b008800890063",
       INIT_3A => X"004f0035003d00390037003b003a003c003d003c00390037003c003e003d003f",
       INIT_3B => X"0043003f003c003b003e003e0040003f003e003c0047006e008e0077004f004a",
       INIT_3C => X"0052003a00420041003f003e003e003e003f003e0041004f004f004c004a004d",
       INIT_3D => X"005400500050004e004c003f003e004100420056007c008d0066004200400045",
       INIT_3E => X"004e0034003a003a003a003a003b0039003a003b003a00450047004700460045",
       INIT_3F => X"004800480049004a0049003f003f0044005a0080008000580042003f00410044",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INIT_40 => X"009500bb00c100cd00ca00b700b500b400b600bd00c100c000c000c000bd00bd",
       INIT_41 => X"00ba00b900bd00c000c100c100c000be00bb00bb00bc00c300ca00d100d400ab",
       INIT_42 => X"009d00cc00d700e300e000be00b300b300b300bb00c300c300bb00be00b400b7",
       INIT_43 => X"00bc00b700b800b700b900bf00bc00bc00be00c200d300e000df00de00e300b7",
       INIT_44 => X"009900c900d500db00df00d500c400b800b100c300d300d400d000d200cc00ca",
       INIT_45 => X"00d100d100d000d100d200d400d000d000d000d500de00df00da00d700e000b8",
       INIT_46 => X"00a600cf00d300de00e200dc00c900830077009e00a600b100b200a700a600ab",
       INIT_47 => X"00b700b200b200ba00b900ba00b400a500cf00e400dc00dd00e000df00e600ba",
       INIT_48 => X"00a700cb00ca00da00e000e100d6008e00990098007800810081007e007c0083",
       INIT_49 => X"008600840082008a00880088008d007b00ba00e300da00d900de00dc00e300b9",
       INIT_4A => X"00a400c900cb00d900dc00da00d100a500c400b5009c00b400b300a000a300ac",
       INIT_4B => X"00bf00c100be00c900bf00c000c600be00d400e100e100e100df00e100e800bc",
       INIT_4C => X"00a400c600c800d900d900d600ac0068009e00a500a600af00a50090009700a0",
       INIT_4D => X"00b200ad00bd00b600aa00b700ad00b900a600b200dc00e200dd00e000e700bc",
       INIT_4E => X"00a900c900c700d800da00cb0092006f00860095009d0090009b008f008f0090",
       INIT_4F => X"0093008e0094008e007f008d008e00b00089009500d100dc00d900dc00e400ba",
       INIT_50 => X"00b100ce00c700d900db00cd00c100c500b800b700bb00b800c000ba00bb00bd",
       INIT_51 => X"00c000c200c200bf00b200ba00bc00c800c100c600d600db00db00dd00e400b9",
       INIT_52 => X"00ba00d400c500d600d700d600dc00d200b900bb00b600ba00b600b400b900ba",
       INIT_53 => X"00c100c600c300b800b500b600b600c600de00de00dd00df00df00de00e300b7",
       INIT_54 => X"00bc00de00c800d800d700d400d600cc00b500b800b600b000b500b800bc00bf",
       INIT_55 => X"00bd00ba00b800b900b600b800ba00c900df00dd00dc00db00db00dc00e300b8",
       INIT_56 => X"00bf00e200cf00e000dc00d100d700de00d900d700d600d700d900db00df00df",
       INIT_57 => X"00df00dd00db00da00d800d600d900db00db00db00d900d600d700db00e300ba",
       INIT_58 => X"00bc00dc00d400ce00b5009900ac00d900e200e100dd00dc00de00df00e100e2",
       INIT_59 => X"00e100dd00dc00da00d900db00dc00da00d900dc00de00e000e000e000e600bb",
       INIT_5A => X"00bd00df00d600c1009d007e00630073009d00c600dd00dd00da00dc00df00e2",
       INIT_5B => X"00e200e000e100df00dc00dd00e000e000df00de00de00de00dd00dd00e200b7",
       INIT_5C => X"00bd00e200de00e900dc00c40092005a0054007100a100ca00da00e000e300e4",
       INIT_5D => X"00e200e100e000dc00d700d700d800d900d800d800d800d800d700da00e100b6",
       INIT_5E => X"00bb00e500e000ea00e100e100da00b300730058006a009100c000dd00e400e1",
       INIT_5F => X"00df00db00da00d900d600d600d900db00db00dd00dc00da00d900dc00e200b7",
       INIT_60 => X"00be00e900de00e900e400e200e000e100b500620050005b006a009200c000d9",
       INIT_61 => X"00e000e100dd00da00d900da00da00d900da00dd00dd00dd00dd00dc00e300bc",
       INIT_62 => X"00bf00ea00dd00e900e700e300e200dd00d500820049004f004b005000640088",
       INIT_63 => X"00ad00c800d700dc00d900d900df00de00dd00dd00db00db00da00db00e300bd",
       INIT_64 => X"00bd00e800d900e400e300e100e200dc00dd0090004a0050004a004c004e004c",
       INIT_65 => X"00530064008100a100b000c900e100e200df00dc00d900d700d700d900e100bb",
       INIT_66 => X"00bb00e800d700e100e000e100e300e200d5007700320038003b0045004d0052",
       INIT_67 => X"005000480042003f0041005b008500a200b800cc00da00df00dd00dd00e300bc",
       INIT_68 => X"00b700e700de00df00df00e600e400e100a20062003c0027003500430044004e",
       INIT_69 => X"005100520053004800390031003f0043004b006d008b00a800c600d700df00c3",
       INIT_6A => X"00b000e200e200de00de00e200e200d4009b008b0096006a003500390033005e",
       INIT_6B => X"009a00a10082004900630072005a00430045008600ab00a900b700c500d000be",
       INIT_6C => X"00af00e100e100df00df00de00de00de00de00e000e400cc009f009f00a000b3",
       INIT_6D => X"00d600dc00cf00a900b200c100c000ad00ab00c300d200d600d800d100d200bd",
       INIT_6E => X"00a600d400d700d100ce00cc00c900c700c700c300c500c200c000c100c200c4",
       INIT_6F => X"00c400c200c400ca00c800c400c800cd00ce00c500c000bf00c500c500c900b5",
       INIT_70 => X"006500780082007800760070006b006a006500620066006300620065006c0080",
       INIT_71 => X"0090009200920093009400960098009e00a400a600a800a800a800a500a70092",
       INIT_72 => X"006f008200860086008a008800890088008400860083007e007f008000830083",
       INIT_73 => X"008a0086007f008100810080007c007e00810082008400840077007300730060",
       INIT_74 => X"0068007100780078007a0076006c00640060005b005500590058005500570056",
       INIT_75 => X"0056004f0046004300420041003f003c003b003c003c003b00360032003f004b",
       INIT_76 => X"003d0037003d0039003a003f003b003600380033002f002f0030003200310032",
       INIT_77 => X"003300370035002f002d002e0032003700360034003400340030003a00680068",
       INIT_78 => X"0044003d0041003c003e003d00370039003d00380037003a003b003800380036",
       INIT_79 => X"0039003b0037003400330033003400340033003500370039004b00710078004b",
       INIT_7A => X"003e0034003b0035003900390034003600360032003000320039003800340035",
       INIT_7B => X"0039003600340033003600370035003000320034003d005f007c0065003e0032",
       INIT_7C => X"003e0035003a0037003b003d003c003c00390037003a004b004c004800440045",
       INIT_7D => X"004b004a004b00490046003a0037003500330045006b007f005b003a00360033",
       INIT_7E => X"004000330033002e0033003800390035003400330032003e0040003e003c0039",
       INIT_7F => X"003c003e00400040004000350034003700460067006900480035003200340032",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
