-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(36-1 downto 0);
        ADDR : in std_logic_vector(9-1 downto 0);
        DO   : out std_logic_vector(36-1 downto 0)
    );
    attribute dont_touch : string;
    attribute dont_touch of bram_single : entity is "true";
   end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(8-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);
    signal bram_di     : std_logic_vector(44-1 downto 0);
    signal bram_do     : std_logic_vector(44-1 downto 0);
    constant bram_par     : std_logic_vector(8-1 downto 0) := "00000000";

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
    bram_di <= bram_par & DI;
    DO <= bram_do(36-1 downto 0);


    MEM_IWGHT_LAYER0_INSTANCE0 : if BRAM_NAME = "iwght_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffec3affffffffffffea99ffffffff0000027e00000000fffff1ebffffffff",
            INIT_01 => X"00000453000000000000077300000000000002fb00000000fffff0f5ffffffff",
            INIT_02 => X"0000017e00000000fffffadbffffffff000031cf00000000000002f800000000",
            INIT_03 => X"0000052800000000000001ec00000000fffffd5bffffffff000017e900000000",
            INIT_04 => X"0000001f000000000000000100000000ffffffe3ffffffff0000000100000000",
            INIT_05 => X"0000002700000000ffffffdeffffffff00000005000000000000000400000000",
            INIT_06 => X"0000002700000000ffffffdcfffffffffffffff2ffffffffffffffd8ffffffff",
            INIT_07 => X"0000000700000000ffffffcefffffffffffffffcfffffffffffffffdffffffff",
            INIT_08 => X"000000290000000000000037000000000000000b00000000ffffffdbffffffff",
            INIT_09 => X"fffffff7ffffffff00000025000000000000002b000000000000003600000000",
            INIT_0A => X"ffffffecffffffff0000000000000000fffffffcffffffff0000000900000000",
            INIT_0B => X"fffffff1ffffffffffffffc3ffffffff0000002600000000ffffffe0ffffffff",
            INIT_0C => X"fffffffaffffffff000000210000000000000014000000000000003d00000000",
            INIT_0D => X"ffffffe7fffffffffffffffcffffffff0000000800000000ffffffbcffffffff",
            INIT_0E => X"fffffff6ffffffffffffffd3ffffffff0000000f000000000000001900000000",
            INIT_0F => X"ffffffefffffffff0000000b00000000fffffffcffffffff0000003800000000",
            INIT_10 => X"00000025000000000000003800000000ffffffd3ffffffffffffffe0ffffffff",
            INIT_11 => X"0000000f000000000000003c000000000000002800000000ffffffdbffffffff",
            INIT_12 => X"000000160000000000000016000000000000002d000000000000003000000000",
            INIT_13 => X"000000180000000000000007000000000000004300000000fffffff3ffffffff",
            INIT_14 => X"fffffff9ffffffff0000000400000000fffffff2fffffffffffffff8ffffffff",
            INIT_15 => X"000000040000000000000014000000000000000500000000ffffffe4ffffffff",
            INIT_16 => X"ffffffc4ffffffffffffffeaffffffff0000000700000000ffffffceffffffff",
            INIT_17 => X"ffffffd2ffffffffffffffdfffffffffffffffffffffffffffffffc0ffffffff",
            INIT_18 => X"00000011000000000000001900000000ffffffdaffffffffffffffdaffffffff",
            INIT_19 => X"0000003800000000fffffff4ffffffff00000013000000000000003700000000",
            INIT_1A => X"0000003400000000000000100000000000000015000000000000001c00000000",
            INIT_1B => X"ffffffe1ffffffff000000320000000000000031000000000000002500000000",
            INIT_1C => X"0000000b00000000ffffffe4ffffffff00000000000000000000001b00000000",
            INIT_1D => X"000000130000000000000036000000000000000f00000000fffffff4ffffffff",
            INIT_1E => X"fffffff3ffffffff000000140000000000000035000000000000000b00000000",
            INIT_1F => X"0000001000000000000000150000000000000035000000000000003100000000",
            INIT_20 => X"00000030000000000000001f000000000000003a00000000ffffffffffffffff",
            INIT_21 => X"fffffff2ffffffff0000001400000000fffffffdffffffffffffffe4ffffffff",
            INIT_22 => X"000000050000000000000009000000000000002200000000ffffffe6ffffffff",
            INIT_23 => X"ffffffe9ffffffff0000001e00000000fffffff5ffffffff0000000100000000",
            INIT_24 => X"ffffffddffffffff0000002900000000fffffff1ffffffffffffffd1ffffffff",
            INIT_25 => X"0000002800000000ffffffd4ffffffffffffffd5fffffffffffffffaffffffff",
            INIT_26 => X"ffffffe1ffffffff0000004400000000ffffffd1ffffffffffffffdbffffffff",
            INIT_27 => X"ffffffd4ffffffff000000110000000000000035000000000000000400000000",
            INIT_28 => X"0000000300000000ffffffeeffffffff0000000d000000000000002b00000000",
            INIT_29 => X"0000002d000000000000000700000000ffffffc2fffffffffffffff5ffffffff",
            INIT_2A => X"ffffffd5ffffffff0000001c000000000000000d00000000ffffffc8ffffffff",
            INIT_2B => X"0000000f00000000ffffffedffffffffffffffe8ffffffff0000003c00000000",
            INIT_2C => X"0000000c000000000000004f00000000ffffffeffffffffffffffff8ffffffff",
            INIT_2D => X"0000000800000000ffffffebffffffffffffffcbffffffffffffffddffffffff",
            INIT_2E => X"0000002800000000ffffffe3ffffffffffffffecffffffff0000000900000000",
            INIT_2F => X"ffffffe7ffffffffffffffb7ffffffff00000008000000000000004200000000",
            INIT_30 => X"00000001000000000000001200000000ffffffcbffffffff0000001000000000",
            INIT_31 => X"ffffffc5fffffffffffffff3ffffffff0000000b000000000000003800000000",
            INIT_32 => X"ffffffe2ffffffff0000002d000000000000001600000000ffffffd5ffffffff",
            INIT_33 => X"0000002800000000ffffffe6ffffffff0000001a000000000000000300000000",
            INIT_34 => X"ffffffe6ffffffff0000001f00000000fffffffaffffffff0000000200000000",
            INIT_35 => X"ffffffdbfffffffffffffffcfffffffffffffffbffffffff0000000400000000",
            INIT_36 => X"00000004000000000000000e00000000ffffffcfffffffff0000001d00000000",
            INIT_37 => X"ffffffd6ffffffff0000003c00000000ffffffeeffffffffffffffbeffffffff",
            INIT_38 => X"0000000400000000ffffffd4ffffffffffffffe6ffffffff0000002d00000000",
            INIT_39 => X"0000001e000000000000002c00000000ffffffcfffffffff0000002d00000000",
            INIT_3A => X"0000002800000000ffffffdeffffffff0000000f000000000000000000000000",
            INIT_3B => X"0000000400000000000000380000000000000034000000000000000400000000",
            INIT_3C => X"0000001f00000000fffffff1ffffffffffffffdaffffffff0000002000000000",
            INIT_3D => X"fffffffbfffffffffffffff4ffffffffffffffedffffffff0000000400000000",
            INIT_3E => X"fffffff2ffffffff000000190000000000000000000000000000000000000000",
            INIT_3F => X"fffffff1ffffffff0000001f00000000ffffffdbffffffffffffffe5ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe0ffffffffffffffd2ffffffff0000000500000000ffffffedffffffff",
            INIT_41 => X"fffffff1fffffffffffffffdffffffffffffffdcffffffff0000000a00000000",
            INIT_42 => X"fffffff3fffffffffffffff2ffffffff0000000e000000000000000300000000",
            INIT_43 => X"fffffff3ffffffffffffffe3ffffffffffffffcfffffffff0000000800000000",
            INIT_44 => X"0000000200000000ffffffd0ffffffffffffffe4ffffffffffffffe0ffffffff",
            INIT_45 => X"0000000a00000000fffffff5ffffffffffffffe0ffffffffffffffe6ffffffff",
            INIT_46 => X"0000001d000000000000000a0000000000000016000000000000001800000000",
            INIT_47 => X"ffffffe2ffffffffffffffe3ffffffff00000019000000000000000c00000000",
            INIT_48 => X"ffffffebffffffff00000006000000000000002200000000ffffffe6ffffffff",
            INIT_49 => X"fffffff6ffffffffffffffdaffffffff0000001400000000ffffffdbffffffff",
            INIT_4A => X"0000000100000000ffffffedffffffffffffffedffffffff0000000600000000",
            INIT_4B => X"ffffffd3ffffffff0000002700000000ffffffedffffffff0000000000000000",
            INIT_4C => X"ffffffccffffffffffffffedffffffff0000002e00000000ffffffdcffffffff",
            INIT_4D => X"ffffffd2ffffffffffffffe4ffffffff0000002d00000000ffffffd5ffffffff",
            INIT_4E => X"ffffffc5fffffffffffffff0fffffffffffffff5ffffffff0000001d00000000",
            INIT_4F => X"0000004200000000fffffffcfffffffffffffffaffffffffffffffe8ffffffff",
            INIT_50 => X"ffffffceffffffffffffffc2ffffffff00000008000000000000002500000000",
            INIT_51 => X"0000001c00000000fffffff0fffffffffffffff3ffffffffffffffdcffffffff",
            INIT_52 => X"ffffffefffffffff00000048000000000000000a00000000ffffffffffffffff",
            INIT_53 => X"fffffff1ffffffff0000001900000000ffffffd6ffffffffffffffe9ffffffff",
            INIT_54 => X"0000000e0000000000000040000000000000003800000000fffffff6ffffffff",
            INIT_55 => X"ffffffdcffffffff0000000e000000000000000600000000ffffffeeffffffff",
            INIT_56 => X"fffffff3ffffffff000000090000000000000003000000000000000500000000",
            INIT_57 => X"00000034000000000000003300000000ffffffdeffffffff0000000300000000",
            INIT_58 => X"0000000300000000fffffffbfffffffffffffff0ffffffff0000002500000000",
            INIT_59 => X"ffffffe7fffffffffffffff3ffffffff00000029000000000000003000000000",
            INIT_5A => X"fffffff9ffffffff0000000b00000000ffffffdfffffffffffffffd2ffffffff",
            INIT_5B => X"ffffffdcffffffff0000000600000000ffffffddffffffffffffffd3ffffffff",
            INIT_5C => X"ffffffe5ffffffffffffffd5ffffffff00000021000000000000000a00000000",
            INIT_5D => X"ffffffd8ffffffffffffffccffffffff0000000300000000ffffffd8ffffffff",
            INIT_5E => X"0000002900000000ffffffe3fffffffffffffff4ffffffff0000000700000000",
            INIT_5F => X"ffffffebfffffffffffffff4fffffffffffffffdffffffff0000002a00000000",
            INIT_60 => X"0000002d000000000000002f000000000000001400000000ffffffdcffffffff",
            INIT_61 => X"0000000700000000fffffff0ffffffff0000002b000000000000003200000000",
            INIT_62 => X"0000000b00000000000000340000000000000015000000000000002700000000",
            INIT_63 => X"00000013000000000000000a00000000fffffff5ffffffff0000004500000000",
            INIT_64 => X"ffffffe8ffffffff0000004400000000ffffffffffffffff0000001300000000",
            INIT_65 => X"0000001800000000ffffffeeffffffffffffffe4fffffffffffffff3ffffffff",
            INIT_66 => X"ffffffccffffffffffffffd8ffffffffffffffd4ffffffff0000001a00000000",
            INIT_67 => X"ffffffecffffffff0000000500000000ffffffe1fffffffffffffff5ffffffff",
            INIT_68 => X"fffffffafffffffffffffffbfffffffffffffff3ffffffff0000000300000000",
            INIT_69 => X"ffffffddffffffffffffffdfffffffff0000001e00000000ffffffdcffffffff",
            INIT_6A => X"00000012000000000000002c00000000fffffffdffffffff0000000800000000",
            INIT_6B => X"00000006000000000000002d0000000000000028000000000000001500000000",
            INIT_6C => X"0000001a000000000000000b00000000ffffffd3ffffffff0000001e00000000",
            INIT_6D => X"00000000000000000000001700000000ffffffd5ffffffff0000002b00000000",
            INIT_6E => X"ffffffc8ffffffff0000001100000000ffffffebffffffffffffffceffffffff",
            INIT_6F => X"ffffffdbffffffffffffffbfffffffff00000006000000000000001a00000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE0 : if BRAM_NAME = "iwght_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00001eac00000000000001350000000000000c2900000000000001eb00000000",
            INIT_01 => X"fffffb4ffffffffffffffb8bffffffff000013af0000000000000c1600000000",
            INIT_02 => X"0000194d00000000fffffb30ffffffff0000044200000000000042b300000000",
            INIT_03 => X"ffffe13affffffff0000044f000000000000165b000000000000090500000000",
            INIT_04 => X"0000000f00000000ffffffe0ffffffff0000000100000000ffffffeaffffffff",
            INIT_05 => X"0000001e0000000000000001000000000000001100000000ffffffdeffffffff",
            INIT_06 => X"000000430000000000000029000000000000000700000000ffffffdcffffffff",
            INIT_07 => X"ffffffefffffffff0000002b0000000000000047000000000000001400000000",
            INIT_08 => X"ffffffd5ffffffff0000000e0000000000000028000000000000004800000000",
            INIT_09 => X"ffffffedffffffffffffffe2ffffffff0000000a000000000000002400000000",
            INIT_0A => X"0000001b00000000ffffffdeffffffff0000000400000000ffffffdbffffffff",
            INIT_0B => X"ffffffdcffffffff00000020000000000000000700000000fffffff1ffffffff",
            INIT_0C => X"fffffffafffffffffffffff4ffffffff0000002c00000000ffffffe8ffffffff",
            INIT_0D => X"fffffff7ffffffff00000007000000000000000600000000fffffff9ffffffff",
            INIT_0E => X"000000000000000000000000000000000000000c00000000ffffffe9ffffffff",
            INIT_0F => X"00000056000000000000007c000000000000006c000000000000000800000000",
            INIT_10 => X"0000006200000000000000530000000000000098000000000000007100000000",
            INIT_11 => X"0000000300000000ffffffe2ffffffff00000022000000000000008d00000000",
            INIT_12 => X"ffffffbeffffffffffffffcbffffffffffffffe3ffffffffffffffc6ffffffff",
            INIT_13 => X"fffffff8ffffffffffffffeaffffffff00000003000000000000000000000000",
            INIT_14 => X"0000006600000000ffffffecffffffff00000032000000000000006800000000",
            INIT_15 => X"00000014000000000000004e000000000000000a000000000000003e00000000",
            INIT_16 => X"fffffff1fffffffffffffff6ffffffffffffffdbffffffff0000001e00000000",
            INIT_17 => X"fffffffcffffffff0000001200000000ffffffe8ffffffffffffffddffffffff",
            INIT_18 => X"fffffffaffffffff0000000000000000fffffff6ffffffff0000001d00000000",
            INIT_19 => X"00000004000000000000001a0000000000000019000000000000001400000000",
            INIT_1A => X"ffffffdcffffffff0000002500000000ffffffbaffffffffffffffeaffffffff",
            INIT_1B => X"0000001e00000000ffffffe8ffffffff00000024000000000000001d00000000",
            INIT_1C => X"ffffffd1ffffffff0000002c00000000ffffffebfffffffffffffffeffffffff",
            INIT_1D => X"ffffffc3ffffffffffffffc2ffffffffffffffecffffffffffffffd0ffffffff",
            INIT_1E => X"ffffffe5ffffffffffffffdefffffffffffffff8ffffffffffffffb8ffffffff",
            INIT_1F => X"000000110000000000000026000000000000001d00000000fffffff2ffffffff",
            INIT_20 => X"ffffffe3ffffffffffffffe9ffffffff00000008000000000000002600000000",
            INIT_21 => X"fffffffffffffffffffffff5ffffffff00000003000000000000002700000000",
            INIT_22 => X"0000001100000000ffffffd9ffffffff00000009000000000000003500000000",
            INIT_23 => X"fffffff5ffffffff0000000700000000ffffffffffffffffffffffe5ffffffff",
            INIT_24 => X"0000002100000000fffffff6fffffffffffffff9ffffffff0000002400000000",
            INIT_25 => X"ffffffdcfffffffffffffffdffffffffffffffefffffffffffffffd5ffffffff",
            INIT_26 => X"0000002200000000fffffff4ffffffffffffffe5ffffffff0000000d00000000",
            INIT_27 => X"00000026000000000000000400000000fffffff1ffffffff0000001c00000000",
            INIT_28 => X"ffffffdaffffffff000000070000000000000005000000000000001900000000",
            INIT_29 => X"ffffffe6ffffffffffffffffffffffffffffffd0ffffffff0000000300000000",
            INIT_2A => X"ffffffe8ffffffffffffffe4fffffffffffffff2fffffffffffffffaffffffff",
            INIT_2B => X"00000001000000000000002c000000000000002600000000ffffffdcffffffff",
            INIT_2C => X"00000055000000000000005900000000ffffffe9fffffffffffffff4ffffffff",
            INIT_2D => X"0000001b00000000fffffffdffffffffffffffebffffffff0000007e00000000",
            INIT_2E => X"0000000e00000000ffffff9fffffffffffffff86ffffffffffffff73ffffffff",
            INIT_2F => X"ffffffeffffffffffffffffffffffffffffffff4ffffffff0000001700000000",
            INIT_30 => X"000000210000000000000005000000000000001100000000ffffffe1ffffffff",
            INIT_31 => X"fffffff9ffffffff000000090000000000000018000000000000001f00000000",
            INIT_32 => X"ffffffe0ffffffffffffffd1ffffffff0000001100000000ffffffdbffffffff",
            INIT_33 => X"000000200000000000000003000000000000002a00000000ffffffd4ffffffff",
            INIT_34 => X"ffffffccffffffffffffffd8ffffffffffffffc2fffffffffffffffaffffffff",
            INIT_35 => X"fffffff5ffffffffffffffc5fffffffffffffff3fffffffffffffffcffffffff",
            INIT_36 => X"00000005000000000000002e0000000000000008000000000000001b00000000",
            INIT_37 => X"0000002d00000000000000390000000000000039000000000000003400000000",
            INIT_38 => X"00000009000000000000000c0000000000000038000000000000002d00000000",
            INIT_39 => X"ffffffcfffffffffffffffaaffffffffffffffd8ffffffff0000000a00000000",
            INIT_3A => X"fffffffdfffffffffffffff0ffffffff00000025000000000000000700000000",
            INIT_3B => X"ffffffdeffffffffffffffecffffffff0000000a00000000ffffffe0ffffffff",
            INIT_3C => X"ffffffceffffffffffffffc7ffffffffffffffefffffffffffffffdcffffffff",
            INIT_3D => X"000000020000000000000000000000000000001000000000fffffffcffffffff",
            INIT_3E => X"00000028000000000000000e000000000000002700000000fffffff0ffffffff",
            INIT_3F => X"fffffff9ffffffff000000060000000000000022000000000000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff6ffffffff0000001b00000000fffffff4ffffffff0000001200000000",
            INIT_41 => X"00000062000000000000004d00000000ffffffecfffffffffffffff1ffffffff",
            INIT_42 => X"000000560000000000000059000000000000001a000000000000005f00000000",
            INIT_43 => X"000000000000000000000007000000000000001700000000fffffff1ffffffff",
            INIT_44 => X"ffffffdbffffffff0000000700000000fffffff7fffffffffffffff4ffffffff",
            INIT_45 => X"0000000600000000fffffffefffffffffffffff1fffffffffffffff9ffffffff",
            INIT_46 => X"0000001c00000000fffffff0ffffffff0000000e00000000fffffff8ffffffff",
            INIT_47 => X"00000061000000000000007100000000ffffffe2fffffffffffffff2ffffffff",
            INIT_48 => X"0000000800000000000000500000000000000001000000000000004f00000000",
            INIT_49 => X"ffffffe8ffffffffffffffdcffffffffffffff8bffffffffffffff9affffffff",
            INIT_4A => X"ffffffdffffffffffffffff4ffffffff00000024000000000000001500000000",
            INIT_4B => X"ffffffe7ffffffffffffffd7ffffffffffffffd0fffffffffffffffcffffffff",
            INIT_4C => X"ffffffdcffffffffffffffdfffffffff0000001c00000000ffffffe4ffffffff",
            INIT_4D => X"00000009000000000000000c00000000ffffffd7fffffffffffffff5ffffffff",
            INIT_4E => X"0000001d000000000000003c000000000000001200000000fffffffeffffffff",
            INIT_4F => X"0000000d00000000000000070000000000000023000000000000002600000000",
            INIT_50 => X"ffffffe6ffffffffffffffcffffffffffffffff1fffffffffffffff6ffffffff",
            INIT_51 => X"ffffffdcfffffffffffffff6ffffffffffffffd4ffffffff0000000200000000",
            INIT_52 => X"000000180000000000000017000000000000000c00000000ffffffd5ffffffff",
            INIT_53 => X"ffffffe4ffffffff0000001300000000ffffffe9ffffffff0000000900000000",
            INIT_54 => X"0000000f0000000000000015000000000000001c00000000ffffffdcffffffff",
            INIT_55 => X"fffffff0ffffffff0000001f000000000000001000000000ffffffe4ffffffff",
            INIT_56 => X"00000005000000000000001200000000ffffffe8ffffffff0000001f00000000",
            INIT_57 => X"000000090000000000000003000000000000000a000000000000000200000000",
            INIT_58 => X"0000000700000000000000050000000000000000000000000000001800000000",
            INIT_59 => X"00000012000000000000001200000000ffffffd2ffffffffffffffddffffffff",
            INIT_5A => X"00000044000000000000001000000000ffffffeaffffffff0000000200000000",
            INIT_5B => X"0000000d00000000fffffffcffffffff00000050000000000000000900000000",
            INIT_5C => X"0000002600000000000000000000000000000009000000000000003900000000",
            INIT_5D => X"ffffffd1ffffffffffffffe3ffffffffffffffdefffffffffffffffcffffffff",
            INIT_5E => X"0000000900000000fffffff0ffffffffffffffe9ffffffffffffffe6ffffffff",
            INIT_5F => X"000000160000000000000013000000000000000a00000000fffffffcffffffff",
            INIT_60 => X"ffffffd0ffffffffffffffcaffffffffffffffd7ffffffff0000000f00000000",
            INIT_61 => X"00000007000000000000001b00000000ffffffb9ffffffffffffffebffffffff",
            INIT_62 => X"0000001500000000fffffffbffffffff0000000800000000ffffffdcffffffff",
            INIT_63 => X"ffffffe3ffffffff00000014000000000000001700000000ffffffeeffffffff",
            INIT_64 => X"0000003d0000000000000028000000000000001e000000000000000500000000",
            INIT_65 => X"000000ab000000000000006b0000000000000078000000000000008b00000000",
            INIT_66 => X"0000005d000000000000003c0000000000000021000000000000008500000000",
            INIT_67 => X"0000001c00000000ffffffe2ffffffff0000001a000000000000001700000000",
            INIT_68 => X"ffffffeafffffffffffffffaffffffff0000000a000000000000003100000000",
            INIT_69 => X"ffffffdafffffffffffffffcffffffff0000000d000000000000002800000000",
            INIT_6A => X"fffffff8ffffffffffffffe6ffffffffffffffddffffffff0000000a00000000",
            INIT_6B => X"fffffff7fffffffffffffffeffffffff0000001d000000000000002100000000",
            INIT_6C => X"0000000000000000ffffffecffffffffffffffbaffffffff0000001d00000000",
            INIT_6D => X"00000003000000000000001e000000000000001100000000ffffffe2ffffffff",
            INIT_6E => X"ffffffffffffffff00000033000000000000000b000000000000000400000000",
            INIT_6F => X"0000000100000000fffffffbffffffff0000002e00000000ffffffe3ffffffff",
            INIT_70 => X"0000000400000000ffffffc6ffffffffffffffe4ffffffffffffffd3ffffffff",
            INIT_71 => X"fffffffaffffffffffffffe8ffffffffffffffd2ffffffffffffffe6ffffffff",
            INIT_72 => X"fffffff3ffffffff0000000500000000ffffffe4fffffffffffffff6ffffffff",
            INIT_73 => X"0000000e000000000000001300000000fffffffeffffffffffffffd7ffffffff",
            INIT_74 => X"00000015000000000000001c0000000000000010000000000000000800000000",
            INIT_75 => X"00000004000000000000002000000000ffffffe7ffffffff0000002800000000",
            INIT_76 => X"00000000000000000000000200000000ffffffc8ffffffffffffffe0ffffffff",
            INIT_77 => X"fffffff9ffffffffffffffefffffffff00000009000000000000000100000000",
            INIT_78 => X"0000001700000000ffffffe7ffffffff00000011000000000000000800000000",
            INIT_79 => X"ffffffebfffffffffffffff9ffffffff00000012000000000000002a00000000",
            INIT_7A => X"00000030000000000000002200000000fffffff0fffffffffffffff1ffffffff",
            INIT_7B => X"0000000800000000ffffffc6ffffffff0000000200000000fffffff8ffffffff",
            INIT_7C => X"000000140000000000000006000000000000001d00000000fffffff6ffffffff",
            INIT_7D => X"fffffff2ffffffff0000000c00000000ffffffceffffffff0000001300000000",
            INIT_7E => X"ffffffeeffffffff00000006000000000000003100000000ffffffe9ffffffff",
            INIT_7F => X"ffffffd1ffffffffffffffe2ffffffffffffffd9fffffffffffffffcffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE1 : if BRAM_NAME = "iwght_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000100000000ffffffd5ffffffffffffffedffffffffffffffd7ffffffff",
            INIT_01 => X"ffffffe7ffffffff00000005000000000000001b000000000000001000000000",
            INIT_02 => X"0000002a000000000000002d000000000000002a000000000000002400000000",
            INIT_03 => X"0000000400000000000000010000000000000010000000000000002700000000",
            INIT_04 => X"ffffffdcffffffffffffffe4ffffffff0000001300000000fffffffbffffffff",
            INIT_05 => X"ffffffe6ffffffff000000060000000000000012000000000000002f00000000",
            INIT_06 => X"00000020000000000000002500000000ffffffedffffffffffffffe5ffffffff",
            INIT_07 => X"0000000d000000000000000b00000000fffffff5ffffffffffffffd7ffffffff",
            INIT_08 => X"ffffffecffffffff0000001200000000ffffffeaffffffff0000000200000000",
            INIT_09 => X"ffffffb2ffffffffffffffbeffffffffffffffa3ffffffffffffff98ffffffff",
            INIT_0A => X"fffffffcffffffffffffffcfffffffffffffffd2ffffffffffffffa1ffffffff",
            INIT_0B => X"0000000100000000000000300000000000000028000000000000001600000000",
            INIT_0C => X"00000048000000000000000a0000000000000013000000000000002500000000",
            INIT_0D => X"ffffffccfffffffffffffff1ffffffffffffffc8ffffffff0000002a00000000",
            INIT_0E => X"ffffffdaffffffffffffffe3ffffffffffffffeeffffffffffffffc2ffffffff",
            INIT_0F => X"00000016000000000000000600000000ffffffd1ffffffffffffffccffffffff",
            INIT_10 => X"00000004000000000000000a0000000000000027000000000000001f00000000",
            INIT_11 => X"0000001700000000ffffffe5ffffffff00000001000000000000000700000000",
            INIT_12 => X"0000001a00000000ffffffebfffffffffffffff9ffffffff0000000e00000000",
            INIT_13 => X"00000032000000000000000f00000000fffffffbffffffff0000002000000000",
            INIT_14 => X"ffffffd8ffffffffffffffe9fffffffffffffff1ffffffffffffffdaffffffff",
            INIT_15 => X"000000220000000000000000000000000000000d00000000ffffffddffffffff",
            INIT_16 => X"00000020000000000000003e000000000000003700000000ffffffecffffffff",
            INIT_17 => X"0000005c0000000000000024000000000000006f000000000000006200000000",
            INIT_18 => X"fffffff3ffffffff000000170000000000000061000000000000006500000000",
            INIT_19 => X"fffffff2ffffffffffffffedfffffffffffffff0ffffffffffffffe9ffffffff",
            INIT_1A => X"ffffffdcffffffffffffffb6fffffffffffffff2ffffffffffffffbdffffffff",
            INIT_1B => X"00000024000000000000000d00000000fffffff7ffffffff0000000b00000000",
            INIT_1C => X"fffffffffffffffffffffffeffffffffffffffe6ffffffff0000001f00000000",
            INIT_1D => X"ffffffedfffffffffffffff0ffffffff00000004000000000000000500000000",
            INIT_1E => X"ffffffe3ffffffff0000001600000000ffffffeaffffffff0000001e00000000",
            INIT_1F => X"0000003200000000000000360000000000000010000000000000001200000000",
            INIT_20 => X"0000004800000000000000270000000000000044000000000000004500000000",
            INIT_21 => X"ffffffd9ffffffffffffffcbffffffff00000039000000000000003d00000000",
            INIT_22 => X"ffffffe5ffffffffffffffe1ffffffff0000002300000000ffffffdeffffffff",
            INIT_23 => X"0000004000000000ffffffcdffffffffffffffb8ffffffff0000000900000000",
            INIT_24 => X"0000007d00000000000000720000000000000049000000000000004f00000000",
            INIT_25 => X"000000350000000000000036000000000000003a000000000000005a00000000",
            INIT_26 => X"0000001a00000000ffffffe0ffffffff00000000000000000000000900000000",
            INIT_27 => X"0000000c0000000000000024000000000000000f000000000000000300000000",
            INIT_28 => X"0000000d000000000000000d0000000000000000000000000000000d00000000",
            INIT_29 => X"ffffffdbffffffff00000015000000000000001b000000000000001e00000000",
            INIT_2A => X"ffffffdafffffffffffffffdffffffffffffffd1ffffffffffffffdfffffffff",
            INIT_2B => X"ffffffe0ffffffff0000000a00000000fffffff6ffffffff0000000300000000",
            INIT_2C => X"ffffffeffffffffffffffff1ffffffffffffffddffffffff0000001100000000",
            INIT_2D => X"ffffffaeffffffffffffffbcffffffffffffffccffffffffffffffbdffffffff",
            INIT_2E => X"ffffffe7ffffffffffffffd7ffffffffffffffe4ffffffffffffffafffffffff",
            INIT_2F => X"000000010000000000000020000000000000002b00000000fffffff2ffffffff",
            INIT_30 => X"00000020000000000000001100000000fffffffcffffffff0000002700000000",
            INIT_31 => X"0000001c00000000ffffffedffffffffffffffd2ffffffff0000001e00000000",
            INIT_32 => X"ffffffdafffffffffffffffefffffffffffffff9ffffffffffffffd0ffffffff",
            INIT_33 => X"00000048000000000000003200000000fffffff8fffffffffffffff0ffffffff",
            INIT_34 => X"ffffffffffffffffffffffe3fffffffffffffffcffffffff0000005d00000000",
            INIT_35 => X"fffffff6fffffffffffffff5ffffffffffffffedfffffffffffffff8ffffffff",
            INIT_36 => X"fffffff2ffffffff00000011000000000000001900000000fffffff3ffffffff",
            INIT_37 => X"fffffff5ffffffff00000019000000000000000900000000fffffff8ffffffff",
            INIT_38 => X"ffffffabffffffff0000000800000000fffffffbffffffff0000002a00000000",
            INIT_39 => X"fffffff2ffffffff0000000000000000ffffffc8ffffffffffffffb4ffffffff",
            INIT_3A => X"ffffffeeffffffffffffffceffffffffffffffc0ffffffffffffffd7ffffffff",
            INIT_3B => X"000000290000000000000001000000000000001800000000ffffffd9ffffffff",
            INIT_3C => X"ffffffd7ffffffff0000000300000000fffffff7fffffffffffffffdffffffff",
            INIT_3D => X"00000006000000000000001900000000ffffffd8ffffffff0000001400000000",
            INIT_3E => X"ffffffe6ffffffff0000000e00000000ffffffe2ffffffff0000002700000000",
            INIT_3F => X"ffffffe1ffffffffffffffaefffffffffffffff9ffffffff0000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffffffffffd4fffffffffffffff5ffffffffffffffeeffffffff",
            INIT_41 => X"ffffffd7ffffffff0000000e00000000ffffffe3ffffffffffffffe4ffffffff",
            INIT_42 => X"0000000800000000fffffff9ffffffff0000000700000000fffffffdffffffff",
            INIT_43 => X"0000000200000000ffffffbdffffffffffffffefffffffffffffffdcffffffff",
            INIT_44 => X"00000012000000000000001400000000ffffffefffffffffffffffbfffffffff",
            INIT_45 => X"0000004c000000000000005100000000fffffffaffffffff0000003700000000",
            INIT_46 => X"0000002300000000000000310000000000000056000000000000005200000000",
            INIT_47 => X"ffffffffffffffff000000260000000000000034000000000000000700000000",
            INIT_48 => X"00000008000000000000000900000000ffffffdaffffffffffffffd5ffffffff",
            INIT_49 => X"000000150000000000000009000000000000000600000000ffffffefffffffff",
            INIT_4A => X"0000000f00000000ffffffe9ffffffff0000000700000000ffffffe3ffffffff",
            INIT_4B => X"00000003000000000000000300000000fffffff8ffffffff0000002a00000000",
            INIT_4C => X"0000001900000000000000310000000000000028000000000000002700000000",
            INIT_4D => X"00000033000000000000003f0000000000000032000000000000002000000000",
            INIT_4E => X"0000000400000000fffffff8ffffffff00000041000000000000000f00000000",
            INIT_4F => X"0000000500000000fffffff4ffffffff0000000400000000ffffffd1ffffffff",
            INIT_50 => X"ffffffc7fffffffffffffff3ffffffff00000009000000000000002500000000",
            INIT_51 => X"0000002400000000fffffffeffffffff00000015000000000000002e00000000",
            INIT_52 => X"0000002800000000fffffffbffffffff0000004d000000000000001b00000000",
            INIT_53 => X"0000000c000000000000000b0000000000000012000000000000001d00000000",
            INIT_54 => X"000000420000000000000030000000000000002b000000000000001900000000",
            INIT_55 => X"ffffffe6ffffffff000000190000000000000018000000000000004400000000",
            INIT_56 => X"ffffffe2ffffffffffffffaaffffffff0000000000000000ffffffd5ffffffff",
            INIT_57 => X"000000000000000000000000000000000000001d00000000ffffffc5ffffffff",
            INIT_58 => X"0000000f00000000ffffffdbffffffffffffffe7fffffffffffffff5ffffffff",
            INIT_59 => X"0000001600000000ffffffd9fffffffffffffffdfffffffffffffff2ffffffff",
            INIT_5A => X"0000000400000000ffffffedffffffff0000000c000000000000000000000000",
            INIT_5B => X"fffffff1fffffffffffffff6ffffffff00000001000000000000000c00000000",
            INIT_5C => X"fffffffaffffffff0000001700000000ffffffe3ffffffffffffffe1ffffffff",
            INIT_5D => X"00000020000000000000001f00000000fffffff6ffffffff0000000f00000000",
            INIT_5E => X"000000180000000000000014000000000000000200000000ffffffeeffffffff",
            INIT_5F => X"0000003a000000000000000a0000000000000021000000000000003b00000000",
            INIT_60 => X"ffffffc2ffffffff00000001000000000000004f000000000000004f00000000",
            INIT_61 => X"ffffffe3ffffffff00000033000000000000000400000000ffffffb2ffffffff",
            INIT_62 => X"fffffffbffffffff000000280000000000000026000000000000004d00000000",
            INIT_63 => X"ffffffe6ffffffff0000000000000000ffffffd4ffffffff0000000100000000",
            INIT_64 => X"0000000000000000000000260000000000000033000000000000001b00000000",
            INIT_65 => X"00000008000000000000000d0000000000000000000000000000000900000000",
            INIT_66 => X"00000021000000000000000400000000fffffff6ffffffff0000001c00000000",
            INIT_67 => X"000000450000000000000043000000000000001c00000000fffffff7ffffffff",
            INIT_68 => X"0000004d00000000000000220000000000000045000000000000002300000000",
            INIT_69 => X"fffffffaffffffffffffffe0ffffffff00000029000000000000006d00000000",
            INIT_6A => X"fffffff6ffffffffffffffd9ffffffffffffffddffffffff0000002500000000",
            INIT_6B => X"ffffffbaffffffff0000000a00000000ffffffa8ffffffffffffffeaffffffff",
            INIT_6C => X"0000000700000000ffffffc0ffffffffffffffefffffffffffffffe2ffffffff",
            INIT_6D => X"0000003e00000000000000120000000000000009000000000000000a00000000",
            INIT_6E => X"00000011000000000000001f0000000000000004000000000000002b00000000",
            INIT_6F => X"0000002d00000000000000340000000000000015000000000000001200000000",
            INIT_70 => X"0000003600000000000000070000000000000039000000000000000d00000000",
            INIT_71 => X"00000018000000000000003e0000000000000042000000000000001f00000000",
            INIT_72 => X"00000010000000000000000c000000000000003f000000000000003e00000000",
            INIT_73 => X"ffffffecffffffffffffffffffffffffffffffe1ffffffff0000000600000000",
            INIT_74 => X"00000034000000000000000f00000000fffffff1ffffffffffffffe5ffffffff",
            INIT_75 => X"0000000b0000000000000008000000000000006c000000000000002600000000",
            INIT_76 => X"0000001e00000000000000000000000000000005000000000000002600000000",
            INIT_77 => X"ffffffd2ffffffffffffff91ffffffffffffffcdffffffffffffffc2ffffffff",
            INIT_78 => X"ffffffb2ffffffffffffffaeffffffffffffffb6ffffffffffffffc2ffffffff",
            INIT_79 => X"0000001000000000ffffffdeffffffffffffffdbffffffffffffffa0ffffffff",
            INIT_7A => X"ffffffeeffffffff0000000a000000000000000400000000ffffffddffffffff",
            INIT_7B => X"ffffffeaffffffffffffffb6fffffffffffffffcffffffff0000000a00000000",
            INIT_7C => X"0000001c000000000000001500000000ffffffe8ffffffffffffffd1ffffffff",
            INIT_7D => X"ffffffe8ffffffff00000069000000000000003e000000000000004100000000",
            INIT_7E => X"0000001b000000000000002000000000ffffffd2ffffffffffffffe3ffffffff",
            INIT_7F => X"00000011000000000000001d000000000000000000000000ffffffeaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE1;


    MEM_IWGHT_LAYER1_INSTANCE2 : if BRAM_NAME = "iwght_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000250000000000000038000000000000001000000000fffffff4ffffffff",
            INIT_01 => X"ffffffddffffffffffffffebffffffff0000001100000000ffffffe7ffffffff",
            INIT_02 => X"ffffffdcfffffffffffffff0ffffffff00000000000000000000000900000000",
            INIT_03 => X"00000038000000000000001f0000000000000029000000000000003700000000",
            INIT_04 => X"0000003a000000000000001c000000000000004f000000000000004700000000",
            INIT_05 => X"0000000b000000000000001b0000000000000016000000000000000e00000000",
            INIT_06 => X"0000000300000000ffffffdcffffffffffffffe8fffffffffffffff1ffffffff",
            INIT_07 => X"fffffff1ffffffffffffffecffffffff00000025000000000000001c00000000",
            INIT_08 => X"ffffffe2fffffffffffffff1fffffffffffffff1ffffffffffffffebffffffff",
            INIT_09 => X"00000004000000000000002f0000000000000010000000000000000f00000000",
            INIT_0A => X"ffffffd5ffffffffffffffdaffffffff0000002000000000ffffffe0ffffffff",
            INIT_0B => X"00000014000000000000000b000000000000001d00000000ffffffebffffffff",
            INIT_0C => X"0000006100000000000000400000000000000037000000000000001c00000000",
            INIT_0D => X"fffffff2ffffffff0000000a0000000000000021000000000000003900000000",
            INIT_0E => X"fffffffdffffffff0000000400000000ffffffdcffffffffffffffc5ffffffff",
            INIT_0F => X"0000004900000000000000000000000000000029000000000000000900000000",
            INIT_10 => X"0000004b000000000000001c0000000000000031000000000000003a00000000",
            INIT_11 => X"000000290000000000000048000000000000002f000000000000005500000000",
            INIT_12 => X"fffffff6ffffffff00000037000000000000002600000000fffffff6ffffffff",
            INIT_13 => X"ffffffcbffffffffffffffddffffffffffffffe9ffffffff0000001c00000000",
            INIT_14 => X"ffffffeaffffffffffffffeaffffffffffffffeaffffffffffffffd9ffffffff",
            INIT_15 => X"00000025000000000000001b0000000000000009000000000000000600000000",
            INIT_16 => X"00000006000000000000000600000000fffffffbffffffff0000002500000000",
            INIT_17 => X"0000001b00000000ffffffe2ffffffffffffffd9fffffffffffffff0ffffffff",
            INIT_18 => X"ffffffb4ffffffff0000000f00000000ffffffe5ffffffff0000000c00000000",
            INIT_19 => X"0000001000000000ffffffe5fffffffffffffffdffffffffffffffc9ffffffff",
            INIT_1A => X"0000001a000000000000000d000000000000001e000000000000000600000000",
            INIT_1B => X"ffffffe9ffffffff0000001200000000fffffff3ffffffff0000003700000000",
            INIT_1C => X"0000000b0000000000000003000000000000000e00000000fffffff3ffffffff",
            INIT_1D => X"000000360000000000000034000000000000001200000000ffffffeeffffffff",
            INIT_1E => X"fffffff3ffffffffffffffffffffffffffffffe1fffffffffffffffdffffffff",
            INIT_1F => X"fffffffcffffffff0000002d00000000ffffffebffffffffffffffefffffffff",
            INIT_20 => X"000000290000000000000011000000000000001e000000000000000000000000",
            INIT_21 => X"0000000b000000000000000c000000000000000b00000000ffffffe8ffffffff",
            INIT_22 => X"ffffffedfffffffffffffff7ffffffff0000001e000000000000002100000000",
            INIT_23 => X"ffffffd9ffffffff0000000c00000000ffffffeeffffffff0000000400000000",
            INIT_24 => X"0000001c00000000ffffffeaffffffffffffffe0fffffffffffffffcffffffff",
            INIT_25 => X"00000000000000000000001900000000ffffffe8fffffffffffffff1ffffffff",
            INIT_26 => X"ffffffd1ffffffffffffffe8ffffffffffffffb8ffffffff0000001200000000",
            INIT_27 => X"ffffffa0ffffffffffffffa9ffffffffffffffb7ffffffffffffffdcffffffff",
            INIT_28 => X"0000001100000000ffffffe3ffffffffffffffa8ffffffffffffffc0ffffffff",
            INIT_29 => X"0000000700000000ffffffeeffffffffffffffa5ffffffff0000000800000000",
            INIT_2A => X"0000000400000000ffffffcaffffffffffffffc7ffffffffffffff82ffffffff",
            INIT_2B => X"fffffff6ffffffff0000003000000000ffffffe3ffffffffffffffdbffffffff",
            INIT_2C => X"ffffffe0ffffffff0000001a0000000000000014000000000000000100000000",
            INIT_2D => X"fffffffcffffffffffffffffffffffff00000015000000000000001600000000",
            INIT_2E => X"fffffff5ffffffffffffffd1fffffffffffffff6ffffffffffffffd5ffffffff",
            INIT_2F => X"ffffffe0ffffffff0000000a000000000000003a00000000ffffffbfffffffff",
            INIT_30 => X"0000003100000000ffffffbffffffffffffffff4ffffffff0000002f00000000",
            INIT_31 => X"fffffff0ffffffff00000012000000000000002f00000000ffffffe7ffffffff",
            INIT_32 => X"ffffffb5fffffffffffffff3ffffffffffffffedffffffff0000000d00000000",
            INIT_33 => X"ffffffe8ffffffffffffffc1ffffffffffffffd9ffffffffffffffd8ffffffff",
            INIT_34 => X"ffffffa7ffffffffffffffecfffffffffffffff2ffffffffffffffdcffffffff",
            INIT_35 => X"ffffffbbffffffffffffffd9ffffffff0000000000000000ffffffe1ffffffff",
            INIT_36 => X"0000000200000000000000320000000000000040000000000000000500000000",
            INIT_37 => X"ffffffd6fffffffffffffffcffffffffffffffe5ffffffff0000000200000000",
            INIT_38 => X"000000290000000000000040000000000000004a00000000ffffffc8ffffffff",
            INIT_39 => X"00000027000000000000004e0000000000000043000000000000005000000000",
            INIT_3A => X"ffffffdefffffffffffffff6ffffffff00000041000000000000004a00000000",
            INIT_3B => X"ffffffe6ffffffff0000001a000000000000001d00000000ffffffe9ffffffff",
            INIT_3C => X"0000000800000000ffffffe9ffffffff0000000d000000000000001100000000",
            INIT_3D => X"0000000e00000000fffffff7ffffffffffffffdaffffffff0000000100000000",
            INIT_3E => X"ffffffcdfffffffffffffff0ffffffff0000000b00000000ffffffb2ffffffff",
            INIT_3F => X"00000007000000000000001b0000000000000048000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff4ffffffff00000012000000000000001a00000000fffffffcffffffff",
            INIT_41 => X"ffffffd0ffffffff0000000400000000fffffffcffffffff0000000b00000000",
            INIT_42 => X"00000020000000000000000400000000ffffffe8ffffffff0000001600000000",
            INIT_43 => X"0000001700000000fffffff0ffffffff0000001e000000000000003000000000",
            INIT_44 => X"ffffffcbffffffffffffffbbffffffffffffffedffffffff0000002500000000",
            INIT_45 => X"fffffff2ffffffffffffffacffffffffffffffe2ffffffffffffffd3ffffffff",
            INIT_46 => X"ffffffd5ffffffff0000001d00000000ffffffe6fffffffffffffff8ffffffff",
            INIT_47 => X"ffffffc7fffffffffffffff3fffffffffffffff5ffffffffffffffddffffffff",
            INIT_48 => X"0000001f00000000000000080000000000000030000000000000001b00000000",
            INIT_49 => X"000000010000000000000016000000000000002b00000000fffffffcffffffff",
            INIT_4A => X"ffffff91ffffffffffffffc0ffffffffffffffe2fffffffffffffff9ffffffff",
            INIT_4B => X"ffffffccffffffffffffffafffffffffffffffa0ffffffffffffffedffffffff",
            INIT_4C => X"ffffffcdffffffffffffffefffffffffffffffadffffffffffffffa5ffffffff",
            INIT_4D => X"ffffffe0fffffffffffffff3ffffffff0000002200000000ffffffefffffffff",
            INIT_4E => X"00000031000000000000000f0000000000000044000000000000002d00000000",
            INIT_4F => X"0000000e00000000000000320000000000000029000000000000000600000000",
            INIT_50 => X"0000001f000000000000000000000000fffffff9fffffffffffffff5ffffffff",
            INIT_51 => X"000000120000000000000011000000000000002c000000000000002300000000",
            INIT_52 => X"0000001b000000000000000a0000000000000000000000000000001d00000000",
            INIT_53 => X"0000000800000000fffffff3fffffffffffffffaffffffffffffffe1ffffffff",
            INIT_54 => X"fffffffafffffffffffffff0ffffffffffffffe3ffffffffffffffd5ffffffff",
            INIT_55 => X"0000000a000000000000001300000000ffffffbeffffffffffffffc0ffffffff",
            INIT_56 => X"ffffffc4ffffffffffffffd2ffffffffffffffecffffffff0000001600000000",
            INIT_57 => X"ffffffc7ffffffffffffffafffffffffffffffa0ffffffffffffffbeffffffff",
            INIT_58 => X"ffffffaaffffffffffffffdfffffffffffffffc8ffffffffffffffbaffffffff",
            INIT_59 => X"ffffffe3ffffffffffffffcbfffffffffffffff5ffffffffffffffd5ffffffff",
            INIT_5A => X"ffffffe2ffffffffffffffe2ffffffff00000012000000000000000300000000",
            INIT_5B => X"00000008000000000000000c00000000ffffffe1ffffffff0000001700000000",
            INIT_5C => X"ffffffd2ffffffffffffffd9fffffffffffffff7ffffffffffffffe7ffffffff",
            INIT_5D => X"0000002900000000ffffffe4fffffffffffffffcfffffffffffffff5ffffffff",
            INIT_5E => X"fffffffafffffffffffffff2ffffffffffffffd7ffffffffffffffe0ffffffff",
            INIT_5F => X"ffffffe8ffffffff0000000c00000000fffffffeffffffff0000002300000000",
            INIT_60 => X"ffffffd0ffffffff00000011000000000000000500000000ffffffd7ffffffff",
            INIT_61 => X"ffffffffffffffffffffffedffffffffffffffceffffffffffffffd7ffffffff",
            INIT_62 => X"ffffffddffffffff00000009000000000000000300000000fffffff0ffffffff",
            INIT_63 => X"0000000b00000000ffffffedffffffffffffffbfffffffffffffffc2ffffffff",
            INIT_64 => X"ffffffd7ffffffff0000000000000000ffffffedffffffffffffffebffffffff",
            INIT_65 => X"00000036000000000000002f000000000000003d00000000ffffffe8ffffffff",
            INIT_66 => X"0000002200000000000000270000000000000000000000000000001900000000",
            INIT_67 => X"ffffffb7ffffffffffffffdbffffffff00000038000000000000003b00000000",
            INIT_68 => X"ffffffe3ffffffff00000009000000000000002e00000000ffffffd3ffffffff",
            INIT_69 => X"ffffffd6ffffffff0000003f000000000000002d000000000000002a00000000",
            INIT_6A => X"ffffffe5ffffffffffffffe6fffffffffffffff6fffffffffffffff6ffffffff",
            INIT_6B => X"0000002500000000ffffffe9ffffffff0000000c000000000000000800000000",
            INIT_6C => X"ffffffe9ffffffff00000024000000000000002d000000000000001800000000",
            INIT_6D => X"ffffffe2ffffffff0000001300000000fffffffcffffffffffffffedffffffff",
            INIT_6E => X"0000000200000000ffffffd9fffffffffffffff7ffffffffffffffdeffffffff",
            INIT_6F => X"0000001e00000000fffffff6ffffffff0000002000000000fffffff2ffffffff",
            INIT_70 => X"fffffffdffffffff0000002400000000fffffffbffffffff0000001000000000",
            INIT_71 => X"0000001200000000000000260000000000000025000000000000001400000000",
            INIT_72 => X"000000190000000000000033000000000000003b000000000000002f00000000",
            INIT_73 => X"ffffffedffffffff00000013000000000000001c000000000000002000000000",
            INIT_74 => X"0000001300000000ffffffdfffffffffffffffdbfffffffffffffffcffffffff",
            INIT_75 => X"0000002d00000000fffffff5ffffffff0000000c000000000000002500000000",
            INIT_76 => X"0000000100000000ffffffd7ffffffffffffffe7fffffffffffffff5ffffffff",
            INIT_77 => X"0000000100000000ffffffffffffffff0000000000000000ffffffdfffffffff",
            INIT_78 => X"00000011000000000000001500000000fffffff0ffffffff0000002100000000",
            INIT_79 => X"00000018000000000000000000000000fffffff1ffffffff0000001800000000",
            INIT_7A => X"00000000000000000000003a000000000000000d000000000000003500000000",
            INIT_7B => X"fffffff0ffffffff0000000f00000000fffffff4ffffffff0000003100000000",
            INIT_7C => X"ffffffffffffffffffffffe1ffffffff0000001f000000000000002000000000",
            INIT_7D => X"fffffffeffffffffffffffeeffffffff0000000d000000000000001000000000",
            INIT_7E => X"fffffff9ffffffff000000240000000000000016000000000000002900000000",
            INIT_7F => X"fffffff1ffffffff00000013000000000000000a000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE2;


    MEM_IWGHT_LAYER1_INSTANCE3 : if BRAM_NAME = "iwght_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffcaffffffffffffffc3ffffffffffffffe8fffffffffffffff1ffffffff",
            INIT_01 => X"0000002b000000000000000800000000fffffff1ffffffff0000000100000000",
            INIT_02 => X"0000001200000000ffffffe6ffffffff0000002900000000ffffffedffffffff",
            INIT_03 => X"0000001400000000ffffffffffffffff00000007000000000000000600000000",
            INIT_04 => X"0000002900000000fffffffcfffffffffffffff8ffffffff0000000800000000",
            INIT_05 => X"0000005f000000000000005c0000000000000053000000000000002e00000000",
            INIT_06 => X"0000003b000000000000000d0000000000000035000000000000006900000000",
            INIT_07 => X"ffffffdbffffffffffffffd1fffffffffffffff6fffffffffffffff2ffffffff",
            INIT_08 => X"ffffffc2fffffffffffffffffffffffffffffff8ffffffffffffffddffffffff",
            INIT_09 => X"00000003000000000000001a00000000ffffffffffffffffffffffd1ffffffff",
            INIT_0A => X"0000000900000000ffffffe8ffffffff00000008000000000000001400000000",
            INIT_0B => X"0000000000000000ffffffdefffffffffffffff6fffffffffffffff3ffffffff",
            INIT_0C => X"0000003b0000000000000010000000000000002300000000ffffffdeffffffff",
            INIT_0D => X"0000002b000000000000001e0000000000000058000000000000005100000000",
            INIT_0E => X"0000000800000000ffffffeafffffffffffffffeffffffff0000001b00000000",
            INIT_0F => X"0000001300000000fffffffbffffffffffffffd9fffffffffffffff8ffffffff",
            INIT_10 => X"0000000e00000000ffffffcbfffffffffffffffffffffffffffffffdffffffff",
            INIT_11 => X"ffffffe0ffffffffffffffdeffffffffffffffc7ffffffffffffffe1ffffffff",
            INIT_12 => X"ffffffebffffffffffffffddffffffffffffffedffffffffffffffe7ffffffff",
            INIT_13 => X"ffffffd5ffffffffffffffe9ffffffffffffffecffffffff0000000500000000",
            INIT_14 => X"0000000b00000000ffffffeeffffffff00000009000000000000000800000000",
            INIT_15 => X"0000002000000000ffffffeeffffffffffffffdfffffffff0000000500000000",
            INIT_16 => X"ffffffe3ffffffff0000000a00000000ffffffecfffffffffffffff9ffffffff",
            INIT_17 => X"000000250000000000000026000000000000001400000000ffffffe8ffffffff",
            INIT_18 => X"fffffff9ffffffff000000200000000000000024000000000000000500000000",
            INIT_19 => X"0000002d0000000000000016000000000000001f000000000000000600000000",
            INIT_1A => X"0000002c000000000000000a0000000000000027000000000000001b00000000",
            INIT_1B => X"fffffffcffffffffffffffeffffffffffffffff0ffffffff0000003200000000",
            INIT_1C => X"fffffff6ffffffffffffffe3ffffffff0000000e00000000fffffff7ffffffff",
            INIT_1D => X"fffffffeffffffffffffffd2ffffffff0000000c00000000ffffffdcffffffff",
            INIT_1E => X"0000002b00000000000000280000000000000047000000000000001400000000",
            INIT_1F => X"00000002000000000000001d000000000000000d00000000ffffffe2ffffffff",
            INIT_20 => X"fffffffeffffffff000000060000000000000001000000000000000e00000000",
            INIT_21 => X"ffffffd4fffffffffffffffbfffffffffffffff0fffffffffffffffbffffffff",
            INIT_22 => X"0000002400000000ffffffffffffffff00000003000000000000002100000000",
            INIT_23 => X"0000000000000000fffffff9ffffffff0000000e000000000000001500000000",
            INIT_24 => X"ffffffd2ffffffffffffffe6fffffffffffffff1fffffffffffffff7ffffffff",
            INIT_25 => X"fffffffbffffffffffffffd2fffffffffffffffaffffffffffffffe7ffffffff",
            INIT_26 => X"0000000d00000000ffffffe1ffffffffffffffb4ffffffffffffffcfffffffff",
            INIT_27 => X"fffffffeffffffff0000001a00000000fffffff4ffffffff0000001900000000",
            INIT_28 => X"fffffff0ffffffff0000001b00000000ffffffd9ffffffffffffffe4ffffffff",
            INIT_29 => X"ffffffb4ffffffffffffff9bffffffffffffffefffffffffffffffc0ffffffff",
            INIT_2A => X"ffffffe0fffffffffffffff0ffffffffffffffc9ffffffffffffffc6ffffffff",
            INIT_2B => X"0000000e0000000000000025000000000000000f000000000000002100000000",
            INIT_2C => X"0000000f00000000000000220000000000000029000000000000003c00000000",
            INIT_2D => X"ffffffc7ffffffffffffffeeffffffffffffffe8ffffffff0000004e00000000",
            INIT_2E => X"ffffffddfffffffffffffff2ffffffffffffffcfffffffffffffffd3ffffffff",
            INIT_2F => X"00000000000000000000001f00000000ffffffccffffffffffffffccffffffff",
            INIT_30 => X"0000000e00000000ffffffeeffffffffffffffeaffffffff0000000700000000",
            INIT_31 => X"fffffff9ffffffffffffffebffffffffffffffecffffffffffffffd9ffffffff",
            INIT_32 => X"000000250000000000000007000000000000003b00000000ffffffffffffffff",
            INIT_33 => X"0000000400000000fffffffbffffffff00000013000000000000000e00000000",
            INIT_34 => X"0000002500000000fffffff5ffffffff0000001000000000ffffffebffffffff",
            INIT_35 => X"fffffffafffffffffffffff7ffffffff0000001a00000000fffffffbffffffff",
            INIT_36 => X"00000021000000000000000d000000000000001a00000000ffffffd9ffffffff",
            INIT_37 => X"ffffffc1ffffffffffffffbcffffffffffffff9fffffffff0000000a00000000",
            INIT_38 => X"ffffffecffffffffffffffe4ffffffff0000001100000000fffffffbffffffff",
            INIT_39 => X"00000030000000000000002300000000fffffff1ffffffffffffffeaffffffff",
            INIT_3A => X"0000002000000000fffffff7ffffffffffffffe9ffffffff0000000600000000",
            INIT_3B => X"00000025000000000000001500000000fffffffdffffffffffffffebffffffff",
            INIT_3C => X"ffffffd9ffffffffffffffebffffffffffffffdbffffffff0000001100000000",
            INIT_3D => X"00000028000000000000001f00000000ffffffe5ffffffffffffffefffffffff",
            INIT_3E => X"ffffffd5ffffffffffffffebffffffff00000028000000000000002c00000000",
            INIT_3F => X"ffffffe4fffffffffffffff3ffffffffffffffd6fffffffffffffff0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001b000000000000000c00000000ffffffd2ffffffffffffffbbffffffff",
            INIT_41 => X"0000002f000000000000001e00000000ffffffd1ffffffffffffffdaffffffff",
            INIT_42 => X"00000050000000000000001b00000000ffffffffffffffff0000001a00000000",
            INIT_43 => X"ffffffd9ffffffff0000003e0000000000000019000000000000000200000000",
            INIT_44 => X"00000020000000000000001700000000fffffff1ffffffffffffffd2ffffffff",
            INIT_45 => X"00000030000000000000001300000000ffffffffffffffffffffffe3ffffffff",
            INIT_46 => X"00000028000000000000003d000000000000001d000000000000000600000000",
            INIT_47 => X"ffffffb4fffffffffffffffafffffffffffffffbffffffff0000000a00000000",
            INIT_48 => X"fffffff7fffffffffffffff9ffffffffffffffe9ffffffffffffffbeffffffff",
            INIT_49 => X"0000000100000000ffffffd9ffffffffffffffd2ffffffffffffffbeffffffff",
            INIT_4A => X"ffffffefffffffff0000002600000000fffffff6ffffffff0000001500000000",
            INIT_4B => X"fffffff4fffffffffffffffeffffffff0000002200000000ffffffe6ffffffff",
            INIT_4C => X"0000003a000000000000001100000000fffffff7fffffffffffffff9ffffffff",
            INIT_4D => X"00000043000000000000005a0000000000000048000000000000003500000000",
            INIT_4E => X"fffffff1ffffffff000000400000000000000040000000000000004400000000",
            INIT_4F => X"000000050000000000000008000000000000002e000000000000002000000000",
            INIT_50 => X"0000000700000000fffffffbfffffffffffffffeffffffff0000000700000000",
            INIT_51 => X"fffffffdfffffffffffffffbffffffffffffffc0ffffffff0000001400000000",
            INIT_52 => X"0000001100000000ffffffe8ffffffff0000001a000000000000001a00000000",
            INIT_53 => X"0000000b00000000ffffffe4ffffffff0000001600000000fffffffaffffffff",
            INIT_54 => X"0000001d0000000000000027000000000000000c000000000000000200000000",
            INIT_55 => X"0000002000000000ffffffcfffffffffffffffe6ffffffff0000000300000000",
            INIT_56 => X"ffffffedffffffff000000150000000000000024000000000000003700000000",
            INIT_57 => X"ffffffbeffffffffffffffc5ffffffffffffffbcffffffff0000002100000000",
            INIT_58 => X"0000002700000000fffffff0ffffffff00000010000000000000003100000000",
            INIT_59 => X"ffffffecfffffffffffffff7ffffffff00000010000000000000001200000000",
            INIT_5A => X"ffffffe7fffffffffffffff3ffffffff0000000100000000fffffff5ffffffff",
            INIT_5B => X"ffffffcdffffffffffffffebffffffffffffffb5ffffffffffffffdbffffffff",
            INIT_5C => X"fffffff9fffffffffffffff8ffffffff0000001000000000ffffffe2ffffffff",
            INIT_5D => X"0000000000000000fffffff1fffffffffffffffdffffffffffffffc2ffffffff",
            INIT_5E => X"0000000300000000ffffffeafffffffffffffff7fffffffffffffff6ffffffff",
            INIT_5F => X"0000001400000000ffffffe8fffffffffffffffbffffffff0000001200000000",
            INIT_60 => X"0000001d0000000000000028000000000000002000000000fffffff3ffffffff",
            INIT_61 => X"00000002000000000000001500000000ffffffe2fffffffffffffff1ffffffff",
            INIT_62 => X"ffffffdeffffffff00000006000000000000000700000000ffffffedffffffff",
            INIT_63 => X"ffffffdfffffffffffffff76ffffffffffffffbfffffffffffffffe1ffffffff",
            INIT_64 => X"ffffffbfffffffffffffffa9ffffffffffffff94ffffffffffffffabffffffff",
            INIT_65 => X"00000006000000000000000800000000ffffffb0ffffffffffffff9dffffffff",
            INIT_66 => X"ffffffeefffffffffffffff6ffffffff00000016000000000000002000000000",
            INIT_67 => X"ffffffd2ffffffffffffffd5ffffffffffffffd9ffffffffffffffe7ffffffff",
            INIT_68 => X"ffffffb1ffffffffffffffaeffffffffffffffcfffffffffffffffc3ffffffff",
            INIT_69 => X"ffffffc5ffffffffffffff99ffffffffffffffa8ffffffffffffffc7ffffffff",
            INIT_6A => X"fffffff1ffffffff0000000700000000fffffff7ffffffff0000000f00000000",
            INIT_6B => X"ffffffe2ffffffff0000001400000000ffffffdbffffffff0000000d00000000",
            INIT_6C => X"ffffffd9ffffffffffffffe1fffffffffffffff8fffffffffffffff2ffffffff",
            INIT_6D => X"0000000500000000ffffffeaffffffffffffffedfffffffffffffffdffffffff",
            INIT_6E => X"0000000600000000fffffff1ffffffffffffffdfffffffff0000000700000000",
            INIT_6F => X"0000001200000000ffffffffffffffffffffffedffffffff0000001400000000",
            INIT_70 => X"ffffffeffffffffffffffffdffffffff0000002a00000000ffffffe1ffffffff",
            INIT_71 => X"0000000000000000fffffffdffffffff0000000d00000000fffffff7ffffffff",
            INIT_72 => X"000000040000000000000000000000000000000000000000fffffffbffffffff",
            INIT_73 => X"00000042000000000000004c0000000000000053000000000000004e00000000",
            INIT_74 => X"00000029000000000000004f0000000000000018000000000000004600000000",
            INIT_75 => X"00000015000000000000003100000000fffffffeffffffff0000006100000000",
            INIT_76 => X"000000110000000000000010000000000000003a000000000000003800000000",
            INIT_77 => X"ffffff9dffffffffffffffaeffffffff00000023000000000000002200000000",
            INIT_78 => X"ffffffcafffffffffffffff9ffffffffffffffd1ffffffffffffffb0ffffffff",
            INIT_79 => X"ffffffeaffffffffffffffc4ffffffffffffffd4ffffffffffffffbfffffffff",
            INIT_7A => X"0000000c000000000000001000000000ffffffe5ffffffff0000002100000000",
            INIT_7B => X"00000032000000000000003400000000ffffffeeffffffffffffffefffffffff",
            INIT_7C => X"fffffff1ffffffff0000000000000000ffffffdeffffffffffffffdaffffffff",
            INIT_7D => X"ffffffe0ffffffff00000000000000000000001f000000000000000b00000000",
            INIT_7E => X"000000000000000000000027000000000000001800000000ffffffedffffffff",
            INIT_7F => X"0000003b000000000000003f00000000fffffff3ffffffff0000002d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE3;


    MEM_IWGHT_LAYER1_INSTANCE4 : if BRAM_NAME = "iwght_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe1ffffffff000000100000000000000013000000000000003100000000",
            INIT_01 => X"ffffffdfffffffffffffffd5ffffffffffffffceffffffff0000000400000000",
            INIT_02 => X"0000000400000000ffffffc6fffffffffffffff8ffffffffffffffe4ffffffff",
            INIT_03 => X"ffffffe3ffffffff000000070000000000000003000000000000001f00000000",
            INIT_04 => X"fffffff8ffffffff000000020000000000000018000000000000001900000000",
            INIT_05 => X"0000001e000000000000002000000000fffffff7fffffffffffffff2ffffffff",
            INIT_06 => X"fffffff8ffffffff00000004000000000000000500000000fffffff3ffffffff",
            INIT_07 => X"0000004b0000000000000053000000000000002900000000fffffffdffffffff",
            INIT_08 => X"0000001e0000000000000064000000000000006e000000000000001e00000000",
            INIT_09 => X"fffffff5ffffffffffffffcdffffffff00000045000000000000004d00000000",
            INIT_0A => X"ffffffe8fffffffffffffff6ffffffffffffffd5ffffffffffffffebffffffff",
            INIT_0B => X"0000004500000000ffffffc6ffffffffffffffcbfffffffffffffff1ffffffff",
            INIT_0C => X"0000002f000000000000003e000000000000005a000000000000005100000000",
            INIT_0D => X"0000005a00000000000000500000000000000015000000000000005f00000000",
            INIT_0E => X"000000210000000000000021000000000000000f000000000000002100000000",
            INIT_0F => X"fffffff2ffffffff00000011000000000000001a000000000000002000000000",
            INIT_10 => X"0000004600000000000000370000000000000021000000000000000700000000",
            INIT_11 => X"0000002300000000000000080000000000000013000000000000004000000000",
            INIT_12 => X"00000001000000000000001100000000ffffffdfffffffff0000000a00000000",
            INIT_13 => X"0000000500000000ffffffe4fffffffffffffffafffffffffffffffdffffffff",
            INIT_14 => X"ffffffeeffffffff0000001500000000ffffffd7ffffffff0000001e00000000",
            INIT_15 => X"ffffffcbffffffffffffffdeffffffffffffffc3ffffffffffffffc5ffffffff",
            INIT_16 => X"ffffffd6ffffffffffffffe8ffffffffffffffddffffffffffffffd2ffffffff",
            INIT_17 => X"fffffff4ffffffffffffffdfffffffffffffffd5fffffffffffffff7ffffffff",
            INIT_18 => X"ffffffe8ffffffffffffffebfffffffffffffffdffffffffffffffedffffffff",
            INIT_19 => X"ffffffc3ffffffffffffffe0fffffffffffffffaffffffffffffffe7ffffffff",
            INIT_1A => X"0000000000000000ffffffd0ffffffffffffffeaffffffff0000001300000000",
            INIT_1B => X"0000000e000000000000001200000000ffffffdbffffffffffffffe9ffffffff",
            INIT_1C => X"fffffff4ffffffff000000060000000000000014000000000000002800000000",
            INIT_1D => X"ffffffeefffffffffffffff0ffffffffffffffc0ffffffffffffffd0ffffffff",
            INIT_1E => X"0000000b000000000000001d000000000000000c00000000fffffff8ffffffff",
            INIT_1F => X"fffffff5ffffffff0000000500000000ffffffefffffffff0000001b00000000",
            INIT_20 => X"0000003d000000000000003a000000000000001a000000000000001e00000000",
            INIT_21 => X"0000001e00000000000000030000000000000020000000000000004800000000",
            INIT_22 => X"ffffffecffffffff00000010000000000000004200000000fffffffdffffffff",
            INIT_23 => X"ffffffeffffffffffffffff3fffffffffffffffdffffffff0000002a00000000",
            INIT_24 => X"ffffffe7ffffffff0000001f00000000ffffffddffffffff0000001a00000000",
            INIT_25 => X"0000001300000000000000110000000000000011000000000000001a00000000",
            INIT_26 => X"ffffffedffffffff000000370000000000000062000000000000004100000000",
            INIT_27 => X"fffffff9ffffffff00000012000000000000001600000000fffffffbffffffff",
            INIT_28 => X"fffffff3ffffffff0000002a0000000000000007000000000000000000000000",
            INIT_29 => X"ffffffe4ffffffff0000001200000000fffffffcffffffff0000000c00000000",
            INIT_2A => X"00000005000000000000000400000000fffffff2ffffffff0000001b00000000",
            INIT_2B => X"fffffff8ffffffff0000002a0000000000000023000000000000001b00000000",
            INIT_2C => X"0000001b0000000000000000000000000000000400000000fffffffbffffffff",
            INIT_2D => X"ffffffe3ffffffffffffffddffffffffffffffdeffffffff0000001500000000",
            INIT_2E => X"ffffff93ffffffffffffff9dfffffffffffffff8ffffffff0000000800000000",
            INIT_2F => X"0000000900000000ffffffa8ffffffffffffffa3ffffffffffffffa4ffffffff",
            INIT_30 => X"fffffffaffffffff000000180000000000000021000000000000000000000000",
            INIT_31 => X"00000004000000000000001c00000000ffffffedffffffff0000000900000000",
            INIT_32 => X"00000005000000000000000d00000000fffffffeffffffffffffffffffffffff",
            INIT_33 => X"0000001b00000000ffffffe5ffffffffffffffeffffffffffffffff8ffffffff",
            INIT_34 => X"0000000f00000000ffffffdffffffffffffffff1fffffffffffffffcffffffff",
            INIT_35 => X"ffffffd6ffffffff0000000000000000fffffff6fffffffffffffff6ffffffff",
            INIT_36 => X"0000000000000000ffffffdfffffffff0000002f000000000000000d00000000",
            INIT_37 => X"fffffffdfffffffffffffffeffffffff0000000c00000000ffffffdaffffffff",
            INIT_38 => X"0000000e00000000ffffffe3fffffffffffffffcffffffff0000001c00000000",
            INIT_39 => X"000000170000000000000024000000000000000d000000000000002500000000",
            INIT_3A => X"fffffffbffffffff0000002400000000fffffffeffffffff0000002400000000",
            INIT_3B => X"ffffffd2ffffffffffffffdbffffffffffffff9cffffffffffffffe0ffffffff",
            INIT_3C => X"ffffffecffffffffffffffcaffffffffffffffbcffffffffffffffd4ffffffff",
            INIT_3D => X"000000490000000000000050000000000000004b00000000ffffffe2ffffffff",
            INIT_3E => X"0000003100000000000000150000000000000034000000000000002300000000",
            INIT_3F => X"ffffffdefffffffffffffff4fffffffffffffffdffffffff0000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001f0000000000000036000000000000000e000000000000001b00000000",
            INIT_41 => X"ffffffd4ffffffff00000017000000000000002c000000000000001600000000",
            INIT_42 => X"00000022000000000000001e00000000ffffffdeffffffffffffffcfffffffff",
            INIT_43 => X"fffffff3ffffffffffffffffffffffff0000002400000000fffffff2ffffffff",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE4;


    MEM_IWGHT_LAYER2_INSTANCE0 : if BRAM_NAME = "iwght_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00001efb00000000fffff7bdfffffffffffffcfcffffffff000004ff00000000",
            INIT_01 => X"ffffe329ffffffff000006b7000000000000245300000000fffff01effffffff",
            INIT_02 => X"0000129b00000000ffffe7e2ffffffff00001b6300000000fffff2c5ffffffff",
            INIT_03 => X"00000806000000000000010d0000000000001bb40000000000000e3d00000000",
            INIT_04 => X"0000002f000000000000001700000000fffffff3ffffffff0000001900000000",
            INIT_05 => X"0000000e00000000000000170000000000000039000000000000002400000000",
            INIT_06 => X"ffffffb8ffffffffffffffdeffffffffffffffebffffffff0000002800000000",
            INIT_07 => X"0000001500000000fffffff1ffffffffffffffa0ffffffffffffffbfffffffff",
            INIT_08 => X"ffffffc7ffffffffffffffc9fffffffffffffff2ffffffffffffffc0ffffffff",
            INIT_09 => X"fffffffaffffffffffffff98ffffffffffffff8affffffffffffffeeffffffff",
            INIT_0A => X"0000003b00000000fffffff8ffffffffffffffb8ffffffffffffffbeffffffff",
            INIT_0B => X"0000004e000000000000006a0000000000000038000000000000005600000000",
            INIT_0C => X"0000004300000000000000450000000000000025000000000000002a00000000",
            INIT_0D => X"0000002700000000ffffffddfffffffffffffffbffffffff0000001900000000",
            INIT_0E => X"0000003700000000000000410000000000000015000000000000001200000000",
            INIT_0F => X"ffffffaaffffffffffffffb3ffffffff00000002000000000000001d00000000",
            INIT_10 => X"00000016000000000000001d00000000fffffff4ffffffff0000000000000000",
            INIT_11 => X"ffffffddffffffff0000000800000000ffffffd9ffffffff0000001600000000",
            INIT_12 => X"0000000300000000ffffffccffffffffffffffd5ffffffff0000000300000000",
            INIT_13 => X"ffffffeeffffffff0000000200000000ffffffd7ffffffffffffffc4ffffffff",
            INIT_14 => X"ffffff9fffffffffffffffbcffffffff00000008000000000000001100000000",
            INIT_15 => X"ffffffbdffffffffffffffa8ffffffffffffffbcffffffffffffffe6ffffffff",
            INIT_16 => X"00000015000000000000000a000000000000001100000000fffffff6ffffffff",
            INIT_17 => X"00000021000000000000003d00000000ffffffcbffffffff0000001400000000",
            INIT_18 => X"000000260000000000000018000000000000001c00000000fffffff9ffffffff",
            INIT_19 => X"0000000e00000000000000090000000000000025000000000000001d00000000",
            INIT_1A => X"ffffffe6fffffffffffffff6ffffffff0000002e000000000000002c00000000",
            INIT_1B => X"ffffffc5ffffffffffffffd7ffffffffffffffc0ffffffffffffffeaffffffff",
            INIT_1C => X"0000001700000000ffffffb8ffffffffffffffb1ffffffffffffffe1ffffffff",
            INIT_1D => X"0000003200000000fffffffaffffffff00000008000000000000002400000000",
            INIT_1E => X"0000001e000000000000001d00000000ffffffecffffffff0000003500000000",
            INIT_1F => X"ffffffd6ffffffffffffffe7ffffffffffffffd0ffffffff0000000200000000",
            INIT_20 => X"ffffff9dffffffffffffffe1ffffffffffffffc4ffffffffffffff95ffffffff",
            INIT_21 => X"fffffff2ffffffff00000026000000000000002c00000000ffffffafffffffff",
            INIT_22 => X"00000004000000000000003a000000000000003e000000000000000c00000000",
            INIT_23 => X"0000001700000000ffffffc8ffffffff0000002f000000000000004200000000",
            INIT_24 => X"fffffff4fffffffffffffff9ffffffffffffffe5ffffffff0000000100000000",
            INIT_25 => X"000000010000000000000012000000000000000e000000000000001300000000",
            INIT_26 => X"ffffffe7ffffffff00000020000000000000000700000000fffffffbffffffff",
            INIT_27 => X"0000001b000000000000002b000000000000002900000000fffffff5ffffffff",
            INIT_28 => X"ffffffdeffffffff0000001000000000fffffffbffffffff0000000b00000000",
            INIT_29 => X"0000002900000000fffffffeffffffff0000000800000000fffffff0ffffffff",
            INIT_2A => X"fffffff3ffffffff000000120000000000000015000000000000001d00000000",
            INIT_2B => X"0000000100000000fffffff6ffffffff0000004c000000000000002600000000",
            INIT_2C => X"000000120000000000000049000000000000000200000000ffffffecffffffff",
            INIT_2D => X"ffffffd5ffffffff000000220000000000000038000000000000000600000000",
            INIT_2E => X"ffffffe4ffffffffffffffd5ffffffffffffffc2ffffffffffffffd3ffffffff",
            INIT_2F => X"0000001b000000000000001f00000000ffffffd7ffffffffffffffbdffffffff",
            INIT_30 => X"00000000000000000000003f0000000000000029000000000000000900000000",
            INIT_31 => X"00000000000000000000001b00000000fffffff4ffffffffffffffcaffffffff",
            INIT_32 => X"0000002f000000000000002a00000000ffffffefffffffff0000000400000000",
            INIT_33 => X"fffffff0ffffffff0000000e00000000fffffff7ffffffff0000001000000000",
            INIT_34 => X"0000001200000000fffffff5ffffffff00000002000000000000000800000000",
            INIT_35 => X"fffffff9ffffffffffffffedffffffffffffffd7ffffffff0000002600000000",
            INIT_36 => X"fffffff2ffffffff00000000000000000000000e00000000fffffff2ffffffff",
            INIT_37 => X"000000420000000000000010000000000000001600000000ffffffe4ffffffff",
            INIT_38 => X"ffffffebffffffff000000020000000000000030000000000000002200000000",
            INIT_39 => X"0000002500000000000000230000000000000009000000000000004300000000",
            INIT_3A => X"00000018000000000000002000000000ffffffe4ffffffffffffffefffffffff",
            INIT_3B => X"ffffffecffffffff0000001400000000ffffffe2ffffffff0000000e00000000",
            INIT_3C => X"00000027000000000000001e000000000000001f000000000000000000000000",
            INIT_3D => X"fffffffaffffffff0000000000000000fffffffafffffffffffffffcffffffff",
            INIT_3E => X"000000150000000000000027000000000000000800000000ffffffe8ffffffff",
            INIT_3F => X"000000310000000000000038000000000000001d00000000fffffffaffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe2ffffffff0000000d000000000000000200000000fffffff0ffffffff",
            INIT_41 => X"ffffffcbfffffffffffffffeffffffffffffffdfffffffffffffffb8ffffffff",
            INIT_42 => X"ffffffe6ffffffffffffffdfffffffff0000000600000000ffffffc9ffffffff",
            INIT_43 => X"0000006000000000000000020000000000000032000000000000004400000000",
            INIT_44 => X"ffffffffffffffff0000003f0000000000000017000000000000003e00000000",
            INIT_45 => X"0000002a0000000000000010000000000000000a000000000000002600000000",
            INIT_46 => X"00000008000000000000002100000000fffffff9ffffffff0000002800000000",
            INIT_47 => X"fffffffdfffffffffffffff8ffffffff00000015000000000000001b00000000",
            INIT_48 => X"0000001600000000ffffffe2ffffffffffffffdbffffffffffffffe5ffffffff",
            INIT_49 => X"00000006000000000000001000000000ffffffe5ffffffff0000000800000000",
            INIT_4A => X"0000000f00000000ffffffe4ffffffff00000014000000000000003d00000000",
            INIT_4B => X"fffffff9fffffffffffffff9ffffffff00000008000000000000001200000000",
            INIT_4C => X"0000000d00000000fffffff1ffffffff0000000b000000000000003000000000",
            INIT_4D => X"fffffff4ffffffff0000000200000000fffffff5ffffffffffffffcaffffffff",
            INIT_4E => X"fffffff7fffffffffffffff7fffffffffffffffcffffffff0000000100000000",
            INIT_4F => X"ffffffe6ffffffff00000040000000000000003c00000000ffffffccffffffff",
            INIT_50 => X"00000007000000000000000d000000000000002f000000000000002700000000",
            INIT_51 => X"0000000000000000000000090000000000000005000000000000002600000000",
            INIT_52 => X"ffffffc8ffffffff0000001d000000000000003000000000fffffffbffffffff",
            INIT_53 => X"fffffff1fffffffffffffffbffffffff0000001100000000fffffff0ffffffff",
            INIT_54 => X"ffffffa6ffffffffffffffcaffffffff0000001500000000fffffff5ffffffff",
            INIT_55 => X"0000000200000000ffffffdfffffffff00000021000000000000002000000000",
            INIT_56 => X"0000000000000000ffffffd8ffffffffffffffcdffffffff0000000000000000",
            INIT_57 => X"ffffffe4ffffffff00000017000000000000000800000000ffffffbeffffffff",
            INIT_58 => X"ffffffdcffffffff0000000d0000000000000009000000000000001100000000",
            INIT_59 => X"fffffff5ffffffff000000160000000000000007000000000000000f00000000",
            INIT_5A => X"ffffffebffffffff00000006000000000000002000000000fffffff0ffffffff",
            INIT_5B => X"ffffffeeffffffffffffffe5ffffffffffffffe9ffffffff0000000c00000000",
            INIT_5C => X"0000003200000000ffffffdeffffffff0000001d000000000000001300000000",
            INIT_5D => X"00000042000000000000000c00000000ffffffe8ffffffff0000001c00000000",
            INIT_5E => X"0000001500000000ffffffbdffffffffffffffefffffffff0000000c00000000",
            INIT_5F => X"0000004b0000000000000036000000000000002500000000ffffffecffffffff",
            INIT_60 => X"00000019000000000000002100000000fffffffeffffffff0000006000000000",
            INIT_61 => X"0000002d00000000ffffffe2ffffffff00000019000000000000002e00000000",
            INIT_62 => X"0000001a00000000fffffff6fffffffffffffffdffffffff0000000600000000",
            INIT_63 => X"fffffff4ffffffff000000020000000000000024000000000000003200000000",
            INIT_64 => X"00000006000000000000003c0000000000000026000000000000002100000000",
            INIT_65 => X"0000000a000000000000000a0000000000000020000000000000002100000000",
            INIT_66 => X"fffffffaffffffffffffffdbffffffff0000000a000000000000000c00000000",
            INIT_67 => X"ffffffffffffffff0000000b0000000000000044000000000000000800000000",
            INIT_68 => X"0000002300000000fffffff5ffffffff0000005d000000000000002d00000000",
            INIT_69 => X"000000050000000000000028000000000000001a000000000000004d00000000",
            INIT_6A => X"ffffffe2ffffffffffffffc2ffffffffffffffe9ffffffff0000001a00000000",
            INIT_6B => X"0000001b000000000000003a00000000ffffffceffffffffffffffd6ffffffff",
            INIT_6C => X"fffffff0ffffffff000000100000000000000028000000000000000500000000",
            INIT_6D => X"0000001700000000ffffffd6ffffffffffffffdaffffffff0000002400000000",
            INIT_6E => X"ffffffe6ffffffff0000001b000000000000001500000000fffffffbffffffff",
            INIT_6F => X"fffffff7fffffffffffffffefffffffffffffff3ffffffffffffffe3ffffffff",
            INIT_70 => X"ffffffcfffffffff00000001000000000000000d00000000ffffffecffffffff",
            INIT_71 => X"0000000400000000fffffffaffffffff00000020000000000000002900000000",
            INIT_72 => X"ffffffd3ffffffffffffffc5ffffffff0000001b000000000000004e00000000",
            INIT_73 => X"0000000b00000000ffffffccffffffffffffffd4ffffffffffffffedffffffff",
            INIT_74 => X"fffffff9ffffffff00000035000000000000002b00000000ffffffe2ffffffff",
            INIT_75 => X"fffffff4fffffffffffffffdfffffffffffffff3ffffffff0000000800000000",
            INIT_76 => X"0000000d0000000000000029000000000000000700000000fffffffdffffffff",
            INIT_77 => X"0000001a000000000000003c0000000000000050000000000000003600000000",
            INIT_78 => X"000000090000000000000013000000000000003b000000000000000b00000000",
            INIT_79 => X"fffffff6ffffffff000000030000000000000014000000000000000500000000",
            INIT_7A => X"0000001c00000000fffffffbffffffff00000019000000000000004d00000000",
            INIT_7B => X"0000007100000000000000590000000000000047000000000000002100000000",
            INIT_7C => X"0000001d00000000fffffffbfffffffffffffff7ffffffff0000002a00000000",
            INIT_7D => X"000000080000000000000019000000000000000d00000000ffffffe2ffffffff",
            INIT_7E => X"ffffffedffffffffffffffe9ffffffffffffffe9ffffffffffffffe9ffffffff",
            INIT_7F => X"fffffff9ffffffffffffffe3fffffffffffffff6ffffffffffffffefffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE0;


    MEM_IWGHT_LAYER2_INSTANCE1 : if BRAM_NAME = "iwght_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffffffffffdaffffffff0000000800000000fffffff7ffffffff",
            INIT_01 => X"0000000700000000000000060000000000000029000000000000000100000000",
            INIT_02 => X"ffffffbfffffffff0000002500000000fffffffcffffffff0000000000000000",
            INIT_03 => X"ffffffcdfffffffffffffff6fffffffffffffffdffffffffffffffc8ffffffff",
            INIT_04 => X"ffffffecffffffffffffffcafffffffffffffff0ffffffffffffffbbffffffff",
            INIT_05 => X"ffffffe2ffffffff00000013000000000000000d000000000000000a00000000",
            INIT_06 => X"ffffffecffffffff00000000000000000000000000000000ffffffdcffffffff",
            INIT_07 => X"0000000400000000ffffffc6fffffffffffffff5ffffffff0000001700000000",
            INIT_08 => X"0000003200000000ffffffdafffffffffffffff9ffffffff0000001e00000000",
            INIT_09 => X"00000036000000000000001d0000000000000036000000000000003700000000",
            INIT_0A => X"fffffffbfffffffffffffff2ffffffff00000013000000000000000900000000",
            INIT_0B => X"0000003900000000ffffffffffffffff00000009000000000000003900000000",
            INIT_0C => X"000000290000000000000029000000000000001c00000000ffffffe5ffffffff",
            INIT_0D => X"0000000f00000000ffffffd7ffffffff0000000d000000000000002800000000",
            INIT_0E => X"0000003b000000000000002100000000ffffffebffffffff0000003800000000",
            INIT_0F => X"00000043000000000000001c00000000fffffff1ffffffff0000002b00000000",
            INIT_10 => X"0000001300000000000000000000000000000009000000000000002200000000",
            INIT_11 => X"ffffffd3ffffffff0000000400000000ffffffd8ffffffff0000001f00000000",
            INIT_12 => X"0000001300000000ffffffeaffffffffffffffdefffffffffffffffdffffffff",
            INIT_13 => X"ffffffcbffffffffffffffcbffffffffffffffd7ffffffff0000000400000000",
            INIT_14 => X"ffffffd1fffffffffffffffdffffffffffffffdaffffffffffffffc0ffffffff",
            INIT_15 => X"00000007000000000000002a00000000ffffffe9ffffffffffffffeaffffffff",
            INIT_16 => X"00000014000000000000002300000000fffffffafffffffffffffff8ffffffff",
            INIT_17 => X"000000210000000000000036000000000000003b000000000000002600000000",
            INIT_18 => X"0000000500000000000000360000000000000045000000000000005300000000",
            INIT_19 => X"0000001d000000000000001d000000000000003600000000ffffffdbffffffff",
            INIT_1A => X"0000000f00000000000000170000000000000032000000000000004800000000",
            INIT_1B => X"fffffff1ffffffff0000002600000000fffffff1ffffffff0000000600000000",
            INIT_1C => X"ffffffeeffffffff00000004000000000000003000000000fffffff4ffffffff",
            INIT_1D => X"0000000200000000fffffff2ffffffffffffffcfffffffffffffffffffffffff",
            INIT_1E => X"ffffffecffffffff00000001000000000000001600000000ffffffeeffffffff",
            INIT_1F => X"0000000c00000000fffffffafffffffffffffff4ffffffff0000001900000000",
            INIT_20 => X"0000001e000000000000001d00000000fffffffefffffffffffffff5ffffffff",
            INIT_21 => X"0000001700000000fffffff9ffffffff00000031000000000000002900000000",
            INIT_22 => X"fffffff0ffffffff00000014000000000000001b000000000000001a00000000",
            INIT_23 => X"fffffff8ffffffff000000330000000000000027000000000000003600000000",
            INIT_24 => X"00000025000000000000003700000000fffffffdffffffff0000003700000000",
            INIT_25 => X"0000004e00000000000000480000000000000027000000000000006000000000",
            INIT_26 => X"fffffff1ffffffff0000001400000000fffffff5ffffffffffffffbcffffffff",
            INIT_27 => X"fffffff3ffffffffffffffb8fffffffffffffffaffffffff0000001a00000000",
            INIT_28 => X"0000002100000000ffffffdefffffffffffffffdffffffff0000001800000000",
            INIT_29 => X"ffffffdffffffffffffffffdffffffff0000001500000000ffffffebffffffff",
            INIT_2A => X"0000000300000000fffffff6ffffffff0000002300000000ffffffdfffffffff",
            INIT_2B => X"00000046000000000000000300000000ffffffd8ffffffff0000000b00000000",
            INIT_2C => X"000000230000000000000036000000000000000c000000000000000b00000000",
            INIT_2D => X"0000000d000000000000003700000000fffffffdffffffffffffffddffffffff",
            INIT_2E => X"0000000500000000fffffff0ffffffff0000001400000000fffffffcffffffff",
            INIT_2F => X"0000002d0000000000000018000000000000002000000000ffffffd6ffffffff",
            INIT_30 => X"0000001f0000000000000028000000000000001b000000000000005500000000",
            INIT_31 => X"0000002e000000000000001a00000000ffffffd1ffffffff0000002100000000",
            INIT_32 => X"ffffffe3ffffffff0000001700000000fffffff8ffffffff0000001100000000",
            INIT_33 => X"ffffffd4fffffffffffffffafffffffffffffff3ffffffffffffffecffffffff",
            INIT_34 => X"0000000c00000000fffffffeffffffffffffffe9fffffffffffffff8ffffffff",
            INIT_35 => X"fffffff2ffffffffffffffe8ffffffffffffffe4ffffffff0000001200000000",
            INIT_36 => X"0000002400000000000000070000000000000006000000000000002600000000",
            INIT_37 => X"0000001b00000000fffffff9ffffffffffffffdbffffffff0000003300000000",
            INIT_38 => X"0000000d00000000000000330000000000000024000000000000001000000000",
            INIT_39 => X"0000003a000000000000002c000000000000004a000000000000006800000000",
            INIT_3A => X"0000001a000000000000000800000000ffffffe0ffffffffffffffffffffffff",
            INIT_3B => X"ffffffdffffffffffffffff8ffffffffffffffbeffffffffffffffeaffffffff",
            INIT_3C => X"0000001d000000000000001600000000ffffffcaffffffffffffffaeffffffff",
            INIT_3D => X"00000010000000000000003c0000000000000002000000000000003800000000",
            INIT_3E => X"00000004000000000000000000000000fffffffcffffffff0000000d00000000",
            INIT_3F => X"fffffff2ffffffffffffffe2ffffffff0000000e00000000fffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002d00000000ffffffffffffffffffffffffffffffff0000001600000000",
            INIT_41 => X"ffffffeeffffffff0000000e0000000000000014000000000000001800000000",
            INIT_42 => X"00000027000000000000002c000000000000000f000000000000003600000000",
            INIT_43 => X"00000010000000000000002d00000000fffffffefffffffffffffffbffffffff",
            INIT_44 => X"0000002b00000000ffffffebffffffff0000001d000000000000000b00000000",
            INIT_45 => X"fffffff2ffffffff00000025000000000000001600000000fffffffcffffffff",
            INIT_46 => X"00000015000000000000001d0000000000000024000000000000002900000000",
            INIT_47 => X"fffffffafffffffffffffff2ffffffff00000000000000000000003e00000000",
            INIT_48 => X"ffffffcafffffffffffffff0ffffffff0000000800000000fffffffeffffffff",
            INIT_49 => X"fffffffaffffffffffffffe0ffffffffffffffdaffffffffffffffa0ffffffff",
            INIT_4A => X"0000000000000000000000140000000000000038000000000000002700000000",
            INIT_4B => X"ffffffdbffffffff00000018000000000000005400000000fffffff3ffffffff",
            INIT_4C => X"ffffffdfffffffffffffffd7fffffffffffffff1ffffffffffffffcdffffffff",
            INIT_4D => X"0000000300000000fffffff7ffffffff0000000600000000ffffffefffffffff",
            INIT_4E => X"000000030000000000000037000000000000000b00000000fffffffaffffffff",
            INIT_4F => X"ffffffdbffffffffffffffe0fffffffffffffff8ffffffffffffffd9ffffffff",
            INIT_50 => X"ffffffebffffffffffffffeeffffffffffffffe1ffffffff0000000400000000",
            INIT_51 => X"000000280000000000000018000000000000001f000000000000000100000000",
            INIT_52 => X"00000035000000000000002e00000000ffffffebffffffff0000000100000000",
            INIT_53 => X"ffffffbeffffffff0000001600000000fffffffdffffffff0000001100000000",
            INIT_54 => X"ffffffcfffffffffffffffe5fffffffffffffff8ffffffffffffffd8ffffffff",
            INIT_55 => X"ffffffe6ffffffff0000000c00000000fffffff7ffffffffffffffedffffffff",
            INIT_56 => X"0000002600000000fffffff4fffffffffffffff3ffffffff0000001500000000",
            INIT_57 => X"000000200000000000000004000000000000001000000000ffffffdeffffffff",
            INIT_58 => X"0000000b0000000000000041000000000000002f000000000000000c00000000",
            INIT_59 => X"ffffffdeffffffff0000001e000000000000001f000000000000000c00000000",
            INIT_5A => X"ffffffcafffffffffffffffbffffffffffffffd3fffffffffffffff8ffffffff",
            INIT_5B => X"0000000900000000ffffffe0ffffffff0000000600000000ffffffd5ffffffff",
            INIT_5C => X"fffffff1ffffffffffffffe2ffffffffffffffe1fffffffffffffff1ffffffff",
            INIT_5D => X"0000001300000000ffffffe8ffffffffffffffe8ffffffffffffffe0ffffffff",
            INIT_5E => X"00000005000000000000000f00000000fffffffaffffffffffffffd0ffffffff",
            INIT_5F => X"00000028000000000000000800000000ffffffe7ffffffff0000001300000000",
            INIT_60 => X"ffffffa6ffffffffffffffc0ffffffff0000002200000000fffffff8ffffffff",
            INIT_61 => X"00000032000000000000000000000000ffffffaefffffffffffffffbffffffff",
            INIT_62 => X"00000026000000000000001e00000000fffffff7ffffffff0000001b00000000",
            INIT_63 => X"0000002b000000000000000d00000000fffffff4ffffffff0000003000000000",
            INIT_64 => X"ffffffe3ffffffff0000000000000000fffffffcffffffff0000000100000000",
            INIT_65 => X"ffffffe9ffffffff0000002f00000000fffffff3ffffffff0000002300000000",
            INIT_66 => X"000000390000000000000009000000000000004a000000000000000d00000000",
            INIT_67 => X"fffffff7fffffffffffffffbffffffffffffffd3ffffffff0000003400000000",
            INIT_68 => X"0000002d00000000000000490000000000000032000000000000002e00000000",
            INIT_69 => X"ffffffd8ffffffffffffffbbffffffff0000000600000000fffffffaffffffff",
            INIT_6A => X"0000000900000000ffffffdcffffffffffffffc2ffffffffffffffffffffffff",
            INIT_6B => X"00000006000000000000001a000000000000001b00000000ffffffe5ffffffff",
            INIT_6C => X"0000001e000000000000001f000000000000000b000000000000000f00000000",
            INIT_6D => X"0000000c000000000000000f000000000000000b000000000000001b00000000",
            INIT_6E => X"0000003600000000ffffffcefffffffffffffff5ffffffff0000004300000000",
            INIT_6F => X"0000000500000000000000190000000000000000000000000000000000000000",
            INIT_70 => X"fffffff3ffffffff0000001e000000000000001700000000ffffffe2ffffffff",
            INIT_71 => X"ffffffb9ffffffff0000003500000000fffffff0ffffffffffffffecffffffff",
            INIT_72 => X"fffffffcffffffffffffffccffffffff0000003000000000ffffffdfffffffff",
            INIT_73 => X"0000000900000000fffffff1ffffffffffffffdcffffffff0000002100000000",
            INIT_74 => X"ffffffebffffffff0000002b00000000fffffff0ffffffffffffffe4ffffffff",
            INIT_75 => X"ffffffd7ffffffffffffffebffffffffffffffedffffffffffffffebffffffff",
            INIT_76 => X"00000009000000000000001a00000000ffffffb8ffffffff0000001b00000000",
            INIT_77 => X"ffffffccffffffffffffffdeffffffffffffffecffffffff0000001800000000",
            INIT_78 => X"fffffff7ffffffff0000000200000000ffffffdeffffffffffffffe3ffffffff",
            INIT_79 => X"fffffffafffffffffffffff9ffffffff0000000900000000ffffffe1ffffffff",
            INIT_7A => X"00000001000000000000000400000000ffffffd2ffffffff0000000600000000",
            INIT_7B => X"00000012000000000000000b000000000000004300000000ffffffeeffffffff",
            INIT_7C => X"0000001a000000000000000c000000000000000b00000000ffffffffffffffff",
            INIT_7D => X"ffffffe3ffffffff0000000b0000000000000031000000000000000500000000",
            INIT_7E => X"ffffffd7ffffffffffffffd5ffffffff0000001700000000ffffffd8ffffffff",
            INIT_7F => X"0000007c00000000fffffffeffffffffffffffc7ffffffff0000004700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE1;


    MEM_IWGHT_LAYER2_INSTANCE2 : if BRAM_NAME = "iwght_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001800000000fffffff2ffffffff0000002000000000ffffffedffffffff",
            INIT_01 => X"0000001000000000fffffff1ffffffffffffffe7ffffffff0000000000000000",
            INIT_02 => X"ffffffefffffffffffffffc8ffffffff00000002000000000000002200000000",
            INIT_03 => X"ffffffbaffffffff0000000e00000000ffffffccffffffffffffffeaffffffff",
            INIT_04 => X"ffffffedffffffffffffffbcffffffffffffffe7ffffffffffffffd0ffffffff",
            INIT_05 => X"ffffffe4ffffffffffffffe3ffffffffffffffe8ffffffff0000000200000000",
            INIT_06 => X"0000001d00000000ffffffe9ffffffffffffffe6ffffffff0000001600000000",
            INIT_07 => X"00000036000000000000002f000000000000000700000000fffffff9ffffffff",
            INIT_08 => X"0000001f000000000000002d00000000ffffffe1ffffffff0000000f00000000",
            INIT_09 => X"0000002800000000ffffffccffffffff0000000f00000000fffffffdffffffff",
            INIT_0A => X"0000003f00000000000000080000000000000003000000000000000700000000",
            INIT_0B => X"ffffffe2ffffffff0000000c0000000000000034000000000000001900000000",
            INIT_0C => X"0000000b000000000000001f000000000000000f000000000000004800000000",
            INIT_0D => X"000000370000000000000023000000000000001500000000fffffff9ffffffff",
            INIT_0E => X"0000002100000000000000210000000000000036000000000000001600000000",
            INIT_0F => X"ffffffd7ffffffff0000002a0000000000000014000000000000001000000000",
            INIT_10 => X"ffffffe6fffffffffffffffdffffffff0000001c00000000ffffffcdffffffff",
            INIT_11 => X"ffffffb7ffffffffffffffd1fffffffffffffff8ffffffffffffffdeffffffff",
            INIT_12 => X"00000000000000000000000b00000000fffffff1ffffffffffffffeeffffffff",
            INIT_13 => X"0000000d00000000fffffff2ffffffff0000004e00000000ffffffe8ffffffff",
            INIT_14 => X"0000001e00000000ffffffeaffffffff00000037000000000000004f00000000",
            INIT_15 => X"ffffffeeffffffff0000001b0000000000000020000000000000001400000000",
            INIT_16 => X"0000000a0000000000000015000000000000003b000000000000002f00000000",
            INIT_17 => X"0000002700000000fffffffaffffffff0000000900000000fffffff4ffffffff",
            INIT_18 => X"0000002000000000fffffffaffffffff0000001e00000000fffffffbffffffff",
            INIT_19 => X"00000026000000000000002d00000000ffffffe1ffffffff0000000600000000",
            INIT_1A => X"ffffffedfffffffffffffff3ffffffff0000000400000000ffffffdfffffffff",
            INIT_1B => X"ffffffdfffffffffffffffecffffffffffffffeaffffffffffffffd9ffffffff",
            INIT_1C => X"ffffffecffffffffffffffcaffffffff0000000f00000000ffffffe7ffffffff",
            INIT_1D => X"ffffffdeffffffffffffffe7fffffffffffffff2ffffffffffffffe5ffffffff",
            INIT_1E => X"ffffffe7ffffffff0000001200000000fffffffafffffffffffffff8ffffffff",
            INIT_1F => X"0000002500000000ffffffffffffffff00000006000000000000002100000000",
            INIT_20 => X"ffffffe0ffffffff0000001c000000000000000000000000ffffffcbffffffff",
            INIT_21 => X"ffffffe7ffffffff0000000e0000000000000014000000000000001700000000",
            INIT_22 => X"0000001b00000000fffffffeffffffff0000002300000000ffffffe8ffffffff",
            INIT_23 => X"000000380000000000000025000000000000003b000000000000001900000000",
            INIT_24 => X"0000002b000000000000001d000000000000000f000000000000002500000000",
            INIT_25 => X"0000000800000000ffffffc9ffffffff0000000e000000000000003d00000000",
            INIT_26 => X"0000004000000000000000180000000000000000000000000000000400000000",
            INIT_27 => X"fffffff8ffffffff0000002d000000000000001f000000000000001100000000",
            INIT_28 => X"ffffffeeffffffff0000001f0000000000000021000000000000002500000000",
            INIT_29 => X"0000003200000000fffffff8ffffffffffffffe6fffffffffffffffbffffffff",
            INIT_2A => X"fffffff4fffffffffffffff6fffffffffffffffbffffffffffffffd6ffffffff",
            INIT_2B => X"ffffffedffffffff0000000e00000000fffffffcffffffffffffffe2ffffffff",
            INIT_2C => X"0000002700000000fffffff4fffffffffffffff3ffffffffffffffefffffffff",
            INIT_2D => X"000000020000000000000038000000000000002200000000ffffffffffffffff",
            INIT_2E => X"0000001800000000fffffff6fffffffffffffff2ffffffffffffffebffffffff",
            INIT_2F => X"ffffffd4ffffffffffffffeeffffffffffffffecffffffff0000002b00000000",
            INIT_30 => X"ffffffdcffffffff0000000300000000ffffffe9ffffffffffffffe5ffffffff",
            INIT_31 => X"00000028000000000000001d000000000000001e00000000fffffff5ffffffff",
            INIT_32 => X"0000000a000000000000000e000000000000001a000000000000001100000000",
            INIT_33 => X"0000004a00000000000000140000000000000000000000000000000200000000",
            INIT_34 => X"0000006b00000000000000230000000000000050000000000000003200000000",
            INIT_35 => X"0000003800000000000000430000000000000009000000000000006e00000000",
            INIT_36 => X"0000004300000000fffffff9ffffffff0000001f000000000000004100000000",
            INIT_37 => X"00000042000000000000000700000000ffffffe0ffffffffffffffe8ffffffff",
            INIT_38 => X"ffffffecffffffffffffffe9ffffffff0000000100000000ffffffecffffffff",
            INIT_39 => X"0000000f00000000ffffffd5ffffffff0000000d000000000000001d00000000",
            INIT_3A => X"0000002d000000000000001e00000000fffffff9ffffffff0000001a00000000",
            INIT_3B => X"00000014000000000000002d0000000000000000000000000000002200000000",
            INIT_3C => X"0000000a00000000ffffffeaffffffff00000010000000000000000700000000",
            INIT_3D => X"0000000c00000000ffffffe6ffffffff0000000900000000ffffffecffffffff",
            INIT_3E => X"0000000a000000000000000600000000fffffff9ffffffff0000000600000000",
            INIT_3F => X"fffffff0ffffffff0000003f0000000000000045000000000000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc0ffffffffffffffcfffffffffffffffffffffffffffffffedffffffff",
            INIT_41 => X"ffffffb3ffffffff0000000300000000ffffffedffffffffffffffbcffffffff",
            INIT_42 => X"0000004000000000ffffffd2ffffffffffffffceffffffff0000000600000000",
            INIT_43 => X"0000000900000000fffffff4fffffffffffffff1ffffffff0000000200000000",
            INIT_44 => X"0000003b00000000fffffffbffffffff00000007000000000000004400000000",
            INIT_45 => X"00000027000000000000002200000000fffffff6ffffffff0000000900000000",
            INIT_46 => X"0000001f000000000000002700000000fffffff4ffffffff0000002000000000",
            INIT_47 => X"00000010000000000000002a000000000000002d000000000000000200000000",
            INIT_48 => X"ffffffd1ffffffff0000000e000000000000001000000000ffffffebffffffff",
            INIT_49 => X"ffffffb5ffffffffffffffc2ffffffffffffffcbffffffffffffffd8ffffffff",
            INIT_4A => X"ffffffd9ffffffffffffffd9ffffffff0000003100000000ffffffd2ffffffff",
            INIT_4B => X"0000000700000000ffffffd7ffffffff00000026000000000000000b00000000",
            INIT_4C => X"0000003400000000000000030000000000000005000000000000000500000000",
            INIT_4D => X"0000000400000000fffffffbffffffff0000000100000000fffffff4ffffffff",
            INIT_4E => X"ffffffc2ffffffffffffffffffffffff0000003b000000000000000500000000",
            INIT_4F => X"0000000c00000000ffffffe3ffffffffffffffdffffffffffffffffcffffffff",
            INIT_50 => X"ffffffdcfffffffffffffff2fffffffffffffffbfffffffffffffff2ffffffff",
            INIT_51 => X"ffffffccffffffff0000000a000000000000002900000000ffffffdbffffffff",
            INIT_52 => X"fffffff5ffffffff0000000e00000000ffffffffffffffffffffffe7ffffffff",
            INIT_53 => X"0000000f00000000000000540000000000000028000000000000002700000000",
            INIT_54 => X"0000000d00000000000000110000000000000030000000000000000e00000000",
            INIT_55 => X"00000017000000000000000b00000000fffffff2ffffffff0000000200000000",
            INIT_56 => X"ffffffe4ffffffff0000001300000000ffffffc9ffffffff0000001200000000",
            INIT_57 => X"000000030000000000000024000000000000001e00000000ffffffe8ffffffff",
            INIT_58 => X"ffffffd0ffffffffffffffebffffffff00000007000000000000000600000000",
            INIT_59 => X"fffffff5ffffffffffffffcfffffffffffffffeeffffffffffffffbdffffffff",
            INIT_5A => X"0000001f00000000ffffffdaffffffffffffffb7ffffffff0000001200000000",
            INIT_5B => X"ffffffd7ffffffff0000000b00000000ffffffdeffffffff0000000a00000000",
            INIT_5C => X"000000240000000000000013000000000000001600000000ffffffefffffffff",
            INIT_5D => X"00000005000000000000001b0000000000000019000000000000000d00000000",
            INIT_5E => X"0000000a000000000000001d000000000000002d00000000ffffffefffffffff",
            INIT_5F => X"00000010000000000000001500000000ffffffedffffffffffffffecffffffff",
            INIT_60 => X"000000040000000000000028000000000000000200000000fffffff5ffffffff",
            INIT_61 => X"0000000b00000000ffffffedffffffff0000002b000000000000001200000000",
            INIT_62 => X"ffffffe8ffffffffffffffe8ffffffff0000000900000000fffffff9ffffffff",
            INIT_63 => X"0000004d0000000000000014000000000000001b000000000000001700000000",
            INIT_64 => X"0000002900000000000000400000000000000007000000000000001100000000",
            INIT_65 => X"ffffffdcfffffffffffffff6ffffffff00000003000000000000005800000000",
            INIT_66 => X"ffffffecffffffffffffffe6ffffffff0000002400000000fffffffeffffffff",
            INIT_67 => X"000000180000000000000016000000000000001900000000fffffffdffffffff",
            INIT_68 => X"0000002c000000000000001b00000000ffffffffffffffff0000003d00000000",
            INIT_69 => X"ffffffdbffffffff0000000100000000ffffffd7ffffffffffffffe6ffffffff",
            INIT_6A => X"fffffffaffffffffffffffcfffffffff0000001e00000000ffffffdcffffffff",
            INIT_6B => X"fffffff2ffffffffffffffe4ffffffffffffffe0ffffffff0000002100000000",
            INIT_6C => X"0000004100000000ffffffe8ffffffff0000004b00000000fffffffdffffffff",
            INIT_6D => X"00000041000000000000005d000000000000001e000000000000004a00000000",
            INIT_6E => X"0000001f00000000000000310000000000000019000000000000004000000000",
            INIT_6F => X"ffffffe6ffffffff0000001f00000000fffffffbffffffff0000003e00000000",
            INIT_70 => X"00000035000000000000003e00000000fffffffbffffffffffffffedffffffff",
            INIT_71 => X"0000002100000000fffffffeffffffff0000002000000000fffffffeffffffff",
            INIT_72 => X"ffffffcfffffffff0000003f000000000000003b000000000000001e00000000",
            INIT_73 => X"ffffffd4ffffffffffffffd9ffffffff0000002e000000000000000100000000",
            INIT_74 => X"000000220000000000000009000000000000000c00000000fffffff4ffffffff",
            INIT_75 => X"0000001600000000fffffff4fffffffffffffff3ffffffffffffffe3ffffffff",
            INIT_76 => X"fffffff6ffffffff0000002c00000000fffffffdffffffff0000001000000000",
            INIT_77 => X"fffffff6ffffffff0000001700000000fffffffbffffffff0000002c00000000",
            INIT_78 => X"fffffff9ffffffffffffffc7ffffffffffffffe6ffffffff0000001b00000000",
            INIT_79 => X"0000001700000000ffffffeeffffffff00000012000000000000000500000000",
            INIT_7A => X"ffffffd4ffffffffffffffe8ffffffff0000002200000000ffffffe1ffffffff",
            INIT_7B => X"0000005200000000ffffffc9ffffffff0000001d000000000000004000000000",
            INIT_7C => X"fffffff2ffffffff00000036000000000000000e000000000000002c00000000",
            INIT_7D => X"00000021000000000000000f00000000ffffffe6ffffffff0000001f00000000",
            INIT_7E => X"ffffffbdffffffffffffffdcffffffff0000001a00000000fffffffdffffffff",
            INIT_7F => X"ffffffbcffffffffffffffaeffffffffffffffc7ffffffffffffffafffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE2;


    MEM_IWGHT_LAYER2_INSTANCE3 : if BRAM_NAME = "iwght_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c000000000000000b00000000fffffff5ffffffffffffff89ffffffff",
            INIT_01 => X"0000001b0000000000000018000000000000000000000000ffffffeaffffffff",
            INIT_02 => X"00000003000000000000000500000000ffffffe2ffffffffffffffeaffffffff",
            INIT_03 => X"fffffff2ffffffff000000070000000000000026000000000000001600000000",
            INIT_04 => X"fffffffcffffffffffffffd7ffffffff00000015000000000000001c00000000",
            INIT_05 => X"ffffffc5ffffffff0000000d00000000fffffff6ffffffffffffffdbffffffff",
            INIT_06 => X"0000002e000000000000002700000000fffffff8ffffffff0000000200000000",
            INIT_07 => X"ffffffe3ffffffff0000000100000000fffffff9fffffffffffffff7ffffffff",
            INIT_08 => X"0000000400000000ffffffd5ffffffff0000001c000000000000001200000000",
            INIT_09 => X"00000023000000000000001e00000000fffffffafffffffffffffff4ffffffff",
            INIT_0A => X"ffffffe0fffffffffffffff8ffffffffffffffe7ffffffffffffffebffffffff",
            INIT_0B => X"0000002400000000000000260000000000000024000000000000002100000000",
            INIT_0C => X"fffffffdffffffff00000026000000000000002000000000fffffff8ffffffff",
            INIT_0D => X"0000001500000000ffffffe9fffffffffffffff4ffffffff0000000300000000",
            INIT_0E => X"0000000e00000000000000200000000000000015000000000000000300000000",
            INIT_0F => X"0000001c0000000000000005000000000000000700000000ffffffe2ffffffff",
            INIT_10 => X"ffffffa0ffffffffffffffcdffffffffffffff98ffffffffffffffc0ffffffff",
            INIT_11 => X"ffffffe7ffffffffffffffdfffffffffffffff96ffffffffffffffa8ffffffff",
            INIT_12 => X"00000013000000000000004300000000fffffff8fffffffffffffff6ffffffff",
            INIT_13 => X"fffffffdffffffff00000012000000000000003c000000000000002e00000000",
            INIT_14 => X"0000002600000000fffffffbfffffffffffffffeffffffff0000001400000000",
            INIT_15 => X"00000040000000000000002c000000000000000d000000000000005400000000",
            INIT_16 => X"0000000f0000000000000022000000000000001700000000ffffffd6ffffffff",
            INIT_17 => X"0000000200000000ffffffd9ffffffff0000000300000000fffffff9ffffffff",
            INIT_18 => X"00000016000000000000001500000000ffffffecfffffffffffffffeffffffff",
            INIT_19 => X"ffffffdaffffffffffffffc9ffffffffffffffccffffffffffffffceffffffff",
            INIT_1A => X"ffffffffffffffff0000002e00000000ffffffdaffffffff0000000000000000",
            INIT_1B => X"0000000800000000ffffffe2ffffffff0000002a00000000fffffff8ffffffff",
            INIT_1C => X"00000006000000000000001300000000fffffff0ffffffff0000000100000000",
            INIT_1D => X"fffffffbffffffff0000002400000000ffffffdcffffffffffffffe6ffffffff",
            INIT_1E => X"0000001b000000000000001a000000000000001a000000000000001500000000",
            INIT_1F => X"ffffffb7fffffffffffffffbffffffff0000000d00000000fffffff7ffffffff",
            INIT_20 => X"00000010000000000000001700000000ffffffecffffffffffffffc6ffffffff",
            INIT_21 => X"fffffffaffffffff00000010000000000000003a000000000000001200000000",
            INIT_22 => X"0000001100000000ffffffd1ffffffffffffffffffffffff0000001d00000000",
            INIT_23 => X"0000002000000000000000510000000000000005000000000000001200000000",
            INIT_24 => X"ffffffffffffffff000000070000000000000024000000000000002300000000",
            INIT_25 => X"0000000000000000ffffffe5ffffffff0000000e000000000000002700000000",
            INIT_26 => X"fffffffcffffffff0000000c000000000000000a000000000000000d00000000",
            INIT_27 => X"fffffffeffffffff0000002c000000000000003600000000ffffffddffffffff",
            INIT_28 => X"ffffffd7fffffffffffffff4ffffffff0000001f000000000000002b00000000",
            INIT_29 => X"00000002000000000000000b000000000000000300000000ffffffeaffffffff",
            INIT_2A => X"0000003f000000000000001700000000fffffff1ffffffff0000002b00000000",
            INIT_2B => X"0000006d0000000000000059000000000000001800000000fffffffbffffffff",
            INIT_2C => X"000000280000000000000028000000000000007c000000000000007200000000",
            INIT_2D => X"000000260000000000000044000000000000003600000000fffffffcffffffff",
            INIT_2E => X"0000000f00000000fffffffbffffffff0000003b000000000000000200000000",
            INIT_2F => X"ffffffbcffffffffffffffc6fffffffffffffff1ffffffffffffffe4ffffffff",
            INIT_30 => X"0000001c00000000ffffffcefffffffffffffffbffffffff0000000100000000",
            INIT_31 => X"000000260000000000000000000000000000001700000000ffffffecffffffff",
            INIT_32 => X"00000003000000000000000c0000000000000005000000000000001c00000000",
            INIT_33 => X"ffffffd7ffffffff0000001400000000ffffffebffffffff0000000a00000000",
            INIT_34 => X"ffffffb7ffffffff00000003000000000000001300000000fffffff4ffffffff",
            INIT_35 => X"ffffffe9ffffffffffffffdaffffffffffffffc3ffffffffffffffc6ffffffff",
            INIT_36 => X"00000009000000000000002b000000000000004700000000ffffffdaffffffff",
            INIT_37 => X"00000031000000000000003e0000000000000030000000000000004100000000",
            INIT_38 => X"0000001f0000000000000014000000000000003a000000000000001f00000000",
            INIT_39 => X"00000032000000000000000200000000fffffff5fffffffffffffffcffffffff",
            INIT_3A => X"ffffffffffffffffffffffe7ffffffff0000001800000000ffffffedffffffff",
            INIT_3B => X"fffffff9ffffffff0000000600000000ffffffd4ffffffffffffffddffffffff",
            INIT_3C => X"00000013000000000000001800000000fffffff0ffffffff0000000600000000",
            INIT_3D => X"ffffffc5ffffffff0000000b000000000000000100000000fffffff8ffffffff",
            INIT_3E => X"ffffffc0ffffffffffffffcdffffffffffffffe1ffffffff0000000a00000000",
            INIT_3F => X"0000000a00000000ffffffefffffffffffffffecffffffffffffffdfffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdbffffffff0000001200000000ffffffe5fffffffffffffffaffffffff",
            INIT_41 => X"fffffff9ffffffff0000001800000000ffffffc0ffffffffffffffe7ffffffff",
            INIT_42 => X"fffffffeffffffff0000002900000000fffffff0ffffffffffffffe3ffffffff",
            INIT_43 => X"00000013000000000000000600000000ffffffccffffffff0000001200000000",
            INIT_44 => X"0000001f00000000fffffff7ffffffff0000001b000000000000000d00000000",
            INIT_45 => X"fffffff2ffffffffffffffe9ffffffff00000030000000000000002600000000",
            INIT_46 => X"00000035000000000000000d00000000fffffff9ffffffff0000001000000000",
            INIT_47 => X"00000037000000000000004a000000000000001a000000000000001300000000",
            INIT_48 => X"0000001c000000000000002d00000000fffffffaffffffff0000003f00000000",
            INIT_49 => X"0000000a000000000000002f0000000000000008000000000000000e00000000",
            INIT_4A => X"0000002700000000000000160000000000000007000000000000000700000000",
            INIT_4B => X"00000035000000000000002a000000000000003a00000000fffffff1ffffffff",
            INIT_4C => X"ffffffdbffffffff0000000c000000000000000f000000000000001d00000000",
            INIT_4D => X"fffffff0ffffffff000000020000000000000000000000000000002000000000",
            INIT_4E => X"ffffffe9ffffffff0000001f00000000ffffffe4ffffffff0000001100000000",
            INIT_4F => X"0000002500000000000000100000000000000037000000000000003300000000",
            INIT_50 => X"0000005500000000000000360000000000000025000000000000005d00000000",
            INIT_51 => X"fffffffcffffffff000000050000000000000023000000000000003b00000000",
            INIT_52 => X"0000000000000000000000110000000000000000000000000000000300000000",
            INIT_53 => X"0000000d000000000000000e000000000000000c000000000000000700000000",
            INIT_54 => X"0000001e00000000ffffffedffffffffffffffe7ffffffff0000002900000000",
            INIT_55 => X"0000000d000000000000000200000000ffffffe5ffffffff0000001100000000",
            INIT_56 => X"0000002600000000ffffffe0ffffffff0000000c000000000000000200000000",
            INIT_57 => X"ffffffd0ffffffff00000006000000000000001600000000ffffffe6ffffffff",
            INIT_58 => X"fffffff7fffffffffffffff0fffffffffffffffffffffffffffffffdffffffff",
            INIT_59 => X"0000003a000000000000001a0000000000000019000000000000001200000000",
            INIT_5A => X"0000003d000000000000000300000000ffffffd7fffffffffffffffdffffffff",
            INIT_5B => X"ffffffd5ffffffffffffffd0ffffffffffffffcfffffffffffffffdcffffffff",
            INIT_5C => X"0000000a00000000ffffffcbffffffffffffffe2fffffffffffffff2ffffffff",
            INIT_5D => X"0000001f00000000ffffffdaffffffffffffffe1ffffffff0000004000000000",
            INIT_5E => X"0000006000000000ffffffe9ffffffff00000011000000000000001000000000",
            INIT_5F => X"0000001a000000000000000100000000ffffffdeffffffff0000002800000000",
            INIT_60 => X"fffffff4ffffffffffffffd9ffffffffffffffedffffffffffffffbbffffffff",
            INIT_61 => X"fffffff9ffffffffffffffdbfffffffffffffffaffffffff0000001b00000000",
            INIT_62 => X"00000016000000000000004a000000000000000e000000000000001000000000",
            INIT_63 => X"00000004000000000000001e00000000fffffffdffffffff0000001b00000000",
            INIT_64 => X"ffffffe1ffffffffffffffccffffffffffffffebffffffffffffffd4ffffffff",
            INIT_65 => X"0000002900000000ffffffe7ffffffffffffffd0ffffffffffffffaeffffffff",
            INIT_66 => X"000000150000000000000019000000000000001f000000000000002100000000",
            INIT_67 => X"ffffffadffffffff0000000c00000000fffffff0ffffffff0000001e00000000",
            INIT_68 => X"ffffffb3ffffffffffffffbdffffffffffffffe8ffffffffffffffd8ffffffff",
            INIT_69 => X"0000000300000000fffffff4ffffffffffffffebffffffffffffffdfffffffff",
            INIT_6A => X"0000001b00000000000000300000000000000024000000000000001300000000",
            INIT_6B => X"0000001900000000000000120000000000000035000000000000001000000000",
            INIT_6C => X"fffffffbffffffff0000002c00000000fffffff8ffffffff0000000200000000",
            INIT_6D => X"00000015000000000000000f0000000000000031000000000000001500000000",
            INIT_6E => X"ffffffe3fffffffffffffff2ffffffff0000001300000000fffffffeffffffff",
            INIT_6F => X"0000001500000000ffffffeaffffffffffffffd0ffffffffffffffe4ffffffff",
            INIT_70 => X"0000004b000000000000001f000000000000002300000000fffffffdffffffff",
            INIT_71 => X"fffffff8ffffffff0000000900000000ffffffdeffffffff0000002b00000000",
            INIT_72 => X"ffffffccffffffff0000000b000000000000000900000000ffffffeeffffffff",
            INIT_73 => X"fffffff7ffffffff0000001f00000000ffffffcafffffffffffffff4ffffffff",
            INIT_74 => X"00000005000000000000001d00000000fffffffcffffffff0000002200000000",
            INIT_75 => X"ffffffe7ffffffff0000001b00000000fffffff6ffffffff0000003a00000000",
            INIT_76 => X"0000001c00000000fffffffeffffffff00000011000000000000001400000000",
            INIT_77 => X"00000011000000000000001600000000ffffffdeffffffffffffffe3ffffffff",
            INIT_78 => X"0000000e00000000ffffffebffffffff0000002400000000ffffffe9ffffffff",
            INIT_79 => X"ffffffd2ffffffff000000040000000000000008000000000000002500000000",
            INIT_7A => X"0000000e00000000ffffffe1ffffffffffffffe1ffffffffffffffd3ffffffff",
            INIT_7B => X"0000002b000000000000000a0000000000000022000000000000000000000000",
            INIT_7C => X"0000003a0000000000000014000000000000004f000000000000000e00000000",
            INIT_7D => X"00000030000000000000004d0000000000000023000000000000002a00000000",
            INIT_7E => X"fffffffaffffffffffffffc7ffffffffffffffe3ffffffff0000001400000000",
            INIT_7F => X"ffffffa8ffffffffffffffbdffffffffffffffe3ffffffffffffffc6ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE3;


    MEM_IWGHT_LAYER2_INSTANCE4 : if BRAM_NAME = "iwght_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003500000000ffffffd4ffffffffffffffdcffffffffffffffd7ffffffff",
            INIT_01 => X"0000000c00000000fffffff9fffffffffffffff9ffffffff0000000600000000",
            INIT_02 => X"0000001400000000ffffffe3ffffffff0000000c000000000000000200000000",
            INIT_03 => X"fffffff4ffffffff00000007000000000000002300000000ffffffffffffffff",
            INIT_04 => X"ffffffe9fffffffffffffffcfffffffffffffff8fffffffffffffff6ffffffff",
            INIT_05 => X"ffffffe1ffffffff0000000e000000000000001500000000ffffffcaffffffff",
            INIT_06 => X"0000003f000000000000000f000000000000001f000000000000002900000000",
            INIT_07 => X"0000000000000000ffffffd2ffffffffffffffd5ffffffff0000002b00000000",
            INIT_08 => X"0000000800000000ffffffddffffffffffffffd1ffffffff0000000a00000000",
            INIT_09 => X"00000008000000000000002500000000ffffffd5fffffffffffffffbffffffff",
            INIT_0A => X"00000004000000000000000d000000000000000f00000000fffffff4ffffffff",
            INIT_0B => X"fffffffafffffffffffffff7ffffffff00000012000000000000000b00000000",
            INIT_0C => X"0000002500000000000000090000000000000004000000000000000700000000",
            INIT_0D => X"ffffffebffffffff000000310000000000000026000000000000000000000000",
            INIT_0E => X"00000009000000000000001400000000ffffffebffffffff0000000400000000",
            INIT_0F => X"000000420000000000000033000000000000004f000000000000002700000000",
            INIT_10 => X"ffffffbeffffffff0000000c0000000000000045000000000000006d00000000",
            INIT_11 => X"ffffffffffffffff0000000f00000000ffffffe8ffffffff0000000a00000000",
            INIT_12 => X"ffffffe3ffffffffffffffeaffffffffffffffecffffffff0000000a00000000",
            INIT_13 => X"ffffffd0ffffffffffffffedffffffffffffffdcffffffff0000000700000000",
            INIT_14 => X"0000002400000000ffffffc6ffffffffffffffdeffffffff0000000900000000",
            INIT_15 => X"ffffffebffffffffffffffebfffffffffffffff0ffffffffffffffdaffffffff",
            INIT_16 => X"ffffffc3fffffffffffffffbffffffffffffffe0ffffffffffffffd1ffffffff",
            INIT_17 => X"ffffffcffffffffffffffff4fffffffffffffff2ffffffffffffffd2ffffffff",
            INIT_18 => X"ffffffc6ffffffffffffffb5ffffffffffffffe9ffffffffffffffb1ffffffff",
            INIT_19 => X"ffffffbcffffffffffffffd4ffffffff0000002500000000ffffffa6ffffffff",
            INIT_1A => X"fffffff7ffffffffffffffcbffffffffffffffbaffffffff0000004000000000",
            INIT_1B => X"00000015000000000000001d000000000000000c00000000fffffff4ffffffff",
            INIT_1C => X"ffffffe7ffffffff0000000d000000000000002900000000ffffffe1ffffffff",
            INIT_1D => X"0000002100000000000000280000000000000003000000000000002b00000000",
            INIT_1E => X"ffffffddffffffff0000003600000000ffffffaaffffffff0000001000000000",
            INIT_1F => X"00000000000000000000000c000000000000001400000000fffffff4ffffffff",
            INIT_20 => X"fffffffcffffffff000000120000000000000023000000000000000f00000000",
            INIT_21 => X"000000060000000000000009000000000000000f000000000000001700000000",
            INIT_22 => X"ffffffc8ffffffffffffffe9ffffffff00000012000000000000000100000000",
            INIT_23 => X"ffffffe0fffffffffffffffbffffffffffffffc8ffffffff0000000800000000",
            INIT_24 => X"000000040000000000000007000000000000001d00000000fffffffbffffffff",
            INIT_25 => X"0000000b0000000000000002000000000000001f00000000ffffffe4ffffffff",
            INIT_26 => X"fffffff8ffffffff00000038000000000000002c000000000000002100000000",
            INIT_27 => X"00000022000000000000001c000000000000001c00000000fffffff3ffffffff",
            INIT_28 => X"0000000800000000fffffffbffffffff0000000100000000fffffffaffffffff",
            INIT_29 => X"0000001000000000ffffffe4ffffffff0000000e000000000000000f00000000",
            INIT_2A => X"000000030000000000000006000000000000001e00000000ffffffe7ffffffff",
            INIT_2B => X"00000049000000000000003c000000000000001b000000000000000800000000",
            INIT_2C => X"0000000e00000000ffffffcdffffffff00000021000000000000004800000000",
            INIT_2D => X"0000001100000000ffffffe5fffffffffffffff0ffffffff0000003800000000",
            INIT_2E => X"ffffffffffffffff0000002c000000000000000900000000ffffffd7ffffffff",
            INIT_2F => X"ffffffd5ffffffff000000120000000000000001000000000000000600000000",
            INIT_30 => X"fffffff8ffffffffffffffebfffffffffffffffbfffffffffffffff3ffffffff",
            INIT_31 => X"0000001400000000fffffffaffffffffffffffbeffffffff0000000700000000",
            INIT_32 => X"0000001b00000000000000350000000000000062000000000000002c00000000",
            INIT_33 => X"000000020000000000000024000000000000003d000000000000004700000000",
            INIT_34 => X"fffffffbffffffffffffffebffffffffffffffccffffffffffffffecffffffff",
            INIT_35 => X"00000029000000000000000000000000fffffff0ffffffffffffffcdffffffff",
            INIT_36 => X"ffffffe5ffffffffffffffb2ffffffffffffffefffffffff0000000c00000000",
            INIT_37 => X"fffffff9ffffffffffffffb7ffffffffffffffd3ffffffffffffffc1ffffffff",
            INIT_38 => X"ffffffdfffffffff000000220000000000000010000000000000001800000000",
            INIT_39 => X"ffffffeaffffffff00000012000000000000000b00000000fffffff4ffffffff",
            INIT_3A => X"ffffffd8fffffffffffffffcffffffff00000003000000000000000d00000000",
            INIT_3B => X"fffffff5ffffffffffffffbcffffffffffffffb4ffffffffffffffddffffffff",
            INIT_3C => X"0000001c000000000000000e00000000ffffffa9ffffffffffffffcaffffffff",
            INIT_3D => X"0000000000000000ffffffc3ffffffffffffffe0ffffffffffffffecffffffff",
            INIT_3E => X"0000001b000000000000000700000000ffffffefffffffff0000000a00000000",
            INIT_3F => X"fffffff0ffffffff0000000500000000fffffff2ffffffff0000000e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000290000000000000006000000000000002b00000000fffffffeffffffff",
            INIT_41 => X"ffffff9ffffffffffffffff8fffffffffffffff7ffffffff0000001300000000",
            INIT_42 => X"ffffffc6ffffffffffffffd3fffffffffffffff5ffffffffffffffdeffffffff",
            INIT_43 => X"fffffffeffffffffffffffeefffffffffffffff6fffffffffffffff6ffffffff",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE4;


    MEM_IWGHT_LAYER3_INSTANCE0 : if BRAM_NAME = "iwght_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000015d0000000000000c87000000000000000600000000ffffdac9ffffffff",
            INIT_01 => X"ffffdf76ffffffff0000271f00000000ffffdba0ffffffff0000263e00000000",
            INIT_02 => X"fffffff7ffffffff0000000e00000000000002c80000000000000d1f00000000",
            INIT_03 => X"ffffffafffffffff0000002b00000000fffffff8ffffffff0000000b00000000",
            INIT_04 => X"0000000100000000ffffffe7ffffffff0000002700000000ffffffdfffffffff",
            INIT_05 => X"fffffff8ffffffff0000001800000000fffffff4fffffffffffffff7ffffffff",
            INIT_06 => X"0000001d000000000000002900000000ffffffd9ffffffff0000001b00000000",
            INIT_07 => X"ffffffb5fffffffffffffff1ffffffff0000002700000000ffffffd8ffffffff",
            INIT_08 => X"ffffffe0ffffffffffffffc9ffffffffffffffeeffffffffffffffeeffffffff",
            INIT_09 => X"0000001000000000ffffffd8ffffffff0000001d00000000ffffffc2ffffffff",
            INIT_0A => X"000000190000000000000009000000000000002f000000000000005700000000",
            INIT_0B => X"ffffffbaffffffff00000013000000000000000900000000ffffffe6ffffffff",
            INIT_0C => X"ffffffe9ffffffffffffffe8ffffffff00000024000000000000006300000000",
            INIT_0D => X"000000160000000000000002000000000000001500000000ffffffccffffffff",
            INIT_0E => X"0000001300000000ffffffb9ffffffffffffffb8ffffffff0000001f00000000",
            INIT_0F => X"ffffffc6ffffffff000000210000000000000032000000000000003200000000",
            INIT_10 => X"0000002800000000fffffff3ffffffff0000000500000000ffffffe4ffffffff",
            INIT_11 => X"ffffffe3ffffffff00000020000000000000001300000000fffffff7ffffffff",
            INIT_12 => X"0000001100000000ffffffedffffffffffffffe3ffffffff0000000900000000",
            INIT_13 => X"0000000500000000fffffff7ffffffffffffffcdffffffffffffffffffffffff",
            INIT_14 => X"ffffffe4ffffffff0000001200000000ffffffe4ffffffff0000000400000000",
            INIT_15 => X"00000000000000000000000e0000000000000040000000000000003600000000",
            INIT_16 => X"ffffffc6ffffffffffffffd9ffffffff0000000800000000ffffffeeffffffff",
            INIT_17 => X"ffffffcbffffffff0000002500000000ffffffe4ffffffff0000000400000000",
            INIT_18 => X"0000004f000000000000001300000000ffffffe5ffffffff0000001d00000000",
            INIT_19 => X"ffffffc0ffffffff0000000f000000000000004500000000ffffffdaffffffff",
            INIT_1A => X"0000000f000000000000002700000000ffffffcbffffffff0000002f00000000",
            INIT_1B => X"ffffffbdfffffffffffffff9ffffffff0000002f00000000fffffff4ffffffff",
            INIT_1C => X"000000140000000000000001000000000000002e00000000ffffffe9ffffffff",
            INIT_1D => X"fffffff0ffffffff00000038000000000000001c00000000fffffffbffffffff",
            INIT_1E => X"00000020000000000000001e0000000000000008000000000000000000000000",
            INIT_1F => X"00000016000000000000000100000000ffffffd0ffffffffffffffe8ffffffff",
            INIT_20 => X"ffffffdffffffffffffffffeffffffff0000000600000000ffffffcdffffffff",
            INIT_21 => X"ffffffabfffffffffffffff4ffffffffffffffe0ffffffffffffffefffffffff",
            INIT_22 => X"0000003b000000000000002c00000000fffffff3ffffffffffffffbbffffffff",
            INIT_23 => X"ffffffe3fffffffffffffff5fffffffffffffff2ffffffff0000000b00000000",
            INIT_24 => X"ffffffebffffffffffffffc7ffffffff0000000200000000ffffffabffffffff",
            INIT_25 => X"ffffffe5ffffffff000000370000000000000011000000000000002200000000",
            INIT_26 => X"0000000700000000ffffffedffffffff0000000b00000000ffffffd4ffffffff",
            INIT_27 => X"ffffffe7ffffffff00000032000000000000003e000000000000003a00000000",
            INIT_28 => X"0000001600000000ffffffd0ffffffff0000002000000000ffffffb4ffffffff",
            INIT_29 => X"00000000000000000000001400000000ffffffb2ffffffff0000002500000000",
            INIT_2A => X"0000001500000000fffffff8fffffffffffffffaffffffffffffffcfffffffff",
            INIT_2B => X"ffffffe0ffffffff00000024000000000000001a000000000000003000000000",
            INIT_2C => X"0000003a000000000000002900000000ffffffbcffffffffffffffd2ffffffff",
            INIT_2D => X"00000006000000000000001800000000ffffffd8ffffffff0000000d00000000",
            INIT_2E => X"ffffffeaffffffffffffffe1ffffffff0000000000000000ffffffe0ffffffff",
            INIT_2F => X"0000000700000000ffffffd7ffffffff00000011000000000000000700000000",
            INIT_30 => X"00000035000000000000001200000000ffffffc5ffffffffffffffd9ffffffff",
            INIT_31 => X"00000021000000000000001e000000000000000e000000000000000700000000",
            INIT_32 => X"0000000a00000000ffffffc5ffffffff0000001d00000000ffffffb6ffffffff",
            INIT_33 => X"ffffffa9ffffffff0000004400000000ffffffd3ffffffff0000000100000000",
            INIT_34 => X"ffffffc6ffffffffffffffc0ffffffff0000003f00000000ffffffa3ffffffff",
            INIT_35 => X"00000006000000000000002b00000000ffffffe5ffffffff0000000500000000",
            INIT_36 => X"0000005000000000fffffffcffffffff0000005400000000ffffffdcffffffff",
            INIT_37 => X"fffffff6ffffffff0000000200000000ffffffbffffffffffffffffbffffffff",
            INIT_38 => X"0000000b00000000ffffffe5ffffffff0000002800000000fffffffcffffffff",
            INIT_39 => X"ffffffdeffffffff0000000e000000000000007500000000fffffffaffffffff",
            INIT_3A => X"0000000400000000ffffffffffffffffffffffeaffffffffffffffc8ffffffff",
            INIT_3B => X"ffffffafffffffff00000000000000000000000900000000ffffffebffffffff",
            INIT_3C => X"fffffff3ffffffff0000003000000000ffffffc9ffffffffffffffbfffffffff",
            INIT_3D => X"00000002000000000000003b000000000000003a00000000fffffff8ffffffff",
            INIT_3E => X"fffffff3ffffffffffffffd7fffffffffffffffaffffffffffffffe0ffffffff",
            INIT_3F => X"ffffffbdfffffffffffffffcffffffff00000007000000000000005b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffceffffffff0000001300000000ffffff94fffffffffffffffdffffffff",
            INIT_41 => X"ffffffe1ffffffff0000000600000000fffffff5ffffffff0000003700000000",
            INIT_42 => X"ffffffeeffffffffffffffddffffffffffffffe2ffffffffffffffa8ffffffff",
            INIT_43 => X"ffffffe6ffffffff0000004e000000000000003a000000000000001200000000",
            INIT_44 => X"ffffffc6ffffffff0000001600000000ffffffcaffffffff0000001100000000",
            INIT_45 => X"ffffffafffffffff0000000700000000fffffff7ffffffff0000000000000000",
            INIT_46 => X"0000001100000000ffffffe2ffffffff00000030000000000000003300000000",
            INIT_47 => X"ffffffc4ffffffff0000001200000000ffffffddfffffffffffffff2ffffffff",
            INIT_48 => X"ffffffbdffffffff0000005400000000ffffffb7fffffffffffffffbffffffff",
            INIT_49 => X"ffffffa5fffffffffffffff1ffffffff0000001400000000fffffffdffffffff",
            INIT_4A => X"00000009000000000000002a00000000ffffffceffffffffffffffc2ffffffff",
            INIT_4B => X"ffffffe2ffffffffffffffeafffffffffffffffbffffffffffffffd4ffffffff",
            INIT_4C => X"0000000900000000000000100000000000000023000000000000001a00000000",
            INIT_4D => X"0000001900000000ffffffe4ffffffffffffffccfffffffffffffff5ffffffff",
            INIT_4E => X"0000000300000000ffffffe6ffffffffffffffd2ffffffff0000001c00000000",
            INIT_4F => X"fffffff1ffffffff00000011000000000000002d00000000ffffffe5ffffffff",
            INIT_50 => X"0000001500000000fffffff6ffffffffffffffe2ffffffff0000003400000000",
            INIT_51 => X"000000300000000000000010000000000000000800000000fffffffaffffffff",
            INIT_52 => X"00000030000000000000002600000000fffffff3ffffffff0000000000000000",
            INIT_53 => X"0000000500000000ffffffd8ffffffff0000002800000000fffffff4ffffffff",
            INIT_54 => X"ffffffe4ffffffffffffffc5ffffffffffffffeeffffffff0000000b00000000",
            INIT_55 => X"0000000200000000ffffffccffffffff0000002f00000000fffffff2ffffffff",
            INIT_56 => X"ffffffddffffffff0000003b0000000000000007000000000000002700000000",
            INIT_57 => X"0000001100000000ffffffe3ffffffff0000000e000000000000001700000000",
            INIT_58 => X"ffffffe9ffffffff0000001000000000fffffff7ffffffff0000001700000000",
            INIT_59 => X"fffffffdffffffff00000026000000000000002300000000ffffffdfffffffff",
            INIT_5A => X"0000000100000000ffffffefffffffff0000001000000000fffffff1ffffffff",
            INIT_5B => X"ffffffdbffffffffffffffe6ffffffff0000000300000000fffffff4ffffffff",
            INIT_5C => X"ffffffe3ffffffffffffffe4fffffffffffffffbffffffff0000001100000000",
            INIT_5D => X"ffffffbeffffffff0000001c00000000ffffffa6ffffffffffffffeeffffffff",
            INIT_5E => X"00000003000000000000000f00000000ffffffb3ffffffff0000001300000000",
            INIT_5F => X"0000003800000000ffffffecfffffffffffffff8ffffffffffffffe5ffffffff",
            INIT_60 => X"0000000d00000000ffffffb2ffffffff00000000000000000000000a00000000",
            INIT_61 => X"ffffffd5ffffffff0000000600000000ffffffccffffffff0000000700000000",
            INIT_62 => X"00000020000000000000002800000000ffffffd7ffffffff0000001500000000",
            INIT_63 => X"0000000a000000000000000b000000000000000600000000ffffffdcffffffff",
            INIT_64 => X"ffffffdeffffffffffffffcaffffffff00000028000000000000005300000000",
            INIT_65 => X"00000042000000000000000e000000000000005400000000ffffffddffffffff",
            INIT_66 => X"0000002000000000fffffff9ffffffff00000015000000000000001100000000",
            INIT_67 => X"0000001900000000fffffff4fffffffffffffff1ffffffffffffffc5ffffffff",
            INIT_68 => X"0000000700000000fffffff4fffffffffffffffafffffffffffffff6ffffffff",
            INIT_69 => X"fffffff7ffffffffffffffd4ffffffffffffffe3ffffffff0000001a00000000",
            INIT_6A => X"0000004c000000000000002000000000ffffffd5ffffffff0000000d00000000",
            INIT_6B => X"ffffffe0ffffffff0000001c0000000000000004000000000000000a00000000",
            INIT_6C => X"0000001e00000000ffffff82ffffffff0000001400000000fffffff8ffffffff",
            INIT_6D => X"0000001a00000000000000210000000000000006000000000000002500000000",
            INIT_6E => X"ffffffb9ffffffff000000170000000000000028000000000000005b00000000",
            INIT_6F => X"fffffffaffffffff00000015000000000000001b00000000fffffff2ffffffff",
            INIT_70 => X"ffffffdcffffffff00000044000000000000002c00000000ffffffdeffffffff",
            INIT_71 => X"ffffffdaffffffff0000000d00000000ffffffdcffffffff0000002800000000",
            INIT_72 => X"ffffffc5fffffffffffffffefffffffffffffff3ffffffff0000000000000000",
            INIT_73 => X"000000010000000000000003000000000000001f000000000000001000000000",
            INIT_74 => X"ffffffe5ffffffff0000003800000000ffffffeefffffffffffffff2ffffffff",
            INIT_75 => X"0000000100000000ffffffd7ffffffff0000000900000000ffffffebffffffff",
            INIT_76 => X"fffffffdffffffff0000000400000000ffffffe6fffffffffffffff3ffffffff",
            INIT_77 => X"0000001e000000000000002c00000000ffffffe6fffffffffffffff2ffffffff",
            INIT_78 => X"0000000800000000fffffffeffffffff00000020000000000000002c00000000",
            INIT_79 => X"fffffffaffffffff0000000000000000ffffffdaffffffffffffffdbffffffff",
            INIT_7A => X"fffffff1ffffffff0000001f00000000ffffffd5ffffffff0000000b00000000",
            INIT_7B => X"ffffffecffffffffffffffa1ffffffffffffffe1ffffffffffffffeeffffffff",
            INIT_7C => X"ffffffe6ffffffff000000290000000000000001000000000000000800000000",
            INIT_7D => X"ffffffe4ffffffffffffffd8ffffffffffffffcfffffffff0000000e00000000",
            INIT_7E => X"ffffffc9ffffffff0000001000000000ffffffe0ffffffff0000000100000000",
            INIT_7F => X"0000003500000000fffffff1ffffffff0000001400000000ffffffcaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE0;


    MEM_IWGHT_LAYER3_INSTANCE1 : if BRAM_NAME = "iwght_layer3_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002c00000000ffffffb7fffffffffffffffbffffffff0000000d00000000",
            INIT_01 => X"fffffff8ffffffffffffffccffffffffffffffd4ffffffff0000001600000000",
            INIT_02 => X"ffffffe0ffffffff000000230000000000000040000000000000003d00000000",
            INIT_03 => X"0000000f00000000ffffffe6ffffffffffffffdffffffffffffffffaffffffff",
            INIT_04 => X"ffffffe5ffffffff0000001b0000000000000029000000000000001300000000",
            INIT_05 => X"0000000400000000fffffffdffffffffffffffc7ffffffffffffffc8ffffffff",
            INIT_06 => X"fffffff8ffffffff0000000b0000000000000011000000000000001000000000",
            INIT_07 => X"fffffff6ffffffff0000001800000000ffffffc5ffffffffffffffd4ffffffff",
            INIT_08 => X"0000000000000000000000030000000000000013000000000000006300000000",
            INIT_09 => X"fffffff2ffffffff000000200000000000000008000000000000000800000000",
            INIT_0A => X"ffffffc4fffffffffffffff4ffffffff0000001100000000ffffffffffffffff",
            INIT_0B => X"fffffffffffffffffffffff2fffffffffffffff4ffffffff0000000a00000000",
            INIT_0C => X"0000002000000000ffffffc4ffffffff00000019000000000000002600000000",
            INIT_0D => X"0000004f000000000000002100000000fffffff4ffffffffffffffe7ffffffff",
            INIT_0E => X"fffffff5ffffffff000000110000000000000032000000000000001b00000000",
            INIT_0F => X"00000008000000000000000100000000ffffffebffffffff0000001200000000",
            INIT_10 => X"fffffffbffffffff0000001c0000000000000037000000000000003f00000000",
            INIT_11 => X"0000003600000000ffffffdfffffffffffffffdaffffffffffffffdeffffffff",
            INIT_12 => X"0000001600000000ffffffe4ffffffffffffffefffffffff0000000b00000000",
            INIT_13 => X"0000003c00000000fffffff1fffffffffffffff0ffffffffffffffd7ffffffff",
            INIT_14 => X"0000000f00000000ffffffdcffffffffffffffefffffffffffffffbeffffffff",
            INIT_15 => X"ffffffefffffffff0000002400000000ffffffd9ffffffffffffffecffffffff",
            INIT_16 => X"00000034000000000000003e00000000fffffffcffffffffffffffc4ffffffff",
            INIT_17 => X"0000002a00000000ffffffbeffffffff0000002800000000ffffffc2ffffffff",
            INIT_18 => X"0000001a00000000ffffffd1ffffffff0000002400000000ffffffb7ffffffff",
            INIT_19 => X"0000000400000000ffffffe9ffffffffffffffe8ffffffff0000001500000000",
            INIT_1A => X"ffffffebfffffffffffffff3ffffffff0000002e00000000fffffff3ffffffff",
            INIT_1B => X"fffffff4ffffffffffffffdaffffffffffffffddffffffffffffffd9ffffffff",
            INIT_1C => X"00000013000000000000000100000000ffffffecffffffffffffffcbffffffff",
            INIT_1D => X"0000001800000000ffffffd8ffffffff0000001b00000000ffffffddffffffff",
            INIT_1E => X"0000004f000000000000000100000000fffffff6ffffffff0000004400000000",
            INIT_1F => X"ffffffdafffffffffffffff2ffffffff0000000f000000000000000e00000000",
            INIT_20 => X"fffffffeffffffff0000001400000000fffffff1fffffffffffffff9ffffffff",
            INIT_21 => X"00000026000000000000002d000000000000000f00000000fffffff1ffffffff",
            INIT_22 => X"ffffffe2ffffffffffffffddffffffff0000002900000000ffffffc1ffffffff",
            INIT_23 => X"0000002f00000000ffffffeeffffffffffffffefffffffffffffffe5ffffffff",
            INIT_24 => X"ffffffbcfffffffffffffffbffffffff00000011000000000000000400000000",
            INIT_25 => X"ffffffe5ffffffffffffffd4ffffffffffffffeffffffffffffffffcffffffff",
            INIT_26 => X"0000003c00000000ffffffefffffffffffffffbbffffffffffffffc3ffffffff",
            INIT_27 => X"000000200000000000000006000000000000001400000000ffffffd3ffffffff",
            INIT_28 => X"ffffffdbffffffffffffffafffffffff00000006000000000000001300000000",
            INIT_29 => X"0000000e00000000fffffff7ffffffff0000001a000000000000000f00000000",
            INIT_2A => X"ffffffedffffffff0000004e00000000ffffffebffffffffffffffebffffffff",
            INIT_2B => X"0000003200000000ffffffdbffffffff0000000b00000000ffffffeaffffffff",
            INIT_2C => X"0000002300000000ffffffddfffffffffffffff3ffffffffffffffc9ffffffff",
            INIT_2D => X"00000012000000000000002a000000000000003b000000000000002700000000",
            INIT_2E => X"ffffffcaffffffff0000001b000000000000000e000000000000000a00000000",
            INIT_2F => X"0000003800000000ffffffd7ffffffff0000001500000000ffffffb0ffffffff",
            INIT_30 => X"ffffffe5ffffffff0000001800000000fffffff3ffffffff0000001f00000000",
            INIT_31 => X"0000002000000000ffffffeaffffffffffffffd3ffffffff0000003a00000000",
            INIT_32 => X"000000110000000000000036000000000000001900000000fffffff2ffffffff",
            INIT_33 => X"00000000000000000000002500000000fffffff0ffffffffffffffd2ffffffff",
            INIT_34 => X"ffffffbdffffffffffffffccffffffff0000001800000000fffffff1ffffffff",
            INIT_35 => X"fffffff0ffffffff0000000000000000ffffffdafffffffffffffffdffffffff",
            INIT_36 => X"ffffffc9ffffffffffffffdcffffffff0000002200000000ffffffd2ffffffff",
            INIT_37 => X"ffffffffffffffff0000001b000000000000002300000000fffffffeffffffff",
            INIT_38 => X"ffffffb4ffffffff0000002c0000000000000004000000000000000f00000000",
            INIT_39 => X"ffffffeeffffffffffffffa7ffffffff0000001100000000ffffffffffffffff",
            INIT_3A => X"ffffffccfffffffffffffffcffffffffffffffa3fffffffffffffff1ffffffff",
            INIT_3B => X"0000000e00000000000000520000000000000002000000000000002b00000000",
            INIT_3C => X"000000090000000000000011000000000000001e000000000000001700000000",
            INIT_3D => X"0000002200000000fffffff1ffffffff00000033000000000000003200000000",
            INIT_3E => X"ffffffe1ffffffff0000000d00000000ffffffbafffffffffffffff3ffffffff",
            INIT_3F => X"000000130000000000000013000000000000000800000000ffffffeaffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff9effffffff0000002c000000000000000d000000000000000e00000000",
            INIT_41 => X"0000001500000000fffffffdffffffff00000020000000000000000000000000",
            INIT_42 => X"ffffffd1ffffffff0000002600000000ffffffecffffffff0000000100000000",
            INIT_43 => X"ffffffd6ffffffffffffffdeffffffff0000000100000000ffffffb8ffffffff",
            INIT_44 => X"ffffffe3ffffffff0000000800000000ffffffdeffffffff0000000100000000",
            INIT_45 => X"ffffffedffffffffffffffb8ffffffffffffffceffffffffffffffc8ffffffff",
            INIT_46 => X"ffffffb5ffffffff0000000100000000ffffffe7ffffffff0000003800000000",
            INIT_47 => X"0000003300000000ffffffbbffffffffffffffe0ffffffffffffffecffffffff",
            INIT_48 => X"00000021000000000000002b0000000000000006000000000000000a00000000",
            INIT_49 => X"ffffffd0ffffffff0000001a00000000ffffffd3ffffffff0000002000000000",
            INIT_4A => X"ffffffd1ffffffff000000070000000000000063000000000000000000000000",
            INIT_4B => X"0000001100000000ffffffb9ffffffffffffffddffffffffffffffd2ffffffff",
            INIT_4C => X"0000000700000000fffffffdffffffff00000013000000000000002c00000000",
            INIT_4D => X"0000000b00000000ffffffaaffffffffffffffcfffffffff0000000c00000000",
            INIT_4E => X"00000004000000000000000e000000000000002100000000fffffffcffffffff",
            INIT_4F => X"ffffffe0ffffffffffffffd5ffffffffffffffefffffffffffffffebffffffff",
            INIT_50 => X"0000001b00000000ffffffe8ffffffff00000013000000000000001600000000",
            INIT_51 => X"fffffff8ffffffff0000001500000000ffffffd6fffffffffffffff5ffffffff",
            INIT_52 => X"ffffffd2ffffffff0000002800000000ffffffe9ffffffff0000004500000000",
            INIT_53 => X"fffffffaffffffffffffffe9ffffffffffffffcfffffffff0000000d00000000",
            INIT_54 => X"ffffffe9ffffffff00000009000000000000004b00000000ffffffe5ffffffff",
            INIT_55 => X"00000049000000000000000700000000ffffffdfffffffff0000003300000000",
            INIT_56 => X"ffffffe7ffffffff0000001300000000fffffff3ffffffffffffffe2ffffffff",
            INIT_57 => X"ffffffebffffffffffffffdafffffffffffffff0ffffffff0000002900000000",
            INIT_58 => X"ffffffe4fffffffffffffffeffffffff00000057000000000000003400000000",
            INIT_59 => X"00000046000000000000001000000000ffffffafffffffff0000000800000000",
            INIT_5A => X"ffffffc5ffffffffffffffffffffffffffffffeeffffffffffffffe4ffffffff",
            INIT_5B => X"fffffff9ffffffffffffffffffffffff0000003a000000000000002d00000000",
            INIT_5C => X"ffffffc9ffffffffffffffeaffffffff00000015000000000000003200000000",
            INIT_5D => X"00000027000000000000001900000000ffffffe6ffffffff0000004b00000000",
            INIT_5E => X"ffffffd1ffffffff00000029000000000000002c00000000ffffff9fffffffff",
            INIT_5F => X"fffffff4ffffffffffffffb2ffffffff0000000300000000ffffffeaffffffff",
            INIT_60 => X"ffffffebffffffffffffffd3ffffffff0000001100000000ffffffb1ffffffff",
            INIT_61 => X"ffffffe3ffffffff000000130000000000000006000000000000000e00000000",
            INIT_62 => X"0000000500000000ffffffe3ffffffff0000000400000000ffffff6cffffffff",
            INIT_63 => X"fffffffaffffffff00000025000000000000001800000000fffffffbffffffff",
            INIT_64 => X"0000002800000000fffffff2ffffffffffffffcefffffffffffffff6ffffffff",
            INIT_65 => X"0000001400000000ffffffc7ffffffffffffffddffffffffffffffe3ffffffff",
            INIT_66 => X"0000000500000000fffffffcffffffff0000006400000000ffffff63ffffffff",
            INIT_67 => X"0000002800000000ffffffabffffffff0000000f000000000000005200000000",
            INIT_68 => X"ffffffc4ffffffff0000001d00000000ffffffe3ffffffffffffffeaffffffff",
            INIT_69 => X"ffffffe1ffffffffffffffd4ffffffff00000003000000000000001000000000",
            INIT_6A => X"00000002000000000000005d00000000ffffff9fffffffffffffffd8ffffffff",
            INIT_6B => X"0000001800000000ffffffc6ffffffff0000006500000000ffffffeaffffffff",
            INIT_6C => X"0000001e00000000ffffffb4ffffffff0000000000000000ffffff82ffffffff",
            INIT_6D => X"0000001c00000000ffffffb4ffffffffffffffe8ffffffffffffffbaffffffff",
            INIT_6E => X"0000002900000000ffffffeeffffffffffffffcfffffffffffffff5cffffffff",
            INIT_6F => X"0000001f0000000000000017000000000000002300000000ffffffe0ffffffff",
            INIT_70 => X"ffffffeefffffffffffffffaffffffff0000000000000000ffffffd1ffffffff",
            INIT_71 => X"0000004000000000ffffffbdffffffffffffff86ffffffffffffffebffffffff",
            INIT_72 => X"fffffffdfffffffffffffffbfffffffffffffff7ffffffff0000001300000000",
            INIT_73 => X"0000003b00000000fffffffaffffffffffffffefffffffff0000002000000000",
            INIT_74 => X"00000021000000000000002a00000000ffffffeefffffffffffffffcffffffff",
            INIT_75 => X"fffffff2fffffffffffffff7ffffffff0000000500000000fffffffbffffffff",
            INIT_76 => X"ffffffefffffffffffffffe3ffffffff0000000500000000ffffffc7ffffffff",
            INIT_77 => X"0000002700000000ffffffffffffffff00000026000000000000004800000000",
            INIT_78 => X"ffffffd3ffffffff0000000100000000ffffffc8ffffffffffffffe3ffffffff",
            INIT_79 => X"00000024000000000000000100000000ffffffe0ffffffff0000003500000000",
            INIT_7A => X"ffffffedffffffffffffffedffffffffffffffe2ffffffffffffffe0ffffffff",
            INIT_7B => X"fffffff7fffffffffffffff1fffffffffffffff7ffffffffffffffbdffffffff",
            INIT_7C => X"fffffffbffffffff00000013000000000000003200000000ffffffe8ffffffff",
            INIT_7D => X"ffffffe6ffffffffffffffd9ffffffffffffffecffffffff0000000700000000",
            INIT_7E => X"00000015000000000000000a00000000ffffffddffffffffffffffe3ffffffff",
            INIT_7F => X"ffffffd9ffffffff0000005b00000000ffffff9efffffffffffffffbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE1;


    MEM_IWGHT_LAYER3_INSTANCE2 : if BRAM_NAME = "iwght_layer3_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000021000000000000000900000000ffffffdaffffffffffffffdeffffffff",
            INIT_01 => X"fffffff2ffffffffffffffebfffffffffffffff1fffffffffffffff4ffffffff",
            INIT_02 => X"0000000800000000ffffffe3ffffffff0000001500000000ffffffe0ffffffff",
            INIT_03 => X"0000001b00000000fffffff3ffffffffffffffdaffffffffffffffe6ffffffff",
            INIT_04 => X"ffffffecffffffff000000060000000000000012000000000000000a00000000",
            INIT_05 => X"ffffffe5fffffffffffffff5ffffffffffffffebffffffffffffffffffffffff",
            INIT_06 => X"0000001900000000fffffffdffffffff0000001c000000000000001b00000000",
            INIT_07 => X"ffffffd2ffffffff0000001000000000ffffff8effffffff0000005a00000000",
            INIT_08 => X"ffffffddffffffff00000006000000000000001100000000fffffffdffffffff",
            INIT_09 => X"ffffffe5ffffffffffffffdaffffffff00000016000000000000002f00000000",
            INIT_0A => X"0000002700000000fffffff9ffffffff0000000f00000000ffffffe5ffffffff",
            INIT_0B => X"000000250000000000000003000000000000004a000000000000000700000000",
            INIT_0C => X"000000140000000000000017000000000000000d000000000000001600000000",
            INIT_0D => X"ffffffdcffffffffffffffcdffffffffffffffb4ffffffff0000002d00000000",
            INIT_0E => X"ffffff9dffffffffffffffe6ffffffff0000001b00000000ffffffdeffffffff",
            INIT_0F => X"ffffffabffffffff0000001600000000ffffffe4ffffffff0000002c00000000",
            INIT_10 => X"00000049000000000000001c000000000000000c00000000ffffffc6ffffffff",
            INIT_11 => X"ffffffdaffffffffffffffd2ffffffffffffffeaffffffff0000005200000000",
            INIT_12 => X"ffffffb8ffffffff0000000f00000000ffffffe9ffffffff0000003a00000000",
            INIT_13 => X"0000001f00000000fffffffafffffffffffffffdfffffffffffffffaffffffff",
            INIT_14 => X"ffffffbeffffffff0000001c00000000fffffffdffffffff0000001b00000000",
            INIT_15 => X"0000001000000000ffffffd7ffffffffffffffd4ffffffff0000001500000000",
            INIT_16 => X"00000037000000000000001900000000ffffffc9ffffffff0000000100000000",
            INIT_17 => X"0000004200000000ffffffb6ffffffff0000001e00000000fffffffaffffffff",
            INIT_18 => X"0000003f00000000ffffffa4ffffffff0000001300000000ffffffb0ffffffff",
            INIT_19 => X"0000000c00000000ffffffe5ffffffffffffffefffffffff0000003700000000",
            INIT_1A => X"fffffff2ffffffff0000000f00000000ffffffd6fffffffffffffff2ffffffff",
            INIT_1B => X"0000004d00000000ffffffc8ffffffff0000000800000000ffffffd3ffffffff",
            INIT_1C => X"ffffffc8ffffffffffffffbfffffffffffffffecffffffffffffffc2ffffffff",
            INIT_1D => X"0000000f00000000ffffffc1ffffffffffffffe0ffffffff0000002c00000000",
            INIT_1E => X"0000002a000000000000004400000000fffffff9ffffffffffffffc3ffffffff",
            INIT_1F => X"fffffff6fffffffffffffffbffffffff0000004e00000000fffffff0ffffffff",
            INIT_20 => X"ffffffcdffffffff0000001000000000fffffff8ffffffffffffff85ffffffff",
            INIT_21 => X"00000002000000000000000100000000ffffffb9ffffffff0000002f00000000",
            INIT_22 => X"00000023000000000000002e000000000000003f00000000ffffffc0ffffffff",
            INIT_23 => X"ffffffe1ffffffff0000000e00000000ffffffd3ffffffffffffffe6ffffffff",
            INIT_24 => X"0000004800000000ffffffd9ffffffff0000000d00000000ffffffe3ffffffff",
            INIT_25 => X"ffffffc4ffffffff00000036000000000000001c00000000ffffffc9ffffffff",
            INIT_26 => X"ffffffd0fffffffffffffffbffffffffffffffeeffffffffffffffdbffffffff",
            INIT_27 => X"0000000400000000fffffffafffffffffffffff4ffffffffffffffdbffffffff",
            INIT_28 => X"0000000000000000ffffffe3ffffffff0000000a000000000000001600000000",
            INIT_29 => X"00000001000000000000000d000000000000002500000000ffffffe4ffffffff",
            INIT_2A => X"0000003000000000000000270000000000000020000000000000000b00000000",
            INIT_2B => X"ffffffb5ffffffff0000001600000000ffffffc1ffffffff0000002200000000",
            INIT_2C => X"0000002000000000ffffff90ffffffff0000002000000000ffffffbfffffffff",
            INIT_2D => X"0000002c00000000fffffffdfffffffffffffff9ffffffff0000000f00000000",
            INIT_2E => X"ffffffbfffffffffffffffedffffffff0000000e00000000ffffffc1ffffffff",
            INIT_2F => X"fffffff0fffffffffffffffbffffffffffffffc1fffffffffffffff3ffffffff",
            INIT_30 => X"0000001900000000fffffff5ffffffff00000002000000000000001800000000",
            INIT_31 => X"fffffffdffffffff0000001b0000000000000024000000000000001f00000000",
            INIT_32 => X"ffffffdbffffffffffffffd8ffffffffffffffddffffffffffffffdeffffffff",
            INIT_33 => X"0000002c00000000fffffff6fffffffffffffff8ffffffff0000003b00000000",
            INIT_34 => X"0000004e0000000000000000000000000000001500000000ffffffd1ffffffff",
            INIT_35 => X"00000010000000000000001a0000000000000023000000000000000d00000000",
            INIT_36 => X"ffffffdafffffffffffffff1ffffffffffffffddffffffffffffffc7ffffffff",
            INIT_37 => X"ffffffedffffffff0000000b00000000ffffffe3ffffffff0000004700000000",
            INIT_38 => X"ffffffedfffffffffffffff7ffffffffffffffecfffffffffffffff1ffffffff",
            INIT_39 => X"fffffff7fffffffffffffff1ffffffff0000001700000000fffffff4ffffffff",
            INIT_3A => X"ffffffeaffffffffffffffaaffffffff0000002600000000ffffffa9ffffffff",
            INIT_3B => X"ffffffe0ffffffffffffffb9ffffffffffffffebffffffff0000001300000000",
            INIT_3C => X"ffffffc5ffffffff0000001d00000000ffffffe2fffffffffffffffeffffffff",
            INIT_3D => X"ffffffc9ffffffff0000003e000000000000001900000000ffffffe6ffffffff",
            INIT_3E => X"0000002600000000fffffff0ffffffffffffffceffffffff0000000500000000",
            INIT_3F => X"ffffffcdfffffffffffffffbffffffff00000011000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004400000000ffffffdfffffffffffffffdeffffffff0000001900000000",
            INIT_41 => X"000000040000000000000047000000000000004400000000ffffff84ffffffff",
            INIT_42 => X"0000003600000000ffffffddffffffff0000003e00000000ffffffb9ffffffff",
            INIT_43 => X"ffffffafffffffffffffffd7ffffffffffffffeeffffffff0000003e00000000",
            INIT_44 => X"0000000200000000fffffff7ffffffffffffffe0ffffffff0000007000000000",
            INIT_45 => X"00000019000000000000002f000000000000001800000000ffffff94ffffffff",
            INIT_46 => X"0000000300000000000000070000000000000034000000000000001000000000",
            INIT_47 => X"ffffffc3ffffffff0000000000000000fffffff8ffffffff0000004900000000",
            INIT_48 => X"0000000400000000fffffffdffffffff0000003900000000fffffffeffffffff",
            INIT_49 => X"fffffff5ffffffff000000190000000000000008000000000000003700000000",
            INIT_4A => X"00000043000000000000001c00000000ffffffd3ffffffff0000005600000000",
            INIT_4B => X"0000000900000000fffffff6fffffffffffffff9ffffffff0000004000000000",
            INIT_4C => X"00000002000000000000002500000000ffffffedffffffff0000001b00000000",
            INIT_4D => X"ffffffdaffffffff0000001f0000000000000024000000000000002000000000",
            INIT_4E => X"0000002e000000000000001500000000ffffffdaffffffff0000005800000000",
            INIT_4F => X"ffffffc6ffffffff0000000a00000000ffffffe7fffffffffffffff5ffffffff",
            INIT_50 => X"0000000500000000fffffff4ffffffff0000000e00000000ffffffe7ffffffff",
            INIT_51 => X"fffffffbffffffff0000001d0000000000000014000000000000002400000000",
            INIT_52 => X"0000001a00000000ffffffcfffffffffffffffddffffffff0000002000000000",
            INIT_53 => X"ffffffd6ffffffff0000004d000000000000000300000000ffffffc4ffffffff",
            INIT_54 => X"0000000b00000000ffffffdbffffffffffffffe9ffffffffffffffa8ffffffff",
            INIT_55 => X"0000001500000000fffffff6ffffffffffffffc9ffffffff0000001300000000",
            INIT_56 => X"00000029000000000000004c00000000ffffffbaffffffffffffffb1ffffffff",
            INIT_57 => X"0000000c00000000fffffff5ffffffff00000035000000000000001000000000",
            INIT_58 => X"ffffffd9ffffffff0000001f000000000000001800000000ffffffd3ffffffff",
            INIT_59 => X"0000002f00000000fffffff2ffffffffffffffcdffffffffffffffffffffffff",
            INIT_5A => X"fffffff1ffffffffffffffedffffffffffffffe8ffffffffffffffd1ffffffff",
            INIT_5B => X"ffffffe9ffffffffffffffe7ffffffffffffffdfffffffff0000002f00000000",
            INIT_5C => X"ffffffe4ffffffff0000001c000000000000000b00000000ffffff71ffffffff",
            INIT_5D => X"ffffffdfffffffff0000001700000000fffffff6ffffffffffffffd6ffffffff",
            INIT_5E => X"0000000c00000000ffffff87ffffffffffffffa6ffffffffffffffceffffffff",
            INIT_5F => X"ffffffe5ffffffff0000003b0000000000000009000000000000000000000000",
            INIT_60 => X"ffffffbeffffffff0000001000000000ffffff89ffffffffffffffc1ffffffff",
            INIT_61 => X"ffffffcfffffffffffffffbfffffffffffffffcbffffffff0000003200000000",
            INIT_62 => X"ffffffdcffffffffffffffd5ffffffffffffffffffffffffffffffaeffffffff",
            INIT_63 => X"fffffff0fffffffffffffff3ffffffff00000014000000000000003700000000",
            INIT_64 => X"ffffffe3ffffffff0000001600000000ffffff9dffffffff0000000a00000000",
            INIT_65 => X"ffffffceffffffff0000001b00000000fffffffaffffffffffffffe3ffffffff",
            INIT_66 => X"ffffffe6ffffffffffffffabffffffffffffffceffffffffffffffd2ffffffff",
            INIT_67 => X"0000000300000000fffffff5ffffffffffffffdaffffffff0000000400000000",
            INIT_68 => X"fffffff3ffffffff0000004800000000ffffff80ffffffff0000000000000000",
            INIT_69 => X"ffffffd5ffffffff000000080000000000000000000000000000003100000000",
            INIT_6A => X"ffffffd6ffffffffffffffbcffffffff",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "ifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE0;


    MEM_IFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "ifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE1;


    MEM_IFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "ifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "ifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE3;


    MEM_IFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "ifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE4;


    MEM_IFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "ifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE0 : if BRAM_NAME = "ifmap_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000d00000000000000000000000000000000000000000000000a00000000",
            INIT_0A => X"0000000000000000000000140000000000000017000000000000002400000000",
            INIT_0B => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002b00000000000000100000000000000016000000000000001200000000",
            INIT_0E => X"00000000000000000000000b000000000000001b000000000000001c00000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000002300000000",
            INIT_10 => X"0000001d0000000000000025000000000000001a000000000000000000000000",
            INIT_11 => X"0000001a00000000000000130000000000000006000000000000001b00000000",
            INIT_12 => X"000000470000000000000000000000000000000a000000000000000b00000000",
            INIT_13 => X"0000003300000000000000220000000000000008000000000000003000000000",
            INIT_14 => X"000000120000000000000011000000000000002e000000000000003c00000000",
            INIT_15 => X"0000000d00000000000000280000000000000040000000000000000000000000",
            INIT_16 => X"00000047000000000000003f0000000000000007000000000000001100000000",
            INIT_17 => X"0000001e00000000000000090000000000000000000000000000000300000000",
            INIT_18 => X"000000150000000000000016000000000000002c000000000000002d00000000",
            INIT_19 => X"0000000f0000000000000014000000000000001d000000000000003a00000000",
            INIT_1A => X"000000130000000000000033000000000000004b000000000000001400000000",
            INIT_1B => X"00000050000000000000001e0000000000000000000000000000000000000000",
            INIT_1C => X"00000039000000000000001c000000000000001a000000000000003200000000",
            INIT_1D => X"0000000b000000000000001f0000000000000011000000000000002000000000",
            INIT_1E => X"00000018000000000000004b0000000000000042000000000000005400000000",
            INIT_1F => X"000000130000000000000019000000000000002d000000000000001c00000000",
            INIT_20 => X"00000028000000000000000f0000000000000017000000000000000200000000",
            INIT_21 => X"0000004e00000000000000000000000000000003000000000000001200000000",
            INIT_22 => X"0000001b00000000000000210000000000000042000000000000004b00000000",
            INIT_23 => X"00000023000000000000001a0000000000000011000000000000002200000000",
            INIT_24 => X"0000000000000000000000030000000000000024000000000000002000000000",
            INIT_25 => X"0000004300000000000000340000000000000000000000000000000000000000",
            INIT_26 => X"0000001400000000000000440000000000000011000000000000004300000000",
            INIT_27 => X"000000170000000000000038000000000000004d000000000000003a00000000",
            INIT_28 => X"0000001400000000000000210000000000000013000000000000000400000000",
            INIT_29 => X"00000034000000000000004f0000000000000042000000000000001400000000",
            INIT_2A => X"00000042000000000000005a0000000000000083000000000000003c00000000",
            INIT_2B => X"0000003700000000000000300000000000000038000000000000003f00000000",
            INIT_2C => X"0000004500000000000000460000000000000041000000000000003d00000000",
            INIT_2D => X"00000065000000000000003c0000000000000045000000000000005000000000",
            INIT_2E => X"0000003a000000000000003d000000000000003b000000000000005900000000",
            INIT_2F => X"0000003e000000000000003b0000000000000037000000000000003700000000",
            INIT_30 => X"000000520000000000000043000000000000004a000000000000004a00000000",
            INIT_31 => X"00000041000000000000006b0000000000000042000000000000004400000000",
            INIT_32 => X"0000003c0000000000000039000000000000003f000000000000003b00000000",
            INIT_33 => X"0000004e000000000000004d000000000000004b000000000000004000000000",
            INIT_34 => X"0000004c000000000000005a000000000000006a000000000000004600000000",
            INIT_35 => X"0000003f000000000000003d0000000000000034000000000000005400000000",
            INIT_36 => X"00000042000000000000003d000000000000003f000000000000004300000000",
            INIT_37 => X"00000056000000000000003c0000000000000042000000000000004700000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000003000000000000000200000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_43 => X"0000003d00000000000000000000000000000001000000000000000a00000000",
            INIT_44 => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_45 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"00000000000000000000002e0000000000000000000000000000002600000000",
            INIT_48 => X"00000000000000000000000c0000000000000000000000000000003d00000000",
            INIT_49 => X"0000000000000000000000410000000000000000000000000000000000000000",
            INIT_4A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000007d000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4F => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_53 => X"0000002a000000000000002c0000000000000000000000000000000700000000",
            INIT_54 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_58 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_59 => X"00000010000000000000000f0000000000000000000000000000000000000000",
            INIT_5A => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5D => X"0000000d0000000000000000000000000000001c000000000000002000000000",
            INIT_5E => X"0000000000000000000000750000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000019000000000000001100000000",
            INIT_60 => X"000000140000000000000013000000000000000e000000000000000000000000",
            INIT_61 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000046000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000002d000000000000001d0000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000900000000000000000000000000000000000000000000000700000000",
            INIT_69 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000060000000000000005c0000000000000000000000000000000000000000",
            INIT_71 => X"0000005a00000000000000610000000000000061000000000000006000000000",
            INIT_72 => X"0000004d00000000000000680000000000000071000000000000006400000000",
            INIT_73 => X"00000050000000000000004a0000000000000043000000000000003d00000000",
            INIT_74 => X"000000630000000000000069000000000000005e000000000000005400000000",
            INIT_75 => X"0000004d00000000000000500000000000000061000000000000006400000000",
            INIT_76 => X"0000000000000000000000180000000000000039000000000000005500000000",
            INIT_77 => X"0000004d000000000000003b000000000000001d000000000000000200000000",
            INIT_78 => X"0000006b000000000000006a000000000000004a000000000000003c00000000",
            INIT_79 => X"0000001b00000000000000370000000000000054000000000000006900000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"00000000000000000000003a0000000000000006000000000000000000000000",
            INIT_7C => X"0000005700000000000000680000000000000058000000000000000a00000000",
            INIT_7D => X"0000000000000000000000000000000000000005000000000000003500000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000001a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE0;


    MEM_IFMAP_LAYER1_INSTANCE1 : if BRAM_NAME = "ifmap_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000038000000000000003b00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000d000000000000004e00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000056000000000000001f0000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000006000000000000000d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000006000000000000001c0000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_0F => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_10 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000c00000000000000000000000000000000000000000000000500000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000004300000000000000260000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000ba00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000bf00000000000000c200000000000000bd00000000000000c100000000",
            INIT_2A => X"000000bb00000000000000c200000000000000c600000000000000bc00000000",
            INIT_2B => X"000000a7000000000000009f00000000000000a500000000000000b500000000",
            INIT_2C => X"000000bd00000000000000b5000000000000009e00000000000000aa00000000",
            INIT_2D => X"000000e300000000000000bf00000000000000c900000000000000c200000000",
            INIT_2E => X"0000008600000000000000ac00000000000000c100000000000000e300000000",
            INIT_2F => X"0000008b000000000000007e000000000000008f00000000000000a100000000",
            INIT_30 => X"000000c0000000000000008800000000000000b600000000000000a300000000",
            INIT_31 => X"000000bf00000000000000ea00000000000000c200000000000000c300000000",
            INIT_32 => X"000000de00000000000000a20000000000000061000000000000007e00000000",
            INIT_33 => X"0000008e000000000000006900000000000000a700000000000000ae00000000",
            INIT_34 => X"000000bf00000000000000c8000000000000006800000000000000c800000000",
            INIT_35 => X"000000a300000000000000d5000000000000009e00000000000000d000000000",
            INIT_36 => X"000000ad00000000000000ef00000000000000a0000000000000009200000000",
            INIT_37 => X"00000103000000000000005e0000000000000062000000000000008e00000000",
            INIT_38 => X"0000014400000000000000b000000000000000f200000000000000ed00000000",
            INIT_39 => X"0000008a00000000000000b50000000000000115000000000000012f00000000",
            INIT_3A => X"0000008c00000000000000ce00000000000000f7000000000000006200000000",
            INIT_3B => X"00000118000000000000011e0000000000000056000000000000007d00000000",
            INIT_3C => X"0000011500000000000000f000000000000000db000000000000010300000000",
            INIT_3D => X"0000007a00000000000000a800000000000000d2000000000000012b00000000",
            INIT_3E => X"00000097000000000000009000000000000000c7000000000000014600000000",
            INIT_3F => X"000000c000000000000001450000000000000113000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000015000000000000000ed00000000000000ac00000000000000c600000000",
            INIT_41 => X"0000012700000000000000be00000000000000cc000000000000010300000000",
            INIT_42 => X"000000a70000000000000096000000000000008c00000000000000ba00000000",
            INIT_43 => X"000000d000000000000000de0000000000000139000000000000013900000000",
            INIT_44 => X"000000de0000000000000146000000000000012400000000000000ac00000000",
            INIT_45 => X"000000c0000000000000010600000000000000cd00000000000000b000000000",
            INIT_46 => X"0000016200000000000000a000000000000000b8000000000000008500000000",
            INIT_47 => X"000000e200000000000000c40000000000000114000000000000014600000000",
            INIT_48 => X"0000009900000000000000bd00000000000000c600000000000000cc00000000",
            INIT_49 => X"00000061000000000000009e00000000000000a800000000000000ec00000000",
            INIT_4A => X"00000149000000000000014900000000000000b7000000000000008400000000",
            INIT_4B => X"000000a800000000000000f500000000000000ca000000000000012a00000000",
            INIT_4C => X"000000b600000000000000d5000000000000011700000000000000b300000000",
            INIT_4D => X"000000b200000000000000610000000000000043000000000000009b00000000",
            INIT_4E => X"0000012e0000000000000146000000000000010900000000000000c800000000",
            INIT_4F => X"0000010f0000000000000109000000000000018d00000000000000d400000000",
            INIT_50 => X"00000058000000000000009100000000000000e9000000000000013700000000",
            INIT_51 => X"000000aa00000000000000ad0000000000000091000000000000006f00000000",
            INIT_52 => X"000001790000000000000128000000000000010e00000000000000cc00000000",
            INIT_53 => X"0000009c00000000000000a300000000000000c700000000000001c800000000",
            INIT_54 => X"00000093000000000000008a0000000000000083000000000000008900000000",
            INIT_55 => X"000000b200000000000000a600000000000000ab000000000000009a00000000",
            INIT_56 => X"000000ff00000000000001c000000000000000e500000000000000b500000000",
            INIT_57 => X"00000087000000000000008c0000000000000097000000000000009500000000",
            INIT_58 => X"000000b400000000000000a1000000000000008f000000000000008500000000",
            INIT_59 => X"0000009500000000000000ae00000000000000b000000000000000aa00000000",
            INIT_5A => X"0000009a00000000000000ac000000000000016a00000000000000bb00000000",
            INIT_5B => X"00000096000000000000008b000000000000008f000000000000009f00000000",
            INIT_5C => X"0000009e000000000000009e00000000000000a300000000000000a200000000",
            INIT_5D => X"000000a3000000000000009500000000000000c100000000000000db00000000",
            INIT_5E => X"0000008f000000000000007c000000000000008b00000000000000ae00000000",
            INIT_5F => X"000000aa00000000000000ad000000000000009d000000000000009200000000",
            INIT_60 => X"000000af00000000000000f300000000000000a7000000000000009000000000",
            INIT_61 => X"0000007b0000000000000078000000000000007e000000000000007600000000",
            INIT_62 => X"0000008500000000000000820000000000000074000000000000007700000000",
            INIT_63 => X"0000006200000000000000620000000000000070000000000000007b00000000",
            INIT_64 => X"000000750000000000000067000000000000006a000000000000006200000000",
            INIT_65 => X"000000770000000000000080000000000000007e000000000000007d00000000",
            INIT_66 => X"0000005f00000000000000790000000000000079000000000000006f00000000",
            INIT_67 => X"0000003f000000000000002e0000000000000026000000000000003400000000",
            INIT_68 => X"00000063000000000000006e0000000000000065000000000000005b00000000",
            INIT_69 => X"00000084000000000000007d0000000000000081000000000000007d00000000",
            INIT_6A => X"00000016000000000000001f0000000000000037000000000000006200000000",
            INIT_6B => X"0000002f00000000000000250000000000000021000000000000003200000000",
            INIT_6C => X"0000007c000000000000001c0000000000000040000000000000005900000000",
            INIT_6D => X"0000004500000000000000420000000000000077000000000000007c00000000",
            INIT_6E => X"0000004100000000000000260000000000000018000000000000002100000000",
            INIT_6F => X"0000003a000000000000001d0000000000000023000000000000003000000000",
            INIT_70 => X"0000005000000000000000740000000000000034000000000000003200000000",
            INIT_71 => X"0000002e000000000000004f0000000000000031000000000000006200000000",
            INIT_72 => X"0000003100000000000000400000000000000000000000000000002100000000",
            INIT_73 => X"000000270000000000000015000000000000001b000000000000001d00000000",
            INIT_74 => X"0000006f000000000000004e0000000000000077000000000000004e00000000",
            INIT_75 => X"000000270000000000000039000000000000005d000000000000005600000000",
            INIT_76 => X"0000002200000000000000360000000000000051000000000000000300000000",
            INIT_77 => X"00000054000000000000001f000000000000000d000000000000001900000000",
            INIT_78 => X"00000040000000000000003d0000000000000075000000000000006900000000",
            INIT_79 => X"0000001300000000000000400000000000000039000000000000007200000000",
            INIT_7A => X"0000001a00000000000000130000000000000029000000000000004f00000000",
            INIT_7B => X"0000002c0000000000000049000000000000002d000000000000002900000000",
            INIT_7C => X"000000500000000000000060000000000000002e000000000000005700000000",
            INIT_7D => X"000000490000000000000031000000000000003c000000000000004300000000",
            INIT_7E => X"00000042000000000000002f000000000000001b000000000000003300000000",
            INIT_7F => X"0000003d000000000000002d0000000000000040000000000000003c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE1;


    MEM_IFMAP_LAYER1_INSTANCE2 : if BRAM_NAME = "ifmap_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003200000000000000450000000000000039000000000000003000000000",
            INIT_01 => X"0000003100000000000000550000000000000036000000000000002800000000",
            INIT_02 => X"0000004b000000000000005f000000000000003c000000000000001100000000",
            INIT_03 => X"00000054000000000000000c0000000000000046000000000000003f00000000",
            INIT_04 => X"000000240000000000000042000000000000001c000000000000001500000000",
            INIT_05 => X"00000017000000000000000a0000000000000029000000000000005000000000",
            INIT_06 => X"000000400000000000000039000000000000006c000000000000004e00000000",
            INIT_07 => X"00000024000000000000003e000000000000000e000000000000004600000000",
            INIT_08 => X"000000010000000000000033000000000000004c000000000000002100000000",
            INIT_09 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000003c0000000000000028000000000000000b000000000000001400000000",
            INIT_0B => X"00000000000000000000001b0000000000000073000000000000003b00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000006e000000000000000f0000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000005000000000000000500000000",
            INIT_1B => X"0000000300000000000000050000000000000008000000000000000400000000",
            INIT_1C => X"0000000c00000000000000060000000000000000000000000000000000000000",
            INIT_1D => X"0000000600000000000000000000000000000000000000000000000100000000",
            INIT_1E => X"00000009000000000000001a0000000000000000000000000000000000000000",
            INIT_1F => X"00000008000000000000000b0000000000000000000000000000000a00000000",
            INIT_20 => X"0000001a00000000000000060000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000012000000000000002b000000000000000000000000",
            INIT_23 => X"0000001f00000000000000110000000000000017000000000000000000000000",
            INIT_24 => X"00000000000000000000005a0000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000016000000000000000e00000000",
            INIT_27 => X"0000001600000000000000220000000000000002000000000000003500000000",
            INIT_28 => X"0000001e00000000000000000000000000000048000000000000000000000000",
            INIT_29 => X"0000003400000000000000060000000000000005000000000000000000000000",
            INIT_2A => X"0000000d0000000000000000000000000000001b000000000000003000000000",
            INIT_2B => X"0000000000000000000000270000000000000004000000000000003300000000",
            INIT_2C => X"00000005000000000000002c0000000000000000000000000000003200000000",
            INIT_2D => X"0000002400000000000000320000000000000006000000000000000000000000",
            INIT_2E => X"00000040000000000000003c0000000000000000000000000000004200000000",
            INIT_2F => X"0000003100000000000000140000000000000018000000000000000000000000",
            INIT_30 => X"00000000000000000000003a0000000000000000000000000000001e00000000",
            INIT_31 => X"000000420000000000000027000000000000000c000000000000000000000000",
            INIT_32 => X"00000000000000000000002d0000000000000045000000000000000000000000",
            INIT_33 => X"0000002200000000000000230000000000000019000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_35 => X"000000000000000000000027000000000000000b000000000000005400000000",
            INIT_36 => X"0000000000000000000000000000000000000036000000000000002900000000",
            INIT_37 => X"0000005d0000000000000000000000000000002d000000000000001200000000",
            INIT_38 => X"0000001800000000000000000000000000000016000000000000000000000000",
            INIT_39 => X"0000000000000000000000120000000000000000000000000000001000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_3B => X"0000000000000000000000650000000000000000000000000000000e00000000",
            INIT_3C => X"0000001500000000000000000000000000000006000000000000002800000000",
            INIT_3D => X"000000000000000000000033000000000000000d000000000000000f00000000",
            INIT_3E => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_3F => X"000000560000000000000000000000000000005a000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003e000000000000000e0000000000000000000000000000001300000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003900000000000000610000000000000000000000000000001300000000",
            INIT_44 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000000b000000000000000500000000",
            INIT_47 => X"000000010000000000000000000000000000007f000000000000000c00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000005100000000000000000000000000000000000000000000001600000000",
            INIT_4B => X"00000000000000000000000b0000000000000000000000000000002100000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000002000000000000000080000000000000000000000000000000100000000",
            INIT_4E => X"0000000b00000000000000010000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000002c000000000000001200000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001e00000000000000040000000000000004000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_5C => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_72 => X"0000000000000000000000070000000000000003000000000000003400000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_75 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_7A => X"0000001900000000000000060000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001c0000000000000031000000000000002a000000000000003f00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7E => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000002d0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE2;


    MEM_IFMAP_LAYER1_INSTANCE3 : if BRAM_NAME = "ifmap_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_06 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000050000000000000011000000000000000900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000004000000000000000200000000",
            INIT_0B => X"0000000200000000000000000000000000000000000000000000000700000000",
            INIT_0C => X"00000007000000000000000b0000000000000003000000000000000000000000",
            INIT_0D => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_0E => X"0000001f00000000000000070000000000000000000000000000000400000000",
            INIT_0F => X"0000001f00000000000000000000000000000001000000000000000000000000",
            INIT_10 => X"0000000f000000000000000b0000000000000000000000000000000000000000",
            INIT_11 => X"0000000100000000000000260000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_13 => X"00000000000000000000002a000000000000000b000000000000000000000000",
            INIT_14 => X"0000001500000000000000040000000000000000000000000000000000000000",
            INIT_15 => X"0000000a00000000000000000000000000000039000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_18 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000003a0000000000000000000000000000000f00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000100000000000000000000000000000000000000000000004b00000000",
            INIT_1C => X"0000000c00000000000000000000000000000009000000000000000000000000",
            INIT_1D => X"0000000000000000000000490000000000000000000000000000000000000000",
            INIT_1E => X"0000008100000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000002f000000000000003a000000000000000000000000",
            INIT_22 => X"0000000000000000000000600000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000c0000000000000003000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000002b000000000000001b00000000",
            INIT_26 => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_28 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_29 => X"0000001800000000000000000000000000000000000000000000000100000000",
            INIT_2A => X"000000110000000000000000000000000000000b000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2C => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_2E => X"0000001400000000000000220000000000000004000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_30 => X"0000001a00000000000000000000000000000000000000000000007200000000",
            INIT_31 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000d0000000000000010000000000000000d00000000",
            INIT_33 => X"0000003a00000000000000000000000000000021000000000000001f00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000045000000000000001a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000050000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_42 => X"0000004600000000000000440000000000000045000000000000003f00000000",
            INIT_43 => X"0000004b00000000000000470000000000000041000000000000004300000000",
            INIT_44 => X"0000002d000000000000002a0000000000000034000000000000004300000000",
            INIT_45 => X"00000043000000000000003b000000000000003d000000000000003500000000",
            INIT_46 => X"0000004400000000000000480000000000000049000000000000004800000000",
            INIT_47 => X"0000002200000000000000380000000000000041000000000000004500000000",
            INIT_48 => X"00000015000000000000000e000000000000000e000000000000001100000000",
            INIT_49 => X"00000025000000000000002b0000000000000038000000000000002700000000",
            INIT_4A => X"0000003100000000000000470000000000000049000000000000004400000000",
            INIT_4B => X"0000000d000000000000000d000000000000000e000000000000002000000000",
            INIT_4C => X"00000010000000000000000f0000000000000011000000000000001500000000",
            INIT_4D => X"0000003c0000000000000019000000000000001c000000000000002900000000",
            INIT_4E => X"00000023000000000000001e000000000000003a000000000000004300000000",
            INIT_4F => X"00000019000000000000000c000000000000000b000000000000001500000000",
            INIT_50 => X"00000019000000000000000c000000000000000a000000000000001100000000",
            INIT_51 => X"0000002e000000000000003a0000000000000022000000000000001600000000",
            INIT_52 => X"000000150000000000000020000000000000002c000000000000003b00000000",
            INIT_53 => X"0000001a000000000000001d0000000000000004000000000000000a00000000",
            INIT_54 => X"00000009000000000000000e000000000000000f000000000000000f00000000",
            INIT_55 => X"00000011000000000000002a000000000000003c000000000000001600000000",
            INIT_56 => X"00000014000000000000001d0000000000000026000000000000001e00000000",
            INIT_57 => X"0000000d000000000000000f000000000000001b000000000000000b00000000",
            INIT_58 => X"00000011000000000000000e0000000000000010000000000000000c00000000",
            INIT_59 => X"0000001b000000000000001b0000000000000036000000000000002300000000",
            INIT_5A => X"0000000700000000000000180000000000000017000000000000001f00000000",
            INIT_5B => X"0000000b00000000000000080000000000000010000000000000001400000000",
            INIT_5C => X"0000001600000000000000110000000000000011000000000000001900000000",
            INIT_5D => X"00000016000000000000001f000000000000001c000000000000002300000000",
            INIT_5E => X"0000001700000000000000170000000000000018000000000000000d00000000",
            INIT_5F => X"0000002700000000000000140000000000000008000000000000000f00000000",
            INIT_60 => X"0000000f000000000000000c000000000000000a000000000000000f00000000",
            INIT_61 => X"0000001200000000000000150000000000000009000000000000001700000000",
            INIT_62 => X"0000000800000000000000120000000000000014000000000000001100000000",
            INIT_63 => X"0000000f000000000000003a0000000000000020000000000000000800000000",
            INIT_64 => X"0000001700000000000000000000000000000011000000000000000e00000000",
            INIT_65 => X"00000015000000000000001b000000000000000c000000000000000f00000000",
            INIT_66 => X"0000001400000000000000000000000000000004000000000000001200000000",
            INIT_67 => X"0000000c00000000000000000000000000000035000000000000002d00000000",
            INIT_68 => X"000000190000000000000023000000000000000c000000000000000e00000000",
            INIT_69 => X"0000000000000000000000060000000000000000000000000000000500000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE3;


    MEM_IFMAP_LAYER1_INSTANCE4 : if BRAM_NAME = "ifmap_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000150000000000000010000000000000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000003000000000000000600000000",
            INIT_27 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_28 => X"0000000400000000000000020000000000000000000000000000000000000000",
            INIT_29 => X"00000009000000000000000a0000000000000006000000000000000400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2B => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_2C => X"0000000600000000000000030000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000030000000000000006000000000000000700000000",
            INIT_2E => X"0000000500000000000000000000000000000003000000000000000300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_30 => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000002000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000004000000000000001c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000003000000000000000a0000000000000004000000000000000000000000",
            INIT_75 => X"000000000000000000000000000000000000000a000000000000000b00000000",
            INIT_76 => X"000000000000000000000000000000000000001a000000000000002500000000",
            INIT_77 => X"0000000a000000000000001e0000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000005f00000000000000000000000000000000000000000000003800000000",
            INIT_7B => X"0000000000000000000000070000000000000001000000000000003600000000",
            INIT_7C => X"0000000a0000000000000016000000000000001e000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000d000000000000001d0000000000000018000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE4;


    MEM_IFMAP_LAYER1_INSTANCE5 : if BRAM_NAME = "ifmap_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000e000000000000002200000000",
            INIT_02 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_04 => X"00000010000000000000000c0000000000000000000000000000000900000000",
            INIT_05 => X"0000001200000000000000180000000000000013000000000000000900000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0A => X"0000000600000000000000070000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0D => X"0000000000000000000000020000000000000002000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000035000000000000000200000000",
            INIT_0F => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000005c0000000000000080000000000000002e00000000",
            INIT_12 => X"00000029000000000000000d0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000013000000000000003400000000",
            INIT_14 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"0000000a00000000000000040000000000000005000000000000000a00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000500000000000000010000000000000002000000000000000500000000",
            INIT_1A => X"0000000000000000000000190000000000000013000000000000000c00000000",
            INIT_1B => X"0000000300000000000000070000000000000023000000000000000000000000",
            INIT_1C => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000700000000000000010000000000000006000000000000001100000000",
            INIT_1E => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000030000000000000009000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000a000000000000001b0000000000000014000000000000000000000000",
            INIT_22 => X"0000000e0000000000000023000000000000002c000000000000000600000000",
            INIT_23 => X"0000003400000000000000340000000000000032000000000000003300000000",
            INIT_24 => X"0000003900000000000000350000000000000030000000000000003700000000",
            INIT_25 => X"000000280000000000000025000000000000002c000000000000003600000000",
            INIT_26 => X"00000037000000000000002f000000000000002d000000000000002900000000",
            INIT_27 => X"0000003700000000000000340000000000000038000000000000003400000000",
            INIT_28 => X"00000020000000000000002a0000000000000029000000000000003400000000",
            INIT_29 => X"0000002100000000000000170000000000000013000000000000001f00000000",
            INIT_2A => X"00000035000000000000001e000000000000002d000000000000002b00000000",
            INIT_2B => X"0000003800000000000000390000000000000037000000000000003600000000",
            INIT_2C => X"000000210000000000000013000000000000001a000000000000001600000000",
            INIT_2D => X"00000021000000000000000f000000000000000a000000000000000100000000",
            INIT_2E => X"00000032000000000000003d0000000000000000000000000000002d00000000",
            INIT_2F => X"000000130000000000000028000000000000002b000000000000003a00000000",
            INIT_30 => X"000000000000000000000023000000000000000f000000000000000600000000",
            INIT_31 => X"00000037000000000000000e0000000000000004000000000000000c00000000",
            INIT_32 => X"0000003e00000000000000210000000000000025000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000a000000000000000f00000000",
            INIT_34 => X"00000000000000000000000b000000000000002b000000000000000900000000",
            INIT_35 => X"0000000000000000000000250000000000000009000000000000001100000000",
            INIT_36 => X"00000018000000000000001d0000000000000012000000000000000e00000000",
            INIT_37 => X"0000000300000000000000070000000000000000000000000000000000000000",
            INIT_38 => X"0000001400000000000000000000000000000000000000000000003b00000000",
            INIT_39 => X"000000040000000000000000000000000000000c000000000000000900000000",
            INIT_3A => X"0000001700000000000000340000000000000018000000000000001900000000",
            INIT_3B => X"0000003900000000000000000000000000000000000000000000000400000000",
            INIT_3C => X"0000001100000000000000130000000000000000000000000000000000000000",
            INIT_3D => X"0000000d00000000000000000000000000000000000000000000000700000000",
            INIT_3E => X"000000000000000000000017000000000000002d000000000000001500000000",
            INIT_3F => X"0000000000000000000000310000000000000000000000000000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000000c0000000000000014000000000000000000000000",
            INIT_41 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000f000000000000000a0000000000000013000000000000000300000000",
            INIT_43 => X"00000000000000000000000e0000000000000020000000000000001b00000000",
            INIT_44 => X"0000000000000000000000300000000000000026000000000000001400000000",
            INIT_45 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_46 => X"0000000500000000000000050000000000000019000000000000000800000000",
            INIT_47 => X"00000020000000000000000e0000000000000002000000000000000400000000",
            INIT_48 => X"0000000000000000000000110000000000000029000000000000003300000000",
            INIT_49 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_4A => X"0000000400000000000000000000000000000000000000000000000700000000",
            INIT_4B => X"00000015000000000000000b0000000000000004000000000000000700000000",
            INIT_4C => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"00000000000000000000000b0000000000000008000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000f0000000000000003000000000000000e000000000000000000000000",
            INIT_66 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_69 => X"0000000600000000000000070000000000000008000000000000000700000000",
            INIT_6A => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_6B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_6D => X"0000000000000000000000050000000000000000000000000000000200000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_70 => X"0000000c00000000000000180000000000000000000000000000000c00000000",
            INIT_71 => X"0000000900000000000000000000000000000005000000000000000200000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_73 => X"0000000f00000000000000000000000000000015000000000000000000000000",
            INIT_74 => X"0000000200000000000000050000000000000017000000000000000000000000",
            INIT_75 => X"0000001800000000000000110000000000000000000000000000000000000000",
            INIT_76 => X"0000000400000000000000000000000000000000000000000000000300000000",
            INIT_77 => X"0000000000000000000000000000000000000015000000000000002500000000",
            INIT_78 => X"000000080000000000000004000000000000000c000000000000000e00000000",
            INIT_79 => X"0000002200000000000000230000000000000023000000000000000000000000",
            INIT_7A => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000001000000000000001700000000",
            INIT_7D => X"0000001000000000000000290000000000000021000000000000001900000000",
            INIT_7E => X"0000000200000000000000000000000000000000000000000000001100000000",
            INIT_7F => X"0000000700000000000000200000000000000007000000000000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE6 : if BRAM_NAME = "ifmap_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000f0000000000000000000000000000002c000000000000001600000000",
            INIT_02 => X"0000002f000000000000003c0000000000000029000000000000000b00000000",
            INIT_03 => X"00000034000000000000001f0000000000000011000000000000001800000000",
            INIT_04 => X"000000320000000000000067000000000000002a000000000000003100000000",
            INIT_05 => X"0000005000000000000000710000000000000010000000000000001100000000",
            INIT_06 => X"0000004500000000000000460000000000000048000000000000004d00000000",
            INIT_07 => X"0000005700000000000000510000000000000053000000000000004f00000000",
            INIT_08 => X"0000000a0000000000000059000000000000006f000000000000005400000000",
            INIT_09 => X"0000004f0000000000000048000000000000004d000000000000004500000000",
            INIT_0A => X"00000052000000000000004a0000000000000049000000000000004900000000",
            INIT_0B => X"0000005400000000000000600000000000000061000000000000005300000000",
            INIT_0C => X"0000006600000000000000440000000000000062000000000000006f00000000",
            INIT_0D => X"0000004b000000000000004b000000000000004a000000000000004100000000",
            INIT_0E => X"0000006700000000000000610000000000000052000000000000004d00000000",
            INIT_0F => X"0000006f000000000000008a000000000000005d000000000000006500000000",
            INIT_10 => X"00000051000000000000005a0000000000000063000000000000006700000000",
            INIT_11 => X"00000048000000000000004b0000000000000056000000000000005300000000",
            INIT_12 => X"000000450000000000000054000000000000005b000000000000004e00000000",
            INIT_13 => X"0000003900000000000000380000000000000071000000000000006d00000000",
            INIT_14 => X"0000003600000000000000340000000000000036000000000000003900000000",
            INIT_15 => X"0000002d0000000000000034000000000000003f000000000000003e00000000",
            INIT_16 => X"00000030000000000000002f0000000000000030000000000000002c00000000",
            INIT_17 => X"0000003b000000000000003b0000000000000036000000000000002c00000000",
            INIT_18 => X"00000029000000000000001c0000000000000036000000000000003900000000",
            INIT_19 => X"00000000000000000000000b000000000000002b000000000000003300000000",
            INIT_1A => X"0000002d0000000000000030000000000000001d000000000000000300000000",
            INIT_1B => X"0000003b000000000000003c0000000000000043000000000000002700000000",
            INIT_1C => X"0000000900000000000000160000000000000028000000000000003c00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1E => X"00000000000000000000002e000000000000001c000000000000000000000000",
            INIT_1F => X"0000002600000000000000370000000000000036000000000000001c00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_22 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000029000000000000002100000000",
            INIT_24 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001f00000000000000000000000000000000000000000000001700000000",
            INIT_27 => X"00000000000000000000000a000000000000001d000000000000002900000000",
            INIT_28 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000019000000000000002a0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000007000000000000001700000000",
            INIT_2C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000f00000000000000090000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_31 => X"000000000000000000000000000000000000000d000000000000000300000000",
            INIT_32 => X"0000000700000000000000020000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_34 => X"0000001200000000000000080000000000000000000000000000001100000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_38 => X"0000001f000000000000001c0000000000000009000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"00000048000000000000004b000000000000004b000000000000004400000000",
            INIT_4D => X"000000470000000000000051000000000000004e000000000000004200000000",
            INIT_4E => X"000000390000000000000033000000000000002e000000000000003700000000",
            INIT_4F => X"000000480000000000000049000000000000003f000000000000004000000000",
            INIT_50 => X"0000001e000000000000004e000000000000004b000000000000004d00000000",
            INIT_51 => X"0000001500000000000000260000000000000034000000000000004c00000000",
            INIT_52 => X"000000350000000000000018000000000000000c000000000000000700000000",
            INIT_53 => X"0000004e0000000000000035000000000000001a000000000000003d00000000",
            INIT_54 => X"000000240000000000000019000000000000004e000000000000004c00000000",
            INIT_55 => X"0000001000000000000000000000000000000023000000000000001800000000",
            INIT_56 => X"0000002a00000000000000220000000000000002000000000000001000000000",
            INIT_57 => X"00000048000000000000004c0000000000000014000000000000000600000000",
            INIT_58 => X"0000001f0000000000000012000000000000002e000000000000002d00000000",
            INIT_59 => X"0000001200000000000000090000000000000019000000000000000800000000",
            INIT_5A => X"0000001f0000000000000020000000000000000f000000000000000a00000000",
            INIT_5B => X"000000110000000000000059000000000000004f000000000000000000000000",
            INIT_5C => X"0000000000000000000000120000000000000010000000000000002c00000000",
            INIT_5D => X"00000006000000000000001a0000000000000015000000000000001f00000000",
            INIT_5E => X"0000000000000000000000330000000000000019000000000000000700000000",
            INIT_5F => X"0000003900000000000000000000000000000033000000000000005600000000",
            INIT_60 => X"0000000e0000000000000000000000000000001a000000000000000400000000",
            INIT_61 => X"0000000b000000000000000c000000000000001a000000000000001400000000",
            INIT_62 => X"0000004100000000000000000000000000000047000000000000001200000000",
            INIT_63 => X"00000003000000000000001b0000000000000000000000000000003100000000",
            INIT_64 => X"0000001700000000000000000000000000000008000000000000001700000000",
            INIT_65 => X"0000001b000000000000000e0000000000000007000000000000001200000000",
            INIT_66 => X"00000020000000000000002f0000000000000000000000000000003100000000",
            INIT_67 => X"00000009000000000000000e000000000000000c000000000000002d00000000",
            INIT_68 => X"0000000e000000000000000f0000000000000002000000000000001c00000000",
            INIT_69 => X"0000001100000000000000350000000000000011000000000000000d00000000",
            INIT_6A => X"0000002c0000000000000001000000000000001c000000000000000000000000",
            INIT_6B => X"0000001e0000000000000000000000000000001b000000000000001100000000",
            INIT_6C => X"0000000a000000000000000a0000000000000019000000000000000000000000",
            INIT_6D => X"000000070000000000000004000000000000003c000000000000002200000000",
            INIT_6E => X"0000002200000000000000250000000000000000000000000000000200000000",
            INIT_6F => X"0000001c000000000000001b0000000000000000000000000000001a00000000",
            INIT_70 => X"0000002300000000000000080000000000000009000000000000000000000000",
            INIT_71 => X"00000000000000000000000d0000000000000000000000000000003900000000",
            INIT_72 => X"00000000000000000000001f0000000000000003000000000000000e00000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000080000000000000000000000000000001c000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE6;


    MEM_IFMAP_LAYER1_INSTANCE7 : if BRAM_NAME = "ifmap_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE7;


    MEM_IFMAP_LAYER2_INSTANCE0 : if BRAM_NAME = "ifmap_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000000000000000000000000000000000001400000000",
            INIT_01 => X"000000d200000000000000360000000000000048000000000000002900000000",
            INIT_02 => X"0000007c00000000000000810000000000000045000000000000002f00000000",
            INIT_03 => X"00000064000000000000009a000000000000009a000000000000008200000000",
            INIT_04 => X"000000c5000000000000012000000000000000b6000000000000000300000000",
            INIT_05 => X"000000480000000000000093000000000000006b000000000000003a00000000",
            INIT_06 => X"0000001d00000000000000a800000000000000a800000000000000aa00000000",
            INIT_07 => X"0000002300000000000000860000000000000118000000000000005500000000",
            INIT_08 => X"0000004c000000000000001a0000000000000052000000000000004f00000000",
            INIT_09 => X"00000032000000000000001200000000000000c100000000000000a400000000",
            INIT_0A => X"0000002a000000000000006a0000000000000004000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000004400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000007500000000000000ba00000000000000a8000000000000008700000000",
            INIT_0E => X"0000003300000000000000bf000000000000005200000000000000d100000000",
            INIT_0F => X"0000000000000000000000560000000000000002000000000000000000000000",
            INIT_10 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_11 => X"000000540000000000000030000000000000001a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000003e00000000000000380000000000000000000000000000000000000000",
            INIT_14 => X"000000550000000000000050000000000000001d000000000000000900000000",
            INIT_15 => X"0000003700000000000000000000000000000000000000000000001600000000",
            INIT_16 => X"0000001a00000000000000130000000000000000000000000000001f00000000",
            INIT_17 => X"0000000400000000000000100000000000000019000000000000001c00000000",
            INIT_18 => X"0000000b00000000000000000000000000000000000000000000000100000000",
            INIT_19 => X"00000039000000000000000e0000000000000000000000000000001400000000",
            INIT_1A => X"0000004e0000000000000023000000000000007d000000000000000700000000",
            INIT_1B => X"0000003200000000000000430000000000000021000000000000004200000000",
            INIT_1C => X"00000068000000000000002c000000000000004b000000000000008500000000",
            INIT_1D => X"00000072000000000000004d0000000000000057000000000000005800000000",
            INIT_1E => X"000000440000000000000033000000000000002b000000000000004700000000",
            INIT_1F => X"0000006b00000000000000020000000000000029000000000000002300000000",
            INIT_20 => X"0000004000000000000000400000000000000057000000000000007c00000000",
            INIT_21 => X"00000085000000000000007d0000000000000000000000000000002b00000000",
            INIT_22 => X"0000001e0000000000000034000000000000002a000000000000001700000000",
            INIT_23 => X"0000000900000000000000110000000000000022000000000000001f00000000",
            INIT_24 => X"0000010700000000000000150000000000000000000000000000000800000000",
            INIT_25 => X"0000009d00000000000000e100000000000000d300000000000000fe00000000",
            INIT_26 => X"0000010e00000000000000ab00000000000000d1000000000000008900000000",
            INIT_27 => X"0000001b0000000000000040000000000000004c000000000000008e00000000",
            INIT_28 => X"0000002d000000000000006e000000000000002a000000000000006700000000",
            INIT_29 => X"0000001f00000000000000230000000000000027000000000000000700000000",
            INIT_2A => X"0000001d00000000000000190000000000000087000000000000000000000000",
            INIT_2B => X"000000000000000000000045000000000000001c000000000000001f00000000",
            INIT_2C => X"0000000f00000000000000000000000000000011000000000000000b00000000",
            INIT_2D => X"000000000000000000000000000000000000004e000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000005b000000000000004b0000000000000029000000000000003900000000",
            INIT_32 => X"00000097000000000000004c000000000000004e000000000000007500000000",
            INIT_33 => X"000000b20000000000000049000000000000005b000000000000007f00000000",
            INIT_34 => X"0000007a00000000000000400000000000000056000000000000002a00000000",
            INIT_35 => X"0000004100000000000001270000000000000039000000000000006400000000",
            INIT_36 => X"000000c30000000000000084000000000000002f000000000000003b00000000",
            INIT_37 => X"0000003d000000000000003b00000000000000bc000000000000004000000000",
            INIT_38 => X"00000051000000000000002100000000000000a5000000000000003900000000",
            INIT_39 => X"0000005200000000000000700000000000000025000000000000004700000000",
            INIT_3A => X"000000000000000000000000000000000000000000000000000000be00000000",
            INIT_3B => X"0000006600000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000002a00000000000000090000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_4B => X"0000004300000000000000120000000000000007000000000000000000000000",
            INIT_4C => X"000000000000000000000073000000000000002c000000000000006d00000000",
            INIT_4D => X"000000c800000000000000640000000000000090000000000000007a00000000",
            INIT_4E => X"000000720000000000000024000000000000009e000000000000007700000000",
            INIT_4F => X"00000049000000000000006b0000000000000026000000000000003c00000000",
            INIT_50 => X"000000960000000000000074000000000000001d000000000000005a00000000",
            INIT_51 => X"00000010000000000000005b000000000000006600000000000000a100000000",
            INIT_52 => X"0000007c00000000000000dd0000000000000025000000000000000000000000",
            INIT_53 => X"0000000b000000000000002e0000000000000035000000000000000000000000",
            INIT_54 => X"0000000b00000000000000040000000000000010000000000000000000000000",
            INIT_55 => X"000000380000000000000038000000000000001d000000000000001c00000000",
            INIT_56 => X"000000680000000000000083000000000000002b000000000000000400000000",
            INIT_57 => X"0000006700000000000000710000000000000060000000000000004300000000",
            INIT_58 => X"0000000000000000000000510000000000000000000000000000003500000000",
            INIT_59 => X"0000000000000000000000500000000000000000000000000000004800000000",
            INIT_5A => X"0000000000000000000000000000000000000081000000000000000000000000",
            INIT_5B => X"0000001500000000000000540000000000000045000000000000000000000000",
            INIT_5C => X"0000000d00000000000000000000000000000007000000000000003b00000000",
            INIT_5D => X"000000310000000000000000000000000000001f000000000000007300000000",
            INIT_5E => X"0000002f000000000000005f000000000000003f000000000000004c00000000",
            INIT_5F => X"000000000000000000000000000000000000002a000000000000000200000000",
            INIT_60 => X"0000001500000000000000620000000000000029000000000000000000000000",
            INIT_61 => X"0000001400000000000000060000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000054000000000000000100000000",
            INIT_64 => X"00000000000000000000005e0000000000000000000000000000000000000000",
            INIT_65 => X"00000000000000000000001f000000000000002d000000000000003400000000",
            INIT_66 => X"0000006b00000000000000000000000000000038000000000000000000000000",
            INIT_67 => X"000000000000000000000037000000000000005f000000000000001e00000000",
            INIT_68 => X"0000000000000000000000350000000000000000000000000000001600000000",
            INIT_69 => X"0000004900000000000000400000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000014000000000000003c000000000000003d00000000",
            INIT_6B => X"00000077000000000000001e00000000000000a9000000000000000000000000",
            INIT_6C => X"0000000000000000000000400000000000000050000000000000005900000000",
            INIT_6D => X"0000003000000000000000520000000000000054000000000000006e00000000",
            INIT_6E => X"0000006a000000000000008b0000000000000065000000000000003e00000000",
            INIT_6F => X"0000001b00000000000000230000000000000028000000000000003800000000",
            INIT_70 => X"0000005200000000000000440000000000000028000000000000000000000000",
            INIT_71 => X"0000009400000000000000130000000000000095000000000000000200000000",
            INIT_72 => X"0000000000000000000000a800000000000000b4000000000000004b00000000",
            INIT_73 => X"0000003700000000000000df0000000000000034000000000000009a00000000",
            INIT_74 => X"0000009b000000000000003600000000000000e0000000000000006400000000",
            INIT_75 => X"0000009d00000000000000470000000000000131000000000000005700000000",
            INIT_76 => X"0000001700000000000000560000000000000070000000000000008f00000000",
            INIT_77 => X"00000110000000000000010a000000000000008000000000000000ea00000000",
            INIT_78 => X"000000ca00000000000000dc000000000000009d00000000000000bf00000000",
            INIT_79 => X"000000f300000000000000f3000000000000010e000000000000010f00000000",
            INIT_7A => X"0000009f000000000000009d000000000000010e00000000000000fe00000000",
            INIT_7B => X"00000027000000000000005e000000000000007c000000000000008600000000",
            INIT_7C => X"000000510000000000000084000000000000005a000000000000005500000000",
            INIT_7D => X"0000001800000000000000260000000000000023000000000000001a00000000",
            INIT_7E => X"00000031000000000000007400000000000000a0000000000000001500000000",
            INIT_7F => X"00000021000000000000000c000000000000002c000000000000001d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE0;


    MEM_IFMAP_LAYER2_INSTANCE1 : if BRAM_NAME = "ifmap_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002300000000000000540000000000000002000000000000002e00000000",
            INIT_01 => X"00000051000000000000003c000000000000001d000000000000003e00000000",
            INIT_02 => X"0000005a000000000000002c0000000000000000000000000000004200000000",
            INIT_03 => X"000000aa00000000000000390000000000000045000000000000000400000000",
            INIT_04 => X"0000000e000000000000000b0000000000000027000000000000005700000000",
            INIT_05 => X"00000024000000000000003c000000000000003b000000000000003300000000",
            INIT_06 => X"0000013f0000000000000031000000000000002b000000000000001600000000",
            INIT_07 => X"000000af0000000000000116000000000000013e000000000000015300000000",
            INIT_08 => X"00000130000000000000010700000000000000f500000000000000c200000000",
            INIT_09 => X"00000084000000000000006c000000000000009600000000000000e900000000",
            INIT_0A => X"000000a100000000000000e800000000000000de000000000000009d00000000",
            INIT_0B => X"0000006f000000000000009a000000000000006d000000000000009100000000",
            INIT_0C => X"0000009100000000000000b500000000000000bf00000000000000a800000000",
            INIT_0D => X"0000006f00000000000000a2000000000000006a000000000000009700000000",
            INIT_0E => X"0000006d000000000000007c0000000000000080000000000000007700000000",
            INIT_0F => X"00000059000000000000000100000000000000ac000000000000001800000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000007400000000000000370000000000000004000000000000003600000000",
            INIT_14 => X"00000000000000000000004b0000000000000019000000000000002600000000",
            INIT_15 => X"0000000100000000000000000000000000000000000000000000001b00000000",
            INIT_16 => X"0000004b000000000000002a0000000000000016000000000000000000000000",
            INIT_17 => X"0000000a00000000000000000000000000000000000000000000004d00000000",
            INIT_18 => X"0000001200000000000000000000000000000000000000000000000a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_1A => X"0000000200000000000000120000000000000000000000000000000000000000",
            INIT_1B => X"0000003e000000000000006c000000000000001e000000000000004300000000",
            INIT_1C => X"0000000f00000000000000110000000000000076000000000000000800000000",
            INIT_1D => X"000000240000000000000000000000000000000a000000000000002900000000",
            INIT_1E => X"0000000c00000000000000030000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_21 => X"0000001000000000000000360000000000000001000000000000000000000000",
            INIT_22 => X"00000012000000000000000b0000000000000035000000000000000600000000",
            INIT_23 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_24 => X"000000000000000000000040000000000000002f000000000000000700000000",
            INIT_25 => X"0000000000000000000000000000000000000020000000000000001a00000000",
            INIT_26 => X"0000006200000000000000000000000000000041000000000000004600000000",
            INIT_27 => X"0000003300000000000000100000000000000032000000000000004000000000",
            INIT_28 => X"0000009d00000000000000240000000000000000000000000000006f00000000",
            INIT_29 => X"0000009500000000000000c4000000000000009e000000000000007c00000000",
            INIT_2A => X"000000ba00000000000000ae000000000000007a000000000000005c00000000",
            INIT_2B => X"00000000000000000000000700000000000000ba00000000000000c500000000",
            INIT_2C => X"0000004c000000000000004f0000000000000041000000000000001f00000000",
            INIT_2D => X"00000062000000000000003e0000000000000064000000000000003000000000",
            INIT_2E => X"0000006c000000000000005b0000000000000080000000000000006500000000",
            INIT_2F => X"000000960000000000000087000000000000006f000000000000006c00000000",
            INIT_30 => X"00000076000000000000003f000000000000008700000000000000c600000000",
            INIT_31 => X"000000960000000000000086000000000000009d000000000000008700000000",
            INIT_32 => X"000000b800000000000000840000000000000024000000000000006d00000000",
            INIT_33 => X"00000040000000000000006d000000000000004f000000000000007000000000",
            INIT_34 => X"00000043000000000000009a000000000000007f000000000000004000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_36 => X"0000000000000000000000000000000000000059000000000000003a00000000",
            INIT_37 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000002f000000000000004f00000000",
            INIT_39 => X"00000019000000000000000c0000000000000000000000000000000000000000",
            INIT_3A => X"0000003e00000000000000140000000000000008000000000000000000000000",
            INIT_3B => X"00000046000000000000002f0000000000000082000000000000000000000000",
            INIT_3C => X"00000001000000000000004c0000000000000021000000000000005200000000",
            INIT_3D => X"000000490000000000000044000000000000000e000000000000007e00000000",
            INIT_3E => X"00000096000000000000000f000000000000002e000000000000002b00000000",
            INIT_3F => X"00000041000000000000003a0000000000000040000000000000005500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a400000000000000ac0000000000000000000000000000000300000000",
            INIT_41 => X"000000a00000000000000083000000000000009200000000000000aa00000000",
            INIT_42 => X"000000c300000000000000d900000000000000e000000000000000ad00000000",
            INIT_43 => X"0000010600000000000000eb00000000000000ce00000000000000c200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE1;


    MEM_IFMAP_LAYER3_INSTANCE0 : if BRAM_NAME = "ifmap_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000099000000000000012d00000000000000f9000000000000014400000000",
            INIT_01 => X"000000f4000000000000004f0000000000000042000000000000009900000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000010c00000000",
            INIT_03 => X"0000006400000000000000000000000000000000000000000000001400000000",
            INIT_04 => X"0000001b0000000000000078000000000000009e00000000000000b300000000",
            INIT_05 => X"0000011b00000000000000990000000000000160000000000000005100000000",
            INIT_06 => X"00000174000000000000008a0000000000000144000000000000014300000000",
            INIT_07 => X"000001260000000000000116000000000000012900000000000001c100000000",
            INIT_08 => X"000000000000000000000000000000000000007e000000000000010d00000000",
            INIT_09 => X"000000eb00000000000000f00000000000000144000000000000019500000000",
            INIT_0A => X"0000000000000000000000490000000000000048000000000000009f00000000",
            INIT_0B => X"00000213000000000000018f00000000000000fa000000000000000600000000",
            INIT_0C => X"0000017a000000000000019a0000000000000215000000000000019200000000",
            INIT_0D => X"0000000d00000000000000540000000000000055000000000000003e00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000015c000000000000000c0000000000000000000000000000000000000000",
            INIT_10 => X"000000dc00000000000000fa000000000000009700000000000000b400000000",
            INIT_11 => X"000001090000000000000152000000000000021d000000000000005600000000",
            INIT_12 => X"00000249000000000000015f0000000000000223000000000000012e00000000",
            INIT_13 => X"000001b30000000000000209000000000000015a000000000000020d00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000018700000000",
            INIT_15 => X"000000170000000000000000000000000000004c000000000000000000000000",
            INIT_16 => X"0000018a00000000000001100000000000000069000000000000007700000000",
            INIT_17 => X"000001840000000000000119000000000000016c000000000000020600000000",
            INIT_18 => X"000000390000000000000014000000000000003a00000000000000fd00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000007900000000000000c40000000000000000000000000000000000000000",
            INIT_1B => X"0000003200000000000000000000000000000000000000000000006600000000",
            INIT_1C => X"0000017e000000000000010c0000000000000056000000000000006500000000",
            INIT_1D => X"00000124000000000000014f00000000000000d7000000000000015b00000000",
            INIT_1E => X"0000013900000000000000f90000000000000116000000000000010100000000",
            INIT_1F => X"00000071000000000000000000000000000000dd00000000000000f000000000",
            INIT_20 => X"0000003700000000000000f300000000000000e800000000000000be00000000",
            INIT_21 => X"000000000000000000000032000000000000006f00000000000001bf00000000",
            INIT_22 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000006600000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "gold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000d00000000000000000000000000000000000000000000000a00000000",
            INIT_0A => X"0000000000000000000000140000000000000017000000000000002400000000",
            INIT_0B => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002b00000000000000100000000000000016000000000000001200000000",
            INIT_0E => X"00000000000000000000000b000000000000001b000000000000001c00000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000002300000000",
            INIT_10 => X"0000001d0000000000000025000000000000001a000000000000000000000000",
            INIT_11 => X"0000001a00000000000000130000000000000006000000000000001b00000000",
            INIT_12 => X"000000470000000000000000000000000000000a000000000000000b00000000",
            INIT_13 => X"0000003300000000000000220000000000000008000000000000003000000000",
            INIT_14 => X"000000120000000000000011000000000000002e000000000000003c00000000",
            INIT_15 => X"0000000d00000000000000280000000000000040000000000000000000000000",
            INIT_16 => X"00000047000000000000003f0000000000000007000000000000001100000000",
            INIT_17 => X"0000001e00000000000000090000000000000000000000000000000300000000",
            INIT_18 => X"000000150000000000000016000000000000002c000000000000002d00000000",
            INIT_19 => X"0000000f0000000000000014000000000000001d000000000000003a00000000",
            INIT_1A => X"000000130000000000000033000000000000004b000000000000001400000000",
            INIT_1B => X"00000050000000000000001e0000000000000000000000000000000000000000",
            INIT_1C => X"00000039000000000000001c000000000000001a000000000000003200000000",
            INIT_1D => X"0000000b000000000000001f0000000000000011000000000000002000000000",
            INIT_1E => X"00000018000000000000004b0000000000000042000000000000005400000000",
            INIT_1F => X"000000130000000000000019000000000000002d000000000000001c00000000",
            INIT_20 => X"00000028000000000000000f0000000000000017000000000000000200000000",
            INIT_21 => X"0000004e00000000000000000000000000000003000000000000001200000000",
            INIT_22 => X"0000001b00000000000000210000000000000042000000000000004b00000000",
            INIT_23 => X"00000023000000000000001a0000000000000011000000000000002200000000",
            INIT_24 => X"0000000000000000000000030000000000000024000000000000002000000000",
            INIT_25 => X"0000004300000000000000340000000000000000000000000000000000000000",
            INIT_26 => X"0000001400000000000000440000000000000011000000000000004300000000",
            INIT_27 => X"000000170000000000000038000000000000004d000000000000003a00000000",
            INIT_28 => X"0000001400000000000000210000000000000013000000000000000400000000",
            INIT_29 => X"00000034000000000000004f0000000000000042000000000000001400000000",
            INIT_2A => X"00000042000000000000005a0000000000000083000000000000003c00000000",
            INIT_2B => X"0000003700000000000000300000000000000038000000000000003f00000000",
            INIT_2C => X"0000004500000000000000460000000000000041000000000000003d00000000",
            INIT_2D => X"00000065000000000000003c0000000000000045000000000000005000000000",
            INIT_2E => X"0000003a000000000000003d000000000000003b000000000000005900000000",
            INIT_2F => X"0000003e000000000000003b0000000000000037000000000000003700000000",
            INIT_30 => X"000000520000000000000043000000000000004a000000000000004a00000000",
            INIT_31 => X"00000041000000000000006b0000000000000042000000000000004400000000",
            INIT_32 => X"0000003c0000000000000039000000000000003f000000000000003b00000000",
            INIT_33 => X"0000004e000000000000004d000000000000004b000000000000004000000000",
            INIT_34 => X"0000004c000000000000005a000000000000006a000000000000004600000000",
            INIT_35 => X"0000003f000000000000003d0000000000000034000000000000005400000000",
            INIT_36 => X"00000042000000000000003d000000000000003f000000000000004300000000",
            INIT_37 => X"00000056000000000000003c0000000000000042000000000000004700000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000003000000000000000200000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_43 => X"0000003d00000000000000000000000000000001000000000000000a00000000",
            INIT_44 => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_45 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"00000000000000000000002e0000000000000000000000000000002600000000",
            INIT_48 => X"00000000000000000000000c0000000000000000000000000000003d00000000",
            INIT_49 => X"0000000000000000000000410000000000000000000000000000000000000000",
            INIT_4A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000007d000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4F => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_53 => X"0000002a000000000000002c0000000000000000000000000000000700000000",
            INIT_54 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_58 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_59 => X"00000010000000000000000f0000000000000000000000000000000000000000",
            INIT_5A => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5D => X"0000000d0000000000000000000000000000001c000000000000002000000000",
            INIT_5E => X"0000000000000000000000750000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000019000000000000001100000000",
            INIT_60 => X"000000140000000000000013000000000000000e000000000000000000000000",
            INIT_61 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000046000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000002d000000000000001d0000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000900000000000000000000000000000000000000000000000700000000",
            INIT_69 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000060000000000000005c0000000000000000000000000000000000000000",
            INIT_71 => X"0000005a00000000000000610000000000000061000000000000006000000000",
            INIT_72 => X"0000004d00000000000000680000000000000071000000000000006400000000",
            INIT_73 => X"00000050000000000000004a0000000000000043000000000000003d00000000",
            INIT_74 => X"000000630000000000000069000000000000005e000000000000005400000000",
            INIT_75 => X"0000004d00000000000000500000000000000061000000000000006400000000",
            INIT_76 => X"0000000000000000000000180000000000000039000000000000005500000000",
            INIT_77 => X"0000004d000000000000003b000000000000001d000000000000000200000000",
            INIT_78 => X"0000006b000000000000006a000000000000004a000000000000003c00000000",
            INIT_79 => X"0000001b00000000000000370000000000000054000000000000006900000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"00000000000000000000003a0000000000000006000000000000000000000000",
            INIT_7C => X"0000005700000000000000680000000000000058000000000000000a00000000",
            INIT_7D => X"0000000000000000000000000000000000000005000000000000003500000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000001a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "gold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000038000000000000003b00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000d000000000000004e00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000056000000000000001f0000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000006000000000000000d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000006000000000000001c0000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_0F => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_10 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000c00000000000000000000000000000000000000000000000500000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000004300000000000000260000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000ba00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000bf00000000000000c200000000000000bd00000000000000c100000000",
            INIT_2A => X"000000bb00000000000000c200000000000000c600000000000000bc00000000",
            INIT_2B => X"000000a7000000000000009f00000000000000a500000000000000b500000000",
            INIT_2C => X"000000bd00000000000000b5000000000000009e00000000000000aa00000000",
            INIT_2D => X"000000e300000000000000bf00000000000000c900000000000000c200000000",
            INIT_2E => X"0000008600000000000000ac00000000000000c100000000000000e300000000",
            INIT_2F => X"0000008b000000000000007e000000000000008f00000000000000a100000000",
            INIT_30 => X"000000c0000000000000008800000000000000b600000000000000a300000000",
            INIT_31 => X"000000bf00000000000000ea00000000000000c200000000000000c300000000",
            INIT_32 => X"000000de00000000000000a20000000000000061000000000000007e00000000",
            INIT_33 => X"0000008e000000000000006900000000000000a700000000000000ae00000000",
            INIT_34 => X"000000bf00000000000000c8000000000000006800000000000000c800000000",
            INIT_35 => X"000000a300000000000000d5000000000000009e00000000000000d000000000",
            INIT_36 => X"000000ad00000000000000ef00000000000000a0000000000000009200000000",
            INIT_37 => X"00000103000000000000005e0000000000000062000000000000008e00000000",
            INIT_38 => X"0000014400000000000000b000000000000000f200000000000000ed00000000",
            INIT_39 => X"0000008a00000000000000b50000000000000115000000000000012f00000000",
            INIT_3A => X"0000008c00000000000000ce00000000000000f7000000000000006200000000",
            INIT_3B => X"00000118000000000000011e0000000000000056000000000000007d00000000",
            INIT_3C => X"0000011500000000000000f000000000000000db000000000000010300000000",
            INIT_3D => X"0000007a00000000000000a800000000000000d2000000000000012b00000000",
            INIT_3E => X"00000097000000000000009000000000000000c7000000000000014600000000",
            INIT_3F => X"000000c000000000000001450000000000000113000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000015000000000000000ed00000000000000ac00000000000000c600000000",
            INIT_41 => X"0000012700000000000000be00000000000000cc000000000000010300000000",
            INIT_42 => X"000000a70000000000000096000000000000008c00000000000000ba00000000",
            INIT_43 => X"000000d000000000000000de0000000000000139000000000000013900000000",
            INIT_44 => X"000000de0000000000000146000000000000012400000000000000ac00000000",
            INIT_45 => X"000000c0000000000000010600000000000000cd00000000000000b000000000",
            INIT_46 => X"0000016200000000000000a000000000000000b8000000000000008500000000",
            INIT_47 => X"000000e200000000000000c40000000000000114000000000000014600000000",
            INIT_48 => X"0000009900000000000000bd00000000000000c600000000000000cc00000000",
            INIT_49 => X"00000061000000000000009e00000000000000a800000000000000ec00000000",
            INIT_4A => X"00000149000000000000014900000000000000b7000000000000008400000000",
            INIT_4B => X"000000a800000000000000f500000000000000ca000000000000012a00000000",
            INIT_4C => X"000000b600000000000000d5000000000000011700000000000000b300000000",
            INIT_4D => X"000000b200000000000000610000000000000043000000000000009b00000000",
            INIT_4E => X"0000012e0000000000000146000000000000010900000000000000c800000000",
            INIT_4F => X"0000010f0000000000000109000000000000018d00000000000000d400000000",
            INIT_50 => X"00000058000000000000009100000000000000e9000000000000013700000000",
            INIT_51 => X"000000aa00000000000000ad0000000000000091000000000000006f00000000",
            INIT_52 => X"000001790000000000000128000000000000010e00000000000000cc00000000",
            INIT_53 => X"0000009c00000000000000a300000000000000c700000000000001c800000000",
            INIT_54 => X"00000093000000000000008a0000000000000083000000000000008900000000",
            INIT_55 => X"000000b200000000000000a600000000000000ab000000000000009a00000000",
            INIT_56 => X"000000ff00000000000001c000000000000000e500000000000000b500000000",
            INIT_57 => X"00000087000000000000008c0000000000000097000000000000009500000000",
            INIT_58 => X"000000b400000000000000a1000000000000008f000000000000008500000000",
            INIT_59 => X"0000009500000000000000ae00000000000000b000000000000000aa00000000",
            INIT_5A => X"0000009a00000000000000ac000000000000016a00000000000000bb00000000",
            INIT_5B => X"00000096000000000000008b000000000000008f000000000000009f00000000",
            INIT_5C => X"0000009e000000000000009e00000000000000a300000000000000a200000000",
            INIT_5D => X"000000a3000000000000009500000000000000c100000000000000db00000000",
            INIT_5E => X"0000008f000000000000007c000000000000008b00000000000000ae00000000",
            INIT_5F => X"000000aa00000000000000ad000000000000009d000000000000009200000000",
            INIT_60 => X"000000af00000000000000f300000000000000a7000000000000009000000000",
            INIT_61 => X"0000007b0000000000000078000000000000007e000000000000007600000000",
            INIT_62 => X"0000008500000000000000820000000000000074000000000000007700000000",
            INIT_63 => X"0000006200000000000000620000000000000070000000000000007b00000000",
            INIT_64 => X"000000750000000000000067000000000000006a000000000000006200000000",
            INIT_65 => X"000000770000000000000080000000000000007e000000000000007d00000000",
            INIT_66 => X"0000005f00000000000000790000000000000079000000000000006f00000000",
            INIT_67 => X"0000003f000000000000002e0000000000000026000000000000003400000000",
            INIT_68 => X"00000063000000000000006e0000000000000065000000000000005b00000000",
            INIT_69 => X"00000084000000000000007d0000000000000081000000000000007d00000000",
            INIT_6A => X"00000016000000000000001f0000000000000037000000000000006200000000",
            INIT_6B => X"0000002f00000000000000250000000000000021000000000000003200000000",
            INIT_6C => X"0000007c000000000000001c0000000000000040000000000000005900000000",
            INIT_6D => X"0000004500000000000000420000000000000077000000000000007c00000000",
            INIT_6E => X"0000004100000000000000260000000000000018000000000000002100000000",
            INIT_6F => X"0000003a000000000000001d0000000000000023000000000000003000000000",
            INIT_70 => X"0000005000000000000000740000000000000034000000000000003200000000",
            INIT_71 => X"0000002e000000000000004f0000000000000031000000000000006200000000",
            INIT_72 => X"0000003100000000000000400000000000000000000000000000002100000000",
            INIT_73 => X"000000270000000000000015000000000000001b000000000000001d00000000",
            INIT_74 => X"0000006f000000000000004e0000000000000077000000000000004e00000000",
            INIT_75 => X"000000270000000000000039000000000000005d000000000000005600000000",
            INIT_76 => X"0000002200000000000000360000000000000051000000000000000300000000",
            INIT_77 => X"00000054000000000000001f000000000000000d000000000000001900000000",
            INIT_78 => X"00000040000000000000003d0000000000000075000000000000006900000000",
            INIT_79 => X"0000001300000000000000400000000000000039000000000000007200000000",
            INIT_7A => X"0000001a00000000000000130000000000000029000000000000004f00000000",
            INIT_7B => X"0000002c0000000000000049000000000000002d000000000000002900000000",
            INIT_7C => X"000000500000000000000060000000000000002e000000000000005700000000",
            INIT_7D => X"000000490000000000000031000000000000003c000000000000004300000000",
            INIT_7E => X"00000042000000000000002f000000000000001b000000000000003300000000",
            INIT_7F => X"0000003d000000000000002d0000000000000040000000000000003c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "gold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003200000000000000450000000000000039000000000000003000000000",
            INIT_01 => X"0000003100000000000000550000000000000036000000000000002800000000",
            INIT_02 => X"0000004b000000000000005f000000000000003c000000000000001100000000",
            INIT_03 => X"00000054000000000000000c0000000000000046000000000000003f00000000",
            INIT_04 => X"000000240000000000000042000000000000001c000000000000001500000000",
            INIT_05 => X"00000017000000000000000a0000000000000029000000000000005000000000",
            INIT_06 => X"000000400000000000000039000000000000006c000000000000004e00000000",
            INIT_07 => X"00000024000000000000003e000000000000000e000000000000004600000000",
            INIT_08 => X"000000010000000000000033000000000000004c000000000000002100000000",
            INIT_09 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000003c0000000000000028000000000000000b000000000000001400000000",
            INIT_0B => X"00000000000000000000001b0000000000000073000000000000003b00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000006e000000000000000f0000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000005000000000000000500000000",
            INIT_1B => X"0000000300000000000000050000000000000008000000000000000400000000",
            INIT_1C => X"0000000c00000000000000060000000000000000000000000000000000000000",
            INIT_1D => X"0000000600000000000000000000000000000000000000000000000100000000",
            INIT_1E => X"00000009000000000000001a0000000000000000000000000000000000000000",
            INIT_1F => X"00000008000000000000000b0000000000000000000000000000000a00000000",
            INIT_20 => X"0000001a00000000000000060000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000012000000000000002b000000000000000000000000",
            INIT_23 => X"0000001f00000000000000110000000000000017000000000000000000000000",
            INIT_24 => X"00000000000000000000005a0000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000016000000000000000e00000000",
            INIT_27 => X"0000001600000000000000220000000000000002000000000000003500000000",
            INIT_28 => X"0000001e00000000000000000000000000000048000000000000000000000000",
            INIT_29 => X"0000003400000000000000060000000000000005000000000000000000000000",
            INIT_2A => X"0000000d0000000000000000000000000000001b000000000000003000000000",
            INIT_2B => X"0000000000000000000000270000000000000004000000000000003300000000",
            INIT_2C => X"00000005000000000000002c0000000000000000000000000000003200000000",
            INIT_2D => X"0000002400000000000000320000000000000006000000000000000000000000",
            INIT_2E => X"00000040000000000000003c0000000000000000000000000000004200000000",
            INIT_2F => X"0000003100000000000000140000000000000018000000000000000000000000",
            INIT_30 => X"00000000000000000000003a0000000000000000000000000000001e00000000",
            INIT_31 => X"000000420000000000000027000000000000000c000000000000000000000000",
            INIT_32 => X"00000000000000000000002d0000000000000045000000000000000000000000",
            INIT_33 => X"0000002200000000000000230000000000000019000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_35 => X"000000000000000000000027000000000000000b000000000000005400000000",
            INIT_36 => X"0000000000000000000000000000000000000036000000000000002900000000",
            INIT_37 => X"0000005d0000000000000000000000000000002d000000000000001200000000",
            INIT_38 => X"0000001800000000000000000000000000000016000000000000000000000000",
            INIT_39 => X"0000000000000000000000120000000000000000000000000000001000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_3B => X"0000000000000000000000650000000000000000000000000000000e00000000",
            INIT_3C => X"0000001500000000000000000000000000000006000000000000002800000000",
            INIT_3D => X"000000000000000000000033000000000000000d000000000000000f00000000",
            INIT_3E => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_3F => X"000000560000000000000000000000000000005a000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003e000000000000000e0000000000000000000000000000001300000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003900000000000000610000000000000000000000000000001300000000",
            INIT_44 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000000b000000000000000500000000",
            INIT_47 => X"000000010000000000000000000000000000007f000000000000000c00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000005100000000000000000000000000000000000000000000001600000000",
            INIT_4B => X"00000000000000000000000b0000000000000000000000000000002100000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000002000000000000000080000000000000000000000000000000100000000",
            INIT_4E => X"0000000b00000000000000010000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000002c000000000000001200000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001e00000000000000040000000000000004000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_5C => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_72 => X"0000000000000000000000070000000000000003000000000000003400000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_75 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_7A => X"0000001900000000000000060000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001c0000000000000031000000000000002a000000000000003f00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7E => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000002d0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE2;


    MEM_GOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "gold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_06 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000050000000000000011000000000000000900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000004000000000000000200000000",
            INIT_0B => X"0000000200000000000000000000000000000000000000000000000700000000",
            INIT_0C => X"00000007000000000000000b0000000000000003000000000000000000000000",
            INIT_0D => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_0E => X"0000001f00000000000000070000000000000000000000000000000400000000",
            INIT_0F => X"0000001f00000000000000000000000000000001000000000000000000000000",
            INIT_10 => X"0000000f000000000000000b0000000000000000000000000000000000000000",
            INIT_11 => X"0000000100000000000000260000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_13 => X"00000000000000000000002a000000000000000b000000000000000000000000",
            INIT_14 => X"0000001500000000000000040000000000000000000000000000000000000000",
            INIT_15 => X"0000000a00000000000000000000000000000039000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_18 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000003a0000000000000000000000000000000f00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000100000000000000000000000000000000000000000000004b00000000",
            INIT_1C => X"0000000c00000000000000000000000000000009000000000000000000000000",
            INIT_1D => X"0000000000000000000000490000000000000000000000000000000000000000",
            INIT_1E => X"0000008100000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000002f000000000000003a000000000000000000000000",
            INIT_22 => X"0000000000000000000000600000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000c0000000000000003000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000002b000000000000001b00000000",
            INIT_26 => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_28 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_29 => X"0000001800000000000000000000000000000000000000000000000100000000",
            INIT_2A => X"000000110000000000000000000000000000000b000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2C => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_2E => X"0000001400000000000000220000000000000004000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_30 => X"0000001a00000000000000000000000000000000000000000000007200000000",
            INIT_31 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000d0000000000000010000000000000000d00000000",
            INIT_33 => X"0000003a00000000000000000000000000000021000000000000001f00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000045000000000000001a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000050000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_42 => X"0000004600000000000000440000000000000045000000000000003f00000000",
            INIT_43 => X"0000004b00000000000000470000000000000041000000000000004300000000",
            INIT_44 => X"0000002d000000000000002a0000000000000034000000000000004300000000",
            INIT_45 => X"00000043000000000000003b000000000000003d000000000000003500000000",
            INIT_46 => X"0000004400000000000000480000000000000049000000000000004800000000",
            INIT_47 => X"0000002200000000000000380000000000000041000000000000004500000000",
            INIT_48 => X"00000015000000000000000e000000000000000e000000000000001100000000",
            INIT_49 => X"00000025000000000000002b0000000000000038000000000000002700000000",
            INIT_4A => X"0000003100000000000000470000000000000049000000000000004400000000",
            INIT_4B => X"0000000d000000000000000d000000000000000e000000000000002000000000",
            INIT_4C => X"00000010000000000000000f0000000000000011000000000000001500000000",
            INIT_4D => X"0000003c0000000000000019000000000000001c000000000000002900000000",
            INIT_4E => X"00000023000000000000001e000000000000003a000000000000004300000000",
            INIT_4F => X"00000019000000000000000c000000000000000b000000000000001500000000",
            INIT_50 => X"00000019000000000000000c000000000000000a000000000000001100000000",
            INIT_51 => X"0000002e000000000000003a0000000000000022000000000000001600000000",
            INIT_52 => X"000000150000000000000020000000000000002c000000000000003b00000000",
            INIT_53 => X"0000001a000000000000001d0000000000000004000000000000000a00000000",
            INIT_54 => X"00000009000000000000000e000000000000000f000000000000000f00000000",
            INIT_55 => X"00000011000000000000002a000000000000003c000000000000001600000000",
            INIT_56 => X"00000014000000000000001d0000000000000026000000000000001e00000000",
            INIT_57 => X"0000000d000000000000000f000000000000001b000000000000000b00000000",
            INIT_58 => X"00000011000000000000000e0000000000000010000000000000000c00000000",
            INIT_59 => X"0000001b000000000000001b0000000000000036000000000000002300000000",
            INIT_5A => X"0000000700000000000000180000000000000017000000000000001f00000000",
            INIT_5B => X"0000000b00000000000000080000000000000010000000000000001400000000",
            INIT_5C => X"0000001600000000000000110000000000000011000000000000001900000000",
            INIT_5D => X"00000016000000000000001f000000000000001c000000000000002300000000",
            INIT_5E => X"0000001700000000000000170000000000000018000000000000000d00000000",
            INIT_5F => X"0000002700000000000000140000000000000008000000000000000f00000000",
            INIT_60 => X"0000000f000000000000000c000000000000000a000000000000000f00000000",
            INIT_61 => X"0000001200000000000000150000000000000009000000000000001700000000",
            INIT_62 => X"0000000800000000000000120000000000000014000000000000001100000000",
            INIT_63 => X"0000000f000000000000003a0000000000000020000000000000000800000000",
            INIT_64 => X"0000001700000000000000000000000000000011000000000000000e00000000",
            INIT_65 => X"00000015000000000000001b000000000000000c000000000000000f00000000",
            INIT_66 => X"0000001400000000000000000000000000000004000000000000001200000000",
            INIT_67 => X"0000000c00000000000000000000000000000035000000000000002d00000000",
            INIT_68 => X"000000190000000000000023000000000000000c000000000000000e00000000",
            INIT_69 => X"0000000000000000000000060000000000000000000000000000000500000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "gold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000150000000000000010000000000000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000003000000000000000600000000",
            INIT_27 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_28 => X"0000000400000000000000020000000000000000000000000000000000000000",
            INIT_29 => X"00000009000000000000000a0000000000000006000000000000000400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2B => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_2C => X"0000000600000000000000030000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000030000000000000006000000000000000700000000",
            INIT_2E => X"0000000500000000000000000000000000000003000000000000000300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_30 => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000002000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000004000000000000001c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000003000000000000000a0000000000000004000000000000000000000000",
            INIT_75 => X"000000000000000000000000000000000000000a000000000000000b00000000",
            INIT_76 => X"000000000000000000000000000000000000001a000000000000002500000000",
            INIT_77 => X"0000000a000000000000001e0000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000005f00000000000000000000000000000000000000000000003800000000",
            INIT_7B => X"0000000000000000000000070000000000000001000000000000003600000000",
            INIT_7C => X"0000000a0000000000000016000000000000001e000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000d000000000000001d0000000000000018000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE4;


    MEM_GOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "gold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000e000000000000002200000000",
            INIT_02 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_04 => X"00000010000000000000000c0000000000000000000000000000000900000000",
            INIT_05 => X"0000001200000000000000180000000000000013000000000000000900000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0A => X"0000000600000000000000070000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0D => X"0000000000000000000000020000000000000002000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000035000000000000000200000000",
            INIT_0F => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000005c0000000000000080000000000000002e00000000",
            INIT_12 => X"00000029000000000000000d0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000013000000000000003400000000",
            INIT_14 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"0000000a00000000000000040000000000000005000000000000000a00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000500000000000000010000000000000002000000000000000500000000",
            INIT_1A => X"0000000000000000000000190000000000000013000000000000000c00000000",
            INIT_1B => X"0000000300000000000000070000000000000023000000000000000000000000",
            INIT_1C => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000700000000000000010000000000000006000000000000001100000000",
            INIT_1E => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000030000000000000009000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000a000000000000001b0000000000000014000000000000000000000000",
            INIT_22 => X"0000000e0000000000000023000000000000002c000000000000000600000000",
            INIT_23 => X"0000003400000000000000340000000000000032000000000000003300000000",
            INIT_24 => X"0000003900000000000000350000000000000030000000000000003700000000",
            INIT_25 => X"000000280000000000000025000000000000002c000000000000003600000000",
            INIT_26 => X"00000037000000000000002f000000000000002d000000000000002900000000",
            INIT_27 => X"0000003700000000000000340000000000000038000000000000003400000000",
            INIT_28 => X"00000020000000000000002a0000000000000029000000000000003400000000",
            INIT_29 => X"0000002100000000000000170000000000000013000000000000001f00000000",
            INIT_2A => X"00000035000000000000001e000000000000002d000000000000002b00000000",
            INIT_2B => X"0000003800000000000000390000000000000037000000000000003600000000",
            INIT_2C => X"000000210000000000000013000000000000001a000000000000001600000000",
            INIT_2D => X"00000021000000000000000f000000000000000a000000000000000100000000",
            INIT_2E => X"00000032000000000000003d0000000000000000000000000000002d00000000",
            INIT_2F => X"000000130000000000000028000000000000002b000000000000003a00000000",
            INIT_30 => X"000000000000000000000023000000000000000f000000000000000600000000",
            INIT_31 => X"00000037000000000000000e0000000000000004000000000000000c00000000",
            INIT_32 => X"0000003e00000000000000210000000000000025000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000a000000000000000f00000000",
            INIT_34 => X"00000000000000000000000b000000000000002b000000000000000900000000",
            INIT_35 => X"0000000000000000000000250000000000000009000000000000001100000000",
            INIT_36 => X"00000018000000000000001d0000000000000012000000000000000e00000000",
            INIT_37 => X"0000000300000000000000070000000000000000000000000000000000000000",
            INIT_38 => X"0000001400000000000000000000000000000000000000000000003b00000000",
            INIT_39 => X"000000040000000000000000000000000000000c000000000000000900000000",
            INIT_3A => X"0000001700000000000000340000000000000018000000000000001900000000",
            INIT_3B => X"0000003900000000000000000000000000000000000000000000000400000000",
            INIT_3C => X"0000001100000000000000130000000000000000000000000000000000000000",
            INIT_3D => X"0000000d00000000000000000000000000000000000000000000000700000000",
            INIT_3E => X"000000000000000000000017000000000000002d000000000000001500000000",
            INIT_3F => X"0000000000000000000000310000000000000000000000000000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000000c0000000000000014000000000000000000000000",
            INIT_41 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000f000000000000000a0000000000000013000000000000000300000000",
            INIT_43 => X"00000000000000000000000e0000000000000020000000000000001b00000000",
            INIT_44 => X"0000000000000000000000300000000000000026000000000000001400000000",
            INIT_45 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_46 => X"0000000500000000000000050000000000000019000000000000000800000000",
            INIT_47 => X"00000020000000000000000e0000000000000002000000000000000400000000",
            INIT_48 => X"0000000000000000000000110000000000000029000000000000003300000000",
            INIT_49 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_4A => X"0000000400000000000000000000000000000000000000000000000700000000",
            INIT_4B => X"00000015000000000000000b0000000000000004000000000000000700000000",
            INIT_4C => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"00000000000000000000000b0000000000000008000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000f0000000000000003000000000000000e000000000000000000000000",
            INIT_66 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_69 => X"0000000600000000000000070000000000000008000000000000000700000000",
            INIT_6A => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_6B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_6D => X"0000000000000000000000050000000000000000000000000000000200000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_70 => X"0000000c00000000000000180000000000000000000000000000000c00000000",
            INIT_71 => X"0000000900000000000000000000000000000005000000000000000200000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_73 => X"0000000f00000000000000000000000000000015000000000000000000000000",
            INIT_74 => X"0000000200000000000000050000000000000017000000000000000000000000",
            INIT_75 => X"0000001800000000000000110000000000000000000000000000000000000000",
            INIT_76 => X"0000000400000000000000000000000000000000000000000000000300000000",
            INIT_77 => X"0000000000000000000000000000000000000015000000000000002500000000",
            INIT_78 => X"000000080000000000000004000000000000000c000000000000000e00000000",
            INIT_79 => X"0000002200000000000000230000000000000023000000000000000000000000",
            INIT_7A => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000001000000000000001700000000",
            INIT_7D => X"0000001000000000000000290000000000000021000000000000001900000000",
            INIT_7E => X"0000000200000000000000000000000000000000000000000000001100000000",
            INIT_7F => X"0000000700000000000000200000000000000007000000000000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE5;


    MEM_GOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "gold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000f0000000000000000000000000000002c000000000000001600000000",
            INIT_02 => X"0000002f000000000000003c0000000000000029000000000000000b00000000",
            INIT_03 => X"00000034000000000000001f0000000000000011000000000000001800000000",
            INIT_04 => X"000000320000000000000067000000000000002a000000000000003100000000",
            INIT_05 => X"0000005000000000000000710000000000000010000000000000001100000000",
            INIT_06 => X"0000004500000000000000460000000000000048000000000000004d00000000",
            INIT_07 => X"0000005700000000000000510000000000000053000000000000004f00000000",
            INIT_08 => X"0000000a0000000000000059000000000000006f000000000000005400000000",
            INIT_09 => X"0000004f0000000000000048000000000000004d000000000000004500000000",
            INIT_0A => X"00000052000000000000004a0000000000000049000000000000004900000000",
            INIT_0B => X"0000005400000000000000600000000000000061000000000000005300000000",
            INIT_0C => X"0000006600000000000000440000000000000062000000000000006f00000000",
            INIT_0D => X"0000004b000000000000004b000000000000004a000000000000004100000000",
            INIT_0E => X"0000006700000000000000610000000000000052000000000000004d00000000",
            INIT_0F => X"0000006f000000000000008a000000000000005d000000000000006500000000",
            INIT_10 => X"00000051000000000000005a0000000000000063000000000000006700000000",
            INIT_11 => X"00000048000000000000004b0000000000000056000000000000005300000000",
            INIT_12 => X"000000450000000000000054000000000000005b000000000000004e00000000",
            INIT_13 => X"0000003900000000000000380000000000000071000000000000006d00000000",
            INIT_14 => X"0000003600000000000000340000000000000036000000000000003900000000",
            INIT_15 => X"0000002d0000000000000034000000000000003f000000000000003e00000000",
            INIT_16 => X"00000030000000000000002f0000000000000030000000000000002c00000000",
            INIT_17 => X"0000003b000000000000003b0000000000000036000000000000002c00000000",
            INIT_18 => X"00000029000000000000001c0000000000000036000000000000003900000000",
            INIT_19 => X"00000000000000000000000b000000000000002b000000000000003300000000",
            INIT_1A => X"0000002d0000000000000030000000000000001d000000000000000300000000",
            INIT_1B => X"0000003b000000000000003c0000000000000043000000000000002700000000",
            INIT_1C => X"0000000900000000000000160000000000000028000000000000003c00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1E => X"00000000000000000000002e000000000000001c000000000000000000000000",
            INIT_1F => X"0000002600000000000000370000000000000036000000000000001c00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_22 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000029000000000000002100000000",
            INIT_24 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001f00000000000000000000000000000000000000000000001700000000",
            INIT_27 => X"00000000000000000000000a000000000000001d000000000000002900000000",
            INIT_28 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000019000000000000002a0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000007000000000000001700000000",
            INIT_2C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000f00000000000000090000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_31 => X"000000000000000000000000000000000000000d000000000000000300000000",
            INIT_32 => X"0000000700000000000000020000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_34 => X"0000001200000000000000080000000000000000000000000000001100000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_38 => X"0000001f000000000000001c0000000000000009000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"00000048000000000000004b000000000000004b000000000000004400000000",
            INIT_4D => X"000000470000000000000051000000000000004e000000000000004200000000",
            INIT_4E => X"000000390000000000000033000000000000002e000000000000003700000000",
            INIT_4F => X"000000480000000000000049000000000000003f000000000000004000000000",
            INIT_50 => X"0000001e000000000000004e000000000000004b000000000000004d00000000",
            INIT_51 => X"0000001500000000000000260000000000000034000000000000004c00000000",
            INIT_52 => X"000000350000000000000018000000000000000c000000000000000700000000",
            INIT_53 => X"0000004e0000000000000035000000000000001a000000000000003d00000000",
            INIT_54 => X"000000240000000000000019000000000000004e000000000000004c00000000",
            INIT_55 => X"0000001000000000000000000000000000000023000000000000001800000000",
            INIT_56 => X"0000002a00000000000000220000000000000002000000000000001000000000",
            INIT_57 => X"00000048000000000000004c0000000000000014000000000000000600000000",
            INIT_58 => X"0000001f0000000000000012000000000000002e000000000000002d00000000",
            INIT_59 => X"0000001200000000000000090000000000000019000000000000000800000000",
            INIT_5A => X"0000001f0000000000000020000000000000000f000000000000000a00000000",
            INIT_5B => X"000000110000000000000059000000000000004f000000000000000000000000",
            INIT_5C => X"0000000000000000000000120000000000000010000000000000002c00000000",
            INIT_5D => X"00000006000000000000001a0000000000000015000000000000001f00000000",
            INIT_5E => X"0000000000000000000000330000000000000019000000000000000700000000",
            INIT_5F => X"0000003900000000000000000000000000000033000000000000005600000000",
            INIT_60 => X"0000000e0000000000000000000000000000001a000000000000000400000000",
            INIT_61 => X"0000000b000000000000000c000000000000001a000000000000001400000000",
            INIT_62 => X"0000004100000000000000000000000000000047000000000000001200000000",
            INIT_63 => X"00000003000000000000001b0000000000000000000000000000003100000000",
            INIT_64 => X"0000001700000000000000000000000000000008000000000000001700000000",
            INIT_65 => X"0000001b000000000000000e0000000000000007000000000000001200000000",
            INIT_66 => X"00000020000000000000002f0000000000000000000000000000003100000000",
            INIT_67 => X"00000009000000000000000e000000000000000c000000000000002d00000000",
            INIT_68 => X"0000000e000000000000000f0000000000000002000000000000001c00000000",
            INIT_69 => X"0000001100000000000000350000000000000011000000000000000d00000000",
            INIT_6A => X"0000002c0000000000000001000000000000001c000000000000000000000000",
            INIT_6B => X"0000001e0000000000000000000000000000001b000000000000001100000000",
            INIT_6C => X"0000000a000000000000000a0000000000000019000000000000000000000000",
            INIT_6D => X"000000070000000000000004000000000000003c000000000000002200000000",
            INIT_6E => X"0000002200000000000000250000000000000000000000000000000200000000",
            INIT_6F => X"0000001c000000000000001b0000000000000000000000000000001a00000000",
            INIT_70 => X"0000002300000000000000080000000000000009000000000000000000000000",
            INIT_71 => X"00000000000000000000000d0000000000000000000000000000003900000000",
            INIT_72 => X"00000000000000000000001f0000000000000003000000000000000e00000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000080000000000000000000000000000001c000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE6;


    MEM_GOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "gold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE7;


    MEM_GOLD_LAYER1_INSTANCE0 : if BRAM_NAME = "gold_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000000000000000000000000000000000001400000000",
            INIT_01 => X"000000d200000000000000360000000000000048000000000000002900000000",
            INIT_02 => X"0000007c00000000000000810000000000000045000000000000002f00000000",
            INIT_03 => X"00000064000000000000009a000000000000009a000000000000008200000000",
            INIT_04 => X"000000c5000000000000012000000000000000b6000000000000000300000000",
            INIT_05 => X"000000480000000000000093000000000000006b000000000000003a00000000",
            INIT_06 => X"0000001d00000000000000a800000000000000a800000000000000aa00000000",
            INIT_07 => X"0000002300000000000000860000000000000118000000000000005500000000",
            INIT_08 => X"0000004c000000000000001a0000000000000052000000000000004f00000000",
            INIT_09 => X"00000032000000000000001200000000000000c100000000000000a400000000",
            INIT_0A => X"0000002a000000000000006a0000000000000004000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000004400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000007500000000000000ba00000000000000a8000000000000008700000000",
            INIT_0E => X"0000003300000000000000bf000000000000005200000000000000d100000000",
            INIT_0F => X"0000000000000000000000560000000000000002000000000000000000000000",
            INIT_10 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_11 => X"000000540000000000000030000000000000001a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000003e00000000000000380000000000000000000000000000000000000000",
            INIT_14 => X"000000550000000000000050000000000000001d000000000000000900000000",
            INIT_15 => X"0000003700000000000000000000000000000000000000000000001600000000",
            INIT_16 => X"0000001a00000000000000130000000000000000000000000000001f00000000",
            INIT_17 => X"0000000400000000000000100000000000000019000000000000001c00000000",
            INIT_18 => X"0000000b00000000000000000000000000000000000000000000000100000000",
            INIT_19 => X"00000039000000000000000e0000000000000000000000000000001400000000",
            INIT_1A => X"0000004e0000000000000023000000000000007d000000000000000700000000",
            INIT_1B => X"0000003200000000000000430000000000000021000000000000004200000000",
            INIT_1C => X"00000068000000000000002c000000000000004b000000000000008500000000",
            INIT_1D => X"00000072000000000000004d0000000000000057000000000000005800000000",
            INIT_1E => X"000000440000000000000033000000000000002b000000000000004700000000",
            INIT_1F => X"0000006b00000000000000020000000000000029000000000000002300000000",
            INIT_20 => X"0000004000000000000000400000000000000057000000000000007c00000000",
            INIT_21 => X"00000085000000000000007d0000000000000000000000000000002b00000000",
            INIT_22 => X"0000001e0000000000000034000000000000002a000000000000001700000000",
            INIT_23 => X"0000000900000000000000110000000000000022000000000000001f00000000",
            INIT_24 => X"0000010700000000000000150000000000000000000000000000000800000000",
            INIT_25 => X"0000009d00000000000000e100000000000000d300000000000000fe00000000",
            INIT_26 => X"0000010e00000000000000ab00000000000000d1000000000000008900000000",
            INIT_27 => X"0000001b0000000000000040000000000000004c000000000000008e00000000",
            INIT_28 => X"0000002d000000000000006e000000000000002a000000000000006700000000",
            INIT_29 => X"0000001f00000000000000230000000000000027000000000000000700000000",
            INIT_2A => X"0000001d00000000000000190000000000000087000000000000000000000000",
            INIT_2B => X"000000000000000000000045000000000000001c000000000000001f00000000",
            INIT_2C => X"0000000f00000000000000000000000000000011000000000000000b00000000",
            INIT_2D => X"000000000000000000000000000000000000004e000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000005b000000000000004b0000000000000029000000000000003900000000",
            INIT_32 => X"00000097000000000000004c000000000000004e000000000000007500000000",
            INIT_33 => X"000000b20000000000000049000000000000005b000000000000007f00000000",
            INIT_34 => X"0000007a00000000000000400000000000000056000000000000002a00000000",
            INIT_35 => X"0000004100000000000001270000000000000039000000000000006400000000",
            INIT_36 => X"000000c30000000000000084000000000000002f000000000000003b00000000",
            INIT_37 => X"0000003d000000000000003b00000000000000bc000000000000004000000000",
            INIT_38 => X"00000051000000000000002100000000000000a5000000000000003900000000",
            INIT_39 => X"0000005200000000000000700000000000000025000000000000004700000000",
            INIT_3A => X"000000000000000000000000000000000000000000000000000000be00000000",
            INIT_3B => X"0000006600000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000002a00000000000000090000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_4B => X"0000004300000000000000120000000000000007000000000000000000000000",
            INIT_4C => X"000000000000000000000073000000000000002c000000000000006d00000000",
            INIT_4D => X"000000c800000000000000640000000000000090000000000000007a00000000",
            INIT_4E => X"000000720000000000000024000000000000009e000000000000007700000000",
            INIT_4F => X"00000049000000000000006b0000000000000026000000000000003c00000000",
            INIT_50 => X"000000960000000000000074000000000000001d000000000000005a00000000",
            INIT_51 => X"00000010000000000000005b000000000000006600000000000000a100000000",
            INIT_52 => X"0000007c00000000000000dd0000000000000025000000000000000000000000",
            INIT_53 => X"0000000b000000000000002e0000000000000035000000000000000000000000",
            INIT_54 => X"0000000b00000000000000040000000000000010000000000000000000000000",
            INIT_55 => X"000000380000000000000038000000000000001d000000000000001c00000000",
            INIT_56 => X"000000680000000000000083000000000000002b000000000000000400000000",
            INIT_57 => X"0000006700000000000000710000000000000060000000000000004300000000",
            INIT_58 => X"0000000000000000000000510000000000000000000000000000003500000000",
            INIT_59 => X"0000000000000000000000500000000000000000000000000000004800000000",
            INIT_5A => X"0000000000000000000000000000000000000081000000000000000000000000",
            INIT_5B => X"0000001500000000000000540000000000000045000000000000000000000000",
            INIT_5C => X"0000000d00000000000000000000000000000007000000000000003b00000000",
            INIT_5D => X"000000310000000000000000000000000000001f000000000000007300000000",
            INIT_5E => X"0000002f000000000000005f000000000000003f000000000000004c00000000",
            INIT_5F => X"000000000000000000000000000000000000002a000000000000000200000000",
            INIT_60 => X"0000001500000000000000620000000000000029000000000000000000000000",
            INIT_61 => X"0000001400000000000000060000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000054000000000000000100000000",
            INIT_64 => X"00000000000000000000005e0000000000000000000000000000000000000000",
            INIT_65 => X"00000000000000000000001f000000000000002d000000000000003400000000",
            INIT_66 => X"0000006b00000000000000000000000000000038000000000000000000000000",
            INIT_67 => X"000000000000000000000037000000000000005f000000000000001e00000000",
            INIT_68 => X"0000000000000000000000350000000000000000000000000000001600000000",
            INIT_69 => X"0000004900000000000000400000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000014000000000000003c000000000000003d00000000",
            INIT_6B => X"00000077000000000000001e00000000000000a9000000000000000000000000",
            INIT_6C => X"0000000000000000000000400000000000000050000000000000005900000000",
            INIT_6D => X"0000003000000000000000520000000000000054000000000000006e00000000",
            INIT_6E => X"0000006a000000000000008b0000000000000065000000000000003e00000000",
            INIT_6F => X"0000001b00000000000000230000000000000028000000000000003800000000",
            INIT_70 => X"0000005200000000000000440000000000000028000000000000000000000000",
            INIT_71 => X"0000009400000000000000130000000000000095000000000000000200000000",
            INIT_72 => X"0000000000000000000000a800000000000000b4000000000000004b00000000",
            INIT_73 => X"0000003700000000000000df0000000000000034000000000000009a00000000",
            INIT_74 => X"0000009b000000000000003600000000000000e0000000000000006400000000",
            INIT_75 => X"0000009d00000000000000470000000000000131000000000000005700000000",
            INIT_76 => X"0000001700000000000000560000000000000070000000000000008f00000000",
            INIT_77 => X"00000110000000000000010a000000000000008000000000000000ea00000000",
            INIT_78 => X"000000ca00000000000000dc000000000000009d00000000000000bf00000000",
            INIT_79 => X"000000f300000000000000f3000000000000010e000000000000010f00000000",
            INIT_7A => X"0000009f000000000000009d000000000000010e00000000000000fe00000000",
            INIT_7B => X"00000027000000000000005e000000000000007c000000000000008600000000",
            INIT_7C => X"000000510000000000000084000000000000005a000000000000005500000000",
            INIT_7D => X"0000001800000000000000260000000000000023000000000000001a00000000",
            INIT_7E => X"00000031000000000000007400000000000000a0000000000000001500000000",
            INIT_7F => X"00000021000000000000000c000000000000002c000000000000001d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE0;


    MEM_GOLD_LAYER1_INSTANCE1 : if BRAM_NAME = "gold_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002300000000000000540000000000000002000000000000002e00000000",
            INIT_01 => X"00000051000000000000003c000000000000001d000000000000003e00000000",
            INIT_02 => X"0000005a000000000000002c0000000000000000000000000000004200000000",
            INIT_03 => X"000000aa00000000000000390000000000000045000000000000000400000000",
            INIT_04 => X"0000000e000000000000000b0000000000000027000000000000005700000000",
            INIT_05 => X"00000024000000000000003c000000000000003b000000000000003300000000",
            INIT_06 => X"0000013f0000000000000031000000000000002b000000000000001600000000",
            INIT_07 => X"000000af0000000000000116000000000000013e000000000000015300000000",
            INIT_08 => X"00000130000000000000010700000000000000f500000000000000c200000000",
            INIT_09 => X"00000084000000000000006c000000000000009600000000000000e900000000",
            INIT_0A => X"000000a100000000000000e800000000000000de000000000000009d00000000",
            INIT_0B => X"0000006f000000000000009a000000000000006d000000000000009100000000",
            INIT_0C => X"0000009100000000000000b500000000000000bf00000000000000a800000000",
            INIT_0D => X"0000006f00000000000000a2000000000000006a000000000000009700000000",
            INIT_0E => X"0000006d000000000000007c0000000000000080000000000000007700000000",
            INIT_0F => X"00000059000000000000000100000000000000ac000000000000001800000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000007400000000000000370000000000000004000000000000003600000000",
            INIT_14 => X"00000000000000000000004b0000000000000019000000000000002600000000",
            INIT_15 => X"0000000100000000000000000000000000000000000000000000001b00000000",
            INIT_16 => X"0000004b000000000000002a0000000000000016000000000000000000000000",
            INIT_17 => X"0000000a00000000000000000000000000000000000000000000004d00000000",
            INIT_18 => X"0000001200000000000000000000000000000000000000000000000a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_1A => X"0000000200000000000000120000000000000000000000000000000000000000",
            INIT_1B => X"0000003e000000000000006c000000000000001e000000000000004300000000",
            INIT_1C => X"0000000f00000000000000110000000000000076000000000000000800000000",
            INIT_1D => X"000000240000000000000000000000000000000a000000000000002900000000",
            INIT_1E => X"0000000c00000000000000030000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_21 => X"0000001000000000000000360000000000000001000000000000000000000000",
            INIT_22 => X"00000012000000000000000b0000000000000035000000000000000600000000",
            INIT_23 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_24 => X"000000000000000000000040000000000000002f000000000000000700000000",
            INIT_25 => X"0000000000000000000000000000000000000020000000000000001a00000000",
            INIT_26 => X"0000006200000000000000000000000000000041000000000000004600000000",
            INIT_27 => X"0000003300000000000000100000000000000032000000000000004000000000",
            INIT_28 => X"0000009d00000000000000240000000000000000000000000000006f00000000",
            INIT_29 => X"0000009500000000000000c4000000000000009e000000000000007c00000000",
            INIT_2A => X"000000ba00000000000000ae000000000000007a000000000000005c00000000",
            INIT_2B => X"00000000000000000000000700000000000000ba00000000000000c500000000",
            INIT_2C => X"0000004c000000000000004f0000000000000041000000000000001f00000000",
            INIT_2D => X"00000062000000000000003e0000000000000064000000000000003000000000",
            INIT_2E => X"0000006c000000000000005b0000000000000080000000000000006500000000",
            INIT_2F => X"000000960000000000000087000000000000006f000000000000006c00000000",
            INIT_30 => X"00000076000000000000003f000000000000008700000000000000c600000000",
            INIT_31 => X"000000960000000000000086000000000000009d000000000000008700000000",
            INIT_32 => X"000000b800000000000000840000000000000024000000000000006d00000000",
            INIT_33 => X"00000040000000000000006d000000000000004f000000000000007000000000",
            INIT_34 => X"00000043000000000000009a000000000000007f000000000000004000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_36 => X"0000000000000000000000000000000000000059000000000000003a00000000",
            INIT_37 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000002f000000000000004f00000000",
            INIT_39 => X"00000019000000000000000c0000000000000000000000000000000000000000",
            INIT_3A => X"0000003e00000000000000140000000000000008000000000000000000000000",
            INIT_3B => X"00000046000000000000002f0000000000000082000000000000000000000000",
            INIT_3C => X"00000001000000000000004c0000000000000021000000000000005200000000",
            INIT_3D => X"000000490000000000000044000000000000000e000000000000007e00000000",
            INIT_3E => X"00000096000000000000000f000000000000002e000000000000002b00000000",
            INIT_3F => X"00000041000000000000003a0000000000000040000000000000005500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a400000000000000ac0000000000000000000000000000000300000000",
            INIT_41 => X"000000a00000000000000083000000000000009200000000000000aa00000000",
            INIT_42 => X"000000c300000000000000d900000000000000e000000000000000ad00000000",
            INIT_43 => X"0000010600000000000000eb00000000000000ce00000000000000c200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE1;


    MEM_GOLD_LAYER2_INSTANCE0 : if BRAM_NAME = "gold_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000099000000000000012d00000000000000f9000000000000014400000000",
            INIT_01 => X"000000f4000000000000004f0000000000000042000000000000009900000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000010c00000000",
            INIT_03 => X"0000006400000000000000000000000000000000000000000000001400000000",
            INIT_04 => X"0000001b0000000000000078000000000000009e00000000000000b300000000",
            INIT_05 => X"0000011b00000000000000990000000000000160000000000000005100000000",
            INIT_06 => X"00000174000000000000008a0000000000000144000000000000014300000000",
            INIT_07 => X"000001260000000000000116000000000000012900000000000001c100000000",
            INIT_08 => X"000000000000000000000000000000000000007e000000000000010d00000000",
            INIT_09 => X"000000eb00000000000000f00000000000000144000000000000019500000000",
            INIT_0A => X"0000000000000000000000490000000000000048000000000000009f00000000",
            INIT_0B => X"00000213000000000000018f00000000000000fa000000000000000600000000",
            INIT_0C => X"0000017a000000000000019a0000000000000215000000000000019200000000",
            INIT_0D => X"0000000d00000000000000540000000000000055000000000000003e00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000015c000000000000000c0000000000000000000000000000000000000000",
            INIT_10 => X"000000dc00000000000000fa000000000000009700000000000000b400000000",
            INIT_11 => X"000001090000000000000152000000000000021d000000000000005600000000",
            INIT_12 => X"00000249000000000000015f0000000000000223000000000000012e00000000",
            INIT_13 => X"000001b30000000000000209000000000000015a000000000000020d00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000018700000000",
            INIT_15 => X"000000170000000000000000000000000000004c000000000000000000000000",
            INIT_16 => X"0000018a00000000000001100000000000000069000000000000007700000000",
            INIT_17 => X"000001840000000000000119000000000000016c000000000000020600000000",
            INIT_18 => X"000000390000000000000014000000000000003a00000000000000fd00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000007900000000000000c40000000000000000000000000000000000000000",
            INIT_1B => X"0000003200000000000000000000000000000000000000000000006600000000",
            INIT_1C => X"0000017e000000000000010c0000000000000056000000000000006500000000",
            INIT_1D => X"00000124000000000000014f00000000000000d7000000000000015b00000000",
            INIT_1E => X"0000013900000000000000f90000000000000116000000000000010100000000",
            INIT_1F => X"00000071000000000000000000000000000000dd00000000000000f000000000",
            INIT_20 => X"0000003700000000000000f300000000000000e800000000000000be00000000",
            INIT_21 => X"000000000000000000000032000000000000006f00000000000001bf00000000",
            INIT_22 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000006600000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE0;


    MEM_GOLD_LAYER3_INSTANCE0 : if BRAM_NAME = "gold_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000065de00000000fffe52cfffffffff0000241000000000ffff1dd9ffffffff",
            INIT_01 => X"fffea670fffffffffffa9f82ffffffffffffbb99fffffffffffedfd3ffffffff",
            INIT_02 => X"fffd3903ffffffffffff4486ffffffff",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER3_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "sampleifmap_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "sampleifmap_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "sampleifmap_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "sampleifmap_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "sampleifmap_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "sampleifmap_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "sampleifmap_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e600000000000000e700000000000000e800000000000000e900000000",
            INIT_05 => X"000000e900000000000000e800000000000000e800000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e800000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ec00000000000000ec00000000000000ed00000000",
            INIT_0D => X"000000ec00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ea00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_15 => X"000000ea00000000000000e700000000000000e700000000000000e300000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000df00000000000000e400000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000cf00000000000000d100000000000000ba00000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000ec00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000cb00000000000000db00000000000000e900000000000000ec00000000",
            INIT_25 => X"000000e600000000000000d600000000000000c300000000000000a300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_28 => X"000000ec00000000000000ec00000000000000ec00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_2A => X"000000ed00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e500000000000000eb00000000000000e800000000000000ea00000000",
            INIT_2C => X"000000ae00000000000000b900000000000000c200000000000000d000000000",
            INIT_2D => X"000000e200000000000000cf00000000000000b800000000000000a500000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e700000000000000e800000000000000e400000000000000e400000000",
            INIT_31 => X"000000ec00000000000000ed00000000000000ed00000000000000ea00000000",
            INIT_32 => X"000000ef00000000000000ef00000000000000ed00000000000000ed00000000",
            INIT_33 => X"000000dd00000000000000e900000000000000e000000000000000e100000000",
            INIT_34 => X"0000009a000000000000009f00000000000000a100000000000000b700000000",
            INIT_35 => X"000000c6000000000000009c000000000000008f000000000000009000000000",
            INIT_36 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_37 => X"000000ef00000000000000ed00000000000000ec00000000000000eb00000000",
            INIT_38 => X"000000e300000000000000e600000000000000e000000000000000d400000000",
            INIT_39 => X"000000ee00000000000000ed00000000000000ea00000000000000e500000000",
            INIT_3A => X"000000f000000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_3B => X"000000d600000000000000e900000000000000db00000000000000c900000000",
            INIT_3C => X"000000ad00000000000000b800000000000000b900000000000000c100000000",
            INIT_3D => X"000000ba00000000000000a2000000000000009f00000000000000a500000000",
            INIT_3E => X"000000e900000000000000e900000000000000ea00000000000000e500000000",
            INIT_3F => X"000000ee00000000000000ed00000000000000ec00000000000000ea00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e100000000000000e100000000000000dd00000000000000d800000000",
            INIT_41 => X"000000ee00000000000000ec00000000000000e700000000000000e300000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_43 => X"000000e600000000000000e900000000000000dc00000000000000c500000000",
            INIT_44 => X"000000d000000000000000db00000000000000d100000000000000d100000000",
            INIT_45 => X"000000da00000000000000d900000000000000d200000000000000d100000000",
            INIT_46 => X"000000e600000000000000e400000000000000e400000000000000e100000000",
            INIT_47 => X"000000ee00000000000000ed00000000000000eb00000000000000e600000000",
            INIT_48 => X"00000088000000000000007c0000000000000077000000000000007600000000",
            INIT_49 => X"000000ed00000000000000eb00000000000000e100000000000000ac00000000",
            INIT_4A => X"000000e900000000000000eb00000000000000eb00000000000000ec00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000e100000000000000e700000000000000e300000000000000e400000000",
            INIT_4D => X"000000b900000000000000c900000000000000d900000000000000e100000000",
            INIT_4E => X"000000ba00000000000000a700000000000000a700000000000000ac00000000",
            INIT_4F => X"000000ee00000000000000ec00000000000000eb00000000000000df00000000",
            INIT_50 => X"0000006f000000000000006c0000000000000067000000000000006d00000000",
            INIT_51 => X"000000e500000000000000e300000000000000de000000000000009200000000",
            INIT_52 => X"000000e600000000000000e700000000000000ea00000000000000ec00000000",
            INIT_53 => X"000000e600000000000000e800000000000000e700000000000000e500000000",
            INIT_54 => X"000000df00000000000000e500000000000000e700000000000000e700000000",
            INIT_55 => X"00000089000000000000009200000000000000a400000000000000bf00000000",
            INIT_56 => X"0000009500000000000000790000000000000080000000000000008600000000",
            INIT_57 => X"000000ed00000000000000eb00000000000000ea00000000000000d800000000",
            INIT_58 => X"000000c800000000000000c700000000000000bc00000000000000c300000000",
            INIT_59 => X"000000d300000000000000d500000000000000df00000000000000d100000000",
            INIT_5A => X"000000d200000000000000db00000000000000dc00000000000000d800000000",
            INIT_5B => X"000000dc00000000000000d800000000000000d300000000000000d100000000",
            INIT_5C => X"000000da00000000000000e100000000000000e200000000000000e100000000",
            INIT_5D => X"000000b200000000000000b500000000000000af00000000000000b700000000",
            INIT_5E => X"000000b9000000000000008e00000000000000aa00000000000000ba00000000",
            INIT_5F => X"000000ec00000000000000ea00000000000000e700000000000000db00000000",
            INIT_60 => X"000000d600000000000000ca00000000000000bf00000000000000c100000000",
            INIT_61 => X"000000ab00000000000000cb00000000000000d600000000000000df00000000",
            INIT_62 => X"0000006200000000000000ae00000000000000cf00000000000000b100000000",
            INIT_63 => X"0000007a000000000000006f0000000000000065000000000000005d00000000",
            INIT_64 => X"000000df00000000000000ca0000000000000099000000000000008900000000",
            INIT_65 => X"000000d900000000000000df00000000000000dc00000000000000da00000000",
            INIT_66 => X"000000de00000000000000c400000000000000d400000000000000dd00000000",
            INIT_67 => X"000000eb00000000000000e800000000000000dd00000000000000db00000000",
            INIT_68 => X"0000007d0000000000000071000000000000006f000000000000007100000000",
            INIT_69 => X"000000be00000000000000bf00000000000000aa000000000000008a00000000",
            INIT_6A => X"00000036000000000000009e00000000000000d800000000000000d000000000",
            INIT_6B => X"0000004200000000000000350000000000000031000000000000002d00000000",
            INIT_6C => X"000000ea00000000000000dd000000000000009f000000000000006600000000",
            INIT_6D => X"000000cf00000000000000df00000000000000e300000000000000e900000000",
            INIT_6E => X"000000c700000000000000d400000000000000d300000000000000ca00000000",
            INIT_6F => X"000000dd00000000000000d300000000000000bc00000000000000b300000000",
            INIT_70 => X"00000044000000000000003f0000000000000045000000000000003d00000000",
            INIT_71 => X"000000c30000000000000097000000000000008b000000000000007b00000000",
            INIT_72 => X"0000006700000000000000a300000000000000ce00000000000000d600000000",
            INIT_73 => X"000000b5000000000000008a0000000000000065000000000000005f00000000",
            INIT_74 => X"000000cd00000000000000db00000000000000dd00000000000000cf00000000",
            INIT_75 => X"000000830000000000000093000000000000009e00000000000000b700000000",
            INIT_76 => X"0000008500000000000000880000000000000082000000000000007d00000000",
            INIT_77 => X"000000c500000000000000b6000000000000008a000000000000008000000000",
            INIT_78 => X"0000007f0000000000000055000000000000003a000000000000002800000000",
            INIT_79 => X"000000a300000000000000770000000000000060000000000000008400000000",
            INIT_7A => X"000000b500000000000000b600000000000000b800000000000000ad00000000",
            INIT_7B => X"000000c800000000000000da00000000000000c600000000000000b700000000",
            INIT_7C => X"000000840000000000000091000000000000009f00000000000000ae00000000",
            INIT_7D => X"00000063000000000000005e0000000000000062000000000000007400000000",
            INIT_7E => X"0000008a000000000000007a000000000000006b000000000000006900000000",
            INIT_7F => X"000000b900000000000000bc000000000000009d000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "sampleifmap_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ce0000000000000086000000000000001a000000000000000d00000000",
            INIT_01 => X"000000ac000000000000008d0000000000000076000000000000008a00000000",
            INIT_02 => X"000000e400000000000000dc00000000000000cf00000000000000b500000000",
            INIT_03 => X"000000b000000000000000e200000000000000e600000000000000e000000000",
            INIT_04 => X"00000091000000000000008e000000000000008a000000000000009000000000",
            INIT_05 => X"0000009a00000000000000950000000000000095000000000000009a00000000",
            INIT_06 => X"000000bb00000000000000ad00000000000000a0000000000000009d00000000",
            INIT_07 => X"0000009d00000000000000a500000000000000b200000000000000be00000000",
            INIT_08 => X"000000e100000000000000c8000000000000003a000000000000000500000000",
            INIT_09 => X"000000e200000000000000d400000000000000c700000000000000c500000000",
            INIT_0A => X"000000e600000000000000e800000000000000e900000000000000e500000000",
            INIT_0B => X"000000d200000000000000dd00000000000000df00000000000000d100000000",
            INIT_0C => X"000000bc00000000000000c100000000000000b400000000000000c600000000",
            INIT_0D => X"000000b800000000000000c000000000000000c200000000000000bd00000000",
            INIT_0E => X"0000009000000000000000a100000000000000ab00000000000000ac00000000",
            INIT_0F => X"0000008a00000000000000800000000000000083000000000000008800000000",
            INIT_10 => X"000000ba00000000000000be0000000000000091000000000000002700000000",
            INIT_11 => X"000000c200000000000000c200000000000000c000000000000000b800000000",
            INIT_12 => X"000000be00000000000000c000000000000000bf00000000000000c200000000",
            INIT_13 => X"00000093000000000000009a00000000000000b400000000000000b100000000",
            INIT_14 => X"000000710000000000000092000000000000009c000000000000009100000000",
            INIT_15 => X"0000006f000000000000007e0000000000000084000000000000007200000000",
            INIT_16 => X"0000005e000000000000005d000000000000005b000000000000005c00000000",
            INIT_17 => X"0000008100000000000000810000000000000079000000000000006900000000",
            INIT_18 => X"00000089000000000000008f00000000000000a2000000000000007a00000000",
            INIT_19 => X"00000082000000000000007f0000000000000080000000000000008300000000",
            INIT_1A => X"00000081000000000000007f0000000000000080000000000000008300000000",
            INIT_1B => X"000000640000000000000068000000000000007c000000000000008100000000",
            INIT_1C => X"0000005e00000000000000700000000000000076000000000000006600000000",
            INIT_1D => X"000000530000000000000057000000000000005e000000000000005e00000000",
            INIT_1E => X"00000065000000000000005d0000000000000053000000000000005000000000",
            INIT_1F => X"0000008200000000000000790000000000000073000000000000006c00000000",
            INIT_20 => X"00000050000000000000004d000000000000004c000000000000004900000000",
            INIT_21 => X"0000005a00000000000000570000000000000057000000000000005400000000",
            INIT_22 => X"00000071000000000000006b0000000000000066000000000000005e00000000",
            INIT_23 => X"0000007800000000000000760000000000000076000000000000007300000000",
            INIT_24 => X"00000064000000000000006a000000000000006e000000000000007300000000",
            INIT_25 => X"00000050000000000000004f0000000000000055000000000000005f00000000",
            INIT_26 => X"000000520000000000000050000000000000004d000000000000005000000000",
            INIT_27 => X"00000088000000000000007d0000000000000071000000000000005c00000000",
            INIT_28 => X"0000001200000000000000090000000000000003000000000000000d00000000",
            INIT_29 => X"0000001600000000000000140000000000000015000000000000001200000000",
            INIT_2A => X"00000030000000000000002a0000000000000022000000000000001a00000000",
            INIT_2B => X"000000460000000000000042000000000000003c000000000000003400000000",
            INIT_2C => X"0000003c00000000000000430000000000000048000000000000004700000000",
            INIT_2D => X"0000003900000000000000350000000000000035000000000000003700000000",
            INIT_2E => X"0000005700000000000000480000000000000039000000000000003900000000",
            INIT_2F => X"0000008900000000000000820000000000000078000000000000006800000000",
            INIT_30 => X"000000200000000000000008000000000000000b000000000000002400000000",
            INIT_31 => X"0000000300000000000000080000000000000016000000000000002400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_33 => X"0000000300000000000000010000000000000005000000000000000600000000",
            INIT_34 => X"0000001500000000000000150000000000000018000000000000000d00000000",
            INIT_35 => X"00000027000000000000001e0000000000000016000000000000001500000000",
            INIT_36 => X"0000007b00000000000000710000000000000055000000000000003900000000",
            INIT_37 => X"000000990000000000000086000000000000007a000000000000007400000000",
            INIT_38 => X"0000001b000000000000000d000000000000001a000000000000002300000000",
            INIT_39 => X"0000001b00000000000000310000000000000046000000000000004700000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000000a000000000000001f0000000000000039000000000000001100000000",
            INIT_3C => X"0000000e00000000000000070000000000000004000000000000000400000000",
            INIT_3D => X"00000056000000000000003e0000000000000029000000000000001900000000",
            INIT_3E => X"0000007200000000000000840000000000000090000000000000007a00000000",
            INIT_3F => X"000000ac00000000000000920000000000000084000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000030000000000000004000000000000000d000000000000001000000000",
            INIT_41 => X"0000002400000000000000360000000000000041000000000000002d00000000",
            INIT_42 => X"0000000000000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"0000008300000000000000a10000000000000076000000000000000700000000",
            INIT_44 => X"0000006d00000000000000690000000000000069000000000000007000000000",
            INIT_45 => X"00000097000000000000009a000000000000008a000000000000007600000000",
            INIT_46 => X"00000078000000000000006a0000000000000069000000000000007f00000000",
            INIT_47 => X"000000b800000000000000a4000000000000008e000000000000008100000000",
            INIT_48 => X"000000000000000000000000000000000000000c000000000000002800000000",
            INIT_49 => X"000000150000000000000020000000000000001e000000000000000c00000000",
            INIT_4A => X"0000000300000000000000020000000000000002000000000000000700000000",
            INIT_4B => X"000000cd00000000000000b60000000000000044000000000000000000000000",
            INIT_4C => X"000000bb00000000000000c300000000000000c200000000000000c400000000",
            INIT_4D => X"00000067000000000000007b000000000000009600000000000000ac00000000",
            INIT_4E => X"00000081000000000000007a0000000000000068000000000000005f00000000",
            INIT_4F => X"000000b900000000000000ab0000000000000098000000000000008400000000",
            INIT_50 => X"000000010000000000000001000000000000001a000000000000004500000000",
            INIT_51 => X"0000000c0000000000000012000000000000000c000000000000000400000000",
            INIT_52 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_53 => X"000000cb00000000000000990000000000000020000000000000000100000000",
            INIT_54 => X"0000009b00000000000000b300000000000000bf00000000000000c300000000",
            INIT_55 => X"0000005e0000000000000051000000000000005b000000000000007700000000",
            INIT_56 => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_57 => X"000000b800000000000000ad00000000000000a2000000000000009000000000",
            INIT_58 => X"000000020000000000000001000000000000002f000000000000005300000000",
            INIT_59 => X"0000000400000000000000070000000000000005000000000000000200000000",
            INIT_5A => X"0000000300000000000000010000000000000001000000000000000100000000",
            INIT_5B => X"000000cd000000000000008e000000000000001b000000000000000100000000",
            INIT_5C => X"00000055000000000000007900000000000000a900000000000000c600000000",
            INIT_5D => X"0000007900000000000000660000000000000055000000000000004a00000000",
            INIT_5E => X"000000840000000000000079000000000000007a000000000000008000000000",
            INIT_5F => X"000000ba00000000000000b000000000000000a5000000000000009300000000",
            INIT_60 => X"0000000300000000000000060000000000000036000000000000005c00000000",
            INIT_61 => X"0000000100000000000000010000000000000001000000000000000200000000",
            INIT_62 => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_63 => X"0000009d0000000000000066000000000000000f000000000000000000000000",
            INIT_64 => X"0000004a0000000000000038000000000000004a000000000000007500000000",
            INIT_65 => X"0000007c000000000000007a0000000000000073000000000000006300000000",
            INIT_66 => X"000000880000000000000080000000000000007d000000000000007b00000000",
            INIT_67 => X"000000bc00000000000000b100000000000000a2000000000000009400000000",
            INIT_68 => X"0000000b0000000000000013000000000000002b000000000000005700000000",
            INIT_69 => X"0000000200000000000000020000000000000005000000000000000800000000",
            INIT_6A => X"0000000200000000000000030000000000000003000000000000000300000000",
            INIT_6B => X"00000047000000000000002a0000000000000004000000000000000000000000",
            INIT_6C => X"0000007100000000000000500000000000000039000000000000003500000000",
            INIT_6D => X"00000074000000000000007b0000000000000086000000000000008400000000",
            INIT_6E => X"0000008f000000000000008b0000000000000083000000000000007800000000",
            INIT_6F => X"000000bc00000000000000b600000000000000a9000000000000009c00000000",
            INIT_70 => X"0000001f0000000000000024000000000000002e000000000000005200000000",
            INIT_71 => X"0000001000000000000000110000000000000016000000000000001b00000000",
            INIT_72 => X"0000001300000000000000140000000000000013000000000000001200000000",
            INIT_73 => X"0000004000000000000000250000000000000017000000000000001300000000",
            INIT_74 => X"0000008000000000000000740000000000000068000000000000005700000000",
            INIT_75 => X"0000007300000000000000750000000000000083000000000000008b00000000",
            INIT_76 => X"00000094000000000000008b0000000000000083000000000000007b00000000",
            INIT_77 => X"000000bb00000000000000b900000000000000ae000000000000009f00000000",
            INIT_78 => X"00000037000000000000003a000000000000003e000000000000005500000000",
            INIT_79 => X"00000030000000000000002e000000000000002f000000000000003300000000",
            INIT_7A => X"0000003700000000000000350000000000000033000000000000003100000000",
            INIT_7B => X"0000006800000000000000510000000000000044000000000000003b00000000",
            INIT_7C => X"0000007f0000000000000085000000000000007f000000000000007400000000",
            INIT_7D => X"0000007a00000000000000720000000000000076000000000000007f00000000",
            INIT_7E => X"00000095000000000000008d0000000000000088000000000000008100000000",
            INIT_7F => X"000000ba00000000000000b400000000000000a8000000000000009e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "sampleifmap_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e900000000000000e900000000000000e700000000000000e700000000",
            INIT_05 => X"000000e900000000000000e800000000000000e700000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e900000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000ea00000000000000ea00000000",
            INIT_0D => X"000000ec00000000000000ec00000000000000ea00000000000000eb00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000eb00000000000000eb00000000000000ea00000000000000e900000000",
            INIT_15 => X"000000ea00000000000000e900000000000000eb00000000000000e600000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e200000000000000e600000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000d200000000000000d800000000000000c000000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000d200000000000000e100000000000000ed00000000000000ee00000000",
            INIT_25 => X"000000e500000000000000da00000000000000cd00000000000000ac00000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e700000000000000ed00000000000000e900000000000000eb00000000",
            INIT_2C => X"000000bc00000000000000c600000000000000cd00000000000000d800000000",
            INIT_2D => X"000000e400000000000000d700000000000000c400000000000000b300000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e400000000000000e600000000000000e300000000000000e500000000",
            INIT_31 => X"000000ed00000000000000ed00000000000000ec00000000000000e800000000",
            INIT_32 => X"000000ed00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_33 => X"000000e200000000000000ed00000000000000e400000000000000e500000000",
            INIT_34 => X"000000b000000000000000b400000000000000b400000000000000c500000000",
            INIT_35 => X"000000ce00000000000000a9000000000000009f00000000000000a300000000",
            INIT_36 => X"000000eb00000000000000ec00000000000000ed00000000000000ee00000000",
            INIT_37 => X"000000ed00000000000000ed00000000000000ee00000000000000ec00000000",
            INIT_38 => X"000000e800000000000000ea00000000000000e600000000000000dc00000000",
            INIT_39 => X"000000ed00000000000000ee00000000000000ed00000000000000ea00000000",
            INIT_3A => X"000000ee00000000000000ec00000000000000ed00000000000000ed00000000",
            INIT_3B => X"000000da00000000000000ec00000000000000de00000000000000cc00000000",
            INIT_3C => X"000000bf00000000000000c900000000000000c900000000000000cc00000000",
            INIT_3D => X"000000c700000000000000b000000000000000ae00000000000000b600000000",
            INIT_3E => X"000000ee00000000000000ee00000000000000ef00000000000000ef00000000",
            INIT_3F => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ef00000000000000ee00000000000000ec00000000000000ea00000000",
            INIT_41 => X"000000ec00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_43 => X"000000e700000000000000ea00000000000000dd00000000000000c600000000",
            INIT_44 => X"000000da00000000000000e400000000000000d800000000000000d500000000",
            INIT_45 => X"000000eb00000000000000e900000000000000e000000000000000dd00000000",
            INIT_46 => X"000000f000000000000000ef00000000000000ee00000000000000f000000000",
            INIT_47 => X"000000ee00000000000000f000000000000000f000000000000000f000000000",
            INIT_48 => X"0000009b000000000000008e000000000000008a000000000000008c00000000",
            INIT_49 => X"000000ea00000000000000ec00000000000000ea00000000000000bc00000000",
            INIT_4A => X"000000ed00000000000000ed00000000000000eb00000000000000e900000000",
            INIT_4B => X"000000ed00000000000000ea00000000000000e400000000000000d800000000",
            INIT_4C => X"000000e800000000000000ec00000000000000e600000000000000e600000000",
            INIT_4D => X"000000cc00000000000000db00000000000000e900000000000000ed00000000",
            INIT_4E => X"000000c700000000000000b400000000000000b300000000000000bd00000000",
            INIT_4F => X"000000f000000000000000f000000000000000f100000000000000eb00000000",
            INIT_50 => X"0000007f000000000000007d0000000000000079000000000000008200000000",
            INIT_51 => X"000000e200000000000000e400000000000000e5000000000000009f00000000",
            INIT_52 => X"000000ed00000000000000ec00000000000000ea00000000000000e800000000",
            INIT_53 => X"000000eb00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_54 => X"000000e800000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_55 => X"0000009c00000000000000a500000000000000b800000000000000ce00000000",
            INIT_56 => X"000000a20000000000000085000000000000008c000000000000009500000000",
            INIT_57 => X"000000f000000000000000f000000000000000f100000000000000e400000000",
            INIT_58 => X"000000d300000000000000d300000000000000ca00000000000000d400000000",
            INIT_59 => X"000000d100000000000000d500000000000000e300000000000000d900000000",
            INIT_5A => X"000000dd00000000000000e200000000000000de00000000000000d500000000",
            INIT_5B => X"000000e500000000000000e100000000000000dd00000000000000db00000000",
            INIT_5C => X"000000e700000000000000ed00000000000000ec00000000000000ea00000000",
            INIT_5D => X"000000c200000000000000c800000000000000c600000000000000cc00000000",
            INIT_5E => X"000000c3000000000000009700000000000000b200000000000000c500000000",
            INIT_5F => X"000000f000000000000000f100000000000000f000000000000000e600000000",
            INIT_60 => X"000000d900000000000000d300000000000000ca00000000000000cf00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000db00000000000000e100000000",
            INIT_62 => X"0000007000000000000000b800000000000000d500000000000000b400000000",
            INIT_63 => X"0000008a00000000000000810000000000000079000000000000007200000000",
            INIT_64 => X"000000ec00000000000000d800000000000000a7000000000000009800000000",
            INIT_65 => X"000000e200000000000000ea00000000000000e900000000000000e800000000",
            INIT_66 => X"000000e600000000000000cb00000000000000db00000000000000e400000000",
            INIT_67 => X"000000f100000000000000ef00000000000000e600000000000000e300000000",
            INIT_68 => X"00000083000000000000007d000000000000007d000000000000008200000000",
            INIT_69 => X"000000c700000000000000c900000000000000b6000000000000009100000000",
            INIT_6A => X"0000004700000000000000ac00000000000000e600000000000000db00000000",
            INIT_6B => X"0000005400000000000000490000000000000049000000000000004600000000",
            INIT_6C => X"000000ef00000000000000e300000000000000a8000000000000007200000000",
            INIT_6D => X"000000d300000000000000e400000000000000e700000000000000ed00000000",
            INIT_6E => X"000000ce00000000000000db00000000000000da00000000000000d000000000",
            INIT_6F => X"000000e700000000000000dd00000000000000c500000000000000ba00000000",
            INIT_70 => X"00000055000000000000004f0000000000000056000000000000005100000000",
            INIT_71 => X"000000c8000000000000009d000000000000009b000000000000008d00000000",
            INIT_72 => X"0000007900000000000000b400000000000000df00000000000000e400000000",
            INIT_73 => X"000000c000000000000000970000000000000075000000000000007000000000",
            INIT_74 => X"000000cb00000000000000db00000000000000de00000000000000d400000000",
            INIT_75 => X"0000008a000000000000009a00000000000000a600000000000000ba00000000",
            INIT_76 => X"0000008e0000000000000092000000000000008b000000000000008500000000",
            INIT_77 => X"000000d400000000000000c50000000000000099000000000000008900000000",
            INIT_78 => X"0000009000000000000000620000000000000046000000000000003500000000",
            INIT_79 => X"0000009e0000000000000073000000000000006b000000000000009700000000",
            INIT_7A => X"000000c100000000000000c200000000000000c200000000000000b400000000",
            INIT_7B => X"000000d200000000000000e400000000000000d100000000000000c200000000",
            INIT_7C => X"00000088000000000000009600000000000000a500000000000000b500000000",
            INIT_7D => X"0000006f000000000000006a000000000000006f000000000000007d00000000",
            INIT_7E => X"0000009700000000000000870000000000000079000000000000007600000000",
            INIT_7F => X"000000cb00000000000000ce00000000000000ae00000000000000a400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "sampleifmap_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000000000008c000000000000001d000000000000000f00000000",
            INIT_01 => X"000000a20000000000000085000000000000007b000000000000009600000000",
            INIT_02 => X"000000ea00000000000000e000000000000000d100000000000000b500000000",
            INIT_03 => X"000000bd00000000000000ee00000000000000f100000000000000ea00000000",
            INIT_04 => X"000000a3000000000000009e000000000000009a000000000000009f00000000",
            INIT_05 => X"000000ab00000000000000a500000000000000a500000000000000ab00000000",
            INIT_06 => X"000000cc00000000000000be00000000000000b100000000000000ae00000000",
            INIT_07 => X"000000af00000000000000b700000000000000c400000000000000cf00000000",
            INIT_08 => X"000000e800000000000000cf000000000000003e000000000000000500000000",
            INIT_09 => X"000000e000000000000000d400000000000000cf00000000000000cd00000000",
            INIT_0A => X"000000ee00000000000000ee00000000000000ec00000000000000e600000000",
            INIT_0B => X"000000e400000000000000ee00000000000000ee00000000000000dd00000000",
            INIT_0C => X"000000d500000000000000d800000000000000c800000000000000d900000000",
            INIT_0D => X"000000cc00000000000000d400000000000000d600000000000000d400000000",
            INIT_0E => X"000000a500000000000000b500000000000000bf00000000000000c100000000",
            INIT_0F => X"0000009a000000000000008f0000000000000092000000000000009c00000000",
            INIT_10 => X"000000c400000000000000cc000000000000009b000000000000002d00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000c500000000",
            INIT_12 => X"000000cf00000000000000cf00000000000000cb00000000000000ce00000000",
            INIT_13 => X"000000a900000000000000b000000000000000c600000000000000c100000000",
            INIT_14 => X"0000008500000000000000a300000000000000ab00000000000000a100000000",
            INIT_15 => X"000000870000000000000096000000000000009d000000000000008900000000",
            INIT_16 => X"0000007400000000000000720000000000000070000000000000007300000000",
            INIT_17 => X"0000008e000000000000008d0000000000000085000000000000007d00000000",
            INIT_18 => X"0000009a00000000000000a000000000000000b3000000000000008700000000",
            INIT_19 => X"0000009600000000000000960000000000000098000000000000009800000000",
            INIT_1A => X"0000009500000000000000930000000000000093000000000000009600000000",
            INIT_1B => X"0000007a000000000000007e0000000000000091000000000000009500000000",
            INIT_1C => X"0000006d00000000000000800000000000000086000000000000007800000000",
            INIT_1D => X"0000006700000000000000700000000000000075000000000000007000000000",
            INIT_1E => X"00000075000000000000006f0000000000000067000000000000006100000000",
            INIT_1F => X"000000900000000000000085000000000000007d000000000000007900000000",
            INIT_20 => X"0000005d000000000000005a000000000000005a000000000000005700000000",
            INIT_21 => X"0000006900000000000000660000000000000066000000000000006200000000",
            INIT_22 => X"00000083000000000000007c0000000000000077000000000000006f00000000",
            INIT_23 => X"0000008500000000000000840000000000000088000000000000008900000000",
            INIT_24 => X"00000077000000000000007f0000000000000085000000000000008800000000",
            INIT_25 => X"0000005c00000000000000610000000000000065000000000000006d00000000",
            INIT_26 => X"0000006200000000000000640000000000000064000000000000005e00000000",
            INIT_27 => X"0000009500000000000000870000000000000077000000000000006800000000",
            INIT_28 => X"0000001a0000000000000010000000000000000b000000000000001900000000",
            INIT_29 => X"0000001e00000000000000190000000000000019000000000000001a00000000",
            INIT_2A => X"0000003b0000000000000033000000000000002b000000000000002400000000",
            INIT_2B => X"0000004f000000000000004d000000000000004b000000000000004500000000",
            INIT_2C => X"0000004800000000000000510000000000000058000000000000005700000000",
            INIT_2D => X"0000004500000000000000450000000000000044000000000000004300000000",
            INIT_2E => X"000000640000000000000059000000000000004e000000000000004700000000",
            INIT_2F => X"000000920000000000000088000000000000007c000000000000007100000000",
            INIT_30 => X"0000002c000000000000000d0000000000000010000000000000002e00000000",
            INIT_31 => X"00000008000000000000000b0000000000000019000000000000002d00000000",
            INIT_32 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_33 => X"0000001700000000000000130000000000000012000000000000000d00000000",
            INIT_34 => X"0000001f00000000000000210000000000000026000000000000001d00000000",
            INIT_35 => X"0000003a0000000000000032000000000000002c000000000000002600000000",
            INIT_36 => X"0000007b0000000000000073000000000000005a000000000000004600000000",
            INIT_37 => X"000000a0000000000000008b000000000000007b000000000000007300000000",
            INIT_38 => X"000000290000000000000013000000000000001b000000000000002900000000",
            INIT_39 => X"0000001f00000000000000320000000000000046000000000000005100000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000002400000000000000320000000000000040000000000000001100000000",
            INIT_3C => X"00000023000000000000001e000000000000001e000000000000001e00000000",
            INIT_3D => X"0000006100000000000000470000000000000037000000000000002b00000000",
            INIT_3E => X"0000006900000000000000780000000000000083000000000000007c00000000",
            INIT_3F => X"000000b300000000000000980000000000000086000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000a000000000000000a000000000000000f00000000",
            INIT_41 => X"00000021000000000000002b0000000000000034000000000000002c00000000",
            INIT_42 => X"0000000100000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"00000080000000000000009e0000000000000075000000000000000800000000",
            INIT_44 => X"0000006900000000000000670000000000000069000000000000007000000000",
            INIT_45 => X"0000007e000000000000007e0000000000000073000000000000006b00000000",
            INIT_46 => X"00000074000000000000005e0000000000000056000000000000006a00000000",
            INIT_47 => X"000000c200000000000000ac0000000000000093000000000000008200000000",
            INIT_48 => X"000000040000000000000003000000000000000a000000000000002800000000",
            INIT_49 => X"0000000a000000000000000c000000000000000c000000000000000600000000",
            INIT_4A => X"0000000200000000000000010000000000000001000000000000000600000000",
            INIT_4B => X"000000820000000000000080000000000000003a000000000000000000000000",
            INIT_4C => X"000000710000000000000077000000000000007b000000000000007f00000000",
            INIT_4D => X"00000042000000000000004b0000000000000060000000000000006e00000000",
            INIT_4E => X"000000840000000000000076000000000000005d000000000000004700000000",
            INIT_4F => X"000000c500000000000000b600000000000000a2000000000000008d00000000",
            INIT_50 => X"000000010000000000000001000000000000001d000000000000004d00000000",
            INIT_51 => X"0000000200000000000000030000000000000002000000000000000100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_53 => X"0000002f000000000000002d000000000000000c000000000000000100000000",
            INIT_54 => X"0000003100000000000000320000000000000030000000000000002e00000000",
            INIT_55 => X"0000004d00000000000000300000000000000026000000000000002a00000000",
            INIT_56 => X"000000870000000000000080000000000000007e000000000000006e00000000",
            INIT_57 => X"000000c600000000000000bb00000000000000b0000000000000009900000000",
            INIT_58 => X"0000000100000000000000010000000000000034000000000000005e00000000",
            INIT_59 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002000000000000000190000000000000003000000000000000200000000",
            INIT_5C => X"0000001d00000000000000190000000000000019000000000000001900000000",
            INIT_5D => X"00000071000000000000005c0000000000000042000000000000002900000000",
            INIT_5E => X"0000008b000000000000007f000000000000007e000000000000007c00000000",
            INIT_5F => X"000000c900000000000000bf00000000000000b3000000000000009d00000000",
            INIT_60 => X"000000020000000000000007000000000000003c000000000000006600000000",
            INIT_61 => X"0000000200000000000000030000000000000003000000000000000200000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000001f00000000000000130000000000000001000000000000000300000000",
            INIT_64 => X"0000003a000000000000001b000000000000000d000000000000001100000000",
            INIT_65 => X"0000007c000000000000007e0000000000000073000000000000005a00000000",
            INIT_66 => X"0000009100000000000000870000000000000082000000000000007b00000000",
            INIT_67 => X"000000ca00000000000000c000000000000000b0000000000000009f00000000",
            INIT_68 => X"0000000c00000000000000170000000000000033000000000000006300000000",
            INIT_69 => X"00000007000000000000000a000000000000000b000000000000000a00000000",
            INIT_6A => X"0000000300000000000000040000000000000004000000000000000400000000",
            INIT_6B => X"00000015000000000000000d0000000000000005000000000000000600000000",
            INIT_6C => X"00000062000000000000004d0000000000000032000000000000001b00000000",
            INIT_6D => X"0000007d000000000000007e000000000000007e000000000000007100000000",
            INIT_6E => X"0000009a0000000000000094000000000000008a000000000000008000000000",
            INIT_6F => X"000000ca00000000000000c500000000000000b800000000000000a800000000",
            INIT_70 => X"00000023000000000000002c0000000000000039000000000000006000000000",
            INIT_71 => X"00000017000000000000001a000000000000001c000000000000001e00000000",
            INIT_72 => X"0000001700000000000000160000000000000015000000000000001500000000",
            INIT_73 => X"000000370000000000000028000000000000001f000000000000001b00000000",
            INIT_74 => X"0000007000000000000000660000000000000058000000000000004600000000",
            INIT_75 => X"0000007f000000000000007a000000000000007a000000000000007900000000",
            INIT_76 => X"000000a00000000000000095000000000000008b000000000000008500000000",
            INIT_77 => X"000000ca00000000000000c800000000000000bd00000000000000ac00000000",
            INIT_78 => X"0000003d0000000000000043000000000000004b000000000000006500000000",
            INIT_79 => X"0000003700000000000000350000000000000035000000000000003800000000",
            INIT_7A => X"0000003e000000000000003a0000000000000038000000000000003700000000",
            INIT_7B => X"0000006000000000000000540000000000000047000000000000004300000000",
            INIT_7C => X"000000790000000000000074000000000000006d000000000000006700000000",
            INIT_7D => X"00000083000000000000007d000000000000007c000000000000007f00000000",
            INIT_7E => X"000000a200000000000000980000000000000091000000000000008800000000",
            INIT_7F => X"000000c800000000000000c300000000000000b700000000000000ab00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "sampleifmap_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_05 => X"000000e600000000000000e800000000000000ea00000000000000ea00000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e700000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ea00000000000000e900000000000000e900000000",
            INIT_0D => X"000000eb00000000000000ed00000000000000ee00000000000000ed00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ec00000000000000ea00000000000000e700000000000000e700000000",
            INIT_15 => X"000000ea00000000000000eb00000000000000ee00000000000000e900000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e700000000000000e800000000000000e700000000000000e600000000",
            INIT_1D => X"000000e600000000000000d500000000000000db00000000000000c500000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000db00000000000000e600000000000000ed00000000000000ec00000000",
            INIT_25 => X"000000e800000000000000dd00000000000000d000000000000000b300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e800000000000000ed00000000000000ea00000000000000ec00000000",
            INIT_2C => X"000000c800000000000000cf00000000000000d200000000000000da00000000",
            INIT_2D => X"000000e800000000000000dc00000000000000ca00000000000000bd00000000",
            INIT_2E => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e600000000000000e700000000000000e400000000000000e500000000",
            INIT_31 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_32 => X"000000ee00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_33 => X"000000e400000000000000ee00000000000000e500000000000000e600000000",
            INIT_34 => X"000000be00000000000000bf00000000000000be00000000000000cc00000000",
            INIT_35 => X"000000d300000000000000b100000000000000ab00000000000000b100000000",
            INIT_36 => X"000000eb00000000000000e900000000000000ea00000000000000ef00000000",
            INIT_37 => X"000000ee00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_38 => X"000000ea00000000000000ee00000000000000e900000000000000de00000000",
            INIT_39 => X"000000ec00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_3A => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_3B => X"000000da00000000000000eb00000000000000dd00000000000000cb00000000",
            INIT_3C => X"000000cb00000000000000d300000000000000d200000000000000d200000000",
            INIT_3D => X"000000cc00000000000000b900000000000000bb00000000000000c400000000",
            INIT_3E => X"000000ee00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_3F => X"000000ee00000000000000ee00000000000000ee00000000000000ee00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f300000000000000f600000000000000f300000000000000f100000000",
            INIT_41 => X"000000eb00000000000000eb00000000000000ed00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ed00000000000000ed00000000",
            INIT_43 => X"000000e500000000000000e700000000000000da00000000000000c400000000",
            INIT_44 => X"000000e300000000000000eb00000000000000de00000000000000d900000000",
            INIT_45 => X"000000f100000000000000f000000000000000eb00000000000000ea00000000",
            INIT_46 => X"000000f000000000000000f000000000000000f000000000000000f300000000",
            INIT_47 => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_48 => X"000000a100000000000000990000000000000094000000000000009500000000",
            INIT_49 => X"000000e800000000000000e900000000000000e900000000000000bf00000000",
            INIT_4A => X"000000eb00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000ef00000000000000f100000000000000eb00000000000000e800000000",
            INIT_4D => X"000000d300000000000000e200000000000000f300000000000000f700000000",
            INIT_4E => X"000000c900000000000000b900000000000000ba00000000000000c300000000",
            INIT_4F => X"000000ef00000000000000ef00000000000000ef00000000000000eb00000000",
            INIT_50 => X"0000008900000000000000890000000000000085000000000000008d00000000",
            INIT_51 => X"000000e000000000000000e100000000000000e700000000000000a500000000",
            INIT_52 => X"000000eb00000000000000ea00000000000000ea00000000000000e900000000",
            INIT_53 => X"000000ec00000000000000ee00000000000000ec00000000000000eb00000000",
            INIT_54 => X"000000ee00000000000000f100000000000000f000000000000000ee00000000",
            INIT_55 => X"000000a300000000000000ac00000000000000bf00000000000000d500000000",
            INIT_56 => X"000000a6000000000000008f0000000000000099000000000000009f00000000",
            INIT_57 => X"000000ef00000000000000ee00000000000000ef00000000000000e500000000",
            INIT_58 => X"000000df00000000000000e000000000000000d700000000000000e000000000",
            INIT_59 => X"000000ce00000000000000d300000000000000e700000000000000e300000000",
            INIT_5A => X"000000db00000000000000e100000000000000de00000000000000d600000000",
            INIT_5B => X"000000e900000000000000e600000000000000e100000000000000df00000000",
            INIT_5C => X"000000ed00000000000000f100000000000000ef00000000000000ed00000000",
            INIT_5D => X"000000ca00000000000000cf00000000000000cb00000000000000d000000000",
            INIT_5E => X"000000ca00000000000000a400000000000000c400000000000000d300000000",
            INIT_5F => X"000000ef00000000000000ef00000000000000ee00000000000000e900000000",
            INIT_60 => X"000000ea00000000000000e000000000000000d900000000000000de00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000e300000000000000f100000000",
            INIT_62 => X"0000007900000000000000bc00000000000000d600000000000000b700000000",
            INIT_63 => X"00000093000000000000008b0000000000000084000000000000007e00000000",
            INIT_64 => X"000000ed00000000000000dc00000000000000ae00000000000000a100000000",
            INIT_65 => X"000000e900000000000000f000000000000000ee00000000000000eb00000000",
            INIT_66 => X"000000ed00000000000000d400000000000000e500000000000000ed00000000",
            INIT_67 => X"000000f200000000000000f200000000000000e900000000000000ea00000000",
            INIT_68 => X"00000097000000000000008d0000000000000093000000000000009800000000",
            INIT_69 => X"000000cc00000000000000cd00000000000000c100000000000000a500000000",
            INIT_6A => X"0000005c00000000000000b700000000000000ea00000000000000e200000000",
            INIT_6B => X"00000062000000000000005a000000000000005b000000000000005b00000000",
            INIT_6C => X"000000f100000000000000e900000000000000b3000000000000008100000000",
            INIT_6D => X"000000d900000000000000e900000000000000ed00000000000000f100000000",
            INIT_6E => X"000000d600000000000000df00000000000000dc00000000000000d400000000",
            INIT_6F => X"000000ea00000000000000e300000000000000cd00000000000000c400000000",
            INIT_70 => X"0000006600000000000000640000000000000072000000000000006c00000000",
            INIT_71 => X"000000cf00000000000000a400000000000000a4000000000000009b00000000",
            INIT_72 => X"0000008a00000000000000be00000000000000e400000000000000ea00000000",
            INIT_73 => X"000000cf00000000000000a80000000000000087000000000000008300000000",
            INIT_74 => X"000000d400000000000000e300000000000000e800000000000000df00000000",
            INIT_75 => X"0000009300000000000000a300000000000000ae00000000000000c300000000",
            INIT_76 => X"0000009700000000000000980000000000000090000000000000008c00000000",
            INIT_77 => X"000000d800000000000000cb00000000000000a0000000000000009300000000",
            INIT_78 => X"000000990000000000000074000000000000005e000000000000004d00000000",
            INIT_79 => X"000000a10000000000000076000000000000006e000000000000009c00000000",
            INIT_7A => X"000000c800000000000000c600000000000000c500000000000000b600000000",
            INIT_7B => X"000000d900000000000000ec00000000000000d900000000000000ca00000000",
            INIT_7C => X"00000095000000000000009f00000000000000ac00000000000000ba00000000",
            INIT_7D => X"0000007b0000000000000076000000000000007b000000000000008a00000000",
            INIT_7E => X"000000a100000000000000910000000000000082000000000000008000000000",
            INIT_7F => X"000000d000000000000000d500000000000000b800000000000000ae00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "sampleifmap_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000dc0000000000000097000000000000002f000000000000002300000000",
            INIT_01 => X"000000a20000000000000086000000000000007b000000000000009600000000",
            INIT_02 => X"000000e900000000000000e100000000000000d300000000000000b400000000",
            INIT_03 => X"000000be00000000000000ee00000000000000f000000000000000e800000000",
            INIT_04 => X"000000b100000000000000aa00000000000000a200000000000000a300000000",
            INIT_05 => X"000000bb00000000000000b600000000000000b600000000000000bb00000000",
            INIT_06 => X"000000d900000000000000cc00000000000000bf00000000000000bd00000000",
            INIT_07 => X"000000b700000000000000c100000000000000d000000000000000da00000000",
            INIT_08 => X"000000ef00000000000000d9000000000000004f000000000000001800000000",
            INIT_09 => X"000000e500000000000000da00000000000000d300000000000000d400000000",
            INIT_0A => X"000000ef00000000000000f500000000000000f600000000000000ed00000000",
            INIT_0B => X"000000ea00000000000000f100000000000000ef00000000000000dc00000000",
            INIT_0C => X"000000e500000000000000e600000000000000d600000000000000e400000000",
            INIT_0D => X"000000e000000000000000e800000000000000ea00000000000000e700000000",
            INIT_0E => X"000000b300000000000000c500000000000000d100000000000000d400000000",
            INIT_0F => X"000000a5000000000000009e00000000000000a100000000000000a900000000",
            INIT_10 => X"000000d800000000000000de00000000000000b3000000000000004700000000",
            INIT_11 => X"000000e300000000000000e600000000000000e500000000000000d900000000",
            INIT_12 => X"000000dd00000000000000e400000000000000e400000000000000e300000000",
            INIT_13 => X"000000bc00000000000000c100000000000000d700000000000000cf00000000",
            INIT_14 => X"0000009c00000000000000ba00000000000000c300000000000000b800000000",
            INIT_15 => X"0000009e00000000000000ad00000000000000b400000000000000a100000000",
            INIT_16 => X"0000008300000000000000850000000000000087000000000000008a00000000",
            INIT_17 => X"0000009c000000000000009e0000000000000097000000000000008c00000000",
            INIT_18 => X"000000bd00000000000000c200000000000000cf00000000000000a100000000",
            INIT_19 => X"000000c100000000000000c000000000000000be00000000000000bb00000000",
            INIT_1A => X"000000bd00000000000000bd00000000000000be00000000000000c000000000",
            INIT_1B => X"0000009a00000000000000a300000000000000ba00000000000000bc00000000",
            INIT_1C => X"0000009100000000000000a300000000000000aa000000000000009a00000000",
            INIT_1D => X"0000008800000000000000900000000000000099000000000000009400000000",
            INIT_1E => X"0000008d000000000000008b0000000000000086000000000000008200000000",
            INIT_1F => X"0000009c00000000000000940000000000000092000000000000009000000000",
            INIT_20 => X"0000007f000000000000007a0000000000000071000000000000006d00000000",
            INIT_21 => X"000000960000000000000093000000000000008e000000000000008600000000",
            INIT_22 => X"000000ac00000000000000a500000000000000a0000000000000009800000000",
            INIT_23 => X"000000af00000000000000b400000000000000ba00000000000000b500000000",
            INIT_24 => X"0000009b00000000000000a300000000000000a800000000000000ac00000000",
            INIT_25 => X"0000007f0000000000000084000000000000008b000000000000009400000000",
            INIT_26 => X"0000007a00000000000000810000000000000085000000000000008100000000",
            INIT_27 => X"0000009c0000000000000092000000000000008a000000000000007e00000000",
            INIT_28 => X"0000003000000000000000230000000000000019000000000000002900000000",
            INIT_29 => X"0000003d000000000000003a0000000000000038000000000000003400000000",
            INIT_2A => X"00000057000000000000004d0000000000000046000000000000003e00000000",
            INIT_2B => X"0000007e000000000000007e0000000000000079000000000000006a00000000",
            INIT_2C => X"000000700000000000000078000000000000007e000000000000007f00000000",
            INIT_2D => X"0000006600000000000000670000000000000068000000000000006a00000000",
            INIT_2E => X"000000770000000000000073000000000000006e000000000000006900000000",
            INIT_2F => X"00000095000000000000008d0000000000000088000000000000008000000000",
            INIT_30 => X"0000003500000000000000130000000000000014000000000000003700000000",
            INIT_31 => X"00000018000000000000001e0000000000000029000000000000003a00000000",
            INIT_32 => X"00000014000000000000000f000000000000000f000000000000001100000000",
            INIT_33 => X"0000003e000000000000003c0000000000000038000000000000002a00000000",
            INIT_34 => X"0000004c000000000000004d0000000000000051000000000000004700000000",
            INIT_35 => X"0000005a0000000000000053000000000000004f000000000000004e00000000",
            INIT_36 => X"0000008a000000000000008a0000000000000076000000000000006500000000",
            INIT_37 => X"0000009e00000000000000890000000000000080000000000000007d00000000",
            INIT_38 => X"000000290000000000000012000000000000001a000000000000002d00000000",
            INIT_39 => X"000000250000000000000039000000000000004c000000000000005400000000",
            INIT_3A => X"000000070000000000000007000000000000000b000000000000001500000000",
            INIT_3B => X"0000003e000000000000004e000000000000005b000000000000002300000000",
            INIT_3C => X"00000045000000000000003f000000000000003e000000000000003c00000000",
            INIT_3D => X"0000007b00000000000000630000000000000053000000000000004a00000000",
            INIT_3E => X"0000007200000000000000870000000000000095000000000000009200000000",
            INIT_3F => X"000000af00000000000000920000000000000085000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000000000080000000000000009000000000000001100000000",
            INIT_41 => X"00000023000000000000002f0000000000000039000000000000002e00000000",
            INIT_42 => X"0000000300000000000000040000000000000007000000000000001400000000",
            INIT_43 => X"0000009400000000000000b30000000000000086000000000000000f00000000",
            INIT_44 => X"0000007f000000000000007c000000000000007d000000000000008300000000",
            INIT_45 => X"0000008d00000000000000900000000000000085000000000000007e00000000",
            INIT_46 => X"000000740000000000000061000000000000005b000000000000007400000000",
            INIT_47 => X"000000be00000000000000a50000000000000090000000000000008100000000",
            INIT_48 => X"0000000400000000000000030000000000000007000000000000002300000000",
            INIT_49 => X"0000000c00000000000000110000000000000011000000000000000700000000",
            INIT_4A => X"0000000300000000000000020000000000000003000000000000000700000000",
            INIT_4B => X"0000009400000000000000920000000000000040000000000000000200000000",
            INIT_4C => X"000000810000000000000089000000000000008d000000000000009000000000",
            INIT_4D => X"000000450000000000000053000000000000006a000000000000007a00000000",
            INIT_4E => X"0000007e00000000000000710000000000000058000000000000004600000000",
            INIT_4F => X"000000c200000000000000b0000000000000009e000000000000008700000000",
            INIT_50 => X"0000000200000000000000010000000000000015000000000000004000000000",
            INIT_51 => X"0000000500000000000000090000000000000005000000000000000000000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000200000000",
            INIT_53 => X"00000044000000000000003b000000000000000b000000000000000100000000",
            INIT_54 => X"0000003b00000000000000430000000000000045000000000000004300000000",
            INIT_55 => X"00000047000000000000002e000000000000002a000000000000003100000000",
            INIT_56 => X"0000008000000000000000780000000000000074000000000000006600000000",
            INIT_57 => X"000000c400000000000000b700000000000000ab000000000000009300000000",
            INIT_58 => X"000000020000000000000001000000000000002b000000000000005200000000",
            INIT_59 => X"0000000200000000000000050000000000000002000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003600000000000000260000000000000002000000000000000000000000",
            INIT_5C => X"000000220000000000000024000000000000002b000000000000002e00000000",
            INIT_5D => X"0000006900000000000000520000000000000038000000000000002700000000",
            INIT_5E => X"0000008300000000000000760000000000000073000000000000007300000000",
            INIT_5F => X"000000c700000000000000bb00000000000000ae000000000000009600000000",
            INIT_60 => X"0000000100000000000000030000000000000032000000000000005d00000000",
            INIT_61 => X"0000000200000000000000030000000000000001000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000002f000000000000001c0000000000000000000000000000000200000000",
            INIT_64 => X"000000370000000000000016000000000000000c000000000000001700000000",
            INIT_65 => X"00000070000000000000006f0000000000000063000000000000005100000000",
            INIT_66 => X"00000089000000000000007e0000000000000077000000000000007100000000",
            INIT_67 => X"000000c900000000000000bc00000000000000ab000000000000009700000000",
            INIT_68 => X"00000004000000000000000b0000000000000025000000000000005900000000",
            INIT_69 => X"0000000200000000000000040000000000000004000000000000000200000000",
            INIT_6A => X"0000000200000000000000010000000000000001000000000000000100000000",
            INIT_6B => X"00000018000000000000000d0000000000000002000000000000000600000000",
            INIT_6C => X"00000052000000000000003e0000000000000029000000000000001900000000",
            INIT_6D => X"0000006f00000000000000700000000000000071000000000000006500000000",
            INIT_6E => X"000000910000000000000089000000000000007e000000000000007300000000",
            INIT_6F => X"000000c900000000000000c100000000000000b300000000000000a100000000",
            INIT_70 => X"0000001100000000000000160000000000000024000000000000005200000000",
            INIT_71 => X"0000000c000000000000000d000000000000000f000000000000000f00000000",
            INIT_72 => X"0000000f000000000000000e000000000000000d000000000000000c00000000",
            INIT_73 => X"0000002d000000000000001b0000000000000015000000000000001400000000",
            INIT_74 => X"0000005800000000000000550000000000000051000000000000004300000000",
            INIT_75 => X"00000070000000000000006b000000000000006e000000000000006900000000",
            INIT_76 => X"00000097000000000000008a000000000000007f000000000000007700000000",
            INIT_77 => X"000000c800000000000000c400000000000000b700000000000000a400000000",
            INIT_78 => X"0000002500000000000000260000000000000030000000000000005300000000",
            INIT_79 => X"0000002600000000000000220000000000000021000000000000002300000000",
            INIT_7A => X"0000002e000000000000002c0000000000000029000000000000002800000000",
            INIT_7B => X"0000004a000000000000003b0000000000000030000000000000002d00000000",
            INIT_7C => X"000000610000000000000061000000000000005c000000000000005300000000",
            INIT_7D => X"00000075000000000000006c000000000000006a000000000000006b00000000",
            INIT_7E => X"00000099000000000000008d0000000000000085000000000000007b00000000",
            INIT_7F => X"000000c700000000000000bf00000000000000b200000000000000a300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "sampleifmap_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000084000000000000008b000000000000009e000000000000009e00000000",
            INIT_01 => X"000000c100000000000000bb00000000000000b600000000000000a600000000",
            INIT_02 => X"000000ce00000000000000d100000000000000cd00000000000000c700000000",
            INIT_03 => X"000000e600000000000000e300000000000000df00000000000000da00000000",
            INIT_04 => X"000000eb00000000000000e700000000000000e200000000000000d500000000",
            INIT_05 => X"000000ea00000000000000ea00000000000000e800000000000000ec00000000",
            INIT_06 => X"000000ee00000000000000e600000000000000e200000000000000ec00000000",
            INIT_07 => X"000000ee00000000000000ed00000000000000e400000000000000e800000000",
            INIT_08 => X"00000089000000000000009700000000000000ac00000000000000aa00000000",
            INIT_09 => X"000000c700000000000000c500000000000000c100000000000000ae00000000",
            INIT_0A => X"000000d200000000000000d900000000000000d700000000000000ce00000000",
            INIT_0B => X"000000ed00000000000000e900000000000000e700000000000000e100000000",
            INIT_0C => X"000000f200000000000000e800000000000000e400000000000000db00000000",
            INIT_0D => X"000000f200000000000000ec00000000000000ea00000000000000f500000000",
            INIT_0E => X"000000f300000000000000eb00000000000000e400000000000000f100000000",
            INIT_0F => X"000000f600000000000000f600000000000000e800000000000000e900000000",
            INIT_10 => X"0000008e000000000000009d00000000000000b000000000000000ae00000000",
            INIT_11 => X"000000c700000000000000ce00000000000000c900000000000000b500000000",
            INIT_12 => X"000000d400000000000000da00000000000000df00000000000000d100000000",
            INIT_13 => X"000000ef00000000000000e600000000000000e600000000000000e000000000",
            INIT_14 => X"000000ef00000000000000e900000000000000e400000000000000dd00000000",
            INIT_15 => X"000000f300000000000000ec00000000000000d500000000000000e800000000",
            INIT_16 => X"000000f800000000000000ee00000000000000e700000000000000f500000000",
            INIT_17 => X"000000f500000000000000fa00000000000000e600000000000000ed00000000",
            INIT_18 => X"0000009300000000000000a000000000000000b200000000000000b400000000",
            INIT_19 => X"000000cf00000000000000d400000000000000cb00000000000000ba00000000",
            INIT_1A => X"000000d600000000000000dd00000000000000e400000000000000d600000000",
            INIT_1B => X"000000f000000000000000df00000000000000e700000000000000dc00000000",
            INIT_1C => X"000000e400000000000000e900000000000000e400000000000000e000000000",
            INIT_1D => X"000000f300000000000000e600000000000000ac00000000000000b100000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f400000000000000f900000000000000e400000000000000ee00000000",
            INIT_20 => X"0000009300000000000000a500000000000000b900000000000000ba00000000",
            INIT_21 => X"000000cf00000000000000d900000000000000cc00000000000000bd00000000",
            INIT_22 => X"000000d600000000000000de00000000000000e700000000000000d300000000",
            INIT_23 => X"000000eb00000000000000d300000000000000e700000000000000da00000000",
            INIT_24 => X"000000d400000000000000e800000000000000e000000000000000e200000000",
            INIT_25 => X"000000ed00000000000000e000000000000000a8000000000000009f00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f200000000000000f800000000000000ea00000000000000e800000000",
            INIT_28 => X"0000008e00000000000000aa00000000000000be00000000000000c100000000",
            INIT_29 => X"000000d300000000000000db00000000000000cb00000000000000bf00000000",
            INIT_2A => X"000000d600000000000000dd00000000000000ea00000000000000d700000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e400000000000000d600000000",
            INIT_2C => X"000000c100000000000000eb00000000000000ce00000000000000cf00000000",
            INIT_2D => X"000000e600000000000000de000000000000009e000000000000007000000000",
            INIT_2E => X"000000f100000000000000e200000000000000e500000000000000f500000000",
            INIT_2F => X"000000eb00000000000000f300000000000000e700000000000000e400000000",
            INIT_30 => X"0000008500000000000000ac00000000000000bf00000000000000c400000000",
            INIT_31 => X"000000d900000000000000de00000000000000ca00000000000000bf00000000",
            INIT_32 => X"000000d600000000000000da00000000000000eb00000000000000df00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e300000000000000d700000000",
            INIT_34 => X"000000bb00000000000000cd00000000000000ba00000000000000bb00000000",
            INIT_35 => X"000000b700000000000000ac0000000000000089000000000000007800000000",
            INIT_36 => X"000000eb00000000000000d800000000000000df00000000000000db00000000",
            INIT_37 => X"000000eb00000000000000f000000000000000e100000000000000e200000000",
            INIT_38 => X"0000008c00000000000000ae00000000000000c500000000000000cc00000000",
            INIT_39 => X"000000e000000000000000e000000000000000da00000000000000cb00000000",
            INIT_3A => X"000000dc00000000000000dc00000000000000ed00000000000000e800000000",
            INIT_3B => X"000000cd00000000000000c900000000000000dd00000000000000dc00000000",
            INIT_3C => X"000000530000000000000064000000000000008a00000000000000ac00000000",
            INIT_3D => X"0000003c0000000000000041000000000000003e000000000000004700000000",
            INIT_3E => X"000000e400000000000000d100000000000000b6000000000000006800000000",
            INIT_3F => X"000000ec00000000000000ef00000000000000d400000000000000da00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000089000000000000009d00000000000000aa00000000000000af00000000",
            INIT_41 => X"000000c500000000000000af00000000000000ba00000000000000b000000000",
            INIT_42 => X"000000d200000000000000ce00000000000000d400000000000000d100000000",
            INIT_43 => X"000000c100000000000000c100000000000000c900000000000000d400000000",
            INIT_44 => X"0000005b00000000000000590000000000000069000000000000008e00000000",
            INIT_45 => X"00000045000000000000005e0000000000000053000000000000005400000000",
            INIT_46 => X"000000b700000000000000a20000000000000079000000000000004e00000000",
            INIT_47 => X"000000c300000000000000cf00000000000000a300000000000000ae00000000",
            INIT_48 => X"0000006800000000000000710000000000000073000000000000007200000000",
            INIT_49 => X"00000080000000000000006f000000000000006b000000000000006900000000",
            INIT_4A => X"0000009b00000000000000970000000000000092000000000000008b00000000",
            INIT_4B => X"0000009600000000000000970000000000000093000000000000009d00000000",
            INIT_4C => X"0000006300000000000000630000000000000064000000000000007600000000",
            INIT_4D => X"0000005300000000000000560000000000000056000000000000005500000000",
            INIT_4E => X"00000099000000000000009a0000000000000080000000000000008b00000000",
            INIT_4F => X"0000007b0000000000000084000000000000006d000000000000007600000000",
            INIT_50 => X"00000044000000000000004b000000000000004c000000000000004200000000",
            INIT_51 => X"0000005a0000000000000054000000000000005a000000000000005300000000",
            INIT_52 => X"000000670000000000000066000000000000006a000000000000005d00000000",
            INIT_53 => X"0000006c0000000000000072000000000000006b000000000000006a00000000",
            INIT_54 => X"00000055000000000000005b000000000000005a000000000000005a00000000",
            INIT_55 => X"00000072000000000000005f0000000000000042000000000000004800000000",
            INIT_56 => X"000000c70000000000000093000000000000006e000000000000008000000000",
            INIT_57 => X"0000005e000000000000005c0000000000000067000000000000007d00000000",
            INIT_58 => X"0000004d000000000000004b0000000000000041000000000000003500000000",
            INIT_59 => X"000000460000000000000055000000000000006a000000000000006f00000000",
            INIT_5A => X"0000005d000000000000005f0000000000000071000000000000005d00000000",
            INIT_5B => X"00000061000000000000006b0000000000000073000000000000006c00000000",
            INIT_5C => X"000000610000000000000062000000000000005f000000000000006200000000",
            INIT_5D => X"000000bb00000000000000950000000000000055000000000000005a00000000",
            INIT_5E => X"000000cc0000000000000070000000000000009200000000000000b300000000",
            INIT_5F => X"000000550000000000000057000000000000005f000000000000009a00000000",
            INIT_60 => X"0000004a000000000000005e0000000000000056000000000000003a00000000",
            INIT_61 => X"00000055000000000000004d0000000000000064000000000000006400000000",
            INIT_62 => X"0000006c000000000000007f0000000000000085000000000000007800000000",
            INIT_63 => X"000000570000000000000062000000000000006e000000000000006900000000",
            INIT_64 => X"0000005f00000000000000570000000000000051000000000000005100000000",
            INIT_65 => X"000000c300000000000000aa0000000000000070000000000000005f00000000",
            INIT_66 => X"000000ad000000000000007f00000000000000c100000000000000d000000000",
            INIT_67 => X"0000004f0000000000000055000000000000005000000000000000b200000000",
            INIT_68 => X"0000004b00000000000000570000000000000059000000000000004a00000000",
            INIT_69 => X"0000005000000000000000470000000000000044000000000000005200000000",
            INIT_6A => X"0000006f00000000000000760000000000000067000000000000005900000000",
            INIT_6B => X"000000620000000000000069000000000000006a000000000000006500000000",
            INIT_6C => X"0000006d00000000000000620000000000000062000000000000006000000000",
            INIT_6D => X"000000b800000000000000b4000000000000008e000000000000007200000000",
            INIT_6E => X"0000008400000000000000a000000000000000c000000000000000bf00000000",
            INIT_6F => X"00000043000000000000003c000000000000005000000000000000aa00000000",
            INIT_70 => X"0000004e0000000000000052000000000000004f000000000000004d00000000",
            INIT_71 => X"0000005600000000000000460000000000000048000000000000004f00000000",
            INIT_72 => X"0000008500000000000000810000000000000079000000000000006d00000000",
            INIT_73 => X"0000008300000000000000870000000000000088000000000000008900000000",
            INIT_74 => X"0000009600000000000000920000000000000094000000000000009200000000",
            INIT_75 => X"000000b500000000000000b300000000000000a3000000000000009400000000",
            INIT_76 => X"0000006500000000000000aa00000000000000b000000000000000b900000000",
            INIT_77 => X"0000003b00000000000000370000000000000049000000000000005a00000000",
            INIT_78 => X"00000068000000000000006a000000000000005e000000000000006000000000",
            INIT_79 => X"0000008a00000000000000840000000000000083000000000000006d00000000",
            INIT_7A => X"0000009a000000000000009b0000000000000098000000000000009000000000",
            INIT_7B => X"00000094000000000000009e000000000000009b000000000000009b00000000",
            INIT_7C => X"00000092000000000000009c000000000000009d000000000000009600000000",
            INIT_7D => X"000000a900000000000000920000000000000082000000000000007700000000",
            INIT_7E => X"0000006900000000000000a700000000000000a800000000000000b100000000",
            INIT_7F => X"0000004800000000000000560000000000000062000000000000004500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "sampleifmap_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008300000000000000730000000000000065000000000000006a00000000",
            INIT_01 => X"0000008f00000000000000900000000000000087000000000000008100000000",
            INIT_02 => X"0000009a000000000000009a0000000000000096000000000000009200000000",
            INIT_03 => X"0000009000000000000000970000000000000099000000000000009a00000000",
            INIT_04 => X"0000007f000000000000008b0000000000000086000000000000008200000000",
            INIT_05 => X"0000009f00000000000000920000000000000075000000000000005e00000000",
            INIT_06 => X"0000008400000000000000a200000000000000a300000000000000a700000000",
            INIT_07 => X"00000069000000000000009a00000000000000c0000000000000009000000000",
            INIT_08 => X"0000006d0000000000000076000000000000006c000000000000005f00000000",
            INIT_09 => X"000000910000000000000081000000000000005d000000000000005f00000000",
            INIT_0A => X"0000009000000000000000960000000000000097000000000000009500000000",
            INIT_0B => X"0000007b000000000000007a000000000000007e000000000000008600000000",
            INIT_0C => X"00000094000000000000009b0000000000000085000000000000007a00000000",
            INIT_0D => X"0000009c00000000000000a20000000000000093000000000000008300000000",
            INIT_0E => X"0000009500000000000000990000000000000097000000000000009d00000000",
            INIT_0F => X"00000094000000000000009d00000000000000a4000000000000009f00000000",
            INIT_10 => X"0000004600000000000000490000000000000059000000000000006600000000",
            INIT_11 => X"0000008c000000000000007b000000000000006f000000000000005600000000",
            INIT_12 => X"0000007500000000000000780000000000000081000000000000008f00000000",
            INIT_13 => X"0000008d0000000000000085000000000000007e000000000000007800000000",
            INIT_14 => X"0000009f0000000000000099000000000000008e000000000000009600000000",
            INIT_15 => X"000000a100000000000000a5000000000000009d000000000000009700000000",
            INIT_16 => X"00000090000000000000009a0000000000000098000000000000009900000000",
            INIT_17 => X"00000095000000000000007d0000000000000079000000000000008300000000",
            INIT_18 => X"0000006e0000000000000047000000000000003d000000000000005600000000",
            INIT_19 => X"0000007b0000000000000082000000000000008a000000000000008000000000",
            INIT_1A => X"000000840000000000000076000000000000006c000000000000007600000000",
            INIT_1B => X"00000099000000000000009c0000000000000098000000000000008f00000000",
            INIT_1C => X"0000009a00000000000000910000000000000089000000000000009500000000",
            INIT_1D => X"000000a400000000000000a0000000000000009a000000000000009900000000",
            INIT_1E => X"00000069000000000000007d0000000000000090000000000000009800000000",
            INIT_1F => X"000000840000000000000056000000000000004b000000000000005c00000000",
            INIT_20 => X"00000072000000000000006b0000000000000067000000000000006800000000",
            INIT_21 => X"00000076000000000000007b0000000000000074000000000000007300000000",
            INIT_22 => X"00000090000000000000008d0000000000000086000000000000007400000000",
            INIT_23 => X"000000750000000000000085000000000000008d000000000000008f00000000",
            INIT_24 => X"0000009600000000000000820000000000000059000000000000006200000000",
            INIT_25 => X"000000910000000000000098000000000000009a000000000000009700000000",
            INIT_26 => X"00000050000000000000005a0000000000000060000000000000007500000000",
            INIT_27 => X"0000004100000000000000490000000000000047000000000000004100000000",
            INIT_28 => X"0000006f000000000000006f000000000000006b000000000000006300000000",
            INIT_29 => X"0000007e000000000000007d0000000000000077000000000000007200000000",
            INIT_2A => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_2B => X"0000003d000000000000005b0000000000000082000000000000008300000000",
            INIT_2C => X"0000009400000000000000730000000000000038000000000000003900000000",
            INIT_2D => X"0000005f00000000000000720000000000000082000000000000008b00000000",
            INIT_2E => X"0000003a00000000000000490000000000000053000000000000005600000000",
            INIT_2F => X"0000001b0000000000000033000000000000004b000000000000003c00000000",
            INIT_30 => X"0000007200000000000000740000000000000068000000000000003e00000000",
            INIT_31 => X"0000005b00000000000000660000000000000075000000000000007400000000",
            INIT_32 => X"00000070000000000000004e0000000000000051000000000000005400000000",
            INIT_33 => X"0000004c00000000000000600000000000000082000000000000008500000000",
            INIT_34 => X"0000006c000000000000006b0000000000000056000000000000005300000000",
            INIT_35 => X"0000005100000000000000530000000000000058000000000000006000000000",
            INIT_36 => X"0000002d0000000000000033000000000000003d000000000000004600000000",
            INIT_37 => X"00000018000000000000001e000000000000002e000000000000003400000000",
            INIT_38 => X"00000069000000000000006a0000000000000060000000000000003900000000",
            INIT_39 => X"0000003500000000000000410000000000000068000000000000006b00000000",
            INIT_3A => X"0000006e00000000000000440000000000000040000000000000003b00000000",
            INIT_3B => X"0000006200000000000000730000000000000085000000000000008700000000",
            INIT_3C => X"00000050000000000000004e000000000000004f000000000000005800000000",
            INIT_3D => X"0000003700000000000000460000000000000050000000000000005100000000",
            INIT_3E => X"00000029000000000000002d0000000000000031000000000000002c00000000",
            INIT_3F => X"00000018000000000000001b000000000000001e000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000068000000000000005a000000000000004100000000",
            INIT_41 => X"00000049000000000000004f000000000000006d000000000000006d00000000",
            INIT_42 => X"0000006a00000000000000620000000000000058000000000000005500000000",
            INIT_43 => X"0000004100000000000000440000000000000053000000000000006200000000",
            INIT_44 => X"000000520000000000000051000000000000004a000000000000004600000000",
            INIT_45 => X"0000002c00000000000000290000000000000033000000000000004800000000",
            INIT_46 => X"0000002300000000000000270000000000000037000000000000003d00000000",
            INIT_47 => X"00000019000000000000001b000000000000001e000000000000002000000000",
            INIT_48 => X"0000006700000000000000690000000000000057000000000000004300000000",
            INIT_49 => X"0000005100000000000000580000000000000063000000000000006600000000",
            INIT_4A => X"00000039000000000000003b0000000000000045000000000000004c00000000",
            INIT_4B => X"000000460000000000000042000000000000003f000000000000003a00000000",
            INIT_4C => X"00000036000000000000003e0000000000000044000000000000004800000000",
            INIT_4D => X"0000002c0000000000000031000000000000002f000000000000002e00000000",
            INIT_4E => X"0000001c000000000000001e000000000000002e000000000000003800000000",
            INIT_4F => X"0000001e00000000000000180000000000000019000000000000001d00000000",
            INIT_50 => X"0000003a0000000000000041000000000000003a000000000000003600000000",
            INIT_51 => X"0000002c000000000000002d0000000000000032000000000000003700000000",
            INIT_52 => X"0000003a00000000000000370000000000000033000000000000002e00000000",
            INIT_53 => X"0000003a000000000000003e0000000000000040000000000000003e00000000",
            INIT_54 => X"0000003000000000000000250000000000000026000000000000003300000000",
            INIT_55 => X"00000026000000000000002a0000000000000030000000000000003100000000",
            INIT_56 => X"0000001c000000000000001b0000000000000020000000000000002900000000",
            INIT_57 => X"0000001f000000000000001c0000000000000019000000000000001b00000000",
            INIT_58 => X"0000001b000000000000001a000000000000001d000000000000001e00000000",
            INIT_59 => X"0000002700000000000000210000000000000020000000000000001f00000000",
            INIT_5A => X"0000003300000000000000350000000000000034000000000000003100000000",
            INIT_5B => X"0000002800000000000000260000000000000028000000000000002e00000000",
            INIT_5C => X"000000370000000000000042000000000000002c000000000000002600000000",
            INIT_5D => X"0000002500000000000000240000000000000025000000000000002900000000",
            INIT_5E => X"0000001b000000000000001a000000000000001b000000000000001f00000000",
            INIT_5F => X"000000170000000000000021000000000000001e000000000000001c00000000",
            INIT_60 => X"0000001c000000000000001b000000000000001f000000000000002100000000",
            INIT_61 => X"00000020000000000000001f000000000000001e000000000000001c00000000",
            INIT_62 => X"0000001e000000000000001e0000000000000021000000000000002300000000",
            INIT_63 => X"0000002d00000000000000290000000000000027000000000000002200000000",
            INIT_64 => X"0000003100000000000000490000000000000034000000000000002a00000000",
            INIT_65 => X"0000002000000000000000260000000000000023000000000000001e00000000",
            INIT_66 => X"0000001d000000000000001b000000000000001a000000000000001b00000000",
            INIT_67 => X"0000000d000000000000001a0000000000000026000000000000001e00000000",
            INIT_68 => X"0000001a000000000000001a000000000000001e000000000000001f00000000",
            INIT_69 => X"0000001b000000000000001a0000000000000019000000000000001900000000",
            INIT_6A => X"0000002800000000000000250000000000000020000000000000001d00000000",
            INIT_6B => X"0000002a00000000000000280000000000000029000000000000002a00000000",
            INIT_6C => X"000000260000000000000040000000000000002e000000000000002700000000",
            INIT_6D => X"0000001d000000000000001e0000000000000024000000000000001c00000000",
            INIT_6E => X"0000001c000000000000001b0000000000000019000000000000001a00000000",
            INIT_6F => X"0000000400000000000000090000000000000025000000000000002100000000",
            INIT_70 => X"0000001c0000000000000019000000000000001b000000000000001700000000",
            INIT_71 => X"0000002500000000000000220000000000000020000000000000001e00000000",
            INIT_72 => X"0000002700000000000000280000000000000027000000000000002700000000",
            INIT_73 => X"00000021000000000000001e0000000000000023000000000000002600000000",
            INIT_74 => X"0000002400000000000000390000000000000024000000000000001c00000000",
            INIT_75 => X"0000001d000000000000001d000000000000001d000000000000001e00000000",
            INIT_76 => X"0000001b00000000000000170000000000000018000000000000001800000000",
            INIT_77 => X"0000000500000000000000040000000000000013000000000000002400000000",
            INIT_78 => X"000000220000000000000020000000000000001e000000000000001c00000000",
            INIT_79 => X"0000002500000000000000230000000000000022000000000000002100000000",
            INIT_7A => X"0000002200000000000000240000000000000026000000000000002600000000",
            INIT_7B => X"0000000c000000000000000f0000000000000018000000000000001e00000000",
            INIT_7C => X"00000020000000000000002d0000000000000013000000000000000800000000",
            INIT_7D => X"0000001c000000000000001b000000000000001b000000000000001900000000",
            INIT_7E => X"0000002200000000000000140000000000000015000000000000001800000000",
            INIT_7F => X"0000000700000000000000040000000000000005000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "sampleifmap_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e00000000000000a600000000000000bb00000000000000be00000000",
            INIT_01 => X"000000d800000000000000d300000000000000d000000000000000c100000000",
            INIT_02 => X"000000da00000000000000de00000000000000dd00000000000000db00000000",
            INIT_03 => X"000000ed00000000000000eb00000000000000e800000000000000e500000000",
            INIT_04 => X"000000ef00000000000000ee00000000000000e900000000000000dc00000000",
            INIT_05 => X"000000f100000000000000f100000000000000ef00000000000000f100000000",
            INIT_06 => X"000000f300000000000000eb00000000000000e700000000000000f200000000",
            INIT_07 => X"000000f100000000000000ef00000000000000e700000000000000ed00000000",
            INIT_08 => X"000000a000000000000000b000000000000000c700000000000000c800000000",
            INIT_09 => X"000000da00000000000000da00000000000000d900000000000000c700000000",
            INIT_0A => X"000000db00000000000000e500000000000000e500000000000000df00000000",
            INIT_0B => X"000000f300000000000000ef00000000000000ee00000000000000e900000000",
            INIT_0C => X"000000f500000000000000ee00000000000000ea00000000000000e100000000",
            INIT_0D => X"000000f500000000000000ef00000000000000ed00000000000000f700000000",
            INIT_0E => X"000000f800000000000000ef00000000000000e900000000000000f500000000",
            INIT_0F => X"000000f700000000000000f600000000000000e800000000000000ec00000000",
            INIT_10 => X"000000a200000000000000b300000000000000c800000000000000c900000000",
            INIT_11 => X"000000d600000000000000df00000000000000dc00000000000000c900000000",
            INIT_12 => X"000000db00000000000000e200000000000000e900000000000000dd00000000",
            INIT_13 => X"000000f400000000000000ea00000000000000ea00000000000000e500000000",
            INIT_14 => X"000000f300000000000000ee00000000000000e900000000000000e200000000",
            INIT_15 => X"000000f100000000000000ea00000000000000d600000000000000eb00000000",
            INIT_16 => X"000000fa00000000000000f000000000000000e900000000000000f700000000",
            INIT_17 => X"000000f400000000000000f900000000000000e500000000000000ee00000000",
            INIT_18 => X"000000a400000000000000b300000000000000c700000000000000cb00000000",
            INIT_19 => X"000000d900000000000000e100000000000000d900000000000000c900000000",
            INIT_1A => X"000000d900000000000000e300000000000000eb00000000000000df00000000",
            INIT_1B => X"000000f400000000000000e200000000000000e800000000000000dd00000000",
            INIT_1C => X"000000eb00000000000000ed00000000000000e700000000000000e400000000",
            INIT_1D => X"000000f100000000000000e400000000000000af00000000000000b800000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f200000000000000f700000000000000e300000000000000ed00000000",
            INIT_20 => X"000000a100000000000000b500000000000000cc00000000000000cf00000000",
            INIT_21 => X"000000d500000000000000e100000000000000d600000000000000c900000000",
            INIT_22 => X"000000d700000000000000e200000000000000ed00000000000000d700000000",
            INIT_23 => X"000000ec00000000000000d400000000000000e500000000000000d900000000",
            INIT_24 => X"000000e100000000000000ec00000000000000e100000000000000e300000000",
            INIT_25 => X"000000ec00000000000000e000000000000000ae00000000000000aa00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000ef00000000000000f500000000000000e700000000000000e700000000",
            INIT_28 => X"0000009a00000000000000b700000000000000cd00000000000000d000000000",
            INIT_29 => X"000000d700000000000000e200000000000000d400000000000000c900000000",
            INIT_2A => X"000000d700000000000000df00000000000000ee00000000000000da00000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e500000000000000d700000000",
            INIT_2C => X"000000cc00000000000000ef00000000000000d000000000000000d100000000",
            INIT_2D => X"000000e900000000000000e300000000000000a7000000000000007c00000000",
            INIT_2E => X"000000ef00000000000000e100000000000000e500000000000000f600000000",
            INIT_2F => X"000000e800000000000000f100000000000000e600000000000000e200000000",
            INIT_30 => X"0000008b00000000000000b300000000000000c700000000000000cc00000000",
            INIT_31 => X"000000d500000000000000dd00000000000000cb00000000000000c200000000",
            INIT_32 => X"000000d400000000000000d800000000000000e900000000000000db00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e600000000000000d800000000",
            INIT_34 => X"000000c000000000000000d400000000000000c000000000000000be00000000",
            INIT_35 => X"000000be00000000000000b70000000000000097000000000000008100000000",
            INIT_36 => X"000000e500000000000000d600000000000000e000000000000000e000000000",
            INIT_37 => X"000000e000000000000000eb00000000000000de00000000000000db00000000",
            INIT_38 => X"0000008a00000000000000af00000000000000c600000000000000cd00000000",
            INIT_39 => X"000000cc00000000000000ce00000000000000cb00000000000000c000000000",
            INIT_3A => X"000000d200000000000000d000000000000000df00000000000000d400000000",
            INIT_3B => X"000000ce00000000000000c700000000000000d800000000000000d500000000",
            INIT_3C => X"0000005d0000000000000071000000000000009500000000000000b200000000",
            INIT_3D => X"0000004500000000000000500000000000000050000000000000005500000000",
            INIT_3E => X"000000de00000000000000ce00000000000000b7000000000000006c00000000",
            INIT_3F => X"000000d400000000000000dd00000000000000c500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000009a00000000000000a800000000000000ad00000000",
            INIT_41 => X"000000b300000000000000a000000000000000ac00000000000000a500000000",
            INIT_42 => X"000000c300000000000000bd00000000000000c200000000000000be00000000",
            INIT_43 => X"000000c600000000000000c100000000000000bf00000000000000c700000000",
            INIT_44 => X"0000006c000000000000006b0000000000000079000000000000009800000000",
            INIT_45 => X"0000004f000000000000006e0000000000000068000000000000006800000000",
            INIT_46 => X"000000af000000000000009f000000000000007a000000000000005200000000",
            INIT_47 => X"000000af00000000000000be000000000000009500000000000000a300000000",
            INIT_48 => X"0000006900000000000000720000000000000074000000000000007300000000",
            INIT_49 => X"0000007f0000000000000070000000000000006e000000000000006d00000000",
            INIT_4A => X"00000093000000000000008c0000000000000088000000000000008700000000",
            INIT_4B => X"000000a1000000000000009e000000000000008f000000000000009700000000",
            INIT_4C => X"0000007800000000000000780000000000000077000000000000008600000000",
            INIT_4D => X"0000005c0000000000000066000000000000006c000000000000006c00000000",
            INIT_4E => X"0000009100000000000000970000000000000080000000000000008f00000000",
            INIT_4F => X"000000780000000000000082000000000000006a000000000000006e00000000",
            INIT_50 => X"0000005200000000000000560000000000000057000000000000004e00000000",
            INIT_51 => X"0000006400000000000000610000000000000069000000000000006300000000",
            INIT_52 => X"0000006f000000000000006a000000000000006d000000000000006500000000",
            INIT_53 => X"0000007f00000000000000840000000000000076000000000000007200000000",
            INIT_54 => X"0000006b000000000000006e000000000000006d000000000000006d00000000",
            INIT_55 => X"00000077000000000000006c0000000000000057000000000000006000000000",
            INIT_56 => X"000000bf0000000000000090000000000000006f000000000000008400000000",
            INIT_57 => X"000000680000000000000066000000000000006f000000000000007800000000",
            INIT_58 => X"00000062000000000000005f0000000000000055000000000000004a00000000",
            INIT_59 => X"000000510000000000000062000000000000007a000000000000008000000000",
            INIT_5A => X"0000007300000000000000710000000000000081000000000000006800000000",
            INIT_5B => X"0000007b0000000000000086000000000000008b000000000000008400000000",
            INIT_5C => X"0000007700000000000000740000000000000073000000000000007800000000",
            INIT_5D => X"000000bd000000000000009e0000000000000068000000000000007100000000",
            INIT_5E => X"000000c5000000000000006d000000000000009400000000000000b700000000",
            INIT_5F => X"0000006300000000000000630000000000000067000000000000009500000000",
            INIT_60 => X"0000005d0000000000000071000000000000006b000000000000005100000000",
            INIT_61 => X"00000066000000000000005d0000000000000073000000000000007500000000",
            INIT_62 => X"0000008300000000000000950000000000000098000000000000008900000000",
            INIT_63 => X"00000071000000000000007d0000000000000088000000000000008200000000",
            INIT_64 => X"0000007b0000000000000072000000000000006c000000000000006c00000000",
            INIT_65 => X"000000c200000000000000af000000000000007f000000000000007600000000",
            INIT_66 => X"000000a2000000000000007600000000000000bd00000000000000ce00000000",
            INIT_67 => X"000000650000000000000062000000000000005000000000000000a700000000",
            INIT_68 => X"0000005d000000000000006a000000000000006e000000000000006100000000",
            INIT_69 => X"0000006400000000000000590000000000000054000000000000006200000000",
            INIT_6A => X"00000086000000000000008a000000000000007b000000000000006e00000000",
            INIT_6B => X"0000007c00000000000000820000000000000083000000000000007e00000000",
            INIT_6C => X"00000087000000000000007e000000000000007f000000000000007b00000000",
            INIT_6D => X"000000b400000000000000b50000000000000099000000000000008600000000",
            INIT_6E => X"0000007a000000000000009700000000000000b700000000000000b800000000",
            INIT_6F => X"000000590000000000000048000000000000004d00000000000000a000000000",
            INIT_70 => X"0000006100000000000000660000000000000065000000000000006600000000",
            INIT_71 => X"0000006b00000000000000580000000000000058000000000000005f00000000",
            INIT_72 => X"0000009e0000000000000097000000000000008e000000000000008200000000",
            INIT_73 => X"0000009d00000000000000a100000000000000a400000000000000a300000000",
            INIT_74 => X"000000a900000000000000aa00000000000000ad00000000000000ab00000000",
            INIT_75 => X"000000ae00000000000000b100000000000000a900000000000000a200000000",
            INIT_76 => X"0000006200000000000000a400000000000000a800000000000000b000000000",
            INIT_77 => X"0000004b000000000000003f0000000000000046000000000000005700000000",
            INIT_78 => X"0000007c000000000000007f0000000000000076000000000000007b00000000",
            INIT_79 => X"000000a000000000000000980000000000000094000000000000007e00000000",
            INIT_7A => X"000000b400000000000000b300000000000000af00000000000000a700000000",
            INIT_7B => X"000000ae00000000000000b900000000000000b800000000000000b700000000",
            INIT_7C => X"000000a000000000000000af00000000000000b200000000000000ad00000000",
            INIT_7D => X"000000a1000000000000008e0000000000000085000000000000008000000000",
            INIT_7E => X"0000006c00000000000000a600000000000000a200000000000000a900000000",
            INIT_7F => X"000000520000000000000059000000000000005f000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "sampleifmap_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000098000000000000008a000000000000007d000000000000008500000000",
            INIT_01 => X"000000a700000000000000a6000000000000009a000000000000009400000000",
            INIT_02 => X"000000b600000000000000b300000000000000ae00000000000000aa00000000",
            INIT_03 => X"000000ab00000000000000b500000000000000b900000000000000b900000000",
            INIT_04 => X"0000008b000000000000009a0000000000000098000000000000009800000000",
            INIT_05 => X"0000009b00000000000000900000000000000078000000000000006600000000",
            INIT_06 => X"0000008800000000000000a300000000000000a200000000000000a500000000",
            INIT_07 => X"0000006c000000000000009900000000000000bb000000000000009100000000",
            INIT_08 => X"00000083000000000000008d0000000000000085000000000000007c00000000",
            INIT_09 => X"000000aa00000000000000980000000000000072000000000000007400000000",
            INIT_0A => X"000000ad00000000000000b000000000000000af00000000000000af00000000",
            INIT_0B => X"00000097000000000000009a00000000000000a000000000000000a700000000",
            INIT_0C => X"000000a000000000000000a80000000000000096000000000000009000000000",
            INIT_0D => X"0000009e00000000000000a50000000000000098000000000000008c00000000",
            INIT_0E => X"00000097000000000000009c000000000000009b00000000000000a300000000",
            INIT_0F => X"000000930000000000000098000000000000009e000000000000009e00000000",
            INIT_10 => X"0000005d00000000000000600000000000000071000000000000008100000000",
            INIT_11 => X"000000a400000000000000940000000000000087000000000000006e00000000",
            INIT_12 => X"000000920000000000000096000000000000009f00000000000000a900000000",
            INIT_13 => X"000000a5000000000000009f0000000000000099000000000000009400000000",
            INIT_14 => X"000000ac00000000000000a800000000000000a000000000000000aa00000000",
            INIT_15 => X"000000a400000000000000a800000000000000a400000000000000a100000000",
            INIT_16 => X"00000092000000000000009e000000000000009e00000000000000a000000000",
            INIT_17 => X"00000096000000000000007d0000000000000079000000000000008400000000",
            INIT_18 => X"0000008700000000000000600000000000000055000000000000007000000000",
            INIT_19 => X"00000093000000000000009c00000000000000a5000000000000009b00000000",
            INIT_1A => X"000000a00000000000000097000000000000008d000000000000008e00000000",
            INIT_1B => X"000000ab00000000000000ae00000000000000ad00000000000000a700000000",
            INIT_1C => X"000000a800000000000000a2000000000000009b00000000000000a700000000",
            INIT_1D => X"000000a600000000000000a300000000000000a100000000000000a300000000",
            INIT_1E => X"0000006f00000000000000820000000000000097000000000000009e00000000",
            INIT_1F => X"0000008a000000000000005c0000000000000052000000000000006200000000",
            INIT_20 => X"0000008f00000000000000870000000000000084000000000000008500000000",
            INIT_21 => X"0000008e0000000000000096000000000000008f000000000000008f00000000",
            INIT_22 => X"000000ab00000000000000a900000000000000a1000000000000008a00000000",
            INIT_23 => X"00000086000000000000009700000000000000a500000000000000a900000000",
            INIT_24 => X"000000a40000000000000094000000000000006b000000000000007400000000",
            INIT_25 => X"00000098000000000000009f00000000000000a300000000000000a300000000",
            INIT_26 => X"0000005b0000000000000066000000000000006c000000000000008000000000",
            INIT_27 => X"000000480000000000000050000000000000004e000000000000004b00000000",
            INIT_28 => X"0000008f0000000000000090000000000000008c000000000000008400000000",
            INIT_29 => X"0000009600000000000000970000000000000093000000000000009000000000",
            INIT_2A => X"0000009a00000000000000940000000000000092000000000000008b00000000",
            INIT_2B => X"0000004e000000000000006e000000000000009c000000000000009f00000000",
            INIT_2C => X"000000a30000000000000084000000000000004a000000000000004b00000000",
            INIT_2D => X"0000006d000000000000007e000000000000008f000000000000009900000000",
            INIT_2E => X"0000004c000000000000005a0000000000000064000000000000006700000000",
            INIT_2F => X"0000002100000000000000390000000000000052000000000000004b00000000",
            INIT_30 => X"0000009200000000000000940000000000000089000000000000005e00000000",
            INIT_31 => X"0000007300000000000000810000000000000091000000000000009200000000",
            INIT_32 => X"0000008700000000000000630000000000000066000000000000006a00000000",
            INIT_33 => X"0000005d0000000000000072000000000000009a000000000000009d00000000",
            INIT_34 => X"0000007c000000000000007d0000000000000068000000000000006500000000",
            INIT_35 => X"000000650000000000000066000000000000006a000000000000007100000000",
            INIT_36 => X"0000003f0000000000000045000000000000004f000000000000005800000000",
            INIT_37 => X"0000001f00000000000000250000000000000035000000000000004300000000",
            INIT_38 => X"000000860000000000000086000000000000007d000000000000005600000000",
            INIT_39 => X"0000004d000000000000005c0000000000000085000000000000008900000000",
            INIT_3A => X"00000083000000000000005c0000000000000059000000000000005200000000",
            INIT_3B => X"0000007300000000000000840000000000000096000000000000009900000000",
            INIT_3C => X"0000006100000000000000600000000000000061000000000000006a00000000",
            INIT_3D => X"0000004f000000000000005f0000000000000065000000000000006300000000",
            INIT_3E => X"00000039000000000000003c0000000000000040000000000000003c00000000",
            INIT_3F => X"0000001f00000000000000220000000000000026000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008300000000000000810000000000000074000000000000005a00000000",
            INIT_41 => X"00000061000000000000006a000000000000008a000000000000008900000000",
            INIT_42 => X"0000007e000000000000007c0000000000000074000000000000006c00000000",
            INIT_43 => X"000000530000000000000054000000000000005f000000000000007100000000",
            INIT_44 => X"000000640000000000000062000000000000005c000000000000005900000000",
            INIT_45 => X"000000450000000000000043000000000000004a000000000000005c00000000",
            INIT_46 => X"0000002e00000000000000330000000000000042000000000000004a00000000",
            INIT_47 => X"0000002000000000000000230000000000000026000000000000002b00000000",
            INIT_48 => X"0000007f00000000000000820000000000000070000000000000005c00000000",
            INIT_49 => X"00000066000000000000006e0000000000000078000000000000007c00000000",
            INIT_4A => X"0000004c0000000000000050000000000000005a000000000000006100000000",
            INIT_4B => X"0000005b00000000000000540000000000000050000000000000004b00000000",
            INIT_4C => X"0000004900000000000000510000000000000059000000000000005f00000000",
            INIT_4D => X"0000003d00000000000000430000000000000041000000000000004100000000",
            INIT_4E => X"00000028000000000000002a000000000000003a000000000000004500000000",
            INIT_4F => X"0000002500000000000000230000000000000028000000000000002a00000000",
            INIT_50 => X"0000004e0000000000000056000000000000004f000000000000004c00000000",
            INIT_51 => X"0000003f00000000000000400000000000000045000000000000004a00000000",
            INIT_52 => X"0000004d000000000000004a0000000000000046000000000000004100000000",
            INIT_53 => X"0000005000000000000000510000000000000052000000000000005100000000",
            INIT_54 => X"000000440000000000000037000000000000003b000000000000004900000000",
            INIT_55 => X"000000320000000000000036000000000000003f000000000000004300000000",
            INIT_56 => X"000000280000000000000028000000000000002d000000000000003600000000",
            INIT_57 => X"0000002500000000000000270000000000000028000000000000002900000000",
            INIT_58 => X"0000002a0000000000000028000000000000002b000000000000002d00000000",
            INIT_59 => X"0000003a00000000000000350000000000000034000000000000003100000000",
            INIT_5A => X"0000004600000000000000480000000000000047000000000000004400000000",
            INIT_5B => X"0000003b000000000000003a000000000000003b000000000000004100000000",
            INIT_5C => X"000000490000000000000055000000000000003f000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000033000000000000003900000000",
            INIT_5E => X"0000002800000000000000270000000000000028000000000000002c00000000",
            INIT_5F => X"0000001d000000000000002a000000000000002a000000000000002900000000",
            INIT_60 => X"0000002600000000000000240000000000000028000000000000002b00000000",
            INIT_61 => X"0000003200000000000000310000000000000030000000000000002c00000000",
            INIT_62 => X"0000003100000000000000310000000000000034000000000000003500000000",
            INIT_63 => X"0000003d000000000000003e000000000000003b000000000000003500000000",
            INIT_64 => X"00000042000000000000005e0000000000000045000000000000003700000000",
            INIT_65 => X"00000028000000000000002f000000000000002e000000000000002c00000000",
            INIT_66 => X"0000002a00000000000000280000000000000027000000000000002700000000",
            INIT_67 => X"000000120000000000000020000000000000002e000000000000002900000000",
            INIT_68 => X"0000002400000000000000230000000000000027000000000000002800000000",
            INIT_69 => X"0000002b00000000000000290000000000000029000000000000002700000000",
            INIT_6A => X"0000003a00000000000000380000000000000033000000000000002e00000000",
            INIT_6B => X"00000037000000000000003c000000000000003d000000000000003d00000000",
            INIT_6C => X"000000360000000000000055000000000000003c000000000000002e00000000",
            INIT_6D => X"000000240000000000000025000000000000002e000000000000002800000000",
            INIT_6E => X"0000002a00000000000000280000000000000026000000000000002600000000",
            INIT_6F => X"00000007000000000000000d0000000000000028000000000000002b00000000",
            INIT_70 => X"0000002800000000000000240000000000000026000000000000002200000000",
            INIT_71 => X"000000330000000000000031000000000000002f000000000000002c00000000",
            INIT_72 => X"00000039000000000000003b0000000000000039000000000000003600000000",
            INIT_73 => X"0000002b00000000000000330000000000000037000000000000003900000000",
            INIT_74 => X"00000032000000000000004e0000000000000030000000000000001f00000000",
            INIT_75 => X"0000002300000000000000230000000000000025000000000000002900000000",
            INIT_76 => X"0000002900000000000000240000000000000025000000000000002500000000",
            INIT_77 => X"0000000700000000000000060000000000000014000000000000002d00000000",
            INIT_78 => X"0000002f000000000000002d000000000000002b000000000000002900000000",
            INIT_79 => X"0000003100000000000000300000000000000030000000000000003000000000",
            INIT_7A => X"0000002d00000000000000310000000000000033000000000000003200000000",
            INIT_7B => X"00000011000000000000001a0000000000000022000000000000002800000000",
            INIT_7C => X"0000002c000000000000003f000000000000001b000000000000000800000000",
            INIT_7D => X"0000002300000000000000220000000000000022000000000000002100000000",
            INIT_7E => X"0000002c00000000000000220000000000000022000000000000002300000000",
            INIT_7F => X"0000000800000000000000050000000000000006000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "sampleifmap_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ba00000000000000c200000000000000da00000000000000de00000000",
            INIT_01 => X"000000f100000000000000ee00000000000000ec00000000000000de00000000",
            INIT_02 => X"000000eb00000000000000f400000000000000f500000000000000f300000000",
            INIT_03 => X"000000f500000000000000f200000000000000f100000000000000f000000000",
            INIT_04 => X"000000f800000000000000f500000000000000f000000000000000e300000000",
            INIT_05 => X"000000f300000000000000f300000000000000f300000000000000f900000000",
            INIT_06 => X"000000f700000000000000ef00000000000000eb00000000000000f500000000",
            INIT_07 => X"000000f600000000000000f300000000000000ea00000000000000f100000000",
            INIT_08 => X"000000b800000000000000c900000000000000e200000000000000e500000000",
            INIT_09 => X"000000ee00000000000000f000000000000000f000000000000000df00000000",
            INIT_0A => X"000000e800000000000000f500000000000000f700000000000000f300000000",
            INIT_0B => X"000000f800000000000000f500000000000000f500000000000000f300000000",
            INIT_0C => X"000000fb00000000000000f300000000000000ef00000000000000e600000000",
            INIT_0D => X"000000f400000000000000ee00000000000000ee00000000000000fb00000000",
            INIT_0E => X"000000fc00000000000000f300000000000000ec00000000000000f800000000",
            INIT_0F => X"000000fb00000000000000fa00000000000000ec00000000000000f000000000",
            INIT_10 => X"000000b500000000000000c700000000000000de00000000000000e100000000",
            INIT_11 => X"000000e400000000000000ef00000000000000ee00000000000000db00000000",
            INIT_12 => X"000000e400000000000000ec00000000000000f400000000000000eb00000000",
            INIT_13 => X"000000f700000000000000ee00000000000000ef00000000000000eb00000000",
            INIT_14 => X"000000f600000000000000f100000000000000ec00000000000000e500000000",
            INIT_15 => X"000000ef00000000000000e800000000000000d700000000000000ec00000000",
            INIT_16 => X"000000fc00000000000000f200000000000000eb00000000000000f800000000",
            INIT_17 => X"000000f700000000000000fb00000000000000e800000000000000f100000000",
            INIT_18 => X"000000b300000000000000c200000000000000d800000000000000de00000000",
            INIT_19 => X"000000e100000000000000eb00000000000000e400000000000000d600000000",
            INIT_1A => X"000000dd00000000000000e600000000000000ef00000000000000e500000000",
            INIT_1B => X"000000f700000000000000e600000000000000ec00000000000000e100000000",
            INIT_1C => X"000000ee00000000000000f000000000000000ea00000000000000e600000000",
            INIT_1D => X"000000f100000000000000e500000000000000b000000000000000ba00000000",
            INIT_1E => X"000000fb00000000000000ef00000000000000e900000000000000f800000000",
            INIT_1F => X"000000f300000000000000f800000000000000e400000000000000ee00000000",
            INIT_20 => X"000000ac00000000000000c100000000000000d900000000000000df00000000",
            INIT_21 => X"000000d900000000000000e700000000000000dd00000000000000d200000000",
            INIT_22 => X"000000d700000000000000e100000000000000eb00000000000000da00000000",
            INIT_23 => X"000000ee00000000000000d600000000000000e800000000000000db00000000",
            INIT_24 => X"000000e400000000000000ee00000000000000e300000000000000e500000000",
            INIT_25 => X"000000ef00000000000000e500000000000000b200000000000000b000000000",
            INIT_26 => X"000000f500000000000000ea00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f000000000000000f600000000000000e800000000000000e700000000",
            INIT_28 => X"000000a400000000000000bf00000000000000d500000000000000dc00000000",
            INIT_29 => X"000000d500000000000000e100000000000000d500000000000000ce00000000",
            INIT_2A => X"000000d600000000000000da00000000000000e600000000000000d600000000",
            INIT_2B => X"000000ce00000000000000c800000000000000e300000000000000d600000000",
            INIT_2C => X"000000cf00000000000000ed00000000000000ce00000000000000d000000000",
            INIT_2D => X"000000e900000000000000e600000000000000ad000000000000008200000000",
            INIT_2E => X"000000e800000000000000db00000000000000e100000000000000f400000000",
            INIT_2F => X"000000e600000000000000f200000000000000e700000000000000dd00000000",
            INIT_30 => X"0000009600000000000000b900000000000000ca00000000000000d400000000",
            INIT_31 => X"000000d000000000000000d900000000000000c900000000000000c400000000",
            INIT_32 => X"000000d300000000000000d000000000000000db00000000000000d300000000",
            INIT_33 => X"000000af00000000000000b900000000000000dd00000000000000d400000000",
            INIT_34 => X"000000c500000000000000d200000000000000bd00000000000000bb00000000",
            INIT_35 => X"000000bb00000000000000b8000000000000009d000000000000008900000000",
            INIT_36 => X"000000da00000000000000ce00000000000000dc00000000000000dd00000000",
            INIT_37 => X"000000d800000000000000e700000000000000db00000000000000d100000000",
            INIT_38 => X"0000009300000000000000b300000000000000c900000000000000d300000000",
            INIT_39 => X"000000cb00000000000000ce00000000000000cc00000000000000c500000000",
            INIT_3A => X"000000cd00000000000000c600000000000000d200000000000000d000000000",
            INIT_3B => X"000000cb00000000000000c000000000000000ce00000000000000ce00000000",
            INIT_3C => X"0000006a000000000000007a000000000000009b00000000000000b300000000",
            INIT_3D => X"000000490000000000000058000000000000005e000000000000006400000000",
            INIT_3E => X"000000d700000000000000ca00000000000000b7000000000000006f00000000",
            INIT_3F => X"000000c100000000000000ce00000000000000b900000000000000c600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000a000000000000000ad00000000000000b300000000",
            INIT_41 => X"000000b300000000000000a100000000000000af00000000000000aa00000000",
            INIT_42 => X"000000bd00000000000000b400000000000000b800000000000000bb00000000",
            INIT_43 => X"000000c400000000000000ba00000000000000b900000000000000c300000000",
            INIT_44 => X"0000008000000000000000800000000000000089000000000000009f00000000",
            INIT_45 => X"0000005a0000000000000080000000000000007e000000000000007e00000000",
            INIT_46 => X"000000ac000000000000009e000000000000007c000000000000005800000000",
            INIT_47 => X"0000009f00000000000000b00000000000000089000000000000009c00000000",
            INIT_48 => X"00000070000000000000007b000000000000007e000000000000007b00000000",
            INIT_49 => X"0000008000000000000000720000000000000072000000000000007200000000",
            INIT_4A => X"0000009000000000000000890000000000000086000000000000008600000000",
            INIT_4B => X"000000a700000000000000a00000000000000092000000000000009800000000",
            INIT_4C => X"0000008c0000000000000090000000000000008b000000000000009300000000",
            INIT_4D => X"0000006800000000000000780000000000000083000000000000008200000000",
            INIT_4E => X"0000008d00000000000000960000000000000083000000000000009500000000",
            INIT_4F => X"0000007500000000000000800000000000000069000000000000006a00000000",
            INIT_50 => X"0000005800000000000000620000000000000066000000000000005900000000",
            INIT_51 => X"0000006a00000000000000680000000000000073000000000000006b00000000",
            INIT_52 => X"0000007300000000000000710000000000000076000000000000006b00000000",
            INIT_53 => X"0000009200000000000000970000000000000086000000000000007b00000000",
            INIT_54 => X"00000078000000000000007f000000000000007f000000000000008000000000",
            INIT_55 => X"00000080000000000000007a0000000000000068000000000000006f00000000",
            INIT_56 => X"000000b6000000000000008b000000000000006e000000000000008600000000",
            INIT_57 => X"00000070000000000000006d0000000000000075000000000000007200000000",
            INIT_58 => X"0000006a000000000000006e0000000000000068000000000000005800000000",
            INIT_59 => X"0000005e00000000000000710000000000000089000000000000008e00000000",
            INIT_5A => X"0000007d000000000000007f0000000000000092000000000000007400000000",
            INIT_5B => X"0000009700000000000000a500000000000000a5000000000000009400000000",
            INIT_5C => X"0000007f000000000000007f0000000000000082000000000000008e00000000",
            INIT_5D => X"000000bf00000000000000a50000000000000072000000000000007b00000000",
            INIT_5E => X"000000b80000000000000064000000000000008e00000000000000b400000000",
            INIT_5F => X"0000006c000000000000006c000000000000006d000000000000008c00000000",
            INIT_60 => X"0000006800000000000000840000000000000082000000000000006400000000",
            INIT_61 => X"00000076000000000000006d0000000000000082000000000000008100000000",
            INIT_62 => X"0000009700000000000000a800000000000000ab000000000000009a00000000",
            INIT_63 => X"0000008b000000000000009a00000000000000a5000000000000009b00000000",
            INIT_64 => X"0000008c0000000000000081000000000000007d000000000000008200000000",
            INIT_65 => X"000000c100000000000000b30000000000000089000000000000008600000000",
            INIT_66 => X"00000098000000000000007000000000000000b900000000000000cb00000000",
            INIT_67 => X"0000006d0000000000000069000000000000005400000000000000a000000000",
            INIT_68 => X"0000006a000000000000007e0000000000000086000000000000007800000000",
            INIT_69 => X"00000079000000000000006c0000000000000065000000000000007100000000",
            INIT_6A => X"0000009f00000000000000a10000000000000091000000000000008300000000",
            INIT_6B => X"00000095000000000000009e00000000000000a1000000000000009900000000",
            INIT_6C => X"0000009b00000000000000910000000000000093000000000000009200000000",
            INIT_6D => X"000000b100000000000000b600000000000000a1000000000000009600000000",
            INIT_6E => X"00000076000000000000009400000000000000b500000000000000b500000000",
            INIT_6F => X"00000060000000000000004e0000000000000050000000000000009d00000000",
            INIT_70 => X"00000072000000000000007d0000000000000080000000000000007f00000000",
            INIT_71 => X"0000008600000000000000730000000000000071000000000000007400000000",
            INIT_72 => X"000000b800000000000000b000000000000000a8000000000000009f00000000",
            INIT_73 => X"000000b900000000000000be00000000000000bf00000000000000be00000000",
            INIT_74 => X"000000b800000000000000be00000000000000c400000000000000c500000000",
            INIT_75 => X"000000a800000000000000af00000000000000ad00000000000000ac00000000",
            INIT_76 => X"0000006300000000000000a300000000000000a500000000000000ab00000000",
            INIT_77 => X"0000005100000000000000430000000000000047000000000000005700000000",
            INIT_78 => X"00000091000000000000009a0000000000000095000000000000009700000000",
            INIT_79 => X"000000c100000000000000b800000000000000b3000000000000009900000000",
            INIT_7A => X"000000d000000000000000cf00000000000000cd00000000000000c900000000",
            INIT_7B => X"000000c800000000000000d400000000000000d200000000000000d100000000",
            INIT_7C => X"000000ab00000000000000c300000000000000c900000000000000c600000000",
            INIT_7D => X"0000009b000000000000008b0000000000000087000000000000008600000000",
            INIT_7E => X"0000007100000000000000a800000000000000a100000000000000a500000000",
            INIT_7F => X"00000056000000000000005a000000000000005c000000000000004900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "sampleifmap_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b000000000000000a7000000000000009f00000000000000a500000000",
            INIT_01 => X"000000c900000000000000c600000000000000b900000000000000af00000000",
            INIT_02 => X"000000d200000000000000d200000000000000d000000000000000cd00000000",
            INIT_03 => X"000000be00000000000000c900000000000000d000000000000000d200000000",
            INIT_04 => X"0000009400000000000000a900000000000000aa00000000000000aa00000000",
            INIT_05 => X"00000099000000000000008e000000000000007a000000000000006c00000000",
            INIT_06 => X"0000008e00000000000000a700000000000000a500000000000000a700000000",
            INIT_07 => X"0000006f000000000000009800000000000000b5000000000000009300000000",
            INIT_08 => X"0000009d00000000000000ae00000000000000aa000000000000009d00000000",
            INIT_09 => X"000000ca00000000000000b6000000000000008f000000000000008d00000000",
            INIT_0A => X"000000ca00000000000000d100000000000000d300000000000000d000000000",
            INIT_0B => X"000000a200000000000000a700000000000000b500000000000000bf00000000",
            INIT_0C => X"000000a900000000000000b200000000000000a0000000000000009b00000000",
            INIT_0D => X"000000a000000000000000a7000000000000009d000000000000009300000000",
            INIT_0E => X"0000009c00000000000000a100000000000000a200000000000000a900000000",
            INIT_0F => X"0000009400000000000000960000000000000096000000000000009e00000000",
            INIT_10 => X"000000790000000000000080000000000000009400000000000000a200000000",
            INIT_11 => X"000000c200000000000000b100000000000000a4000000000000008a00000000",
            INIT_12 => X"000000ab00000000000000b200000000000000bc00000000000000c700000000",
            INIT_13 => X"000000b000000000000000ac00000000000000ac00000000000000aa00000000",
            INIT_14 => X"000000b500000000000000b000000000000000a800000000000000b400000000",
            INIT_15 => X"000000ac00000000000000af00000000000000ad00000000000000aa00000000",
            INIT_16 => X"0000009600000000000000a300000000000000a500000000000000a800000000",
            INIT_17 => X"00000099000000000000007d0000000000000076000000000000008500000000",
            INIT_18 => X"000000a6000000000000007f0000000000000075000000000000008f00000000",
            INIT_19 => X"000000b000000000000000ba00000000000000c500000000000000bc00000000",
            INIT_1A => X"000000b200000000000000ab00000000000000a300000000000000a900000000",
            INIT_1B => X"000000ba00000000000000bf00000000000000be00000000000000b900000000",
            INIT_1C => X"000000b100000000000000ac00000000000000a500000000000000b400000000",
            INIT_1D => X"000000b200000000000000af00000000000000ac00000000000000ad00000000",
            INIT_1E => X"000000740000000000000088000000000000009c00000000000000a400000000",
            INIT_1F => X"0000009000000000000000620000000000000057000000000000006700000000",
            INIT_20 => X"000000b000000000000000a800000000000000a500000000000000a600000000",
            INIT_21 => X"000000aa00000000000000b300000000000000ae00000000000000b000000000",
            INIT_22 => X"000000bd00000000000000be00000000000000b800000000000000a400000000",
            INIT_23 => X"0000009600000000000000a800000000000000b500000000000000b900000000",
            INIT_24 => X"000000ad000000000000009d0000000000000076000000000000008100000000",
            INIT_25 => X"000000a200000000000000ab00000000000000ad00000000000000ad00000000",
            INIT_26 => X"0000005f000000000000006a0000000000000070000000000000008500000000",
            INIT_27 => X"0000004e00000000000000560000000000000054000000000000005000000000",
            INIT_28 => X"000000af00000000000000b100000000000000ac00000000000000a500000000",
            INIT_29 => X"000000b000000000000000b300000000000000b000000000000000ae00000000",
            INIT_2A => X"000000ad00000000000000ab00000000000000ab00000000000000a400000000",
            INIT_2B => X"0000005e000000000000007e00000000000000ab00000000000000af00000000",
            INIT_2C => X"000000ac000000000000008e0000000000000055000000000000005800000000",
            INIT_2D => X"000000750000000000000088000000000000009800000000000000a200000000",
            INIT_2E => X"00000050000000000000005e0000000000000068000000000000006c00000000",
            INIT_2F => X"00000027000000000000003f0000000000000058000000000000004f00000000",
            INIT_30 => X"000000af00000000000000b200000000000000a6000000000000007c00000000",
            INIT_31 => X"0000008b000000000000009a00000000000000ad00000000000000af00000000",
            INIT_32 => X"0000009a000000000000007a000000000000007e000000000000008200000000",
            INIT_33 => X"0000006c000000000000008300000000000000a900000000000000ae00000000",
            INIT_34 => X"0000008500000000000000860000000000000072000000000000007200000000",
            INIT_35 => X"0000006c000000000000006d0000000000000071000000000000007900000000",
            INIT_36 => X"00000045000000000000004b0000000000000056000000000000005f00000000",
            INIT_37 => X"00000026000000000000002b000000000000003b000000000000004900000000",
            INIT_38 => X"0000009f00000000000000a00000000000000096000000000000006f00000000",
            INIT_39 => X"000000640000000000000074000000000000009e00000000000000a300000000",
            INIT_3A => X"0000009700000000000000730000000000000070000000000000006800000000",
            INIT_3B => X"00000083000000000000009500000000000000a800000000000000ac00000000",
            INIT_3C => X"0000006a000000000000006a000000000000006b000000000000007700000000",
            INIT_3D => X"000000540000000000000064000000000000006c000000000000006a00000000",
            INIT_3E => X"0000004100000000000000440000000000000049000000000000004500000000",
            INIT_3F => X"000000250000000000000028000000000000002c000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009a0000000000000097000000000000008a000000000000007100000000",
            INIT_41 => X"00000077000000000000008000000000000000a200000000000000a100000000",
            INIT_42 => X"0000009200000000000000900000000000000088000000000000008100000000",
            INIT_43 => X"0000006200000000000000650000000000000072000000000000008400000000",
            INIT_44 => X"0000006c000000000000006d0000000000000067000000000000006500000000",
            INIT_45 => X"0000004b00000000000000480000000000000050000000000000006300000000",
            INIT_46 => X"0000003a000000000000003d000000000000004d000000000000005500000000",
            INIT_47 => X"000000270000000000000029000000000000002d000000000000003400000000",
            INIT_48 => X"00000097000000000000009a0000000000000088000000000000007400000000",
            INIT_49 => X"0000007c0000000000000084000000000000008f000000000000009400000000",
            INIT_4A => X"00000057000000000000005b0000000000000067000000000000007600000000",
            INIT_4B => X"000000650000000000000063000000000000005b000000000000005600000000",
            INIT_4C => X"00000052000000000000005e0000000000000063000000000000006500000000",
            INIT_4D => X"00000045000000000000004a0000000000000048000000000000004800000000",
            INIT_4E => X"0000003200000000000000340000000000000044000000000000004e00000000",
            INIT_4F => X"00000030000000000000002f0000000000000030000000000000003300000000",
            INIT_50 => X"00000063000000000000006a0000000000000064000000000000006000000000",
            INIT_51 => X"0000005100000000000000520000000000000056000000000000005c00000000",
            INIT_52 => X"000000540000000000000051000000000000004f000000000000005200000000",
            INIT_53 => X"00000058000000000000005e000000000000005b000000000000005700000000",
            INIT_54 => X"0000004c00000000000000440000000000000044000000000000004d00000000",
            INIT_55 => X"0000003b00000000000000400000000000000048000000000000004a00000000",
            INIT_56 => X"0000003200000000000000310000000000000036000000000000003f00000000",
            INIT_57 => X"0000003000000000000000340000000000000030000000000000003100000000",
            INIT_58 => X"0000003700000000000000360000000000000039000000000000003b00000000",
            INIT_59 => X"00000044000000000000003e000000000000003d000000000000003c00000000",
            INIT_5A => X"0000004d000000000000004f000000000000004f000000000000004e00000000",
            INIT_5B => X"0000004200000000000000450000000000000044000000000000004800000000",
            INIT_5C => X"0000005200000000000000610000000000000047000000000000003d00000000",
            INIT_5D => X"000000390000000000000038000000000000003c000000000000004100000000",
            INIT_5E => X"0000003100000000000000300000000000000031000000000000003500000000",
            INIT_5F => X"0000002300000000000000320000000000000032000000000000003200000000",
            INIT_60 => X"0000002d000000000000002c0000000000000030000000000000003200000000",
            INIT_61 => X"0000003700000000000000350000000000000035000000000000003100000000",
            INIT_62 => X"000000380000000000000038000000000000003b000000000000003a00000000",
            INIT_63 => X"0000004400000000000000470000000000000042000000000000003c00000000",
            INIT_64 => X"0000004b0000000000000068000000000000004b000000000000003b00000000",
            INIT_65 => X"00000033000000000000003a0000000000000038000000000000003500000000",
            INIT_66 => X"0000003300000000000000310000000000000030000000000000003100000000",
            INIT_67 => X"0000001400000000000000250000000000000035000000000000003200000000",
            INIT_68 => X"000000290000000000000028000000000000002c000000000000002d00000000",
            INIT_69 => X"00000030000000000000002e000000000000002e000000000000002c00000000",
            INIT_6A => X"00000041000000000000003f0000000000000039000000000000003300000000",
            INIT_6B => X"0000003d00000000000000440000000000000044000000000000004400000000",
            INIT_6C => X"0000003f000000000000005d0000000000000042000000000000003200000000",
            INIT_6D => X"0000002f00000000000000300000000000000038000000000000003100000000",
            INIT_6E => X"000000330000000000000031000000000000002f000000000000002f00000000",
            INIT_6F => X"00000005000000000000000e000000000000002e000000000000003400000000",
            INIT_70 => X"0000002d0000000000000029000000000000002b000000000000002700000000",
            INIT_71 => X"0000003b00000000000000380000000000000036000000000000003200000000",
            INIT_72 => X"0000004000000000000000420000000000000040000000000000003e00000000",
            INIT_73 => X"00000031000000000000003a000000000000003d000000000000004000000000",
            INIT_74 => X"0000003b00000000000000550000000000000035000000000000002400000000",
            INIT_75 => X"0000002f000000000000002f0000000000000030000000000000003200000000",
            INIT_76 => X"00000032000000000000002d000000000000002e000000000000002e00000000",
            INIT_77 => X"0000000300000000000000030000000000000018000000000000003600000000",
            INIT_78 => X"0000003600000000000000340000000000000032000000000000002f00000000",
            INIT_79 => X"0000003a00000000000000380000000000000038000000000000003800000000",
            INIT_7A => X"0000003200000000000000350000000000000037000000000000003a00000000",
            INIT_7B => X"00000014000000000000001e0000000000000027000000000000002d00000000",
            INIT_7C => X"0000003600000000000000480000000000000021000000000000000b00000000",
            INIT_7D => X"0000002e000000000000002d000000000000002d000000000000002c00000000",
            INIT_7E => X"00000034000000000000002b000000000000002c000000000000002c00000000",
            INIT_7F => X"0000000700000000000000030000000000000008000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "sampleifmap_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be00000000000000b000000000000000a7000000000000009b00000000",
            INIT_01 => X"000000a600000000000000a800000000000000a600000000000000b100000000",
            INIT_02 => X"000000bb00000000000000bb00000000000000b300000000000000aa00000000",
            INIT_03 => X"000000b800000000000000b800000000000000bb00000000000000bb00000000",
            INIT_04 => X"000000ba00000000000000b800000000000000b400000000000000b600000000",
            INIT_05 => X"000000bd00000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000c000000000000000ca00000000000000c900000000000000c900000000",
            INIT_08 => X"000000bb00000000000000ab00000000000000a3000000000000009900000000",
            INIT_09 => X"0000009f000000000000009a000000000000009b00000000000000b300000000",
            INIT_0A => X"000000af00000000000000ab00000000000000a5000000000000009f00000000",
            INIT_0B => X"000000a500000000000000a200000000000000ab00000000000000a900000000",
            INIT_0C => X"000000a500000000000000a600000000000000a400000000000000aa00000000",
            INIT_0D => X"000000a800000000000000a900000000000000ad00000000000000a700000000",
            INIT_0E => X"000000ca00000000000000be00000000000000ad00000000000000a900000000",
            INIT_0F => X"000000bd00000000000000cb00000000000000ca00000000000000cc00000000",
            INIT_10 => X"000000b800000000000000a800000000000000a0000000000000009b00000000",
            INIT_11 => X"000000bc00000000000000b000000000000000ae00000000000000bb00000000",
            INIT_12 => X"000000be00000000000000b100000000000000b300000000000000b600000000",
            INIT_13 => X"000000b900000000000000bc00000000000000c200000000000000c000000000",
            INIT_14 => X"000000c200000000000000c100000000000000c200000000000000c100000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c500000000000000c300000000",
            INIT_16 => X"000000cf00000000000000ce00000000000000c500000000000000bf00000000",
            INIT_17 => X"000000bd00000000000000cc00000000000000ce00000000000000d000000000",
            INIT_18 => X"000000b100000000000000a6000000000000009d000000000000009700000000",
            INIT_19 => X"000000c500000000000000c700000000000000b900000000000000b400000000",
            INIT_1A => X"000000c600000000000000cd00000000000000cc00000000000000b600000000",
            INIT_1B => X"000000cb00000000000000c400000000000000c500000000000000d200000000",
            INIT_1C => X"000000cb00000000000000d200000000000000cf00000000000000cd00000000",
            INIT_1D => X"000000cc00000000000000c500000000000000d200000000000000cf00000000",
            INIT_1E => X"000000c900000000000000cc00000000000000c600000000000000d000000000",
            INIT_1F => X"000000c000000000000000ce00000000000000cf00000000000000d100000000",
            INIT_20 => X"000000ae00000000000000a8000000000000009e000000000000009700000000",
            INIT_21 => X"000000c400000000000000bf00000000000000b500000000000000b100000000",
            INIT_22 => X"000000b900000000000000bd00000000000000c200000000000000b700000000",
            INIT_23 => X"000000ca00000000000000b900000000000000b900000000000000c400000000",
            INIT_24 => X"000000c000000000000000c800000000000000c700000000000000c700000000",
            INIT_25 => X"000000bc00000000000000be00000000000000c700000000000000c300000000",
            INIT_26 => X"000000c400000000000000c900000000000000c700000000000000c900000000",
            INIT_27 => X"000000c400000000000000cf00000000000000cc00000000000000ce00000000",
            INIT_28 => X"000000ae00000000000000a7000000000000009c000000000000009400000000",
            INIT_29 => X"000000c300000000000000c400000000000000ae00000000000000ab00000000",
            INIT_2A => X"000000b800000000000000bd00000000000000be00000000000000c000000000",
            INIT_2B => X"000000bf00000000000000bd00000000000000bd00000000000000bb00000000",
            INIT_2C => X"000000c600000000000000bb00000000000000c300000000000000be00000000",
            INIT_2D => X"000000c100000000000000c000000000000000bc00000000000000c000000000",
            INIT_2E => X"000000d100000000000000cb00000000000000ce00000000000000cd00000000",
            INIT_2F => X"000000c400000000000000d100000000000000d000000000000000d400000000",
            INIT_30 => X"000000ae00000000000000a50000000000000099000000000000009400000000",
            INIT_31 => X"000000c300000000000000cb00000000000000b000000000000000a800000000",
            INIT_32 => X"000000be00000000000000bb00000000000000bc00000000000000bc00000000",
            INIT_33 => X"000000c300000000000000c500000000000000c200000000000000b600000000",
            INIT_34 => X"000000cd00000000000000c800000000000000c100000000000000c400000000",
            INIT_35 => X"000000c900000000000000c500000000000000c500000000000000c600000000",
            INIT_36 => X"000000c300000000000000c600000000000000c800000000000000c500000000",
            INIT_37 => X"000000c300000000000000cf00000000000000cb00000000000000c500000000",
            INIT_38 => X"000000ac00000000000000a3000000000000009b000000000000009900000000",
            INIT_39 => X"000000d100000000000000c700000000000000bc00000000000000ac00000000",
            INIT_3A => X"000000bf00000000000000bd00000000000000be00000000000000c400000000",
            INIT_3B => X"000000c400000000000000bb00000000000000bc00000000000000c100000000",
            INIT_3C => X"000000ce00000000000000c400000000000000c200000000000000ca00000000",
            INIT_3D => X"000000c800000000000000c400000000000000c900000000000000c200000000",
            INIT_3E => X"000000c900000000000000c800000000000000bb00000000000000b500000000",
            INIT_3F => X"000000bd00000000000000c700000000000000c400000000000000c800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000a3000000000000009f00000000000000a000000000",
            INIT_41 => X"000000be00000000000000b000000000000000b000000000000000ae00000000",
            INIT_42 => X"000000b000000000000000b000000000000000af00000000000000b400000000",
            INIT_43 => X"000000b600000000000000ac00000000000000aa00000000000000b500000000",
            INIT_44 => X"000000bb00000000000000b500000000000000b200000000000000bb00000000",
            INIT_45 => X"000000bb00000000000000b400000000000000bc00000000000000b100000000",
            INIT_46 => X"000000bc00000000000000bc00000000000000c400000000000000c700000000",
            INIT_47 => X"000000b800000000000000c200000000000000c000000000000000c500000000",
            INIT_48 => X"000000ac00000000000000a200000000000000a700000000000000ab00000000",
            INIT_49 => X"000000b000000000000000b400000000000000ab00000000000000aa00000000",
            INIT_4A => X"0000009c0000000000000096000000000000009c000000000000009b00000000",
            INIT_4B => X"0000009e00000000000000990000000000000092000000000000009600000000",
            INIT_4C => X"0000009d00000000000000a400000000000000a600000000000000a600000000",
            INIT_4D => X"000000a6000000000000009c00000000000000a2000000000000009d00000000",
            INIT_4E => X"000000bd00000000000000bc00000000000000c700000000000000c800000000",
            INIT_4F => X"000000b600000000000000c200000000000000c100000000000000c500000000",
            INIT_50 => X"000000b000000000000000a800000000000000b400000000000000af00000000",
            INIT_51 => X"000000ae00000000000000b600000000000000b100000000000000ad00000000",
            INIT_52 => X"0000009a000000000000009f00000000000000a0000000000000009c00000000",
            INIT_53 => X"000000ad00000000000000a800000000000000a3000000000000009f00000000",
            INIT_54 => X"000000a200000000000000a000000000000000a400000000000000aa00000000",
            INIT_55 => X"000000ac00000000000000a700000000000000a800000000000000a000000000",
            INIT_56 => X"000000c400000000000000c400000000000000c300000000000000c200000000",
            INIT_57 => X"000000b700000000000000c100000000000000bf00000000000000c500000000",
            INIT_58 => X"000000bb00000000000000b200000000000000bb00000000000000b500000000",
            INIT_59 => X"000000b600000000000000ae00000000000000aa00000000000000b700000000",
            INIT_5A => X"000000b500000000000000b400000000000000b300000000000000b300000000",
            INIT_5B => X"000000c100000000000000c100000000000000bb00000000000000b800000000",
            INIT_5C => X"000000b900000000000000bc00000000000000c000000000000000c100000000",
            INIT_5D => X"000000c000000000000000c000000000000000ba00000000000000b800000000",
            INIT_5E => X"000000bd00000000000000c000000000000000bc00000000000000bb00000000",
            INIT_5F => X"000000ba00000000000000c400000000000000bf00000000000000be00000000",
            INIT_60 => X"000000ab00000000000000ba00000000000000be00000000000000b900000000",
            INIT_61 => X"000000c100000000000000950000000000000084000000000000009900000000",
            INIT_62 => X"000000bc00000000000000ba00000000000000bf00000000000000c600000000",
            INIT_63 => X"000000c400000000000000c300000000000000c100000000000000bf00000000",
            INIT_64 => X"000000bc00000000000000be00000000000000c000000000000000c300000000",
            INIT_65 => X"000000bf00000000000000c000000000000000be00000000000000bc00000000",
            INIT_66 => X"000000c500000000000000c300000000000000c100000000000000bf00000000",
            INIT_67 => X"000000c100000000000000cc00000000000000ca00000000000000ca00000000",
            INIT_68 => X"0000009e00000000000000bc00000000000000c200000000000000ba00000000",
            INIT_69 => X"0000006d000000000000005e0000000000000074000000000000008400000000",
            INIT_6A => X"000000c200000000000000c200000000000000b1000000000000009100000000",
            INIT_6B => X"000000c700000000000000c400000000000000c100000000000000bf00000000",
            INIT_6C => X"000000c600000000000000c800000000000000c700000000000000c700000000",
            INIT_6D => X"000000c600000000000000c700000000000000c400000000000000c400000000",
            INIT_6E => X"000000c400000000000000c400000000000000c400000000000000c500000000",
            INIT_6F => X"000000b900000000000000c600000000000000c500000000000000c600000000",
            INIT_70 => X"000000c600000000000000c400000000000000c500000000000000ba00000000",
            INIT_71 => X"0000005c000000000000008d00000000000000b800000000000000c200000000",
            INIT_72 => X"000000b3000000000000008e0000000000000068000000000000005400000000",
            INIT_73 => X"000000cc00000000000000cc00000000000000c900000000000000c300000000",
            INIT_74 => X"000000c700000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_75 => X"000000bf00000000000000c200000000000000c200000000000000c200000000",
            INIT_76 => X"000000be00000000000000be00000000000000be00000000000000bd00000000",
            INIT_77 => X"000000b500000000000000c000000000000000be00000000000000bf00000000",
            INIT_78 => X"000000c800000000000000c600000000000000c700000000000000b800000000",
            INIT_79 => X"000000b100000000000000c900000000000000c800000000000000c500000000",
            INIT_7A => X"00000080000000000000005d0000000000000054000000000000007500000000",
            INIT_7B => X"000000cd00000000000000d000000000000000ca00000000000000ad00000000",
            INIT_7C => X"000000c700000000000000c700000000000000c800000000000000ca00000000",
            INIT_7D => X"000000c300000000000000c500000000000000c400000000000000c300000000",
            INIT_7E => X"000000bf00000000000000c200000000000000c300000000000000c100000000",
            INIT_7F => X"000000b200000000000000be00000000000000bd00000000000000bf00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "sampleifmap_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d000000000000000cb00000000000000c900000000000000b900000000",
            INIT_01 => X"000000d600000000000000d000000000000000ce00000000000000cd00000000",
            INIT_02 => X"0000005b000000000000004c000000000000005c00000000000000af00000000",
            INIT_03 => X"000000cb00000000000000b5000000000000008c000000000000006900000000",
            INIT_04 => X"000000c200000000000000c500000000000000ca00000000000000ce00000000",
            INIT_05 => X"000000c200000000000000c200000000000000c200000000000000c100000000",
            INIT_06 => X"000000bf00000000000000c100000000000000c300000000000000c200000000",
            INIT_07 => X"000000b400000000000000be00000000000000be00000000000000c100000000",
            INIT_08 => X"000000d600000000000000cf00000000000000cc00000000000000bb00000000",
            INIT_09 => X"000000d000000000000000d300000000000000d400000000000000d400000000",
            INIT_0A => X"000000570000000000000047000000000000007c00000000000000cb00000000",
            INIT_0B => X"0000008400000000000000630000000000000054000000000000005400000000",
            INIT_0C => X"000000cb00000000000000cb00000000000000be00000000000000a700000000",
            INIT_0D => X"000000c400000000000000c500000000000000c000000000000000c300000000",
            INIT_0E => X"000000bf00000000000000c000000000000000c200000000000000c200000000",
            INIT_0F => X"000000b700000000000000c000000000000000bf00000000000000c100000000",
            INIT_10 => X"000000d600000000000000cf00000000000000cf00000000000000be00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000d400000000",
            INIT_12 => X"000000570000000000000048000000000000008900000000000000d300000000",
            INIT_13 => X"0000005300000000000000560000000000000054000000000000005300000000",
            INIT_14 => X"0000009b0000000000000083000000000000006b000000000000005900000000",
            INIT_15 => X"000000cc00000000000000cb00000000000000b600000000000000a300000000",
            INIT_16 => X"000000bf00000000000000c200000000000000c600000000000000ca00000000",
            INIT_17 => X"000000b600000000000000bf00000000000000c000000000000000c100000000",
            INIT_18 => X"000000d700000000000000d100000000000000d200000000000000bf00000000",
            INIT_19 => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1A => X"0000003a000000000000002f000000000000007100000000000000cc00000000",
            INIT_1B => X"0000005d0000000000000057000000000000004c000000000000003f00000000",
            INIT_1C => X"0000003e00000000000000460000000000000050000000000000005a00000000",
            INIT_1D => X"0000009f000000000000007a000000000000004d000000000000003a00000000",
            INIT_1E => X"000000c800000000000000c900000000000000c200000000000000b400000000",
            INIT_1F => X"000000b900000000000000c400000000000000c400000000000000c800000000",
            INIT_20 => X"000000d300000000000000cf00000000000000d000000000000000bf00000000",
            INIT_21 => X"000000d400000000000000d100000000000000d200000000000000d100000000",
            INIT_22 => X"0000002500000000000000410000000000000065000000000000009d00000000",
            INIT_23 => X"00000058000000000000004a0000000000000044000000000000003300000000",
            INIT_24 => X"0000004900000000000000550000000000000056000000000000005b00000000",
            INIT_25 => X"00000048000000000000003e000000000000002e000000000000003700000000",
            INIT_26 => X"0000009e0000000000000085000000000000006b000000000000004e00000000",
            INIT_27 => X"000000ba00000000000000c400000000000000c300000000000000b800000000",
            INIT_28 => X"000000d100000000000000cb00000000000000ca00000000000000ba00000000",
            INIT_29 => X"000000c800000000000000d100000000000000ce00000000000000cf00000000",
            INIT_2A => X"000000640000000000000097000000000000008c000000000000009500000000",
            INIT_2B => X"0000006000000000000000320000000000000035000000000000002d00000000",
            INIT_2C => X"00000048000000000000008000000000000000a0000000000000009c00000000",
            INIT_2D => X"0000004200000000000000590000000000000070000000000000006200000000",
            INIT_2E => X"000000a300000000000000a60000000000000083000000000000004300000000",
            INIT_2F => X"000000b200000000000000bc00000000000000b700000000000000ad00000000",
            INIT_30 => X"000000d200000000000000ca00000000000000c900000000000000b900000000",
            INIT_31 => X"000000d100000000000000d100000000000000d000000000000000d200000000",
            INIT_32 => X"000000bd00000000000000d700000000000000d300000000000000d200000000",
            INIT_33 => X"000000a800000000000000940000000000000092000000000000009000000000",
            INIT_34 => X"0000009a00000000000000c000000000000000ce00000000000000ca00000000",
            INIT_35 => X"0000009f00000000000000b100000000000000b200000000000000a300000000",
            INIT_36 => X"000000c200000000000000bf00000000000000b2000000000000009c00000000",
            INIT_37 => X"000000b000000000000000bc00000000000000c100000000000000c400000000",
            INIT_38 => X"000000c400000000000000c000000000000000bc00000000000000b000000000",
            INIT_39 => X"000000b700000000000000b900000000000000bc00000000000000c000000000",
            INIT_3A => X"000000ad00000000000000b300000000000000b200000000000000b600000000",
            INIT_3B => X"000000ad00000000000000ab00000000000000aa00000000000000aa00000000",
            INIT_3C => X"000000a700000000000000a100000000000000a000000000000000a900000000",
            INIT_3D => X"000000aa00000000000000a500000000000000a100000000000000a500000000",
            INIT_3E => X"00000096000000000000009800000000000000a000000000000000aa00000000",
            INIT_3F => X"0000009c00000000000000a400000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b000000000000006e0000000000000063000000000000007200000000",
            INIT_41 => X"0000005d000000000000005e0000000000000061000000000000006600000000",
            INIT_42 => X"0000005000000000000000580000000000000055000000000000005800000000",
            INIT_43 => X"000000650000000000000053000000000000004e000000000000004d00000000",
            INIT_44 => X"0000006b000000000000006a000000000000006c000000000000007100000000",
            INIT_45 => X"00000071000000000000006f000000000000006e000000000000006c00000000",
            INIT_46 => X"0000007700000000000000780000000000000077000000000000007500000000",
            INIT_47 => X"0000007c000000000000007a0000000000000079000000000000007800000000",
            INIT_48 => X"000000750000000000000071000000000000006d000000000000007a00000000",
            INIT_49 => X"0000007100000000000000720000000000000070000000000000007300000000",
            INIT_4A => X"0000006d000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006c000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006b00000000000000690000000000000070000000000000007300000000",
            INIT_4D => X"000000680000000000000065000000000000006a000000000000006c00000000",
            INIT_4E => X"0000006d000000000000006d000000000000006b000000000000006a00000000",
            INIT_4F => X"00000065000000000000005e0000000000000066000000000000006700000000",
            INIT_50 => X"00000070000000000000006b0000000000000061000000000000007800000000",
            INIT_51 => X"0000005e00000000000000620000000000000068000000000000006d00000000",
            INIT_52 => X"000000560000000000000058000000000000005d000000000000005e00000000",
            INIT_53 => X"0000004e0000000000000050000000000000004f000000000000005200000000",
            INIT_54 => X"000000450000000000000048000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000042000000000000004300000000",
            INIT_56 => X"0000004000000000000000420000000000000041000000000000004000000000",
            INIT_57 => X"0000004d0000000000000035000000000000003f000000000000004300000000",
            INIT_58 => X"0000004500000000000000410000000000000037000000000000005b00000000",
            INIT_59 => X"0000003d000000000000003f0000000000000042000000000000004200000000",
            INIT_5A => X"00000039000000000000003c0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003a00000000000000400000000000000042000000000000003f00000000",
            INIT_5D => X"0000003c000000000000003b0000000000000039000000000000003800000000",
            INIT_5E => X"0000003900000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000005c000000000000004b0000000000000031000000000000003400000000",
            INIT_60 => X"000000440000000000000042000000000000003c000000000000005d00000000",
            INIT_61 => X"0000004100000000000000400000000000000043000000000000004300000000",
            INIT_62 => X"0000003b000000000000003e0000000000000041000000000000004500000000",
            INIT_63 => X"0000003d000000000000003c000000000000003b000000000000003b00000000",
            INIT_64 => X"00000038000000000000003a000000000000003f000000000000004000000000",
            INIT_65 => X"0000003800000000000000380000000000000037000000000000003700000000",
            INIT_66 => X"000000350000000000000038000000000000003a000000000000003900000000",
            INIT_67 => X"000000510000000000000061000000000000005d000000000000004100000000",
            INIT_68 => X"00000039000000000000003d0000000000000039000000000000005900000000",
            INIT_69 => X"0000003b0000000000000039000000000000003b000000000000003900000000",
            INIT_6A => X"000000360000000000000038000000000000003a000000000000003c00000000",
            INIT_6B => X"0000003d000000000000003b000000000000003d000000000000003c00000000",
            INIT_6C => X"00000039000000000000003a000000000000003d000000000000004100000000",
            INIT_6D => X"0000003d000000000000003d000000000000003c000000000000003c00000000",
            INIT_6E => X"000000460000000000000039000000000000003e000000000000004200000000",
            INIT_6F => X"00000043000000000000003b0000000000000059000000000000006100000000",
            INIT_70 => X"0000003e000000000000003f000000000000003c000000000000005900000000",
            INIT_71 => X"0000003f000000000000003e000000000000003e000000000000003e00000000",
            INIT_72 => X"000000520000000000000041000000000000003d000000000000003e00000000",
            INIT_73 => X"00000051000000000000004e0000000000000051000000000000005400000000",
            INIT_74 => X"0000005300000000000000550000000000000054000000000000005800000000",
            INIT_75 => X"0000004000000000000000420000000000000043000000000000005000000000",
            INIT_76 => X"0000006700000000000000560000000000000038000000000000003400000000",
            INIT_77 => X"0000004b000000000000003d0000000000000039000000000000004c00000000",
            INIT_78 => X"0000003c000000000000003d000000000000003c000000000000005c00000000",
            INIT_79 => X"0000004100000000000000430000000000000042000000000000003f00000000",
            INIT_7A => X"0000004800000000000000410000000000000043000000000000004200000000",
            INIT_7B => X"0000004600000000000000480000000000000049000000000000004900000000",
            INIT_7C => X"0000004b000000000000004b000000000000004a000000000000004900000000",
            INIT_7D => X"0000003e00000000000000400000000000000040000000000000004b00000000",
            INIT_7E => X"0000004000000000000000580000000000000056000000000000004100000000",
            INIT_7F => X"000000490000000000000040000000000000003c000000000000003900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "sampleifmap_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c000000000000000b300000000000000b0000000000000009c00000000",
            INIT_01 => X"000000ad00000000000000ad00000000000000ab00000000000000b900000000",
            INIT_02 => X"000000b800000000000000b600000000000000b300000000000000af00000000",
            INIT_03 => X"000000b500000000000000b600000000000000b800000000000000b900000000",
            INIT_04 => X"000000b900000000000000b700000000000000b300000000000000b300000000",
            INIT_05 => X"000000bd00000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000b700000000000000ca00000000000000c400000000000000c500000000",
            INIT_08 => X"000000c300000000000000b800000000000000b3000000000000009b00000000",
            INIT_09 => X"000000a4000000000000009f00000000000000a200000000000000be00000000",
            INIT_0A => X"000000b000000000000000a900000000000000a500000000000000a300000000",
            INIT_0B => X"000000a700000000000000a400000000000000ae00000000000000ab00000000",
            INIT_0C => X"000000a600000000000000a800000000000000a600000000000000ac00000000",
            INIT_0D => X"000000a900000000000000ab00000000000000af00000000000000a900000000",
            INIT_0E => X"000000cc00000000000000bf00000000000000ae00000000000000aa00000000",
            INIT_0F => X"000000be00000000000000d700000000000000d000000000000000ce00000000",
            INIT_10 => X"000000c400000000000000b900000000000000b2000000000000009a00000000",
            INIT_11 => X"000000a800000000000000b200000000000000c100000000000000cb00000000",
            INIT_12 => X"000000c400000000000000be00000000000000af00000000000000a000000000",
            INIT_13 => X"000000bc00000000000000be00000000000000c500000000000000c300000000",
            INIT_14 => X"000000c300000000000000c200000000000000c300000000000000c400000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c600000000000000c400000000",
            INIT_16 => X"000000cd00000000000000cd00000000000000c400000000000000c000000000",
            INIT_17 => X"000000bf00000000000000d700000000000000d000000000000000ce00000000",
            INIT_18 => X"000000c300000000000000bc00000000000000b2000000000000009a00000000",
            INIT_19 => X"0000008000000000000000bc00000000000000c500000000000000ca00000000",
            INIT_1A => X"0000009b000000000000009a0000000000000098000000000000006c00000000",
            INIT_1B => X"0000009400000000000000950000000000000095000000000000009e00000000",
            INIT_1C => X"000000ad00000000000000a300000000000000a100000000000000a700000000",
            INIT_1D => X"0000009f00000000000000ae00000000000000a300000000000000a800000000",
            INIT_1E => X"000000ce00000000000000cc00000000000000d000000000000000bc00000000",
            INIT_1F => X"000000bc00000000000000d400000000000000cd00000000000000cc00000000",
            INIT_20 => X"000000bf00000000000000bb00000000000000b1000000000000009a00000000",
            INIT_21 => X"0000007e00000000000000bd00000000000000c400000000000000c600000000",
            INIT_22 => X"0000006b000000000000006a000000000000008b000000000000008000000000",
            INIT_23 => X"0000007100000000000000760000000000000078000000000000007300000000",
            INIT_24 => X"0000007e00000000000000720000000000000072000000000000007700000000",
            INIT_25 => X"0000007000000000000000880000000000000070000000000000007600000000",
            INIT_26 => X"000000ce00000000000000c900000000000000cb00000000000000a000000000",
            INIT_27 => X"000000be00000000000000d600000000000000cd00000000000000ce00000000",
            INIT_28 => X"000000bd00000000000000bb00000000000000ae000000000000009700000000",
            INIT_29 => X"0000009300000000000000b700000000000000c800000000000000c500000000",
            INIT_2A => X"000000a5000000000000009100000000000000a800000000000000a900000000",
            INIT_2B => X"0000009d0000000000000095000000000000009200000000000000aa00000000",
            INIT_2C => X"000000bd00000000000000b000000000000000b200000000000000b400000000",
            INIT_2D => X"000000b100000000000000bc00000000000000b300000000000000b000000000",
            INIT_2E => X"000000d000000000000000cf00000000000000d000000000000000c400000000",
            INIT_2F => X"000000be00000000000000d800000000000000d100000000000000d000000000",
            INIT_30 => X"000000bd00000000000000b900000000000000ac000000000000009800000000",
            INIT_31 => X"00000060000000000000009300000000000000c600000000000000c200000000",
            INIT_32 => X"0000009800000000000000900000000000000097000000000000009500000000",
            INIT_33 => X"0000008b00000000000000800000000000000079000000000000009800000000",
            INIT_34 => X"000000a200000000000000aa0000000000000097000000000000009c00000000",
            INIT_35 => X"000000a4000000000000009600000000000000ad000000000000009600000000",
            INIT_36 => X"000000d200000000000000cc00000000000000a6000000000000009c00000000",
            INIT_37 => X"000000bc00000000000000d400000000000000cf00000000000000d300000000",
            INIT_38 => X"000000bb00000000000000b600000000000000ac000000000000009b00000000",
            INIT_39 => X"00000065000000000000007700000000000000b500000000000000c200000000",
            INIT_3A => X"0000007800000000000000830000000000000083000000000000007b00000000",
            INIT_3B => X"0000007f00000000000000870000000000000087000000000000009200000000",
            INIT_3C => X"0000007b0000000000000083000000000000007b000000000000007b00000000",
            INIT_3D => X"0000009f000000000000007b0000000000000084000000000000006d00000000",
            INIT_3E => X"000000c700000000000000bf0000000000000084000000000000007b00000000",
            INIT_3F => X"000000ba00000000000000d000000000000000c900000000000000c900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b900000000000000b400000000000000af00000000000000a100000000",
            INIT_41 => X"000000af00000000000000ab00000000000000ba00000000000000c000000000",
            INIT_42 => X"000000a600000000000000ac00000000000000a500000000000000a200000000",
            INIT_43 => X"000000aa00000000000000ad00000000000000ac00000000000000af00000000",
            INIT_44 => X"000000af00000000000000b200000000000000b200000000000000ac00000000",
            INIT_45 => X"000000be00000000000000b200000000000000ac00000000000000a300000000",
            INIT_46 => X"000000cd00000000000000c800000000000000b000000000000000ac00000000",
            INIT_47 => X"000000b900000000000000d100000000000000c900000000000000c800000000",
            INIT_48 => X"000000ba00000000000000b400000000000000b700000000000000ac00000000",
            INIT_49 => X"000000b700000000000000c200000000000000c000000000000000be00000000",
            INIT_4A => X"000000a300000000000000a200000000000000a500000000000000a000000000",
            INIT_4B => X"000000a200000000000000a4000000000000009e000000000000009f00000000",
            INIT_4C => X"000000a200000000000000ac00000000000000ae00000000000000a700000000",
            INIT_4D => X"000000b600000000000000a500000000000000a300000000000000a000000000",
            INIT_4E => X"000000cd00000000000000ca00000000000000c600000000000000c800000000",
            INIT_4F => X"000000b800000000000000d000000000000000ca00000000000000ca00000000",
            INIT_50 => X"000000be00000000000000ba00000000000000c400000000000000b100000000",
            INIT_51 => X"000000b700000000000000c100000000000000c100000000000000c000000000",
            INIT_52 => X"0000009f00000000000000a500000000000000a700000000000000a300000000",
            INIT_53 => X"000000ac00000000000000aa00000000000000a600000000000000a400000000",
            INIT_54 => X"000000ab00000000000000a600000000000000a600000000000000a800000000",
            INIT_55 => X"000000b200000000000000ab00000000000000ad00000000000000a800000000",
            INIT_56 => X"000000c700000000000000c700000000000000c600000000000000c700000000",
            INIT_57 => X"000000b800000000000000d000000000000000c800000000000000c800000000",
            INIT_58 => X"000000c800000000000000c300000000000000cc00000000000000b700000000",
            INIT_59 => X"000000c600000000000000be00000000000000bb00000000000000c900000000",
            INIT_5A => X"000000c100000000000000c100000000000000c100000000000000c200000000",
            INIT_5B => X"000000c600000000000000c600000000000000c200000000000000c100000000",
            INIT_5C => X"000000c600000000000000c300000000000000c300000000000000c600000000",
            INIT_5D => X"000000c500000000000000c400000000000000c400000000000000c500000000",
            INIT_5E => X"000000c900000000000000c900000000000000cb00000000000000c900000000",
            INIT_5F => X"000000bb00000000000000d100000000000000c800000000000000ca00000000",
            INIT_60 => X"000000b200000000000000c600000000000000cd00000000000000b900000000",
            INIT_61 => X"000000c4000000000000009a000000000000008d00000000000000a600000000",
            INIT_62 => X"000000c500000000000000c700000000000000ca00000000000000ca00000000",
            INIT_63 => X"000000ca00000000000000c900000000000000c700000000000000c500000000",
            INIT_64 => X"000000c400000000000000c600000000000000c700000000000000c900000000",
            INIT_65 => X"000000c600000000000000c700000000000000c600000000000000c400000000",
            INIT_66 => X"000000ce00000000000000cb00000000000000ca00000000000000c700000000",
            INIT_67 => X"000000bd00000000000000d400000000000000ce00000000000000cf00000000",
            INIT_68 => X"000000a500000000000000c800000000000000d000000000000000ba00000000",
            INIT_69 => X"0000006b000000000000005f000000000000007c000000000000009000000000",
            INIT_6A => X"000000c700000000000000c700000000000000b3000000000000008f00000000",
            INIT_6B => X"000000cc00000000000000c900000000000000c600000000000000c500000000",
            INIT_6C => X"000000cc00000000000000ce00000000000000cd00000000000000cc00000000",
            INIT_6D => X"000000cd00000000000000cd00000000000000c900000000000000c900000000",
            INIT_6E => X"000000cb00000000000000cb00000000000000cb00000000000000cc00000000",
            INIT_6F => X"000000b700000000000000cf00000000000000ca00000000000000ca00000000",
            INIT_70 => X"000000cc00000000000000d000000000000000d400000000000000ba00000000",
            INIT_71 => X"0000005b000000000000008f00000000000000c100000000000000ce00000000",
            INIT_72 => X"000000b5000000000000008e0000000000000065000000000000005100000000",
            INIT_73 => X"000000cf00000000000000cf00000000000000cc00000000000000c600000000",
            INIT_74 => X"000000ca00000000000000cf00000000000000cf00000000000000cf00000000",
            INIT_75 => X"000000c500000000000000c600000000000000c500000000000000c500000000",
            INIT_76 => X"000000c500000000000000c500000000000000c500000000000000c500000000",
            INIT_77 => X"000000b500000000000000cc00000000000000c500000000000000c400000000",
            INIT_78 => X"000000ce00000000000000d200000000000000d600000000000000b800000000",
            INIT_79 => X"000000b300000000000000cf00000000000000d400000000000000d100000000",
            INIT_7A => X"00000080000000000000005d0000000000000053000000000000007400000000",
            INIT_7B => X"000000ce00000000000000d200000000000000cb00000000000000ae00000000",
            INIT_7C => X"000000c900000000000000ca00000000000000ca00000000000000cc00000000",
            INIT_7D => X"000000c900000000000000c900000000000000c700000000000000c600000000",
            INIT_7E => X"000000c700000000000000c900000000000000ca00000000000000c800000000",
            INIT_7F => X"000000b400000000000000cb00000000000000c600000000000000c600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "sampleifmap_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d500000000000000d600000000000000d700000000000000ba00000000",
            INIT_01 => X"000000d900000000000000d400000000000000d600000000000000d600000000",
            INIT_02 => X"000000560000000000000049000000000000005b00000000000000af00000000",
            INIT_03 => X"000000cc00000000000000b5000000000000008a000000000000006500000000",
            INIT_04 => X"000000c600000000000000c700000000000000cb00000000000000d000000000",
            INIT_05 => X"000000c800000000000000c900000000000000c900000000000000c700000000",
            INIT_06 => X"000000c900000000000000c900000000000000ca00000000000000c800000000",
            INIT_07 => X"000000b600000000000000cc00000000000000c800000000000000ca00000000",
            INIT_08 => X"000000d900000000000000d800000000000000d800000000000000bb00000000",
            INIT_09 => X"000000d300000000000000d600000000000000d900000000000000db00000000",
            INIT_0A => X"000000520000000000000044000000000000007b00000000000000cc00000000",
            INIT_0B => X"0000008200000000000000610000000000000051000000000000004f00000000",
            INIT_0C => X"000000ca00000000000000c900000000000000bc00000000000000a500000000",
            INIT_0D => X"000000c600000000000000c700000000000000c100000000000000c400000000",
            INIT_0E => X"000000c800000000000000c800000000000000c700000000000000c600000000",
            INIT_0F => X"000000b600000000000000cc00000000000000c700000000000000c900000000",
            INIT_10 => X"000000d600000000000000d500000000000000d900000000000000bc00000000",
            INIT_11 => X"000000d200000000000000d600000000000000d800000000000000d800000000",
            INIT_12 => X"000000530000000000000046000000000000008800000000000000d400000000",
            INIT_13 => X"0000004d00000000000000500000000000000050000000000000004e00000000",
            INIT_14 => X"00000097000000000000007e0000000000000066000000000000005300000000",
            INIT_15 => X"000000cc00000000000000c900000000000000b2000000000000009f00000000",
            INIT_16 => X"000000c600000000000000c800000000000000c900000000000000cb00000000",
            INIT_17 => X"000000b400000000000000c900000000000000c500000000000000c700000000",
            INIT_18 => X"000000d500000000000000d600000000000000da00000000000000bb00000000",
            INIT_19 => X"000000d800000000000000d700000000000000d800000000000000d700000000",
            INIT_1A => X"00000037000000000000002d000000000000007000000000000000cc00000000",
            INIT_1B => X"00000051000000000000004d0000000000000045000000000000003a00000000",
            INIT_1C => X"0000003e0000000000000046000000000000004d000000000000005000000000",
            INIT_1D => X"000000a0000000000000007c000000000000004f000000000000003b00000000",
            INIT_1E => X"000000cd00000000000000cd00000000000000c400000000000000b500000000",
            INIT_1F => X"000000b400000000000000ca00000000000000c800000000000000cb00000000",
            INIT_20 => X"000000d100000000000000d200000000000000d800000000000000bc00000000",
            INIT_21 => X"000000d400000000000000d400000000000000d600000000000000d300000000",
            INIT_22 => X"00000021000000000000003a000000000000005f000000000000009a00000000",
            INIT_23 => X"0000004d0000000000000041000000000000003e000000000000003000000000",
            INIT_24 => X"0000004800000000000000540000000000000054000000000000005200000000",
            INIT_25 => X"00000048000000000000003f000000000000002f000000000000003800000000",
            INIT_26 => X"0000009e0000000000000084000000000000006b000000000000004e00000000",
            INIT_27 => X"000000b600000000000000ca00000000000000c100000000000000b500000000",
            INIT_28 => X"000000cf00000000000000ce00000000000000d200000000000000b800000000",
            INIT_29 => X"000000c800000000000000d400000000000000d300000000000000d100000000",
            INIT_2A => X"00000061000000000000008f0000000000000085000000000000009100000000",
            INIT_2B => X"0000005a000000000000002e0000000000000032000000000000002d00000000",
            INIT_2C => X"00000047000000000000007f000000000000009e000000000000009600000000",
            INIT_2D => X"0000004100000000000000580000000000000070000000000000006100000000",
            INIT_2E => X"000000a200000000000000a50000000000000082000000000000004300000000",
            INIT_2F => X"000000b000000000000000c500000000000000b500000000000000a800000000",
            INIT_30 => X"000000d000000000000000cd00000000000000d200000000000000b700000000",
            INIT_31 => X"000000d200000000000000d500000000000000d400000000000000d300000000",
            INIT_32 => X"000000bf00000000000000d400000000000000d100000000000000d100000000",
            INIT_33 => X"000000a600000000000000930000000000000093000000000000009400000000",
            INIT_34 => X"0000009d00000000000000c300000000000000d000000000000000c800000000",
            INIT_35 => X"000000a200000000000000b400000000000000b500000000000000a600000000",
            INIT_36 => X"000000c500000000000000c100000000000000b4000000000000009f00000000",
            INIT_37 => X"000000b100000000000000c700000000000000c100000000000000c300000000",
            INIT_38 => X"000000c200000000000000c300000000000000c400000000000000ae00000000",
            INIT_39 => X"000000b900000000000000bb00000000000000be00000000000000c200000000",
            INIT_3A => X"000000b500000000000000b700000000000000b500000000000000b800000000",
            INIT_3B => X"000000ad00000000000000ae00000000000000b000000000000000b200000000",
            INIT_3C => X"000000ac00000000000000a600000000000000a400000000000000aa00000000",
            INIT_3D => X"000000b000000000000000aa00000000000000a600000000000000aa00000000",
            INIT_3E => X"0000009b000000000000009d00000000000000a500000000000000af00000000",
            INIT_3F => X"0000009e00000000000000af00000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000070000000000000006c000000000000007000000000",
            INIT_41 => X"0000006000000000000000610000000000000064000000000000006700000000",
            INIT_42 => X"00000057000000000000005e000000000000005a000000000000005c00000000",
            INIT_43 => X"0000006700000000000000570000000000000053000000000000005400000000",
            INIT_44 => X"00000070000000000000006f0000000000000070000000000000007300000000",
            INIT_45 => X"0000007600000000000000740000000000000073000000000000007100000000",
            INIT_46 => X"0000007b000000000000007c000000000000007b000000000000007a00000000",
            INIT_47 => X"0000007c0000000000000084000000000000007a000000000000007900000000",
            INIT_48 => X"0000007000000000000000710000000000000073000000000000007500000000",
            INIT_49 => X"000000710000000000000071000000000000006f000000000000007100000000",
            INIT_4A => X"0000006e000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006b000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006e000000000000006c0000000000000073000000000000007300000000",
            INIT_4D => X"0000006b0000000000000068000000000000006d000000000000006f00000000",
            INIT_4E => X"000000700000000000000070000000000000006e000000000000006d00000000",
            INIT_4F => X"000000650000000000000062000000000000005f000000000000006400000000",
            INIT_50 => X"0000006a00000000000000690000000000000066000000000000007100000000",
            INIT_51 => X"0000005d00000000000000610000000000000066000000000000006a00000000",
            INIT_52 => X"000000550000000000000059000000000000005e000000000000005f00000000",
            INIT_53 => X"0000004e000000000000004f000000000000004e000000000000005200000000",
            INIT_54 => X"000000440000000000000047000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000041000000000000004300000000",
            INIT_56 => X"0000004100000000000000420000000000000042000000000000004100000000",
            INIT_57 => X"0000006400000000000000470000000000000037000000000000003c00000000",
            INIT_58 => X"000000400000000000000041000000000000003c000000000000005400000000",
            INIT_59 => X"0000003c000000000000003e0000000000000040000000000000004000000000",
            INIT_5A => X"00000038000000000000003d0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003b00000000000000410000000000000043000000000000004000000000",
            INIT_5D => X"0000003c000000000000003b000000000000003a000000000000003800000000",
            INIT_5E => X"0000003800000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000008000000000000000750000000000000048000000000000003800000000",
            INIT_60 => X"0000003e000000000000003f000000000000003b000000000000005300000000",
            INIT_61 => X"0000003f000000000000003d0000000000000041000000000000003f00000000",
            INIT_62 => X"00000039000000000000003c000000000000003e000000000000004300000000",
            INIT_63 => X"0000003d000000000000003c000000000000003a000000000000003a00000000",
            INIT_64 => X"0000003e00000000000000400000000000000044000000000000004100000000",
            INIT_65 => X"0000003d000000000000003e000000000000003c000000000000003d00000000",
            INIT_66 => X"00000041000000000000003d000000000000003a000000000000003a00000000",
            INIT_67 => X"0000006300000000000000890000000000000088000000000000005b00000000",
            INIT_68 => X"00000039000000000000003d0000000000000035000000000000004f00000000",
            INIT_69 => X"0000003c000000000000003a000000000000003b000000000000003700000000",
            INIT_6A => X"000000370000000000000039000000000000003c000000000000003d00000000",
            INIT_6B => X"0000003f000000000000003d000000000000003e000000000000003c00000000",
            INIT_6C => X"0000003b000000000000003c000000000000003f000000000000004300000000",
            INIT_6D => X"0000003f0000000000000040000000000000003e000000000000003e00000000",
            INIT_6E => X"0000006e0000000000000047000000000000003c000000000000003e00000000",
            INIT_6F => X"0000004a000000000000004f0000000000000077000000000000008e00000000",
            INIT_70 => X"000000410000000000000042000000000000003a000000000000005200000000",
            INIT_71 => X"0000003e000000000000003e000000000000003e000000000000003f00000000",
            INIT_72 => X"0000004f0000000000000041000000000000003e000000000000003f00000000",
            INIT_73 => X"0000004d000000000000004a000000000000004c000000000000004f00000000",
            INIT_74 => X"0000004e00000000000000500000000000000050000000000000005400000000",
            INIT_75 => X"00000041000000000000003e000000000000003f000000000000004c00000000",
            INIT_76 => X"0000008d000000000000007c0000000000000056000000000000004200000000",
            INIT_77 => X"0000004500000000000000400000000000000042000000000000006600000000",
            INIT_78 => X"0000003a000000000000003a0000000000000034000000000000004e00000000",
            INIT_79 => X"00000039000000000000003b000000000000003a000000000000003a00000000",
            INIT_7A => X"00000045000000000000003a000000000000003b000000000000003a00000000",
            INIT_7B => X"0000004500000000000000460000000000000047000000000000004700000000",
            INIT_7C => X"0000004a00000000000000490000000000000048000000000000004800000000",
            INIT_7D => X"00000044000000000000003f000000000000003f000000000000004900000000",
            INIT_7E => X"0000005800000000000000800000000000000080000000000000005a00000000",
            INIT_7F => X"000000440000000000000041000000000000003f000000000000004200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "sampleifmap_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cd00000000000000c100000000000000bb000000000000009500000000",
            INIT_01 => X"000000b400000000000000b500000000000000b700000000000000ca00000000",
            INIT_02 => X"000000c000000000000000c100000000000000bd00000000000000b600000000",
            INIT_03 => X"000000bd00000000000000bd00000000000000c000000000000000c000000000",
            INIT_04 => X"000000c000000000000000bd00000000000000b900000000000000ba00000000",
            INIT_05 => X"000000be00000000000000c000000000000000c100000000000000c100000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000ab00000000000000d400000000000000d100000000000000ca00000000",
            INIT_08 => X"000000e300000000000000d700000000000000cc000000000000009d00000000",
            INIT_09 => X"000000b300000000000000b300000000000000be00000000000000e000000000",
            INIT_0A => X"000000c300000000000000c300000000000000bb00000000000000b300000000",
            INIT_0B => X"000000b700000000000000b400000000000000be00000000000000bb00000000",
            INIT_0C => X"000000b700000000000000b800000000000000b700000000000000bc00000000",
            INIT_0D => X"000000bc00000000000000bc00000000000000bf00000000000000b900000000",
            INIT_0E => X"000000e000000000000000d300000000000000c200000000000000be00000000",
            INIT_0F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_10 => X"000000db00000000000000d500000000000000c9000000000000009900000000",
            INIT_11 => X"000000b800000000000000c400000000000000d500000000000000df00000000",
            INIT_12 => X"000000d400000000000000d300000000000000c300000000000000b100000000",
            INIT_13 => X"000000ca00000000000000cc00000000000000d200000000000000d000000000",
            INIT_14 => X"000000d100000000000000d000000000000000d100000000000000d100000000",
            INIT_15 => X"000000d000000000000000d000000000000000d400000000000000d200000000",
            INIT_16 => X"000000df00000000000000de00000000000000d500000000000000d000000000",
            INIT_17 => X"000000b800000000000000e000000000000000d700000000000000da00000000",
            INIT_18 => X"000000de00000000000000d300000000000000cf00000000000000a600000000",
            INIT_19 => X"0000008300000000000000c900000000000000dc00000000000000e200000000",
            INIT_1A => X"000000b100000000000000a6000000000000009e000000000000007700000000",
            INIT_1B => X"000000ab00000000000000a600000000000000a700000000000000b200000000",
            INIT_1C => X"000000ba00000000000000b200000000000000b200000000000000b700000000",
            INIT_1D => X"000000a500000000000000b400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000dd00000000000000dc00000000000000e400000000000000cf00000000",
            INIT_1F => X"000000ba00000000000000e600000000000000df00000000000000e000000000",
            INIT_20 => X"000000da00000000000000ca00000000000000cb00000000000000a700000000",
            INIT_21 => X"0000008e00000000000000d600000000000000e100000000000000e000000000",
            INIT_22 => X"0000008100000000000000780000000000000098000000000000009900000000",
            INIT_23 => X"00000083000000000000007c000000000000007e000000000000008100000000",
            INIT_24 => X"0000008a00000000000000820000000000000084000000000000008600000000",
            INIT_25 => X"0000007b000000000000008d0000000000000088000000000000008800000000",
            INIT_26 => X"000000d900000000000000da00000000000000e300000000000000ba00000000",
            INIT_27 => X"000000b900000000000000e300000000000000dc00000000000000de00000000",
            INIT_28 => X"000000d900000000000000cb00000000000000c900000000000000a400000000",
            INIT_29 => X"000000a500000000000000d100000000000000da00000000000000dc00000000",
            INIT_2A => X"000000b4000000000000009c00000000000000b500000000000000c400000000",
            INIT_2B => X"000000ac00000000000000a300000000000000a000000000000000b300000000",
            INIT_2C => X"000000c900000000000000be00000000000000c100000000000000bf00000000",
            INIT_2D => X"000000be00000000000000c600000000000000c000000000000000bf00000000",
            INIT_2E => X"000000e100000000000000e100000000000000e100000000000000d400000000",
            INIT_2F => X"000000bc00000000000000e800000000000000e100000000000000df00000000",
            INIT_30 => X"000000d900000000000000c800000000000000c600000000000000a400000000",
            INIT_31 => X"0000006800000000000000ac00000000000000d600000000000000d900000000",
            INIT_32 => X"000000af00000000000000a600000000000000a5000000000000009e00000000",
            INIT_33 => X"000000a00000000000000097000000000000009000000000000000a500000000",
            INIT_34 => X"000000b600000000000000bd00000000000000ad00000000000000b200000000",
            INIT_35 => X"000000b900000000000000ad00000000000000b700000000000000aa00000000",
            INIT_36 => X"000000e200000000000000dc00000000000000b200000000000000a600000000",
            INIT_37 => X"000000bc00000000000000e700000000000000e000000000000000dd00000000",
            INIT_38 => X"000000d800000000000000c700000000000000c900000000000000a900000000",
            INIT_39 => X"0000006f000000000000009200000000000000cb00000000000000da00000000",
            INIT_3A => X"00000090000000000000009d0000000000000095000000000000008600000000",
            INIT_3B => X"00000090000000000000008f000000000000008f000000000000009b00000000",
            INIT_3C => X"0000008e0000000000000094000000000000008e000000000000009300000000",
            INIT_3D => X"000000b0000000000000008e000000000000008d000000000000007f00000000",
            INIT_3E => X"000000dc00000000000000d10000000000000095000000000000008900000000",
            INIT_3F => X"000000ba00000000000000e400000000000000dc00000000000000d900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d900000000000000c700000000000000ce00000000000000b100000000",
            INIT_41 => X"000000c500000000000000c100000000000000cd00000000000000db00000000",
            INIT_42 => X"000000b800000000000000bb00000000000000b700000000000000b800000000",
            INIT_43 => X"000000bd00000000000000bb00000000000000ba00000000000000c000000000",
            INIT_44 => X"000000bf00000000000000c200000000000000c200000000000000c000000000",
            INIT_45 => X"000000c800000000000000bc00000000000000ba00000000000000b200000000",
            INIT_46 => X"000000db00000000000000d600000000000000c600000000000000c100000000",
            INIT_47 => X"000000b900000000000000e400000000000000dd00000000000000db00000000",
            INIT_48 => X"000000d600000000000000c500000000000000d400000000000000ba00000000",
            INIT_49 => X"000000d200000000000000dc00000000000000d600000000000000d700000000",
            INIT_4A => X"000000ba00000000000000b600000000000000bb00000000000000b900000000",
            INIT_4B => X"000000ba00000000000000b900000000000000b400000000000000b600000000",
            INIT_4C => X"000000b800000000000000c300000000000000c600000000000000c100000000",
            INIT_4D => X"000000c600000000000000b600000000000000b600000000000000b500000000",
            INIT_4E => X"000000df00000000000000dd00000000000000de00000000000000de00000000",
            INIT_4F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_50 => X"000000d800000000000000c800000000000000de00000000000000bc00000000",
            INIT_51 => X"000000cc00000000000000d600000000000000d400000000000000d700000000",
            INIT_52 => X"000000b000000000000000b600000000000000b800000000000000b500000000",
            INIT_53 => X"000000bf00000000000000bc00000000000000b800000000000000b500000000",
            INIT_54 => X"000000b900000000000000b800000000000000ba00000000000000bd00000000",
            INIT_55 => X"000000c900000000000000ba00000000000000b800000000000000b600000000",
            INIT_56 => X"000000db00000000000000dc00000000000000dd00000000000000df00000000",
            INIT_57 => X"000000b800000000000000e300000000000000dc00000000000000db00000000",
            INIT_58 => X"000000e000000000000000cf00000000000000e200000000000000bf00000000",
            INIT_59 => X"000000de00000000000000d700000000000000d100000000000000dc00000000",
            INIT_5A => X"000000d700000000000000d600000000000000d700000000000000d900000000",
            INIT_5B => X"000000df00000000000000df00000000000000db00000000000000d900000000",
            INIT_5C => X"000000da00000000000000db00000000000000dd00000000000000df00000000",
            INIT_5D => X"000000db00000000000000d900000000000000d600000000000000d800000000",
            INIT_5E => X"000000d600000000000000d900000000000000db00000000000000db00000000",
            INIT_5F => X"000000ba00000000000000e300000000000000db00000000000000d700000000",
            INIT_60 => X"000000ce00000000000000d400000000000000dc00000000000000bc00000000",
            INIT_61 => X"000000d900000000000000ac000000000000009900000000000000b500000000",
            INIT_62 => X"000000dc00000000000000dd00000000000000e100000000000000e200000000",
            INIT_63 => X"000000e200000000000000e100000000000000df00000000000000de00000000",
            INIT_64 => X"000000da00000000000000dc00000000000000dd00000000000000e100000000",
            INIT_65 => X"000000da00000000000000dc00000000000000db00000000000000d900000000",
            INIT_66 => X"000000e000000000000000de00000000000000dc00000000000000d900000000",
            INIT_67 => X"000000bb00000000000000e600000000000000e000000000000000e000000000",
            INIT_68 => X"000000c100000000000000d600000000000000df00000000000000bd00000000",
            INIT_69 => X"000000730000000000000063000000000000007e000000000000009d00000000",
            INIT_6A => X"000000dd00000000000000dd00000000000000c6000000000000009d00000000",
            INIT_6B => X"000000e200000000000000df00000000000000dc00000000000000da00000000",
            INIT_6C => X"000000df00000000000000e100000000000000e000000000000000e200000000",
            INIT_6D => X"000000e000000000000000e000000000000000dd00000000000000dc00000000",
            INIT_6E => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_6F => X"000000b700000000000000e200000000000000dd00000000000000dd00000000",
            INIT_70 => X"000000e900000000000000de00000000000000e200000000000000bd00000000",
            INIT_71 => X"0000005a000000000000009200000000000000c400000000000000dc00000000",
            INIT_72 => X"000000ca00000000000000a10000000000000071000000000000005400000000",
            INIT_73 => X"000000e400000000000000e300000000000000e000000000000000da00000000",
            INIT_74 => X"000000dc00000000000000e000000000000000e100000000000000e200000000",
            INIT_75 => X"000000d900000000000000d800000000000000d700000000000000d700000000",
            INIT_76 => X"000000d800000000000000d800000000000000d800000000000000d800000000",
            INIT_77 => X"000000b600000000000000e100000000000000da00000000000000d700000000",
            INIT_78 => X"000000ea00000000000000e000000000000000e500000000000000bb00000000",
            INIT_79 => X"000000b300000000000000da00000000000000e100000000000000e100000000",
            INIT_7A => X"00000091000000000000006a0000000000000058000000000000007300000000",
            INIT_7B => X"000000e100000000000000e400000000000000dd00000000000000c000000000",
            INIT_7C => X"000000d900000000000000da00000000000000db00000000000000df00000000",
            INIT_7D => X"000000db00000000000000d900000000000000d600000000000000d600000000",
            INIT_7E => X"000000da00000000000000dc00000000000000dd00000000000000db00000000",
            INIT_7F => X"000000b700000000000000e200000000000000dc00000000000000d900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "sampleifmap_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e900000000000000de00000000000000e900000000000000be00000000",
            INIT_01 => X"000000e100000000000000e000000000000000e200000000000000e400000000",
            INIT_02 => X"0000005b0000000000000050000000000000006200000000000000b500000000",
            INIT_03 => X"000000d900000000000000c00000000000000092000000000000006a00000000",
            INIT_04 => X"000000da00000000000000dd00000000000000e100000000000000e000000000",
            INIT_05 => X"000000d900000000000000da00000000000000da00000000000000d900000000",
            INIT_06 => X"000000dd00000000000000dd00000000000000dd00000000000000da00000000",
            INIT_07 => X"000000bc00000000000000e300000000000000dc00000000000000dd00000000",
            INIT_08 => X"000000e900000000000000dd00000000000000ea00000000000000bf00000000",
            INIT_09 => X"000000dd00000000000000e200000000000000e300000000000000e700000000",
            INIT_0A => X"0000004f0000000000000049000000000000008200000000000000d500000000",
            INIT_0B => X"0000008800000000000000640000000000000050000000000000004b00000000",
            INIT_0C => X"000000dc00000000000000d700000000000000c800000000000000ad00000000",
            INIT_0D => X"000000de00000000000000df00000000000000d900000000000000d900000000",
            INIT_0E => X"000000db00000000000000db00000000000000dd00000000000000dd00000000",
            INIT_0F => X"000000bd00000000000000e300000000000000db00000000000000da00000000",
            INIT_10 => X"000000e400000000000000d900000000000000e800000000000000bd00000000",
            INIT_11 => X"000000dc00000000000000e200000000000000e100000000000000e300000000",
            INIT_12 => X"00000050000000000000004a000000000000009000000000000000dd00000000",
            INIT_13 => X"0000004c000000000000004e000000000000004c000000000000004a00000000",
            INIT_14 => X"000000a100000000000000810000000000000064000000000000005300000000",
            INIT_15 => X"000000e200000000000000e100000000000000c900000000000000b000000000",
            INIT_16 => X"000000d700000000000000d900000000000000dc00000000000000df00000000",
            INIT_17 => X"000000bb00000000000000e100000000000000d900000000000000d700000000",
            INIT_18 => X"000000e100000000000000d700000000000000e800000000000000bb00000000",
            INIT_19 => X"000000e200000000000000e300000000000000e100000000000000e000000000",
            INIT_1A => X"000000380000000000000032000000000000007700000000000000d500000000",
            INIT_1B => X"00000052000000000000004d0000000000000045000000000000003b00000000",
            INIT_1C => X"0000003f00000000000000420000000000000048000000000000005000000000",
            INIT_1D => X"000000a20000000000000085000000000000005b000000000000004100000000",
            INIT_1E => X"000000df00000000000000da00000000000000cc00000000000000b800000000",
            INIT_1F => X"000000bc00000000000000e300000000000000dd00000000000000dd00000000",
            INIT_20 => X"000000df00000000000000de00000000000000e700000000000000b700000000",
            INIT_21 => X"000000e100000000000000e400000000000000e600000000000000df00000000",
            INIT_22 => X"00000027000000000000003c000000000000006200000000000000a200000000",
            INIT_23 => X"0000004e00000000000000440000000000000043000000000000003500000000",
            INIT_24 => X"0000004800000000000000530000000000000052000000000000005100000000",
            INIT_25 => X"00000043000000000000003f0000000000000031000000000000003900000000",
            INIT_26 => X"000000a8000000000000008b000000000000006d000000000000004b00000000",
            INIT_27 => X"000000c300000000000000df00000000000000d700000000000000c600000000",
            INIT_28 => X"000000de00000000000000e200000000000000e200000000000000b000000000",
            INIT_29 => X"000000d400000000000000e200000000000000e200000000000000de00000000",
            INIT_2A => X"0000006a0000000000000096000000000000008b000000000000009b00000000",
            INIT_2B => X"0000005e00000000000000330000000000000039000000000000003500000000",
            INIT_2C => X"00000049000000000000008200000000000000a1000000000000009a00000000",
            INIT_2D => X"00000043000000000000005a0000000000000072000000000000006300000000",
            INIT_2E => X"000000a900000000000000ab0000000000000086000000000000004500000000",
            INIT_2F => X"000000be00000000000000d000000000000000c500000000000000b700000000",
            INIT_30 => X"000000df00000000000000e100000000000000e100000000000000af00000000",
            INIT_31 => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_32 => X"000000cc00000000000000e400000000000000e000000000000000de00000000",
            INIT_33 => X"000000b300000000000000a0000000000000009f000000000000009f00000000",
            INIT_34 => X"000000a900000000000000cf00000000000000dc00000000000000d600000000",
            INIT_35 => X"000000ad00000000000000c000000000000000c100000000000000b200000000",
            INIT_36 => X"000000d600000000000000d200000000000000c300000000000000ab00000000",
            INIT_37 => X"000000bd00000000000000d200000000000000d100000000000000d800000000",
            INIT_38 => X"000000d100000000000000d700000000000000d400000000000000a600000000",
            INIT_39 => X"000000c700000000000000c900000000000000cc00000000000000ce00000000",
            INIT_3A => X"000000c200000000000000c500000000000000c300000000000000c700000000",
            INIT_3B => X"000000c400000000000000c200000000000000c100000000000000c000000000",
            INIT_3C => X"000000ca00000000000000c400000000000000c200000000000000c400000000",
            INIT_3D => X"000000cd00000000000000c800000000000000c400000000000000c800000000",
            INIT_3E => X"000000bf00000000000000c000000000000000c500000000000000ce00000000",
            INIT_3F => X"000000b500000000000000c900000000000000c500000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000820000000000000078000000000000006500000000",
            INIT_41 => X"0000006a000000000000006b0000000000000070000000000000007600000000",
            INIT_42 => X"0000006300000000000000660000000000000062000000000000006500000000",
            INIT_43 => X"00000080000000000000006c0000000000000065000000000000006200000000",
            INIT_44 => X"0000009300000000000000920000000000000092000000000000009000000000",
            INIT_45 => X"0000009e00000000000000980000000000000096000000000000009400000000",
            INIT_46 => X"000000a800000000000000a800000000000000a600000000000000a400000000",
            INIT_47 => X"0000009200000000000000a700000000000000a500000000000000a800000000",
            INIT_48 => X"0000008600000000000000860000000000000082000000000000006f00000000",
            INIT_49 => X"0000008800000000000000890000000000000088000000000000008a00000000",
            INIT_4A => X"0000007e00000000000000830000000000000086000000000000008400000000",
            INIT_4B => X"0000008300000000000000830000000000000080000000000000007f00000000",
            INIT_4C => X"00000081000000000000007f0000000000000086000000000000008a00000000",
            INIT_4D => X"0000007e000000000000007c0000000000000080000000000000008100000000",
            INIT_4E => X"0000008400000000000000840000000000000082000000000000008100000000",
            INIT_4F => X"0000006000000000000000730000000000000073000000000000007700000000",
            INIT_50 => X"0000007800000000000000780000000000000071000000000000006800000000",
            INIT_51 => X"00000064000000000000006c0000000000000076000000000000007a00000000",
            INIT_52 => X"000000590000000000000055000000000000005b000000000000006000000000",
            INIT_53 => X"0000005600000000000000570000000000000055000000000000005800000000",
            INIT_54 => X"000000430000000000000046000000000000004f000000000000005600000000",
            INIT_55 => X"0000003c000000000000003f0000000000000041000000000000004200000000",
            INIT_56 => X"0000003b000000000000003c000000000000003c000000000000003b00000000",
            INIT_57 => X"0000004b000000000000003f0000000000000032000000000000003600000000",
            INIT_58 => X"00000039000000000000003d0000000000000037000000000000003d00000000",
            INIT_59 => X"00000036000000000000003b000000000000003f000000000000003a00000000",
            INIT_5A => X"0000002f000000000000002f0000000000000033000000000000003800000000",
            INIT_5B => X"0000003200000000000000310000000000000032000000000000003000000000",
            INIT_5C => X"0000002f00000000000000350000000000000037000000000000003300000000",
            INIT_5D => X"000000370000000000000032000000000000002e000000000000002d00000000",
            INIT_5E => X"0000003400000000000000340000000000000034000000000000003600000000",
            INIT_5F => X"000000680000000000000068000000000000003a000000000000003000000000",
            INIT_60 => X"0000003c0000000000000041000000000000003d000000000000004400000000",
            INIT_61 => X"000000390000000000000037000000000000003d000000000000003e00000000",
            INIT_62 => X"0000003a00000000000000370000000000000038000000000000003d00000000",
            INIT_63 => X"0000003600000000000000380000000000000038000000000000003b00000000",
            INIT_64 => X"000000340000000000000037000000000000003b000000000000003900000000",
            INIT_65 => X"0000003400000000000000340000000000000033000000000000003300000000",
            INIT_66 => X"0000003900000000000000370000000000000035000000000000003300000000",
            INIT_67 => X"0000004b00000000000000780000000000000071000000000000004b00000000",
            INIT_68 => X"00000035000000000000003b0000000000000034000000000000003e00000000",
            INIT_69 => X"0000003600000000000000340000000000000039000000000000003900000000",
            INIT_6A => X"0000003200000000000000300000000000000032000000000000003600000000",
            INIT_6B => X"0000003500000000000000340000000000000038000000000000003900000000",
            INIT_6C => X"0000003300000000000000340000000000000036000000000000003900000000",
            INIT_6D => X"0000003000000000000000350000000000000037000000000000003600000000",
            INIT_6E => X"0000005f000000000000003d0000000000000034000000000000003200000000",
            INIT_6F => X"00000032000000000000003e0000000000000065000000000000007c00000000",
            INIT_70 => X"00000037000000000000003a0000000000000035000000000000003e00000000",
            INIT_71 => X"0000003c000000000000003c000000000000003d000000000000003b00000000",
            INIT_72 => X"0000004b000000000000003a0000000000000037000000000000003900000000",
            INIT_73 => X"0000004500000000000000440000000000000048000000000000004c00000000",
            INIT_74 => X"00000049000000000000004b000000000000004a000000000000004b00000000",
            INIT_75 => X"000000350000000000000037000000000000003a000000000000004600000000",
            INIT_76 => X"0000007f000000000000006b0000000000000045000000000000003300000000",
            INIT_77 => X"000000330000000000000036000000000000003a000000000000005b00000000",
            INIT_78 => X"0000002e00000000000000330000000000000033000000000000004000000000",
            INIT_79 => X"0000003500000000000000390000000000000038000000000000003300000000",
            INIT_7A => X"0000003e00000000000000320000000000000033000000000000003400000000",
            INIT_7B => X"00000039000000000000003c000000000000003e000000000000004000000000",
            INIT_7C => X"000000400000000000000040000000000000003e000000000000003c00000000",
            INIT_7D => X"0000003700000000000000340000000000000035000000000000004000000000",
            INIT_7E => X"0000004800000000000000690000000000000067000000000000004600000000",
            INIT_7F => X"0000003200000000000000340000000000000032000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "sampleifmap_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000300000000000000046000000000000004100000000",
            INIT_01 => X"0000002d000000000000002c0000000000000028000000000000001700000000",
            INIT_02 => X"0000000f000000000000000a0000000000000028000000000000002d00000000",
            INIT_03 => X"0000003000000000000000330000000000000035000000000000002c00000000",
            INIT_04 => X"0000005b000000000000005d000000000000005a000000000000004100000000",
            INIT_05 => X"00000037000000000000003c0000000000000051000000000000005f00000000",
            INIT_06 => X"000000440000000000000029000000000000006f000000000000007000000000",
            INIT_07 => X"0000004300000000000000360000000000000033000000000000004d00000000",
            INIT_08 => X"0000001e000000000000003c000000000000004f000000000000004500000000",
            INIT_09 => X"0000003100000000000000310000000000000041000000000000002900000000",
            INIT_0A => X"0000001900000000000000070000000000000023000000000000003100000000",
            INIT_0B => X"0000003100000000000000370000000000000045000000000000004100000000",
            INIT_0C => X"0000005000000000000000530000000000000055000000000000004d00000000",
            INIT_0D => X"0000003b00000000000000370000000000000051000000000000005700000000",
            INIT_0E => X"0000002f000000000000001f0000000000000079000000000000008300000000",
            INIT_0F => X"0000003d00000000000000410000000000000036000000000000003800000000",
            INIT_10 => X"0000002900000000000000480000000000000054000000000000004900000000",
            INIT_11 => X"000000360000000000000032000000000000004a000000000000004000000000",
            INIT_12 => X"00000024000000000000000b0000000000000020000000000000003600000000",
            INIT_13 => X"00000027000000000000002f0000000000000043000000000000003c00000000",
            INIT_14 => X"0000003e000000000000003b000000000000004d000000000000004b00000000",
            INIT_15 => X"0000003f00000000000000300000000000000055000000000000005300000000",
            INIT_16 => X"0000002900000000000000170000000000000080000000000000008b00000000",
            INIT_17 => X"000000300000000000000049000000000000004e000000000000004600000000",
            INIT_18 => X"000000360000000000000050000000000000004b000000000000005800000000",
            INIT_19 => X"0000003f00000000000000370000000000000044000000000000005000000000",
            INIT_1A => X"000000250000000000000011000000000000001c000000000000003a00000000",
            INIT_1B => X"0000002700000000000000280000000000000033000000000000002b00000000",
            INIT_1C => X"00000046000000000000004b0000000000000062000000000000005500000000",
            INIT_1D => X"0000004400000000000000320000000000000054000000000000005600000000",
            INIT_1E => X"0000004b000000000000002f0000000000000089000000000000008e00000000",
            INIT_1F => X"000000260000000000000041000000000000005d000000000000006400000000",
            INIT_20 => X"00000042000000000000006f0000000000000059000000000000005f00000000",
            INIT_21 => X"00000044000000000000003d000000000000003d000000000000005100000000",
            INIT_22 => X"00000016000000000000000f0000000000000016000000000000003e00000000",
            INIT_23 => X"0000003f00000000000000330000000000000023000000000000001f00000000",
            INIT_24 => X"000000470000000000000048000000000000004b000000000000004800000000",
            INIT_25 => X"0000004e00000000000000330000000000000053000000000000004d00000000",
            INIT_26 => X"000000570000000000000057000000000000009c000000000000009500000000",
            INIT_27 => X"00000058000000000000004b000000000000005f000000000000006300000000",
            INIT_28 => X"0000004d00000000000000520000000000000053000000000000005200000000",
            INIT_29 => X"000000390000000000000040000000000000003a000000000000004700000000",
            INIT_2A => X"0000001c00000000000000110000000000000014000000000000003b00000000",
            INIT_2B => X"000000470000000000000047000000000000003d000000000000003200000000",
            INIT_2C => X"0000003800000000000000440000000000000043000000000000004500000000",
            INIT_2D => X"0000004e00000000000000460000000000000053000000000000002900000000",
            INIT_2E => X"00000059000000000000006200000000000000ac000000000000009c00000000",
            INIT_2F => X"000000630000000000000070000000000000006f000000000000005e00000000",
            INIT_30 => X"0000003b00000000000000200000000000000040000000000000004500000000",
            INIT_31 => X"000000310000000000000049000000000000004a000000000000004800000000",
            INIT_32 => X"0000003e000000000000001d0000000000000012000000000000003100000000",
            INIT_33 => X"0000003f00000000000000560000000000000055000000000000005200000000",
            INIT_34 => X"0000002b000000000000005f0000000000000034000000000000002200000000",
            INIT_35 => X"0000004e0000000000000055000000000000005e000000000000001900000000",
            INIT_36 => X"0000006b000000000000006d00000000000000b400000000000000a600000000",
            INIT_37 => X"0000002f00000000000000560000000000000083000000000000006c00000000",
            INIT_38 => X"0000004600000000000000190000000000000035000000000000003b00000000",
            INIT_39 => X"0000003d0000000000000050000000000000004e000000000000005100000000",
            INIT_3A => X"0000005e0000000000000035000000000000000a000000000000002800000000",
            INIT_3B => X"00000019000000000000004b0000000000000058000000000000005700000000",
            INIT_3C => X"00000039000000000000005c000000000000002d000000000000000d00000000",
            INIT_3D => X"0000006200000000000000590000000000000065000000000000003200000000",
            INIT_3E => X"0000007c000000000000007800000000000000b3000000000000009000000000",
            INIT_3F => X"0000001800000000000000340000000000000080000000000000007c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000660000000000000031000000000000002f000000000000004400000000",
            INIT_41 => X"0000004f000000000000003f0000000000000059000000000000007700000000",
            INIT_42 => X"0000006000000000000000510000000000000022000000000000004200000000",
            INIT_43 => X"0000000e0000000000000029000000000000005a000000000000005900000000",
            INIT_44 => X"000000470000000000000043000000000000005c000000000000003400000000",
            INIT_45 => X"00000073000000000000006e0000000000000071000000000000006f00000000",
            INIT_46 => X"0000007f0000000000000079000000000000009c000000000000008800000000",
            INIT_47 => X"00000016000000000000001f0000000000000073000000000000007c00000000",
            INIT_48 => X"0000007200000000000000370000000000000035000000000000004d00000000",
            INIT_49 => X"000000370000000000000041000000000000007b000000000000008000000000",
            INIT_4A => X"0000006e000000000000006f0000000000000052000000000000004f00000000",
            INIT_4B => X"0000002500000000000000140000000000000045000000000000006a00000000",
            INIT_4C => X"0000006100000000000000530000000000000069000000000000005c00000000",
            INIT_4D => X"0000005c00000000000000730000000000000078000000000000007600000000",
            INIT_4E => X"0000007f000000000000007d0000000000000093000000000000009000000000",
            INIT_4F => X"00000017000000000000000e000000000000005f000000000000007700000000",
            INIT_50 => X"000000700000000000000036000000000000003a000000000000005500000000",
            INIT_51 => X"0000003100000000000000640000000000000084000000000000008100000000",
            INIT_52 => X"0000006d00000000000000680000000000000054000000000000002700000000",
            INIT_53 => X"00000053000000000000003f000000000000005d000000000000007d00000000",
            INIT_54 => X"0000006e0000000000000068000000000000005e000000000000006100000000",
            INIT_55 => X"000000390000000000000055000000000000007f000000000000006d00000000",
            INIT_56 => X"0000007c000000000000007b0000000000000096000000000000009800000000",
            INIT_57 => X"00000015000000000000000c000000000000005d000000000000007200000000",
            INIT_58 => X"0000006b00000000000000320000000000000035000000000000006c00000000",
            INIT_59 => X"0000004b00000000000000800000000000000083000000000000007e00000000",
            INIT_5A => X"0000006b0000000000000055000000000000005b000000000000003300000000",
            INIT_5B => X"000000930000000000000081000000000000006e000000000000008a00000000",
            INIT_5C => X"0000007700000000000000710000000000000078000000000000008400000000",
            INIT_5D => X"0000005d000000000000005a0000000000000073000000000000007500000000",
            INIT_5E => X"0000007d0000000000000071000000000000008d00000000000000a000000000",
            INIT_5F => X"00000009000000000000000e0000000000000065000000000000007900000000",
            INIT_60 => X"0000005c000000000000002b000000000000002a000000000000006000000000",
            INIT_61 => X"0000007700000000000000820000000000000080000000000000006a00000000",
            INIT_62 => X"000000890000000000000072000000000000007b000000000000007800000000",
            INIT_63 => X"000000840000000000000069000000000000006e000000000000009400000000",
            INIT_64 => X"0000008600000000000000800000000000000087000000000000009200000000",
            INIT_65 => X"00000077000000000000007e0000000000000078000000000000008c00000000",
            INIT_66 => X"0000006a00000000000000630000000000000091000000000000009800000000",
            INIT_67 => X"0000002800000000000000120000000000000063000000000000008200000000",
            INIT_68 => X"00000059000000000000003b0000000000000042000000000000006100000000",
            INIT_69 => X"000000880000000000000085000000000000006f000000000000006400000000",
            INIT_6A => X"000000910000000000000096000000000000008c000000000000009300000000",
            INIT_6B => X"0000007f00000000000000830000000000000088000000000000008e00000000",
            INIT_6C => X"000000930000000000000088000000000000007b000000000000007d00000000",
            INIT_6D => X"00000088000000000000009c000000000000008e000000000000009700000000",
            INIT_6E => X"00000070000000000000006d0000000000000090000000000000009200000000",
            INIT_6F => X"000000530000000000000032000000000000005c000000000000008200000000",
            INIT_70 => X"0000005f000000000000004b0000000000000048000000000000006900000000",
            INIT_71 => X"000000850000000000000085000000000000005e000000000000006800000000",
            INIT_72 => X"0000008500000000000000800000000000000087000000000000008f00000000",
            INIT_73 => X"0000009800000000000000a00000000000000096000000000000009300000000",
            INIT_74 => X"0000008700000000000000840000000000000090000000000000009100000000",
            INIT_75 => X"000000a500000000000000a2000000000000008a000000000000008a00000000",
            INIT_76 => X"00000077000000000000007e000000000000007f00000000000000a300000000",
            INIT_77 => X"0000004d000000000000003b000000000000005f000000000000007600000000",
            INIT_78 => X"0000005b00000000000000440000000000000044000000000000005e00000000",
            INIT_79 => X"00000083000000000000007b0000000000000062000000000000006500000000",
            INIT_7A => X"0000004f000000000000008a00000000000000c1000000000000009300000000",
            INIT_7B => X"000000a200000000000000930000000000000093000000000000007c00000000",
            INIT_7C => X"00000090000000000000009800000000000000ab00000000000000b400000000",
            INIT_7D => X"000000b300000000000000940000000000000079000000000000009000000000",
            INIT_7E => X"0000007b000000000000008000000000000000a000000000000000b400000000",
            INIT_7F => X"00000054000000000000001a000000000000003f000000000000007000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "sampleifmap_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000004a000000000000004f000000000000005800000000",
            INIT_01 => X"0000008100000000000000780000000000000078000000000000006e00000000",
            INIT_02 => X"0000005700000000000000c000000000000000b8000000000000007800000000",
            INIT_03 => X"000000a600000000000000a4000000000000009c000000000000007200000000",
            INIT_04 => X"000000b600000000000000b700000000000000a1000000000000009a00000000",
            INIT_05 => X"0000008f000000000000009400000000000000ad00000000000000bb00000000",
            INIT_06 => X"0000007c000000000000008e00000000000000c300000000000000b500000000",
            INIT_07 => X"000000760000000000000029000000000000002c000000000000006b00000000",
            INIT_08 => X"0000006000000000000000670000000000000059000000000000005b00000000",
            INIT_09 => X"0000006a000000000000006f0000000000000064000000000000007400000000",
            INIT_0A => X"000000a800000000000000bb0000000000000080000000000000007200000000",
            INIT_0B => X"000000ac00000000000000ac0000000000000099000000000000008c00000000",
            INIT_0C => X"000000a3000000000000009d00000000000000a400000000000000a700000000",
            INIT_0D => X"0000009c00000000000000ab00000000000000a500000000000000a100000000",
            INIT_0E => X"0000007200000000000000a7000000000000009100000000000000a100000000",
            INIT_0F => X"0000005e000000000000002a000000000000004a000000000000006a00000000",
            INIT_10 => X"0000007a00000000000000780000000000000061000000000000006500000000",
            INIT_11 => X"0000005b000000000000005f000000000000004e000000000000007200000000",
            INIT_12 => X"000000cc0000000000000081000000000000006e000000000000007300000000",
            INIT_13 => X"0000009900000000000000a0000000000000008900000000000000a700000000",
            INIT_14 => X"000000b200000000000000aa00000000000000ba00000000000000b300000000",
            INIT_15 => X"000000a500000000000000a2000000000000009c00000000000000b300000000",
            INIT_16 => X"000000480000000000000068000000000000008c000000000000009c00000000",
            INIT_17 => X"0000007200000000000000460000000000000059000000000000005400000000",
            INIT_18 => X"00000060000000000000007a000000000000006b000000000000006e00000000",
            INIT_19 => X"000000640000000000000048000000000000004c000000000000005a00000000",
            INIT_1A => X"0000008c0000000000000057000000000000007f000000000000006d00000000",
            INIT_1B => X"000000b400000000000000a6000000000000009f00000000000000bd00000000",
            INIT_1C => X"000000bc00000000000000be00000000000000ad00000000000000ae00000000",
            INIT_1D => X"000000a100000000000000a2000000000000009900000000000000a200000000",
            INIT_1E => X"0000004a000000000000004b0000000000000095000000000000009900000000",
            INIT_1F => X"0000008a0000000000000070000000000000003e000000000000004200000000",
            INIT_20 => X"0000004e0000000000000059000000000000006a000000000000007700000000",
            INIT_21 => X"00000067000000000000003c0000000000000047000000000000005900000000",
            INIT_22 => X"000000420000000000000072000000000000005f000000000000004b00000000",
            INIT_23 => X"000000be00000000000000ae00000000000000b5000000000000007f00000000",
            INIT_24 => X"000000c100000000000000b800000000000000ab00000000000000ba00000000",
            INIT_25 => X"000000a500000000000000ab00000000000000a000000000000000a400000000",
            INIT_26 => X"0000005c0000000000000068000000000000008b000000000000009200000000",
            INIT_27 => X"000000730000000000000070000000000000005e000000000000004d00000000",
            INIT_28 => X"00000067000000000000003a000000000000005e000000000000007e00000000",
            INIT_29 => X"0000005f0000000000000048000000000000004c000000000000006a00000000",
            INIT_2A => X"0000006300000000000000780000000000000041000000000000005e00000000",
            INIT_2B => X"000000bc00000000000000c400000000000000a1000000000000005b00000000",
            INIT_2C => X"000000a700000000000000a700000000000000c100000000000000b600000000",
            INIT_2D => X"000000a1000000000000009a00000000000000a000000000000000aa00000000",
            INIT_2E => X"00000051000000000000006e000000000000008a000000000000009100000000",
            INIT_2F => X"00000064000000000000006d0000000000000088000000000000006900000000",
            INIT_30 => X"0000006800000000000000460000000000000052000000000000006f00000000",
            INIT_31 => X"000000540000000000000045000000000000005e000000000000007100000000",
            INIT_32 => X"0000007d0000000000000055000000000000006d000000000000007400000000",
            INIT_33 => X"000000c800000000000000ba000000000000009b000000000000007f00000000",
            INIT_34 => X"0000009d00000000000000b100000000000000bb00000000000000bb00000000",
            INIT_35 => X"000000a600000000000000a400000000000000a2000000000000009400000000",
            INIT_36 => X"000000610000000000000079000000000000009500000000000000a200000000",
            INIT_37 => X"0000006100000000000000610000000000000073000000000000007800000000",
            INIT_38 => X"000000b4000000000000008c000000000000005c000000000000006500000000",
            INIT_39 => X"0000004c0000000000000055000000000000007b000000000000009700000000",
            INIT_3A => X"00000054000000000000005a000000000000007c000000000000006700000000",
            INIT_3B => X"000000c800000000000000ad00000000000000af000000000000009200000000",
            INIT_3C => X"0000009f00000000000000ad00000000000000ad00000000000000bc00000000",
            INIT_3D => X"000000ad00000000000000a300000000000000ac000000000000009f00000000",
            INIT_3E => X"000000830000000000000083000000000000008b00000000000000a400000000",
            INIT_3F => X"000000600000000000000064000000000000005f000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000c00000000000000090000000000000007700000000",
            INIT_41 => X"0000006c000000000000007f000000000000009d00000000000000c200000000",
            INIT_42 => X"0000006f000000000000006a000000000000005e000000000000006a00000000",
            INIT_43 => X"000000c500000000000000b000000000000000af000000000000007c00000000",
            INIT_44 => X"000000a500000000000000b000000000000000aa00000000000000b800000000",
            INIT_45 => X"000000a300000000000000af00000000000000c5000000000000009c00000000",
            INIT_46 => X"00000065000000000000007a0000000000000083000000000000009300000000",
            INIT_47 => X"00000066000000000000006b0000000000000060000000000000006400000000",
            INIT_48 => X"000000a9000000000000008a0000000000000074000000000000006e00000000",
            INIT_49 => X"0000008800000000000000a000000000000000c400000000000000c500000000",
            INIT_4A => X"0000008a000000000000005c0000000000000063000000000000008100000000",
            INIT_4B => X"000000a900000000000000b4000000000000009f000000000000009200000000",
            INIT_4C => X"000000b200000000000000af000000000000008d000000000000008e00000000",
            INIT_4D => X"0000009700000000000000b300000000000000bc00000000000000a600000000",
            INIT_4E => X"0000003a0000000000000070000000000000009a000000000000008f00000000",
            INIT_4F => X"0000004900000000000000660000000000000065000000000000005b00000000",
            INIT_50 => X"0000006b000000000000004a0000000000000057000000000000005b00000000",
            INIT_51 => X"000000a300000000000000bf00000000000000b900000000000000a500000000",
            INIT_52 => X"00000066000000000000006a0000000000000080000000000000008600000000",
            INIT_53 => X"0000007400000000000000920000000000000084000000000000007600000000",
            INIT_54 => X"000000b600000000000000a10000000000000063000000000000004d00000000",
            INIT_55 => X"000000a700000000000000ad000000000000009f00000000000000b700000000",
            INIT_56 => X"0000002b000000000000005e0000000000000087000000000000009c00000000",
            INIT_57 => X"0000004d0000000000000044000000000000005c000000000000005b00000000",
            INIT_58 => X"0000002c0000000000000032000000000000005f000000000000005100000000",
            INIT_59 => X"000000bb00000000000000a60000000000000094000000000000005f00000000",
            INIT_5A => X"00000072000000000000007e000000000000009000000000000000ae00000000",
            INIT_5B => X"0000006b00000000000000770000000000000072000000000000006800000000",
            INIT_5C => X"000000b6000000000000009d0000000000000052000000000000005100000000",
            INIT_5D => X"0000009600000000000000a900000000000000b200000000000000a900000000",
            INIT_5E => X"0000003f000000000000002c000000000000006c000000000000009800000000",
            INIT_5F => X"0000005600000000000000500000000000000045000000000000006100000000",
            INIT_60 => X"000000150000000000000034000000000000005f000000000000005a00000000",
            INIT_61 => X"000000b00000000000000092000000000000006d000000000000001c00000000",
            INIT_62 => X"0000007f000000000000008e00000000000000b500000000000000ca00000000",
            INIT_63 => X"0000008200000000000000720000000000000077000000000000007800000000",
            INIT_64 => X"000000a900000000000000900000000000000076000000000000008100000000",
            INIT_65 => X"0000009800000000000000b400000000000000ad000000000000009f00000000",
            INIT_66 => X"00000055000000000000002c0000000000000044000000000000007700000000",
            INIT_67 => X"0000006a00000000000000a70000000000000072000000000000003300000000",
            INIT_68 => X"000000340000000000000039000000000000005b000000000000005f00000000",
            INIT_69 => X"0000009c00000000000000770000000000000031000000000000001800000000",
            INIT_6A => X"0000009b00000000000000ba00000000000000cb00000000000000bb00000000",
            INIT_6B => X"0000007500000000000000740000000000000085000000000000008d00000000",
            INIT_6C => X"00000099000000000000008b0000000000000077000000000000006d00000000",
            INIT_6D => X"0000007d000000000000009c00000000000000a7000000000000009f00000000",
            INIT_6E => X"0000004000000000000000440000000000000041000000000000006500000000",
            INIT_6F => X"0000007a00000000000000aa0000000000000090000000000000003700000000",
            INIT_70 => X"000000490000000000000020000000000000004b000000000000005e00000000",
            INIT_71 => X"0000007300000000000000360000000000000021000000000000002e00000000",
            INIT_72 => X"000000c200000000000000c300000000000000b0000000000000009600000000",
            INIT_73 => X"000000920000000000000088000000000000009b00000000000000b100000000",
            INIT_74 => X"00000077000000000000005e0000000000000065000000000000008b00000000",
            INIT_75 => X"000000690000000000000060000000000000005f000000000000006500000000",
            INIT_76 => X"0000006d000000000000006b0000000000000076000000000000008300000000",
            INIT_77 => X"0000006a000000000000009a000000000000008f000000000000008000000000",
            INIT_78 => X"0000004c00000000000000180000000000000023000000000000004e00000000",
            INIT_79 => X"0000003b000000000000001b0000000000000028000000000000004100000000",
            INIT_7A => X"000000b000000000000000960000000000000088000000000000007800000000",
            INIT_7B => X"000000ba00000000000000a500000000000000b700000000000000c000000000",
            INIT_7C => X"00000056000000000000006b00000000000000aa00000000000000cf00000000",
            INIT_7D => X"0000008c00000000000000700000000000000055000000000000004200000000",
            INIT_7E => X"000000890000000000000089000000000000009500000000000000a900000000",
            INIT_7F => X"00000080000000000000009a000000000000008f000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "sampleifmap_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000000000400000000000000051000000000000004400000000",
            INIT_01 => X"00000050000000000000004b0000000000000039000000000000002100000000",
            INIT_02 => X"0000002200000000000000140000000000000046000000000000005300000000",
            INIT_03 => X"000000420000000000000046000000000000004b000000000000004700000000",
            INIT_04 => X"00000079000000000000007c0000000000000078000000000000005700000000",
            INIT_05 => X"000000520000000000000054000000000000006c000000000000007e00000000",
            INIT_06 => X"0000005b000000000000003b0000000000000081000000000000008800000000",
            INIT_07 => X"00000057000000000000004c0000000000000043000000000000006000000000",
            INIT_08 => X"0000002f000000000000004a0000000000000066000000000000005000000000",
            INIT_09 => X"000000540000000000000054000000000000005c000000000000003800000000",
            INIT_0A => X"000000300000000000000012000000000000003e000000000000005800000000",
            INIT_0B => X"00000049000000000000004d000000000000005c000000000000005d00000000",
            INIT_0C => X"0000006a000000000000006f0000000000000075000000000000006b00000000",
            INIT_0D => X"00000053000000000000004d000000000000006c000000000000007500000000",
            INIT_0E => X"00000041000000000000002d000000000000008b000000000000009700000000",
            INIT_0F => X"00000051000000000000005a0000000000000042000000000000004700000000",
            INIT_10 => X"000000380000000000000058000000000000006d000000000000005f00000000",
            INIT_11 => X"0000005a00000000000000560000000000000069000000000000005400000000",
            INIT_12 => X"0000003c00000000000000140000000000000035000000000000005c00000000",
            INIT_13 => X"0000003c00000000000000420000000000000058000000000000005900000000",
            INIT_14 => X"00000054000000000000004e0000000000000066000000000000006700000000",
            INIT_15 => X"0000005600000000000000420000000000000072000000000000007200000000",
            INIT_16 => X"000000370000000000000023000000000000008f000000000000009e00000000",
            INIT_17 => X"0000003b00000000000000620000000000000062000000000000005400000000",
            INIT_18 => X"0000004900000000000000640000000000000064000000000000007400000000",
            INIT_19 => X"0000006000000000000000580000000000000066000000000000006d00000000",
            INIT_1A => X"00000038000000000000001a000000000000002d000000000000005e00000000",
            INIT_1B => X"0000003700000000000000360000000000000043000000000000004100000000",
            INIT_1C => X"0000006200000000000000610000000000000075000000000000006a00000000",
            INIT_1D => X"0000005b00000000000000450000000000000072000000000000007600000000",
            INIT_1E => X"0000005d0000000000000040000000000000009600000000000000a000000000",
            INIT_1F => X"00000032000000000000005e000000000000007e000000000000007800000000",
            INIT_20 => X"0000005d00000000000000800000000000000068000000000000007800000000",
            INIT_21 => X"0000005e000000000000005a000000000000005e000000000000007200000000",
            INIT_22 => X"00000024000000000000001a0000000000000027000000000000005d00000000",
            INIT_23 => X"0000005600000000000000490000000000000037000000000000002f00000000",
            INIT_24 => X"00000065000000000000006b0000000000000071000000000000006900000000",
            INIT_25 => X"00000067000000000000004a000000000000006d000000000000006700000000",
            INIT_26 => X"00000074000000000000007000000000000000ac00000000000000a200000000",
            INIT_27 => X"0000006c00000000000000670000000000000084000000000000008100000000",
            INIT_28 => X"0000006200000000000000620000000000000066000000000000006900000000",
            INIT_29 => X"0000004e000000000000005b0000000000000059000000000000005f00000000",
            INIT_2A => X"0000002b000000000000001b0000000000000023000000000000005800000000",
            INIT_2B => X"0000006c000000000000006a000000000000005d000000000000004d00000000",
            INIT_2C => X"0000004e00000000000000640000000000000065000000000000006700000000",
            INIT_2D => X"000000660000000000000062000000000000006e000000000000003900000000",
            INIT_2E => X"0000007f000000000000008200000000000000ba00000000000000a700000000",
            INIT_2F => X"0000007800000000000000840000000000000090000000000000008100000000",
            INIT_30 => X"0000004f00000000000000300000000000000060000000000000005e00000000",
            INIT_31 => X"0000003f000000000000005d0000000000000064000000000000005a00000000",
            INIT_32 => X"0000005a0000000000000026000000000000001d000000000000004a00000000",
            INIT_33 => X"0000006300000000000000820000000000000081000000000000007e00000000",
            INIT_34 => X"0000003900000000000000730000000000000047000000000000003a00000000",
            INIT_35 => X"0000006a0000000000000071000000000000007b000000000000002500000000",
            INIT_36 => X"0000008c000000000000008d00000000000000c100000000000000b700000000",
            INIT_37 => X"0000003b000000000000006500000000000000a0000000000000008900000000",
            INIT_38 => X"00000069000000000000002f0000000000000054000000000000005600000000",
            INIT_39 => X"00000047000000000000005e0000000000000061000000000000006700000000",
            INIT_3A => X"0000008b00000000000000490000000000000014000000000000003800000000",
            INIT_3B => X"000000290000000000000072000000000000008c000000000000008a00000000",
            INIT_3C => X"0000004f00000000000000730000000000000041000000000000001a00000000",
            INIT_3D => X"0000008c0000000000000078000000000000007d000000000000003b00000000",
            INIT_3E => X"00000094000000000000009600000000000000c300000000000000b000000000",
            INIT_3F => X"00000018000000000000003f000000000000009b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c000000000000004a000000000000004e000000000000006200000000",
            INIT_41 => X"0000005c00000000000000500000000000000072000000000000009500000000",
            INIT_42 => X"000000900000000000000071000000000000002c000000000000004700000000",
            INIT_43 => X"00000017000000000000003f0000000000000086000000000000008800000000",
            INIT_44 => X"00000056000000000000005e000000000000007c000000000000004500000000",
            INIT_45 => X"000000a5000000000000009b000000000000008b000000000000007000000000",
            INIT_46 => X"00000096000000000000009600000000000000b100000000000000aa00000000",
            INIT_47 => X"000000160000000000000029000000000000008e000000000000009200000000",
            INIT_48 => X"00000094000000000000004e0000000000000051000000000000007400000000",
            INIT_49 => X"000000450000000000000054000000000000009b00000000000000a300000000",
            INIT_4A => X"0000008e0000000000000089000000000000005a000000000000005100000000",
            INIT_4B => X"000000380000000000000021000000000000005d000000000000008a00000000",
            INIT_4C => X"000000800000000000000073000000000000008f000000000000007c00000000",
            INIT_4D => X"00000081000000000000009c000000000000009c000000000000009700000000",
            INIT_4E => X"0000009a000000000000009800000000000000ad00000000000000a700000000",
            INIT_4F => X"0000001800000000000000160000000000000079000000000000009400000000",
            INIT_50 => X"000000910000000000000049000000000000004f000000000000007800000000",
            INIT_51 => X"00000041000000000000007f00000000000000a600000000000000a500000000",
            INIT_52 => X"0000007f000000000000008e0000000000000072000000000000003600000000",
            INIT_53 => X"0000006c0000000000000047000000000000005d000000000000007e00000000",
            INIT_54 => X"000000a100000000000000920000000000000085000000000000008700000000",
            INIT_55 => X"00000057000000000000007500000000000000a5000000000000009c00000000",
            INIT_56 => X"0000009c000000000000009700000000000000af00000000000000a900000000",
            INIT_57 => X"0000001700000000000000130000000000000074000000000000009100000000",
            INIT_58 => X"0000008a00000000000000420000000000000045000000000000007b00000000",
            INIT_59 => X"0000005f00000000000000a500000000000000a800000000000000a100000000",
            INIT_5A => X"00000070000000000000008a000000000000008c000000000000004b00000000",
            INIT_5B => X"000000a200000000000000880000000000000066000000000000006d00000000",
            INIT_5C => X"000000870000000000000097000000000000009a000000000000009900000000",
            INIT_5D => X"0000008800000000000000760000000000000085000000000000007c00000000",
            INIT_5E => X"0000009d000000000000009200000000000000aa00000000000000bd00000000",
            INIT_5F => X"0000000b00000000000000140000000000000077000000000000009400000000",
            INIT_60 => X"00000079000000000000003c0000000000000039000000000000006a00000000",
            INIT_61 => X"0000009800000000000000ad00000000000000a4000000000000008700000000",
            INIT_62 => X"00000076000000000000007f0000000000000093000000000000009000000000",
            INIT_63 => X"0000008b0000000000000066000000000000005c000000000000007300000000",
            INIT_64 => X"000000740000000000000085000000000000008a000000000000008d00000000",
            INIT_65 => X"000000880000000000000077000000000000006b000000000000007800000000",
            INIT_66 => X"00000091000000000000008700000000000000ae00000000000000b000000000",
            INIT_67 => X"0000002b000000000000001a000000000000007200000000000000a100000000",
            INIT_68 => X"00000074000000000000004e0000000000000055000000000000007400000000",
            INIT_69 => X"000000ab00000000000000ac000000000000008c000000000000007f00000000",
            INIT_6A => X"000000780000000000000082000000000000007c000000000000009900000000",
            INIT_6B => X"0000006e00000000000000710000000000000076000000000000007700000000",
            INIT_6C => X"0000007d0000000000000077000000000000006c000000000000006900000000",
            INIT_6D => X"000000750000000000000081000000000000007a000000000000008300000000",
            INIT_6E => X"0000009a000000000000008d00000000000000a2000000000000009000000000",
            INIT_6F => X"0000005f0000000000000041000000000000007000000000000000a600000000",
            INIT_70 => X"0000007800000000000000630000000000000060000000000000008400000000",
            INIT_71 => X"000000a800000000000000a50000000000000072000000000000008200000000",
            INIT_72 => X"000000700000000000000068000000000000006b000000000000008b00000000",
            INIT_73 => X"00000084000000000000008e0000000000000081000000000000007c00000000",
            INIT_74 => X"0000006f000000000000006b0000000000000077000000000000007a00000000",
            INIT_75 => X"00000090000000000000008d0000000000000076000000000000007300000000",
            INIT_76 => X"0000009f0000000000000092000000000000007b000000000000008e00000000",
            INIT_77 => X"0000005e00000000000000480000000000000070000000000000009d00000000",
            INIT_78 => X"00000076000000000000005d000000000000005a000000000000007900000000",
            INIT_79 => X"000000a60000000000000097000000000000007c000000000000007f00000000",
            INIT_7A => X"00000045000000000000007900000000000000ab000000000000009900000000",
            INIT_7B => X"0000008b000000000000007b000000000000007c000000000000006b00000000",
            INIT_7C => X"0000007700000000000000800000000000000090000000000000009b00000000",
            INIT_7D => X"000000a700000000000000830000000000000067000000000000007a00000000",
            INIT_7E => X"000000a00000000000000080000000000000008c000000000000009f00000000",
            INIT_7F => X"000000680000000000000022000000000000004b000000000000009500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "sampleifmap_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e00000000000000640000000000000064000000000000007000000000",
            INIT_01 => X"000000a300000000000000950000000000000098000000000000008d00000000",
            INIT_02 => X"0000004700000000000000a600000000000000a3000000000000008a00000000",
            INIT_03 => X"0000008d000000000000008b0000000000000085000000000000006400000000",
            INIT_04 => X"0000009e00000000000000a00000000000000088000000000000008100000000",
            INIT_05 => X"0000007e000000000000007d000000000000009700000000000000a300000000",
            INIT_06 => X"0000008f000000000000007a00000000000000b100000000000000a900000000",
            INIT_07 => X"0000008b0000000000000033000000000000003d000000000000008f00000000",
            INIT_08 => X"0000008100000000000000830000000000000070000000000000007000000000",
            INIT_09 => X"000000890000000000000090000000000000007c000000000000009300000000",
            INIT_0A => X"0000009900000000000000a80000000000000079000000000000008f00000000",
            INIT_0B => X"000000930000000000000092000000000000007f000000000000007a00000000",
            INIT_0C => X"0000008a0000000000000084000000000000008b000000000000008d00000000",
            INIT_0D => X"000000860000000000000099000000000000008f000000000000008600000000",
            INIT_0E => X"0000007a00000000000000920000000000000082000000000000009100000000",
            INIT_0F => X"0000006f000000000000003a0000000000000064000000000000008600000000",
            INIT_10 => X"0000008e00000000000000950000000000000076000000000000007900000000",
            INIT_11 => X"00000076000000000000007b0000000000000061000000000000008d00000000",
            INIT_12 => X"000000bb0000000000000079000000000000007e000000000000008f00000000",
            INIT_13 => X"000000820000000000000088000000000000006e000000000000009100000000",
            INIT_14 => X"0000009a000000000000009400000000000000a1000000000000009a00000000",
            INIT_15 => X"0000009100000000000000960000000000000086000000000000009700000000",
            INIT_16 => X"000000570000000000000061000000000000007b000000000000008600000000",
            INIT_17 => X"0000008600000000000000610000000000000077000000000000006700000000",
            INIT_18 => X"0000006f00000000000000970000000000000087000000000000008800000000",
            INIT_19 => X"0000007d000000000000005d0000000000000065000000000000007a00000000",
            INIT_1A => X"0000007d00000000000000600000000000000099000000000000008600000000",
            INIT_1B => X"000000a00000000000000092000000000000008800000000000000a900000000",
            INIT_1C => X"000000a700000000000000a60000000000000094000000000000009600000000",
            INIT_1D => X"0000009100000000000000900000000000000080000000000000008d00000000",
            INIT_1E => X"0000005e000000000000004b0000000000000082000000000000008400000000",
            INIT_1F => X"000000a900000000000000950000000000000057000000000000005300000000",
            INIT_20 => X"0000005e0000000000000070000000000000008c000000000000009400000000",
            INIT_21 => X"0000008200000000000000540000000000000068000000000000007900000000",
            INIT_22 => X"0000004a000000000000008d0000000000000074000000000000006600000000",
            INIT_23 => X"000000aa000000000000009b00000000000000a3000000000000007600000000",
            INIT_24 => X"000000a7000000000000009d000000000000009500000000000000a500000000",
            INIT_25 => X"0000009100000000000000930000000000000089000000000000009200000000",
            INIT_26 => X"00000071000000000000006d000000000000007c000000000000007f00000000",
            INIT_27 => X"000000a1000000000000009c0000000000000077000000000000006000000000",
            INIT_28 => X"0000007d00000000000000480000000000000077000000000000009800000000",
            INIT_29 => X"0000007900000000000000630000000000000065000000000000008100000000",
            INIT_2A => X"0000007d000000000000009a000000000000005b000000000000007800000000",
            INIT_2B => X"000000a900000000000000b50000000000000096000000000000005d00000000",
            INIT_2C => X"0000008f000000000000009100000000000000ad00000000000000a200000000",
            INIT_2D => X"0000008b00000000000000810000000000000087000000000000008f00000000",
            INIT_2E => X"0000006600000000000000750000000000000078000000000000007d00000000",
            INIT_2F => X"00000099000000000000009a00000000000000ab000000000000008100000000",
            INIT_30 => X"0000007b00000000000000520000000000000068000000000000008800000000",
            INIT_31 => X"0000007300000000000000620000000000000076000000000000008800000000",
            INIT_32 => X"000000940000000000000075000000000000008d000000000000009600000000",
            INIT_33 => X"000000b300000000000000ad0000000000000095000000000000008100000000",
            INIT_34 => X"0000008f000000000000009f00000000000000a800000000000000a500000000",
            INIT_35 => X"0000008d000000000000008c000000000000008b000000000000007e00000000",
            INIT_36 => X"0000006d000000000000007a0000000000000085000000000000008800000000",
            INIT_37 => X"00000095000000000000009600000000000000a4000000000000009800000000",
            INIT_38 => X"000000bf0000000000000096000000000000006f000000000000007d00000000",
            INIT_39 => X"0000006f0000000000000079000000000000009e00000000000000ac00000000",
            INIT_3A => X"0000006900000000000000730000000000000099000000000000009100000000",
            INIT_3B => X"000000ac000000000000009a00000000000000a1000000000000009400000000",
            INIT_3C => X"0000008d000000000000009c000000000000009b00000000000000a100000000",
            INIT_3D => X"0000008f00000000000000880000000000000093000000000000008900000000",
            INIT_3E => X"00000086000000000000007b000000000000008c000000000000008900000000",
            INIT_3F => X"00000095000000000000009e0000000000000095000000000000009c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000dc00000000000000c800000000000000a2000000000000009500000000",
            INIT_41 => X"0000009300000000000000aa00000000000000bd00000000000000d100000000",
            INIT_42 => X"00000088000000000000007d000000000000007a000000000000009100000000",
            INIT_43 => X"000000a40000000000000096000000000000009f000000000000008b00000000",
            INIT_44 => X"0000008e000000000000009f000000000000009b000000000000009b00000000",
            INIT_45 => X"00000088000000000000009300000000000000a9000000000000008500000000",
            INIT_46 => X"00000072000000000000006b000000000000007e000000000000007f00000000",
            INIT_47 => X"0000009c00000000000000a0000000000000008f000000000000009a00000000",
            INIT_48 => X"000000be000000000000009d0000000000000089000000000000008b00000000",
            INIT_49 => X"000000b000000000000000bf00000000000000d700000000000000d500000000",
            INIT_4A => X"000000a30000000000000075000000000000008400000000000000a900000000",
            INIT_4B => X"0000008f000000000000009a000000000000009700000000000000ad00000000",
            INIT_4C => X"0000009800000000000000990000000000000081000000000000007c00000000",
            INIT_4D => X"0000007c000000000000009500000000000000a3000000000000009100000000",
            INIT_4E => X"0000004a00000000000000600000000000000083000000000000007700000000",
            INIT_4F => X"0000007800000000000000970000000000000095000000000000009100000000",
            INIT_50 => X"000000860000000000000061000000000000006f000000000000007300000000",
            INIT_51 => X"000000c100000000000000d300000000000000cf00000000000000bf00000000",
            INIT_52 => X"0000007f000000000000009100000000000000ad00000000000000b100000000",
            INIT_53 => X"000000680000000000000086000000000000008f000000000000009000000000",
            INIT_54 => X"0000009b000000000000008b000000000000005c000000000000004900000000",
            INIT_55 => X"0000008e0000000000000094000000000000008a00000000000000a100000000",
            INIT_56 => X"0000003c00000000000000550000000000000075000000000000008300000000",
            INIT_57 => X"0000006d000000000000006f0000000000000091000000000000009200000000",
            INIT_58 => X"0000004000000000000000410000000000000072000000000000006a00000000",
            INIT_59 => X"000000d500000000000000c300000000000000b2000000000000007800000000",
            INIT_5A => X"0000009900000000000000ad00000000000000b900000000000000ca00000000",
            INIT_5B => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_5C => X"0000009a000000000000008e0000000000000060000000000000006c00000000",
            INIT_5D => X"0000007f000000000000009500000000000000a1000000000000009000000000",
            INIT_5E => X"0000006100000000000000310000000000000062000000000000008300000000",
            INIT_5F => X"000000750000000000000076000000000000006c000000000000009300000000",
            INIT_60 => X"00000026000000000000003e0000000000000070000000000000007400000000",
            INIT_61 => X"000000c700000000000000b40000000000000087000000000000002900000000",
            INIT_62 => X"000000b200000000000000b700000000000000cc00000000000000d400000000",
            INIT_63 => X"000000a1000000000000009e00000000000000a400000000000000ab00000000",
            INIT_64 => X"0000008d0000000000000087000000000000008b000000000000009d00000000",
            INIT_65 => X"0000007e000000000000009c0000000000000099000000000000008700000000",
            INIT_66 => X"0000007c000000000000003b0000000000000042000000000000006700000000",
            INIT_67 => X"0000008300000000000000c50000000000000088000000000000005400000000",
            INIT_68 => X"0000004e000000000000004f000000000000007b000000000000007f00000000",
            INIT_69 => X"000000bf00000000000000950000000000000042000000000000002500000000",
            INIT_6A => X"000000c200000000000000d600000000000000db00000000000000d000000000",
            INIT_6B => X"0000009f00000000000000a500000000000000b400000000000000b800000000",
            INIT_6C => X"00000083000000000000007b000000000000007d000000000000008700000000",
            INIT_6D => X"0000007200000000000000870000000000000093000000000000008a00000000",
            INIT_6E => X"0000005b0000000000000055000000000000004f000000000000006c00000000",
            INIT_6F => X"0000008f00000000000000c900000000000000ac000000000000004e00000000",
            INIT_70 => X"0000006b00000000000000340000000000000068000000000000007d00000000",
            INIT_71 => X"00000097000000000000004e0000000000000030000000000000004300000000",
            INIT_72 => X"000000da00000000000000d900000000000000cb00000000000000bd00000000",
            INIT_73 => X"000000b600000000000000b400000000000000c300000000000000cd00000000",
            INIT_74 => X"0000007a000000000000005e000000000000007400000000000000a500000000",
            INIT_75 => X"0000006f00000000000000590000000000000059000000000000006100000000",
            INIT_76 => X"000000860000000000000082000000000000008a000000000000009600000000",
            INIT_77 => X"0000008100000000000000bc00000000000000b5000000000000009f00000000",
            INIT_78 => X"0000007300000000000000280000000000000033000000000000006600000000",
            INIT_79 => X"0000004e0000000000000029000000000000003a000000000000006000000000",
            INIT_7A => X"000000cf00000000000000b900000000000000b500000000000000a000000000",
            INIT_7B => X"000000ce00000000000000c400000000000000d200000000000000da00000000",
            INIT_7C => X"00000071000000000000007c00000000000000b400000000000000d600000000",
            INIT_7D => X"000000a000000000000000840000000000000066000000000000005600000000",
            INIT_7E => X"000000a700000000000000a700000000000000a700000000000000ba00000000",
            INIT_7F => X"0000009c00000000000000b900000000000000b300000000000000b400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "sampleifmap_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000002e0000000000000040000000000000003200000000",
            INIT_01 => X"0000003900000000000000370000000000000024000000000000001600000000",
            INIT_02 => X"00000012000000000000000c0000000000000036000000000000003b00000000",
            INIT_03 => X"000000320000000000000031000000000000002c000000000000002b00000000",
            INIT_04 => X"0000004d0000000000000051000000000000004d000000000000003a00000000",
            INIT_05 => X"000000390000000000000038000000000000004e000000000000005300000000",
            INIT_06 => X"0000003a000000000000001f000000000000005d000000000000006100000000",
            INIT_07 => X"0000004200000000000000350000000000000029000000000000004100000000",
            INIT_08 => X"0000001d00000000000000390000000000000051000000000000003a00000000",
            INIT_09 => X"0000003c000000000000003b000000000000003d000000000000002300000000",
            INIT_0A => X"0000001b0000000000000007000000000000002f000000000000004000000000",
            INIT_0B => X"0000002f000000000000003b000000000000003e000000000000003800000000",
            INIT_0C => X"00000044000000000000004a000000000000004a000000000000004400000000",
            INIT_0D => X"0000003c00000000000000330000000000000051000000000000004e00000000",
            INIT_0E => X"0000002700000000000000150000000000000060000000000000006f00000000",
            INIT_0F => X"000000420000000000000045000000000000002c000000000000002d00000000",
            INIT_10 => X"0000002300000000000000460000000000000057000000000000004800000000",
            INIT_11 => X"00000041000000000000003c0000000000000048000000000000003500000000",
            INIT_12 => X"0000002300000000000000070000000000000026000000000000004500000000",
            INIT_13 => X"0000002100000000000000300000000000000041000000000000003400000000",
            INIT_14 => X"0000003700000000000000320000000000000042000000000000004300000000",
            INIT_15 => X"0000003e000000000000002d0000000000000052000000000000004d00000000",
            INIT_16 => X"0000002600000000000000100000000000000063000000000000007400000000",
            INIT_17 => X"00000033000000000000004d000000000000004b000000000000003f00000000",
            INIT_18 => X"0000002f0000000000000050000000000000004c000000000000005e00000000",
            INIT_19 => X"0000004a00000000000000410000000000000048000000000000004700000000",
            INIT_1A => X"00000022000000000000000c000000000000001e000000000000004800000000",
            INIT_1B => X"0000001e00000000000000230000000000000034000000000000002800000000",
            INIT_1C => X"0000004500000000000000440000000000000057000000000000004b00000000",
            INIT_1D => X"00000043000000000000002e000000000000004d000000000000005100000000",
            INIT_1E => X"00000049000000000000002a000000000000006b000000000000007700000000",
            INIT_1F => X"0000002200000000000000440000000000000060000000000000005f00000000",
            INIT_20 => X"0000003c000000000000006a000000000000004f000000000000006100000000",
            INIT_21 => X"0000004c00000000000000480000000000000044000000000000004b00000000",
            INIT_22 => X"00000011000000000000000c0000000000000018000000000000004900000000",
            INIT_23 => X"0000003b00000000000000330000000000000025000000000000001c00000000",
            INIT_24 => X"00000047000000000000004b000000000000004f000000000000004800000000",
            INIT_25 => X"0000004d000000000000002d0000000000000049000000000000004700000000",
            INIT_26 => X"0000005500000000000000520000000000000081000000000000008000000000",
            INIT_27 => X"0000005000000000000000490000000000000061000000000000005e00000000",
            INIT_28 => X"00000043000000000000004b000000000000004d000000000000005200000000",
            INIT_29 => X"0000003d000000000000004d0000000000000045000000000000003d00000000",
            INIT_2A => X"00000016000000000000000d0000000000000013000000000000004300000000",
            INIT_2B => X"000000490000000000000047000000000000003b000000000000002c00000000",
            INIT_2C => X"0000003500000000000000490000000000000048000000000000004800000000",
            INIT_2D => X"0000004d000000000000003e0000000000000049000000000000002200000000",
            INIT_2E => X"0000005b00000000000000600000000000000093000000000000008800000000",
            INIT_2F => X"0000005c0000000000000068000000000000006e000000000000005c00000000",
            INIT_30 => X"0000003300000000000000190000000000000046000000000000004800000000",
            INIT_31 => X"00000032000000000000004f000000000000004f000000000000003e00000000",
            INIT_32 => X"000000360000000000000018000000000000000f000000000000003800000000",
            INIT_33 => X"0000003e000000000000004d000000000000004b000000000000004900000000",
            INIT_34 => X"0000002a00000000000000600000000000000033000000000000002200000000",
            INIT_35 => X"0000004a00000000000000480000000000000058000000000000001600000000",
            INIT_36 => X"0000006c000000000000006800000000000000a1000000000000009500000000",
            INIT_37 => X"0000002b00000000000000510000000000000083000000000000006b00000000",
            INIT_38 => X"000000460000000000000015000000000000003b000000000000003f00000000",
            INIT_39 => X"0000003a000000000000004b0000000000000048000000000000004d00000000",
            INIT_3A => X"00000051000000000000002f0000000000000008000000000000002900000000",
            INIT_3B => X"00000012000000000000003e000000000000004b000000000000004b00000000",
            INIT_3C => X"0000004000000000000000590000000000000027000000000000000600000000",
            INIT_3D => X"000000530000000000000048000000000000005e000000000000002a00000000",
            INIT_3E => X"00000078000000000000007200000000000000a2000000000000008300000000",
            INIT_3F => X"0000001500000000000000340000000000000085000000000000007600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006800000000000000310000000000000035000000000000004900000000",
            INIT_41 => X"0000004600000000000000390000000000000058000000000000007900000000",
            INIT_42 => X"0000005300000000000000470000000000000017000000000000003300000000",
            INIT_43 => X"000000070000000000000022000000000000004f000000000000004e00000000",
            INIT_44 => X"0000003e000000000000003c0000000000000051000000000000002800000000",
            INIT_45 => X"0000005d000000000000005b0000000000000063000000000000005000000000",
            INIT_46 => X"000000790000000000000078000000000000008d000000000000007300000000",
            INIT_47 => X"000000140000000000000021000000000000007c000000000000007900000000",
            INIT_48 => X"000000760000000000000038000000000000003a000000000000005600000000",
            INIT_49 => X"000000330000000000000040000000000000007f000000000000008300000000",
            INIT_4A => X"0000006300000000000000610000000000000040000000000000003b00000000",
            INIT_4B => X"0000001c000000000000000d000000000000003a000000000000005e00000000",
            INIT_4C => X"000000500000000000000049000000000000005d000000000000005300000000",
            INIT_4D => X"0000004a000000000000005f0000000000000069000000000000006200000000",
            INIT_4E => X"0000007e00000000000000770000000000000084000000000000007400000000",
            INIT_4F => X"00000017000000000000000d0000000000000065000000000000007f00000000",
            INIT_50 => X"000000740000000000000035000000000000003b000000000000005b00000000",
            INIT_51 => X"0000003000000000000000670000000000000087000000000000008400000000",
            INIT_52 => X"000000610000000000000060000000000000004b000000000000002000000000",
            INIT_53 => X"000000490000000000000032000000000000004a000000000000006600000000",
            INIT_54 => X"0000006100000000000000590000000000000052000000000000005a00000000",
            INIT_55 => X"000000310000000000000047000000000000006c000000000000006200000000",
            INIT_56 => X"0000008a0000000000000077000000000000007c000000000000007700000000",
            INIT_57 => X"00000014000000000000000a000000000000005b000000000000007b00000000",
            INIT_58 => X"0000006e000000000000002f0000000000000033000000000000006500000000",
            INIT_59 => X"0000004800000000000000870000000000000087000000000000008100000000",
            INIT_5A => X"0000004f00000000000000520000000000000054000000000000002e00000000",
            INIT_5B => X"0000008700000000000000750000000000000056000000000000005e00000000",
            INIT_5C => X"0000005e000000000000005d0000000000000066000000000000007800000000",
            INIT_5D => X"00000058000000000000004a0000000000000058000000000000005c00000000",
            INIT_5E => X"0000008d00000000000000760000000000000073000000000000008400000000",
            INIT_5F => X"00000007000000000000000b000000000000005b000000000000007700000000",
            INIT_60 => X"0000006000000000000000280000000000000028000000000000005800000000",
            INIT_61 => X"00000077000000000000008b0000000000000083000000000000006b00000000",
            INIT_62 => X"0000005900000000000000570000000000000066000000000000006b00000000",
            INIT_63 => X"0000006c0000000000000051000000000000004a000000000000005f00000000",
            INIT_64 => X"0000005d0000000000000064000000000000006e000000000000007600000000",
            INIT_65 => X"0000005f00000000000000570000000000000055000000000000006600000000",
            INIT_66 => X"0000007100000000000000650000000000000078000000000000007c00000000",
            INIT_67 => X"00000020000000000000000f0000000000000059000000000000007b00000000",
            INIT_68 => X"0000005c0000000000000037000000000000003f000000000000005f00000000",
            INIT_69 => X"00000089000000000000008b000000000000006e000000000000006400000000",
            INIT_6A => X"0000005c00000000000000650000000000000061000000000000007b00000000",
            INIT_6B => X"0000005600000000000000560000000000000058000000000000005a00000000",
            INIT_6C => X"0000006c00000000000000640000000000000058000000000000005500000000",
            INIT_6D => X"0000005f000000000000006e000000000000006c000000000000007200000000",
            INIT_6E => X"00000073000000000000006b0000000000000075000000000000006d00000000",
            INIT_6F => X"0000004c00000000000000310000000000000058000000000000008000000000",
            INIT_70 => X"0000006000000000000000470000000000000045000000000000006a00000000",
            INIT_71 => X"0000008700000000000000860000000000000056000000000000006800000000",
            INIT_72 => X"0000005800000000000000510000000000000057000000000000007400000000",
            INIT_73 => X"0000006a000000000000006e0000000000000060000000000000006000000000",
            INIT_74 => X"0000005c0000000000000057000000000000005f000000000000006200000000",
            INIT_75 => X"00000080000000000000007f000000000000006b000000000000006100000000",
            INIT_76 => X"000000770000000000000074000000000000005e000000000000007a00000000",
            INIT_77 => X"000000460000000000000035000000000000005c000000000000007a00000000",
            INIT_78 => X"0000005c00000000000000400000000000000040000000000000006000000000",
            INIT_79 => X"000000850000000000000079000000000000005f000000000000006700000000",
            INIT_7A => X"0000003300000000000000640000000000000096000000000000008100000000",
            INIT_7B => X"0000007100000000000000620000000000000065000000000000005800000000",
            INIT_7C => X"0000005f00000000000000650000000000000077000000000000008300000000",
            INIT_7D => X"0000009800000000000000710000000000000053000000000000006000000000",
            INIT_7E => X"0000007c00000000000000620000000000000078000000000000009400000000",
            INIT_7F => X"00000048000000000000000d0000000000000039000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "sampleifmap_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005a0000000000000047000000000000004c000000000000005700000000",
            INIT_01 => X"000000820000000000000078000000000000007c000000000000007300000000",
            INIT_02 => X"0000003a0000000000000096000000000000008e000000000000006e00000000",
            INIT_03 => X"0000007800000000000000770000000000000074000000000000005400000000",
            INIT_04 => X"0000008600000000000000850000000000000071000000000000006c00000000",
            INIT_05 => X"0000006e0000000000000067000000000000007e000000000000008900000000",
            INIT_06 => X"00000072000000000000006300000000000000a3000000000000009f00000000",
            INIT_07 => X"0000006b0000000000000021000000000000002a000000000000007500000000",
            INIT_08 => X"0000005d00000000000000640000000000000058000000000000005600000000",
            INIT_09 => X"0000006900000000000000750000000000000063000000000000007500000000",
            INIT_0A => X"0000008b000000000000009b0000000000000066000000000000006e00000000",
            INIT_0B => X"000000810000000000000081000000000000006f000000000000006b00000000",
            INIT_0C => X"00000076000000000000006d0000000000000077000000000000007c00000000",
            INIT_0D => X"00000071000000000000007c0000000000000076000000000000007100000000",
            INIT_0E => X"0000006300000000000000830000000000000075000000000000008300000000",
            INIT_0F => X"0000005700000000000000270000000000000048000000000000006900000000",
            INIT_10 => X"0000007300000000000000780000000000000060000000000000005f00000000",
            INIT_11 => X"0000005600000000000000630000000000000047000000000000006d00000000",
            INIT_12 => X"000000b0000000000000006a0000000000000063000000000000006c00000000",
            INIT_13 => X"00000075000000000000007b000000000000005e000000000000008200000000",
            INIT_14 => X"000000880000000000000081000000000000008d000000000000008900000000",
            INIT_15 => X"000000790000000000000078000000000000006f000000000000008300000000",
            INIT_16 => X"000000430000000000000050000000000000006b000000000000007500000000",
            INIT_17 => X"0000006e00000000000000430000000000000051000000000000004800000000",
            INIT_18 => X"00000057000000000000007d0000000000000070000000000000006d00000000",
            INIT_19 => X"0000005e00000000000000470000000000000048000000000000005800000000",
            INIT_1A => X"0000007300000000000000490000000000000079000000000000006400000000",
            INIT_1B => X"0000009400000000000000870000000000000076000000000000009800000000",
            INIT_1C => X"0000009500000000000000940000000000000082000000000000008500000000",
            INIT_1D => X"0000007a00000000000000790000000000000071000000000000007d00000000",
            INIT_1E => X"0000004e000000000000003a0000000000000071000000000000007200000000",
            INIT_1F => X"0000008a00000000000000730000000000000038000000000000003d00000000",
            INIT_20 => X"0000004300000000000000590000000000000074000000000000007700000000",
            INIT_21 => X"00000066000000000000003c0000000000000048000000000000005800000000",
            INIT_22 => X"00000037000000000000006d0000000000000057000000000000004800000000",
            INIT_23 => X"0000009c000000000000008d0000000000000092000000000000006500000000",
            INIT_24 => X"00000098000000000000008c0000000000000088000000000000009800000000",
            INIT_25 => X"0000007c000000000000007f000000000000007b000000000000008600000000",
            INIT_26 => X"00000062000000000000005d0000000000000069000000000000006d00000000",
            INIT_27 => X"00000077000000000000007a0000000000000062000000000000004d00000000",
            INIT_28 => X"0000005d00000000000000320000000000000061000000000000007e00000000",
            INIT_29 => X"00000060000000000000004b0000000000000046000000000000006000000000",
            INIT_2A => X"000000610000000000000076000000000000003b000000000000005a00000000",
            INIT_2B => X"0000009700000000000000a20000000000000083000000000000004900000000",
            INIT_2C => X"0000007f000000000000008400000000000000a3000000000000009600000000",
            INIT_2D => X"00000075000000000000006e0000000000000076000000000000007d00000000",
            INIT_2E => X"0000004f000000000000005e0000000000000066000000000000006900000000",
            INIT_2F => X"0000006a0000000000000070000000000000008e000000000000006b00000000",
            INIT_30 => X"0000005900000000000000370000000000000051000000000000007000000000",
            INIT_31 => X"000000590000000000000045000000000000004e000000000000005c00000000",
            INIT_32 => X"000000760000000000000053000000000000006b000000000000007700000000",
            INIT_33 => X"0000009c0000000000000097000000000000007d000000000000006b00000000",
            INIT_34 => X"0000007e0000000000000094000000000000009b000000000000009400000000",
            INIT_35 => X"000000750000000000000078000000000000007b000000000000006c00000000",
            INIT_36 => X"0000005600000000000000540000000000000066000000000000007200000000",
            INIT_37 => X"0000006900000000000000630000000000000079000000000000008100000000",
            INIT_38 => X"0000009a00000000000000780000000000000056000000000000006200000000",
            INIT_39 => X"0000004e0000000000000045000000000000005f000000000000007700000000",
            INIT_3A => X"0000004e0000000000000057000000000000007e000000000000007300000000",
            INIT_3B => X"000000960000000000000084000000000000008b000000000000007d00000000",
            INIT_3C => X"0000007e0000000000000092000000000000008e000000000000008d00000000",
            INIT_3D => X"0000007b00000000000000760000000000000084000000000000007900000000",
            INIT_3E => X"0000006f00000000000000520000000000000058000000000000007300000000",
            INIT_3F => X"00000067000000000000006a0000000000000065000000000000007900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a70000000000000088000000000000007400000000",
            INIT_41 => X"0000005c00000000000000600000000000000077000000000000009f00000000",
            INIT_42 => X"0000006f0000000000000066000000000000005a000000000000006600000000",
            INIT_43 => X"0000008f00000000000000830000000000000088000000000000007000000000",
            INIT_44 => X"000000800000000000000096000000000000008e000000000000008600000000",
            INIT_45 => X"000000770000000000000084000000000000009c000000000000007500000000",
            INIT_46 => X"00000053000000000000004e0000000000000059000000000000006600000000",
            INIT_47 => X"0000006c00000000000000710000000000000060000000000000006a00000000",
            INIT_48 => X"000000920000000000000071000000000000006d000000000000006c00000000",
            INIT_49 => X"00000069000000000000007b000000000000009e00000000000000a600000000",
            INIT_4A => X"0000008c00000000000000550000000000000052000000000000006600000000",
            INIT_4B => X"0000007b0000000000000086000000000000007e000000000000009100000000",
            INIT_4C => X"00000089000000000000008a0000000000000073000000000000006800000000",
            INIT_4D => X"0000006a000000000000008a0000000000000096000000000000008300000000",
            INIT_4E => X"0000002d000000000000004a000000000000006f000000000000006100000000",
            INIT_4F => X"0000004b00000000000000690000000000000065000000000000006000000000",
            INIT_50 => X"0000005600000000000000370000000000000055000000000000005800000000",
            INIT_51 => X"0000007e00000000000000970000000000000097000000000000008b00000000",
            INIT_52 => X"0000005700000000000000570000000000000068000000000000006800000000",
            INIT_53 => X"00000052000000000000006e000000000000006e000000000000006f00000000",
            INIT_54 => X"0000008c0000000000000079000000000000004b000000000000003500000000",
            INIT_55 => X"0000007a00000000000000810000000000000078000000000000009100000000",
            INIT_56 => X"00000020000000000000003e0000000000000062000000000000007400000000",
            INIT_57 => X"0000004000000000000000410000000000000062000000000000006100000000",
            INIT_58 => X"000000200000000000000022000000000000005c000000000000005200000000",
            INIT_59 => X"0000009c00000000000000860000000000000075000000000000004b00000000",
            INIT_5A => X"000000570000000000000062000000000000006d000000000000008d00000000",
            INIT_5B => X"0000005f000000000000005b000000000000005a000000000000005200000000",
            INIT_5C => X"0000008b00000000000000790000000000000046000000000000005200000000",
            INIT_5D => X"0000006b0000000000000080000000000000008f000000000000008100000000",
            INIT_5E => X"0000003f000000000000001d000000000000004e000000000000007100000000",
            INIT_5F => X"0000004200000000000000470000000000000047000000000000006300000000",
            INIT_60 => X"0000000d00000000000000230000000000000056000000000000005a00000000",
            INIT_61 => X"000000940000000000000072000000000000004e000000000000000f00000000",
            INIT_62 => X"00000062000000000000006f000000000000008b00000000000000a200000000",
            INIT_63 => X"000000710000000000000056000000000000005b000000000000006100000000",
            INIT_64 => X"0000007e0000000000000073000000000000006a000000000000007800000000",
            INIT_65 => X"0000006a00000000000000870000000000000087000000000000007600000000",
            INIT_66 => X"0000005b0000000000000026000000000000002a000000000000004f00000000",
            INIT_67 => X"0000005300000000000000990000000000000060000000000000002c00000000",
            INIT_68 => X"00000025000000000000002d0000000000000056000000000000005c00000000",
            INIT_69 => X"0000007a0000000000000057000000000000001f000000000000000d00000000",
            INIT_6A => X"0000007a000000000000009e00000000000000ad000000000000009600000000",
            INIT_6B => X"0000005c000000000000005d0000000000000072000000000000007500000000",
            INIT_6C => X"0000007100000000000000670000000000000055000000000000004d00000000",
            INIT_6D => X"0000005b00000000000000730000000000000085000000000000007e00000000",
            INIT_6E => X"0000003c000000000000003b0000000000000032000000000000004e00000000",
            INIT_6F => X"000000620000000000000086000000000000006c000000000000002a00000000",
            INIT_70 => X"0000003800000000000000180000000000000047000000000000005200000000",
            INIT_71 => X"0000005400000000000000230000000000000017000000000000002400000000",
            INIT_72 => X"000000a500000000000000a50000000000000092000000000000007600000000",
            INIT_73 => X"00000079000000000000006f0000000000000082000000000000009600000000",
            INIT_74 => X"00000062000000000000003f0000000000000042000000000000006c00000000",
            INIT_75 => X"0000005600000000000000460000000000000045000000000000004e00000000",
            INIT_76 => X"000000620000000000000060000000000000006c000000000000007500000000",
            INIT_77 => X"00000059000000000000007b0000000000000074000000000000007800000000",
            INIT_78 => X"000000400000000000000011000000000000001b000000000000004100000000",
            INIT_79 => X"00000025000000000000000f000000000000001d000000000000003400000000",
            INIT_7A => X"0000009600000000000000740000000000000064000000000000005900000000",
            INIT_7B => X"0000009c0000000000000088000000000000009800000000000000aa00000000",
            INIT_7C => X"0000004a0000000000000045000000000000007900000000000000a600000000",
            INIT_7D => X"0000007f00000000000000660000000000000047000000000000002f00000000",
            INIT_7E => X"000000820000000000000083000000000000008b000000000000009c00000000",
            INIT_7F => X"0000007500000000000000920000000000000088000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "sampleifmap_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000058000000000000004d000000000000008b00000000000000b300000000",
            INIT_01 => X"00000097000000000000009c000000000000009d000000000000008d00000000",
            INIT_02 => X"000000970000000000000090000000000000009e000000000000009c00000000",
            INIT_03 => X"0000007600000000000000790000000000000088000000000000009700000000",
            INIT_04 => X"000000540000000000000054000000000000006c000000000000007e00000000",
            INIT_05 => X"00000053000000000000005e0000000000000062000000000000006200000000",
            INIT_06 => X"0000006000000000000000540000000000000056000000000000005a00000000",
            INIT_07 => X"0000004d000000000000004c0000000000000057000000000000007500000000",
            INIT_08 => X"000000920000000000000080000000000000008500000000000000b800000000",
            INIT_09 => X"000000a7000000000000009e000000000000009f000000000000009f00000000",
            INIT_0A => X"0000009a000000000000009900000000000000a200000000000000a500000000",
            INIT_0B => X"0000007d00000000000000880000000000000096000000000000009600000000",
            INIT_0C => X"00000052000000000000005a000000000000006d000000000000008100000000",
            INIT_0D => X"00000058000000000000005e0000000000000062000000000000005d00000000",
            INIT_0E => X"0000006a000000000000005b000000000000004c000000000000004e00000000",
            INIT_0F => X"0000005a000000000000005b0000000000000062000000000000007600000000",
            INIT_10 => X"000000aa00000000000000b0000000000000009800000000000000b400000000",
            INIT_11 => X"000000a4000000000000009b000000000000009800000000000000a400000000",
            INIT_12 => X"0000009f00000000000000a200000000000000aa00000000000000a200000000",
            INIT_13 => X"0000008c00000000000000920000000000000097000000000000009c00000000",
            INIT_14 => X"000000470000000000000058000000000000007c000000000000009200000000",
            INIT_15 => X"0000006b00000000000000670000000000000062000000000000005500000000",
            INIT_16 => X"0000006f000000000000006f000000000000006d000000000000006500000000",
            INIT_17 => X"0000005f000000000000005d0000000000000065000000000000006f00000000",
            INIT_18 => X"000000b500000000000000b800000000000000ae00000000000000af00000000",
            INIT_19 => X"000000a300000000000000a4000000000000009800000000000000a800000000",
            INIT_1A => X"000000a800000000000000a700000000000000b300000000000000a600000000",
            INIT_1B => X"000000a4000000000000009f00000000000000a200000000000000ae00000000",
            INIT_1C => X"0000003a00000000000000590000000000000089000000000000009700000000",
            INIT_1D => X"0000006b0000000000000063000000000000005a000000000000004800000000",
            INIT_1E => X"00000079000000000000007d0000000000000080000000000000007500000000",
            INIT_1F => X"0000006f000000000000006d0000000000000061000000000000006900000000",
            INIT_20 => X"000000ac00000000000000a700000000000000ae00000000000000af00000000",
            INIT_21 => X"000000af00000000000000b000000000000000a100000000000000a200000000",
            INIT_22 => X"000000b400000000000000b300000000000000b200000000000000b200000000",
            INIT_23 => X"000000a400000000000000a000000000000000a800000000000000b000000000",
            INIT_24 => X"000000450000000000000078000000000000009c00000000000000ad00000000",
            INIT_25 => X"0000005e0000000000000063000000000000005a000000000000004200000000",
            INIT_26 => X"0000007b000000000000007f000000000000007c000000000000006900000000",
            INIT_27 => X"0000007400000000000000710000000000000068000000000000007000000000",
            INIT_28 => X"000000aa000000000000009000000000000000ae00000000000000b500000000",
            INIT_29 => X"000000b300000000000000b000000000000000a600000000000000a900000000",
            INIT_2A => X"000000b500000000000000b400000000000000b400000000000000b400000000",
            INIT_2B => X"00000096000000000000009f00000000000000ae00000000000000b000000000",
            INIT_2C => X"00000074000000000000009b00000000000000af00000000000000b500000000",
            INIT_2D => X"000000700000000000000083000000000000007d000000000000006000000000",
            INIT_2E => X"00000079000000000000007a0000000000000078000000000000007500000000",
            INIT_2F => X"0000007c00000000000000760000000000000078000000000000007900000000",
            INIT_30 => X"000000b2000000000000008a000000000000009c00000000000000c000000000",
            INIT_31 => X"000000af00000000000000b000000000000000ae00000000000000af00000000",
            INIT_32 => X"000000b800000000000000ba00000000000000b400000000000000b800000000",
            INIT_33 => X"0000009900000000000000ad00000000000000bb00000000000000bb00000000",
            INIT_34 => X"000000a700000000000000ad00000000000000ad00000000000000a600000000",
            INIT_35 => X"0000007900000000000000940000000000000095000000000000009600000000",
            INIT_36 => X"0000006f000000000000006d0000000000000075000000000000007300000000",
            INIT_37 => X"00000080000000000000007b000000000000007a000000000000007800000000",
            INIT_38 => X"000000ab000000000000009c000000000000007d00000000000000b900000000",
            INIT_39 => X"000000b800000000000000af00000000000000af00000000000000ad00000000",
            INIT_3A => X"000000c200000000000000c100000000000000b700000000000000bc00000000",
            INIT_3B => X"000000a600000000000000b800000000000000b900000000000000bd00000000",
            INIT_3C => X"000000b000000000000000b100000000000000ac00000000000000a400000000",
            INIT_3D => X"0000007a000000000000008f000000000000008900000000000000aa00000000",
            INIT_3E => X"000000670000000000000060000000000000006e000000000000006b00000000",
            INIT_3F => X"0000007d000000000000007b0000000000000076000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a0000000000000009f0000000000000095000000000000009b00000000",
            INIT_41 => X"000000b400000000000000b200000000000000ad00000000000000ac00000000",
            INIT_42 => X"000000bf00000000000000ba00000000000000ba00000000000000bb00000000",
            INIT_43 => X"000000a000000000000000ac00000000000000af00000000000000bb00000000",
            INIT_44 => X"000000b000000000000000a60000000000000097000000000000009a00000000",
            INIT_45 => X"0000008500000000000000a6000000000000009b00000000000000b700000000",
            INIT_46 => X"0000007700000000000000700000000000000068000000000000006800000000",
            INIT_47 => X"0000007d000000000000007a000000000000007a000000000000007600000000",
            INIT_48 => X"000000a900000000000000930000000000000098000000000000009a00000000",
            INIT_49 => X"000000aa00000000000000b700000000000000b200000000000000b200000000",
            INIT_4A => X"000000c100000000000000c600000000000000bc00000000000000b000000000",
            INIT_4B => X"000000a900000000000000a500000000000000a700000000000000ae00000000",
            INIT_4C => X"000000a90000000000000092000000000000008c000000000000009d00000000",
            INIT_4D => X"0000008d00000000000000ab00000000000000a000000000000000b300000000",
            INIT_4E => X"0000007700000000000000750000000000000068000000000000005f00000000",
            INIT_4F => X"0000007d0000000000000076000000000000007b000000000000007400000000",
            INIT_50 => X"000000b1000000000000009f0000000000000070000000000000008600000000",
            INIT_51 => X"000000ba00000000000000b800000000000000b800000000000000ae00000000",
            INIT_52 => X"000000b000000000000000bf00000000000000c200000000000000ba00000000",
            INIT_53 => X"000000bb00000000000000a7000000000000009e000000000000009b00000000",
            INIT_54 => X"000000970000000000000086000000000000009300000000000000ae00000000",
            INIT_55 => X"0000007c000000000000009b000000000000009c00000000000000a000000000",
            INIT_56 => X"0000006600000000000000690000000000000066000000000000004a00000000",
            INIT_57 => X"0000007f000000000000007b0000000000000075000000000000006b00000000",
            INIT_58 => X"0000009d00000000000000ae000000000000005b000000000000004100000000",
            INIT_59 => X"000000be00000000000000bf00000000000000b1000000000000009300000000",
            INIT_5A => X"000000b000000000000000ac00000000000000b000000000000000bc00000000",
            INIT_5B => X"000000a3000000000000009400000000000000ae00000000000000b800000000",
            INIT_5C => X"000000950000000000000085000000000000009a00000000000000b000000000",
            INIT_5D => X"0000005000000000000000830000000000000095000000000000009800000000",
            INIT_5E => X"0000006600000000000000670000000000000061000000000000004200000000",
            INIT_5F => X"0000007d00000000000000780000000000000071000000000000006700000000",
            INIT_60 => X"000000b100000000000000bf000000000000005c000000000000001500000000",
            INIT_61 => X"000000b600000000000000bd00000000000000ca00000000000000bc00000000",
            INIT_62 => X"000000bc00000000000000a5000000000000009c00000000000000b300000000",
            INIT_63 => X"00000072000000000000009800000000000000ae00000000000000c800000000",
            INIT_64 => X"000000890000000000000078000000000000007f000000000000005f00000000",
            INIT_65 => X"0000004e00000000000000720000000000000088000000000000009700000000",
            INIT_66 => X"0000006200000000000000590000000000000049000000000000004000000000",
            INIT_67 => X"0000007600000000000000750000000000000071000000000000006200000000",
            INIT_68 => X"000000ad00000000000000a80000000000000063000000000000002c00000000",
            INIT_69 => X"000000bb00000000000000bc00000000000000c300000000000000c800000000",
            INIT_6A => X"000000c200000000000000b4000000000000009500000000000000a500000000",
            INIT_6B => X"0000009a00000000000000a800000000000000a800000000000000b900000000",
            INIT_6C => X"0000008a00000000000000910000000000000092000000000000006b00000000",
            INIT_6D => X"000000480000000000000064000000000000007f000000000000009c00000000",
            INIT_6E => X"0000006000000000000000530000000000000040000000000000003900000000",
            INIT_6F => X"0000006f000000000000006c000000000000006a000000000000006200000000",
            INIT_70 => X"0000009f00000000000000750000000000000076000000000000006900000000",
            INIT_71 => X"000000bb00000000000000b400000000000000be00000000000000c400000000",
            INIT_72 => X"000000c100000000000000c600000000000000ad00000000000000ad00000000",
            INIT_73 => X"000000bc00000000000000b400000000000000a500000000000000ab00000000",
            INIT_74 => X"000000b300000000000000ad00000000000000bb00000000000000ae00000000",
            INIT_75 => X"000000480000000000000069000000000000008000000000000000a000000000",
            INIT_76 => X"0000006c00000000000000570000000000000045000000000000004300000000",
            INIT_77 => X"0000006600000000000000610000000000000064000000000000006300000000",
            INIT_78 => X"0000009d00000000000000680000000000000071000000000000008a00000000",
            INIT_79 => X"000000a800000000000000b400000000000000c400000000000000c600000000",
            INIT_7A => X"000000cd00000000000000cb00000000000000bf00000000000000b400000000",
            INIT_7B => X"000000c800000000000000c400000000000000bf00000000000000d200000000",
            INIT_7C => X"000000be00000000000000bc00000000000000bb00000000000000c000000000",
            INIT_7D => X"000000500000000000000071000000000000009900000000000000a800000000",
            INIT_7E => X"0000008700000000000000600000000000000040000000000000004600000000",
            INIT_7F => X"00000062000000000000005a000000000000005a000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "sampleifmap_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000930000000000000073000000000000008a000000000000009600000000",
            INIT_01 => X"0000009600000000000000b000000000000000bb00000000000000be00000000",
            INIT_02 => X"000000c600000000000000d300000000000000c700000000000000ab00000000",
            INIT_03 => X"000000cb00000000000000be00000000000000c200000000000000d300000000",
            INIT_04 => X"000000bd00000000000000b800000000000000ba00000000000000bf00000000",
            INIT_05 => X"00000046000000000000006400000000000000a600000000000000be00000000",
            INIT_06 => X"0000008f000000000000006a0000000000000038000000000000002f00000000",
            INIT_07 => X"0000005e000000000000004a000000000000005c000000000000009500000000",
            INIT_08 => X"000000a50000000000000092000000000000009b000000000000009b00000000",
            INIT_09 => X"0000009100000000000000bf00000000000000c000000000000000bd00000000",
            INIT_0A => X"0000009500000000000000a900000000000000d2000000000000009c00000000",
            INIT_0B => X"000000a800000000000000b200000000000000c200000000000000c000000000",
            INIT_0C => X"000000a700000000000000aa00000000000000b500000000000000a900000000",
            INIT_0D => X"0000002b00000000000000430000000000000075000000000000009a00000000",
            INIT_0E => X"0000008f00000000000000680000000000000031000000000000002200000000",
            INIT_0F => X"00000050000000000000003f000000000000006a000000000000009c00000000",
            INIT_10 => X"000000a6000000000000008a00000000000000a200000000000000a500000000",
            INIT_11 => X"0000008900000000000000ba00000000000000be00000000000000c400000000",
            INIT_12 => X"000000a9000000000000009d00000000000000c9000000000000007400000000",
            INIT_13 => X"0000008f000000000000008000000000000000b600000000000000d200000000",
            INIT_14 => X"00000061000000000000007f0000000000000093000000000000007c00000000",
            INIT_15 => X"00000033000000000000002f0000000000000038000000000000005200000000",
            INIT_16 => X"0000009d00000000000000690000000000000040000000000000002b00000000",
            INIT_17 => X"000000410000000000000039000000000000007b000000000000009d00000000",
            INIT_18 => X"0000009e0000000000000078000000000000009600000000000000a900000000",
            INIT_19 => X"0000009800000000000000be00000000000000be00000000000000be00000000",
            INIT_1A => X"000000b900000000000000bc0000000000000099000000000000003c00000000",
            INIT_1B => X"000000ce000000000000009000000000000000a500000000000000c300000000",
            INIT_1C => X"0000003d0000000000000065000000000000008900000000000000b100000000",
            INIT_1D => X"0000005000000000000000470000000000000033000000000000003700000000",
            INIT_1E => X"000000a0000000000000006e000000000000004a000000000000003700000000",
            INIT_1F => X"000000320000000000000036000000000000008e00000000000000b000000000",
            INIT_20 => X"000000a6000000000000009600000000000000a000000000000000aa00000000",
            INIT_21 => X"0000009a00000000000000ba00000000000000bc00000000000000ba00000000",
            INIT_22 => X"00000092000000000000007e0000000000000031000000000000002000000000",
            INIT_23 => X"000000c0000000000000008c000000000000008c000000000000009b00000000",
            INIT_24 => X"0000003e0000000000000061000000000000009c00000000000000cc00000000",
            INIT_25 => X"0000005700000000000000520000000000000049000000000000004900000000",
            INIT_26 => X"000000a6000000000000006b000000000000003e000000000000003a00000000",
            INIT_27 => X"00000033000000000000004800000000000000a700000000000000bc00000000",
            INIT_28 => X"0000009c000000000000009700000000000000ab00000000000000b200000000",
            INIT_29 => X"0000007c00000000000000a300000000000000b200000000000000b500000000",
            INIT_2A => X"000000370000000000000028000000000000001d000000000000002400000000",
            INIT_2B => X"0000008200000000000000650000000000000063000000000000004e00000000",
            INIT_2C => X"00000037000000000000005f000000000000007b000000000000009000000000",
            INIT_2D => X"00000055000000000000003c0000000000000033000000000000003400000000",
            INIT_2E => X"000000990000000000000066000000000000004d000000000000004e00000000",
            INIT_2F => X"00000037000000000000005900000000000000b100000000000000bb00000000",
            INIT_30 => X"00000098000000000000009200000000000000ab00000000000000b500000000",
            INIT_31 => X"00000069000000000000009500000000000000a700000000000000a900000000",
            INIT_32 => X"0000002e0000000000000042000000000000005e000000000000004f00000000",
            INIT_33 => X"00000078000000000000005c0000000000000047000000000000002f00000000",
            INIT_34 => X"0000002900000000000000380000000000000037000000000000005a00000000",
            INIT_35 => X"00000037000000000000001e0000000000000022000000000000002300000000",
            INIT_36 => X"0000007700000000000000610000000000000056000000000000005200000000",
            INIT_37 => X"0000003c000000000000006a00000000000000ae00000000000000ad00000000",
            INIT_38 => X"000000a3000000000000009e000000000000009c00000000000000b100000000",
            INIT_39 => X"00000089000000000000009400000000000000a0000000000000009c00000000",
            INIT_3A => X"0000006b00000000000000660000000000000076000000000000008f00000000",
            INIT_3B => X"00000067000000000000007d000000000000006d000000000000006e00000000",
            INIT_3C => X"0000001300000000000000100000000000000011000000000000002f00000000",
            INIT_3D => X"00000013000000000000000e000000000000001c000000000000001800000000",
            INIT_3E => X"0000006300000000000000600000000000000041000000000000002b00000000",
            INIT_3F => X"00000043000000000000008500000000000000ad000000000000008c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a7000000000000008b000000000000009e00000000",
            INIT_41 => X"000000c000000000000000ab000000000000008c000000000000009700000000",
            INIT_42 => X"000000880000000000000085000000000000007400000000000000ac00000000",
            INIT_43 => X"00000065000000000000007f000000000000008d000000000000009200000000",
            INIT_44 => X"0000001900000000000000200000000000000025000000000000004100000000",
            INIT_45 => X"0000000f000000000000000a0000000000000011000000000000001800000000",
            INIT_46 => X"0000004e00000000000000610000000000000042000000000000001400000000",
            INIT_47 => X"00000069000000000000009c0000000000000094000000000000006200000000",
            INIT_48 => X"000000ab00000000000000ae00000000000000a400000000000000a000000000",
            INIT_49 => X"000000b100000000000000940000000000000088000000000000009e00000000",
            INIT_4A => X"0000009700000000000000a9000000000000009300000000000000b800000000",
            INIT_4B => X"0000007d000000000000008e000000000000008b000000000000007f00000000",
            INIT_4C => X"0000002b000000000000003f000000000000004d000000000000006700000000",
            INIT_4D => X"0000001a00000000000000110000000000000018000000000000002100000000",
            INIT_4E => X"000000320000000000000048000000000000003e000000000000001f00000000",
            INIT_4F => X"000000880000000000000078000000000000005a000000000000004800000000",
            INIT_50 => X"000000a700000000000000a700000000000000a300000000000000a000000000",
            INIT_51 => X"00000078000000000000008c00000000000000a800000000000000b100000000",
            INIT_52 => X"000000820000000000000076000000000000008f00000000000000ab00000000",
            INIT_53 => X"0000009100000000000000a6000000000000009c000000000000007b00000000",
            INIT_54 => X"0000004e000000000000005b0000000000000069000000000000007c00000000",
            INIT_55 => X"0000004300000000000000380000000000000042000000000000004c00000000",
            INIT_56 => X"0000004900000000000000410000000000000041000000000000004600000000",
            INIT_57 => X"0000006a0000000000000051000000000000007b000000000000006400000000",
            INIT_58 => X"00000093000000000000008c000000000000009f000000000000009c00000000",
            INIT_59 => X"0000007b000000000000009900000000000000aa00000000000000b400000000",
            INIT_5A => X"0000007e0000000000000073000000000000009c000000000000008b00000000",
            INIT_5B => X"000000a200000000000000a8000000000000009e000000000000008300000000",
            INIT_5C => X"00000078000000000000007b0000000000000077000000000000007f00000000",
            INIT_5D => X"0000007700000000000000690000000000000068000000000000007000000000",
            INIT_5E => X"0000006d00000000000000680000000000000069000000000000007400000000",
            INIT_5F => X"00000068000000000000005c0000000000000086000000000000007a00000000",
            INIT_60 => X"0000008b000000000000007b000000000000009e00000000000000a400000000",
            INIT_61 => X"0000008c000000000000008d000000000000009c00000000000000ad00000000",
            INIT_62 => X"000000a100000000000000820000000000000079000000000000008d00000000",
            INIT_63 => X"000000a800000000000000a6000000000000009d000000000000009700000000",
            INIT_64 => X"00000084000000000000008f000000000000008a000000000000009000000000",
            INIT_65 => X"00000094000000000000008a0000000000000085000000000000008100000000",
            INIT_66 => X"0000008400000000000000860000000000000089000000000000008f00000000",
            INIT_67 => X"0000009300000000000000730000000000000064000000000000007800000000",
            INIT_68 => X"000000a800000000000000900000000000000095000000000000008e00000000",
            INIT_69 => X"0000009e000000000000009e00000000000000a100000000000000a700000000",
            INIT_6A => X"000000a90000000000000097000000000000009000000000000000a500000000",
            INIT_6B => X"000000a2000000000000009e00000000000000a000000000000000a100000000",
            INIT_6C => X"0000007f00000000000000890000000000000091000000000000009900000000",
            INIT_6D => X"0000009e00000000000000960000000000000095000000000000008d00000000",
            INIT_6E => X"0000008f00000000000000940000000000000096000000000000009f00000000",
            INIT_6F => X"0000009f000000000000008b0000000000000077000000000000007b00000000",
            INIT_70 => X"000000b900000000000000b300000000000000a6000000000000009800000000",
            INIT_71 => X"000000a800000000000000aa00000000000000a700000000000000a700000000",
            INIT_72 => X"000000b200000000000000ad00000000000000a400000000000000a700000000",
            INIT_73 => X"000000850000000000000089000000000000009d00000000000000a900000000",
            INIT_74 => X"00000088000000000000008c000000000000008f000000000000009200000000",
            INIT_75 => X"0000009d00000000000000980000000000000097000000000000008c00000000",
            INIT_76 => X"000000900000000000000099000000000000009c00000000000000a600000000",
            INIT_77 => X"0000009900000000000000900000000000000083000000000000008500000000",
            INIT_78 => X"000000ab00000000000000b700000000000000b2000000000000009f00000000",
            INIT_79 => X"0000009f0000000000000091000000000000007d000000000000008b00000000",
            INIT_7A => X"0000009c0000000000000095000000000000008b00000000000000a200000000",
            INIT_7B => X"0000007300000000000000830000000000000098000000000000009e00000000",
            INIT_7C => X"0000008f0000000000000094000000000000008e000000000000008400000000",
            INIT_7D => X"000000a1000000000000009c000000000000009d000000000000009000000000",
            INIT_7E => X"0000009c0000000000000094000000000000009f00000000000000a700000000",
            INIT_7F => X"0000009800000000000000990000000000000096000000000000009c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "sampleifmap_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000310000000000000060000000000000007600000000",
            INIT_01 => X"000000530000000000000054000000000000005f000000000000006000000000",
            INIT_02 => X"0000005a00000000000000530000000000000061000000000000005f00000000",
            INIT_03 => X"0000004f000000000000004b0000000000000052000000000000005c00000000",
            INIT_04 => X"00000032000000000000003b0000000000000050000000000000005b00000000",
            INIT_05 => X"0000003300000000000000380000000000000038000000000000003700000000",
            INIT_06 => X"0000003a00000000000000330000000000000038000000000000003c00000000",
            INIT_07 => X"0000002f000000000000002f0000000000000035000000000000004c00000000",
            INIT_08 => X"0000006900000000000000590000000000000058000000000000008200000000",
            INIT_09 => X"00000068000000000000005d0000000000000060000000000000006c00000000",
            INIT_0A => X"0000005b000000000000005a0000000000000062000000000000006500000000",
            INIT_0B => X"00000048000000000000004f0000000000000057000000000000005400000000",
            INIT_0C => X"00000032000000000000003d0000000000000048000000000000005200000000",
            INIT_0D => X"0000003300000000000000370000000000000038000000000000003700000000",
            INIT_0E => X"0000004100000000000000350000000000000028000000000000002b00000000",
            INIT_0F => X"00000039000000000000003a000000000000003d000000000000004b00000000",
            INIT_10 => X"0000007a00000000000000810000000000000068000000000000008400000000",
            INIT_11 => X"0000006a000000000000005f0000000000000059000000000000006c00000000",
            INIT_12 => X"0000005e00000000000000620000000000000069000000000000006200000000",
            INIT_13 => X"0000004c000000000000004f0000000000000050000000000000005500000000",
            INIT_14 => X"0000002a0000000000000036000000000000004c000000000000005500000000",
            INIT_15 => X"00000042000000000000003f000000000000003a000000000000003300000000",
            INIT_16 => X"0000004200000000000000430000000000000042000000000000003c00000000",
            INIT_17 => X"000000390000000000000038000000000000003e000000000000004300000000",
            INIT_18 => X"000000840000000000000088000000000000007f000000000000008100000000",
            INIT_19 => X"000000690000000000000068000000000000005a000000000000007000000000",
            INIT_1A => X"0000006600000000000000650000000000000071000000000000006500000000",
            INIT_1B => X"0000005d0000000000000057000000000000005a000000000000006700000000",
            INIT_1C => X"0000001f0000000000000033000000000000004e000000000000004f00000000",
            INIT_1D => X"0000003e00000000000000390000000000000033000000000000002a00000000",
            INIT_1E => X"0000004a000000000000004b000000000000004d000000000000004600000000",
            INIT_1F => X"0000004500000000000000430000000000000037000000000000003c00000000",
            INIT_20 => X"0000007f0000000000000079000000000000007f000000000000008000000000",
            INIT_21 => X"0000007200000000000000720000000000000063000000000000006d00000000",
            INIT_22 => X"000000710000000000000070000000000000006f000000000000006f00000000",
            INIT_23 => X"0000005c00000000000000590000000000000063000000000000006c00000000",
            INIT_24 => X"0000002c000000000000004e0000000000000059000000000000005e00000000",
            INIT_25 => X"0000002e00000000000000380000000000000034000000000000002700000000",
            INIT_26 => X"0000004900000000000000470000000000000043000000000000003500000000",
            INIT_27 => X"000000470000000000000045000000000000003b000000000000004200000000",
            INIT_28 => X"0000007f00000000000000680000000000000083000000000000008900000000",
            INIT_29 => X"000000740000000000000071000000000000006a000000000000007600000000",
            INIT_2A => X"0000007100000000000000740000000000000075000000000000007300000000",
            INIT_2B => X"00000054000000000000005a0000000000000069000000000000006d00000000",
            INIT_2C => X"0000004f00000000000000670000000000000068000000000000006a00000000",
            INIT_2D => X"0000003d0000000000000052000000000000004d000000000000003a00000000",
            INIT_2E => X"000000460000000000000043000000000000003f000000000000003e00000000",
            INIT_2F => X"0000004b00000000000000460000000000000048000000000000004900000000",
            INIT_30 => X"0000008700000000000000660000000000000077000000000000009800000000",
            INIT_31 => X"0000006f00000000000000730000000000000075000000000000007a00000000",
            INIT_32 => X"00000070000000000000007c000000000000007b000000000000007900000000",
            INIT_33 => X"0000005c00000000000000660000000000000071000000000000007300000000",
            INIT_34 => X"0000006e000000000000006d0000000000000065000000000000006400000000",
            INIT_35 => X"00000043000000000000005b0000000000000057000000000000005c00000000",
            INIT_36 => X"0000003b00000000000000380000000000000040000000000000003e00000000",
            INIT_37 => X"0000004e000000000000004a0000000000000048000000000000004500000000",
            INIT_38 => X"0000007e00000000000000780000000000000059000000000000009300000000",
            INIT_39 => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_3A => X"00000073000000000000007c000000000000007a000000000000008000000000",
            INIT_3B => X"00000064000000000000006c000000000000006d000000000000007300000000",
            INIT_3C => X"0000006a000000000000006d0000000000000068000000000000006500000000",
            INIT_3D => X"000000480000000000000057000000000000004b000000000000006600000000",
            INIT_3E => X"00000035000000000000002e000000000000003c000000000000003b00000000",
            INIT_3F => X"0000004b00000000000000490000000000000044000000000000004200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000720000000000000078000000000000006f000000000000007600000000",
            INIT_41 => X"0000007700000000000000750000000000000074000000000000007700000000",
            INIT_42 => X"0000006d000000000000006f000000000000007a000000000000008000000000",
            INIT_43 => X"0000005e00000000000000610000000000000067000000000000007300000000",
            INIT_44 => X"0000006400000000000000610000000000000059000000000000005e00000000",
            INIT_45 => X"000000590000000000000072000000000000005f000000000000006d00000000",
            INIT_46 => X"000000470000000000000040000000000000003a000000000000003e00000000",
            INIT_47 => X"0000004b00000000000000480000000000000048000000000000004600000000",
            INIT_48 => X"0000007800000000000000690000000000000071000000000000007700000000",
            INIT_49 => X"0000006f000000000000007b000000000000007a000000000000007c00000000",
            INIT_4A => X"00000079000000000000007d000000000000007b000000000000007600000000",
            INIT_4B => X"0000006f0000000000000065000000000000006d000000000000007600000000",
            INIT_4C => X"0000006000000000000000520000000000000055000000000000006900000000",
            INIT_4D => X"00000067000000000000007a0000000000000064000000000000006a00000000",
            INIT_4E => X"000000490000000000000047000000000000003e000000000000003d00000000",
            INIT_4F => X"0000004b0000000000000044000000000000004b000000000000004700000000",
            INIT_50 => X"0000007e00000000000000720000000000000048000000000000006400000000",
            INIT_51 => X"0000007e000000000000007c000000000000007f000000000000007800000000",
            INIT_52 => X"0000007b00000000000000800000000000000081000000000000007f00000000",
            INIT_53 => X"0000009000000000000000780000000000000077000000000000007900000000",
            INIT_54 => X"00000058000000000000004f0000000000000063000000000000008300000000",
            INIT_55 => X"0000005b000000000000006c0000000000000061000000000000005f00000000",
            INIT_56 => X"0000003b000000000000003d000000000000003e000000000000002e00000000",
            INIT_57 => X"0000004c00000000000000490000000000000046000000000000004000000000",
            INIT_58 => X"00000069000000000000007f0000000000000034000000000000002200000000",
            INIT_59 => X"000000830000000000000084000000000000007a000000000000005d00000000",
            INIT_5A => X"0000008c00000000000000780000000000000073000000000000008100000000",
            INIT_5B => X"000000850000000000000074000000000000009700000000000000a600000000",
            INIT_5C => X"000000610000000000000056000000000000006e000000000000008d00000000",
            INIT_5D => X"000000310000000000000056000000000000005c000000000000006000000000",
            INIT_5E => X"0000003c000000000000003e000000000000003c000000000000002a00000000",
            INIT_5F => X"0000004a00000000000000450000000000000042000000000000003e00000000",
            INIT_60 => X"0000007d000000000000008e0000000000000040000000000000000400000000",
            INIT_61 => X"00000084000000000000008c000000000000009a000000000000008c00000000",
            INIT_62 => X"0000009c000000000000007b000000000000006b000000000000007f00000000",
            INIT_63 => X"000000530000000000000077000000000000009300000000000000b200000000",
            INIT_64 => X"000000640000000000000053000000000000005b000000000000004000000000",
            INIT_65 => X"00000031000000000000004d000000000000005c000000000000006f00000000",
            INIT_66 => X"000000390000000000000037000000000000002f000000000000002900000000",
            INIT_67 => X"0000004400000000000000420000000000000043000000000000003b00000000",
            INIT_68 => X"0000007b000000000000007a0000000000000048000000000000001800000000",
            INIT_69 => X"0000008d000000000000008f0000000000000096000000000000009c00000000",
            INIT_6A => X"000000a0000000000000008f000000000000006a000000000000007700000000",
            INIT_6B => X"0000007700000000000000800000000000000081000000000000009700000000",
            INIT_6C => X"0000006d00000000000000730000000000000074000000000000004d00000000",
            INIT_6D => X"0000002d0000000000000044000000000000005a000000000000007b00000000",
            INIT_6E => X"000000370000000000000033000000000000002b000000000000002300000000",
            INIT_6F => X"0000003e000000000000003a000000000000003e000000000000003b00000000",
            INIT_70 => X"00000070000000000000004a0000000000000052000000000000004500000000",
            INIT_71 => X"0000008f00000000000000860000000000000091000000000000009600000000",
            INIT_72 => X"0000009c00000000000000a10000000000000084000000000000008300000000",
            INIT_73 => X"0000009700000000000000850000000000000072000000000000007d00000000",
            INIT_74 => X"00000098000000000000009200000000000000a0000000000000009100000000",
            INIT_75 => X"0000002f000000000000004b000000000000005d000000000000008100000000",
            INIT_76 => X"0000004400000000000000380000000000000030000000000000002f00000000",
            INIT_77 => X"000000390000000000000036000000000000003c000000000000003c00000000",
            INIT_78 => X"00000070000000000000003b0000000000000041000000000000005700000000",
            INIT_79 => X"0000007d00000000000000860000000000000096000000000000009800000000",
            INIT_7A => X"000000a500000000000000a7000000000000009b000000000000008f00000000",
            INIT_7B => X"000000a0000000000000008f0000000000000084000000000000009b00000000",
            INIT_7C => X"000000a1000000000000009f000000000000009e00000000000000a200000000",
            INIT_7D => X"0000003900000000000000540000000000000078000000000000008900000000",
            INIT_7E => X"0000005f0000000000000040000000000000002b000000000000003300000000",
            INIT_7F => X"0000003900000000000000360000000000000037000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "sampleifmap_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000660000000000000040000000000000004e000000000000005800000000",
            INIT_01 => X"0000006c0000000000000081000000000000008d000000000000009000000000",
            INIT_02 => X"0000009d00000000000000af00000000000000a5000000000000008b00000000",
            INIT_03 => X"0000009f00000000000000860000000000000086000000000000009e00000000",
            INIT_04 => X"0000009800000000000000930000000000000094000000000000009a00000000",
            INIT_05 => X"0000003100000000000000490000000000000087000000000000009a00000000",
            INIT_06 => X"00000067000000000000004b0000000000000023000000000000001e00000000",
            INIT_07 => X"00000039000000000000002c000000000000003d000000000000006f00000000",
            INIT_08 => X"0000007400000000000000570000000000000057000000000000005600000000",
            INIT_09 => X"0000006900000000000000910000000000000093000000000000008f00000000",
            INIT_0A => X"0000006c000000000000008500000000000000b3000000000000008000000000",
            INIT_0B => X"00000079000000000000007a000000000000008b000000000000009100000000",
            INIT_0C => X"00000079000000000000007c0000000000000087000000000000007d00000000",
            INIT_0D => X"00000018000000000000002a0000000000000058000000000000007200000000",
            INIT_0E => X"000000660000000000000049000000000000001d000000000000001300000000",
            INIT_0F => X"0000002e00000000000000270000000000000050000000000000007500000000",
            INIT_10 => X"00000076000000000000004d000000000000005c000000000000005c00000000",
            INIT_11 => X"0000006200000000000000910000000000000099000000000000009c00000000",
            INIT_12 => X"0000007a000000000000007400000000000000aa000000000000005c00000000",
            INIT_13 => X"00000062000000000000004b000000000000008300000000000000a500000000",
            INIT_14 => X"0000004000000000000000550000000000000061000000000000004c00000000",
            INIT_15 => X"0000001b0000000000000011000000000000001b000000000000003600000000",
            INIT_16 => X"0000007500000000000000450000000000000028000000000000001a00000000",
            INIT_17 => X"0000002800000000000000240000000000000064000000000000007f00000000",
            INIT_18 => X"0000006e000000000000003c0000000000000054000000000000005e00000000",
            INIT_19 => X"00000073000000000000009b00000000000000a3000000000000009c00000000",
            INIT_1A => X"000000890000000000000094000000000000007c000000000000002700000000",
            INIT_1B => X"0000009c00000000000000570000000000000071000000000000009500000000",
            INIT_1C => X"00000027000000000000003d0000000000000050000000000000007800000000",
            INIT_1D => X"0000002e00000000000000220000000000000018000000000000002700000000",
            INIT_1E => X"000000780000000000000045000000000000002d000000000000001f00000000",
            INIT_1F => X"000000200000000000000022000000000000007b000000000000009900000000",
            INIT_20 => X"000000720000000000000059000000000000005d000000000000006100000000",
            INIT_21 => X"00000075000000000000009800000000000000a2000000000000009600000000",
            INIT_22 => X"000000740000000000000064000000000000001d000000000000000d00000000",
            INIT_23 => X"0000007c00000000000000490000000000000056000000000000007300000000",
            INIT_24 => X"0000001b000000000000002f000000000000005b000000000000008600000000",
            INIT_25 => X"0000003200000000000000310000000000000032000000000000003100000000",
            INIT_26 => X"0000007d0000000000000042000000000000001e000000000000001900000000",
            INIT_27 => X"000000200000000000000038000000000000009600000000000000a200000000",
            INIT_28 => X"0000006300000000000000570000000000000068000000000000006a00000000",
            INIT_29 => X"0000005700000000000000810000000000000096000000000000008d00000000",
            INIT_2A => X"000000250000000000000016000000000000000b000000000000000f00000000",
            INIT_2B => X"0000003e00000000000000290000000000000039000000000000003600000000",
            INIT_2C => X"0000001a00000000000000360000000000000048000000000000005300000000",
            INIT_2D => X"0000003300000000000000220000000000000023000000000000002000000000",
            INIT_2E => X"00000070000000000000003e000000000000002b000000000000002800000000",
            INIT_2F => X"0000001f000000000000004a000000000000009e000000000000009b00000000",
            INIT_30 => X"0000005a000000000000004f0000000000000068000000000000007000000000",
            INIT_31 => X"0000004200000000000000730000000000000089000000000000007b00000000",
            INIT_32 => X"0000001700000000000000280000000000000042000000000000002f00000000",
            INIT_33 => X"00000045000000000000002c0000000000000026000000000000001b00000000",
            INIT_34 => X"0000001d0000000000000026000000000000001f000000000000003600000000",
            INIT_35 => X"0000001f000000000000000f0000000000000016000000000000001900000000",
            INIT_36 => X"0000004e000000000000003a0000000000000033000000000000003100000000",
            INIT_37 => X"0000001f00000000000000570000000000000094000000000000008600000000",
            INIT_38 => X"0000006000000000000000590000000000000058000000000000006d00000000",
            INIT_39 => X"0000005e00000000000000730000000000000081000000000000006900000000",
            INIT_3A => X"0000003c00000000000000360000000000000047000000000000006100000000",
            INIT_3B => X"0000003c000000000000004b000000000000003e000000000000004200000000",
            INIT_3C => X"0000000e0000000000000009000000000000000a000000000000001a00000000",
            INIT_3D => X"0000000c000000000000000b0000000000000013000000000000001100000000",
            INIT_3E => X"0000003b000000000000003a000000000000001f000000000000001700000000",
            INIT_3F => X"0000002300000000000000690000000000000088000000000000005e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007000000000000000600000000000000046000000000000005b00000000",
            INIT_41 => X"0000009300000000000000890000000000000068000000000000006000000000",
            INIT_42 => X"000000430000000000000045000000000000003a000000000000007500000000",
            INIT_43 => X"00000035000000000000003f0000000000000045000000000000004a00000000",
            INIT_44 => X"0000000d00000000000000130000000000000019000000000000002900000000",
            INIT_45 => X"00000012000000000000000d0000000000000009000000000000000c00000000",
            INIT_46 => X"00000027000000000000003e0000000000000024000000000000000c00000000",
            INIT_47 => X"0000004700000000000000790000000000000068000000000000003400000000",
            INIT_48 => X"000000620000000000000062000000000000005c000000000000005b00000000",
            INIT_49 => X"0000008600000000000000690000000000000056000000000000006100000000",
            INIT_4A => X"00000061000000000000007c000000000000006b000000000000008e00000000",
            INIT_4B => X"00000049000000000000004e0000000000000049000000000000004400000000",
            INIT_4C => X"0000001c0000000000000026000000000000002b000000000000003e00000000",
            INIT_4D => X"00000014000000000000000b000000000000000e000000000000001600000000",
            INIT_4E => X"000000140000000000000030000000000000002a000000000000001400000000",
            INIT_4F => X"0000006400000000000000580000000000000038000000000000002500000000",
            INIT_50 => X"000000620000000000000061000000000000005e000000000000005b00000000",
            INIT_51 => X"0000004c000000000000005b000000000000006f000000000000007100000000",
            INIT_52 => X"000000510000000000000050000000000000006e000000000000008400000000",
            INIT_53 => X"000000540000000000000063000000000000005f000000000000004700000000",
            INIT_54 => X"000000330000000000000038000000000000003d000000000000004800000000",
            INIT_55 => X"0000002b0000000000000020000000000000002b000000000000003500000000",
            INIT_56 => X"0000002800000000000000250000000000000028000000000000002e00000000",
            INIT_57 => X"000000420000000000000030000000000000005a000000000000004000000000",
            INIT_58 => X"0000005200000000000000500000000000000060000000000000005700000000",
            INIT_59 => X"000000480000000000000062000000000000006d000000000000007100000000",
            INIT_5A => X"0000004600000000000000450000000000000073000000000000005c00000000",
            INIT_5B => X"000000580000000000000060000000000000005e000000000000004a00000000",
            INIT_5C => X"0000004a000000000000004c0000000000000047000000000000004500000000",
            INIT_5D => X"0000004b000000000000003d000000000000003c000000000000004200000000",
            INIT_5E => X"00000041000000000000003f0000000000000040000000000000004900000000",
            INIT_5F => X"0000003a0000000000000036000000000000005e000000000000004c00000000",
            INIT_60 => X"0000004c00000000000000430000000000000061000000000000006000000000",
            INIT_61 => X"00000050000000000000004e000000000000005a000000000000006900000000",
            INIT_62 => X"00000062000000000000004c0000000000000048000000000000005700000000",
            INIT_63 => X"0000005a000000000000005d000000000000005c000000000000005700000000",
            INIT_64 => X"0000004600000000000000550000000000000054000000000000004f00000000",
            INIT_65 => X"00000057000000000000004d0000000000000048000000000000004200000000",
            INIT_66 => X"0000004f00000000000000500000000000000052000000000000005300000000",
            INIT_67 => X"0000005e00000000000000460000000000000035000000000000004300000000",
            INIT_68 => X"0000006500000000000000510000000000000054000000000000004900000000",
            INIT_69 => X"0000005b0000000000000058000000000000005b000000000000006100000000",
            INIT_6A => X"00000063000000000000005b0000000000000059000000000000006900000000",
            INIT_6B => X"0000005a000000000000005d000000000000005d000000000000005900000000",
            INIT_6C => X"0000003c00000000000000490000000000000055000000000000005800000000",
            INIT_6D => X"0000005b00000000000000540000000000000052000000000000004900000000",
            INIT_6E => X"0000005500000000000000570000000000000056000000000000005d00000000",
            INIT_6F => X"0000006400000000000000570000000000000044000000000000004300000000",
            INIT_70 => X"00000071000000000000006a0000000000000060000000000000005300000000",
            INIT_71 => X"0000005f0000000000000060000000000000005f000000000000006000000000",
            INIT_72 => X"00000068000000000000006d0000000000000069000000000000006600000000",
            INIT_73 => X"0000004a0000000000000052000000000000005a000000000000005b00000000",
            INIT_74 => X"0000004a000000000000004d000000000000004e000000000000005200000000",
            INIT_75 => X"0000005c00000000000000570000000000000055000000000000004d00000000",
            INIT_76 => X"00000054000000000000005a0000000000000059000000000000006400000000",
            INIT_77 => X"0000005a0000000000000057000000000000004d000000000000004e00000000",
            INIT_78 => X"000000680000000000000071000000000000006b000000000000005c00000000",
            INIT_79 => X"0000005c000000000000004d0000000000000042000000000000005200000000",
            INIT_7A => X"0000005a000000000000005b0000000000000051000000000000005f00000000",
            INIT_7B => X"0000003d000000000000004d000000000000005b000000000000005800000000",
            INIT_7C => X"000000520000000000000056000000000000004d000000000000004600000000",
            INIT_7D => X"00000060000000000000005b000000000000005c000000000000005300000000",
            INIT_7E => X"0000005b0000000000000057000000000000005c000000000000006500000000",
            INIT_7F => X"00000057000000000000005b000000000000005a000000000000005c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "sampleifmap_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000001a000000000000003d000000000000005300000000",
            INIT_01 => X"00000036000000000000003a0000000000000043000000000000004100000000",
            INIT_02 => X"0000003b00000000000000340000000000000041000000000000003f00000000",
            INIT_03 => X"00000034000000000000002e0000000000000035000000000000003e00000000",
            INIT_04 => X"00000027000000000000002b0000000000000041000000000000004700000000",
            INIT_05 => X"00000026000000000000002d000000000000002f000000000000002f00000000",
            INIT_06 => X"00000032000000000000002a000000000000002d000000000000002f00000000",
            INIT_07 => X"000000290000000000000029000000000000002e000000000000004500000000",
            INIT_08 => X"00000046000000000000003a0000000000000035000000000000006100000000",
            INIT_09 => X"0000004d00000000000000440000000000000043000000000000004600000000",
            INIT_0A => X"0000003900000000000000380000000000000041000000000000004400000000",
            INIT_0B => X"0000002e00000000000000320000000000000039000000000000003400000000",
            INIT_0C => X"00000026000000000000002b0000000000000034000000000000003c00000000",
            INIT_0D => X"00000028000000000000002c000000000000002f000000000000002f00000000",
            INIT_0E => X"00000038000000000000002b000000000000001e000000000000002000000000",
            INIT_0F => X"0000003100000000000000330000000000000035000000000000004300000000",
            INIT_10 => X"00000051000000000000005c0000000000000047000000000000006400000000",
            INIT_11 => X"0000004e00000000000000440000000000000039000000000000004400000000",
            INIT_12 => X"0000003b000000000000003f0000000000000047000000000000004000000000",
            INIT_13 => X"0000003000000000000000310000000000000030000000000000003400000000",
            INIT_14 => X"0000001e00000000000000210000000000000032000000000000003b00000000",
            INIT_15 => X"0000003800000000000000350000000000000030000000000000002b00000000",
            INIT_16 => X"0000003800000000000000390000000000000038000000000000003300000000",
            INIT_17 => X"00000031000000000000002f0000000000000035000000000000003900000000",
            INIT_18 => X"000000590000000000000061000000000000005f000000000000006000000000",
            INIT_19 => X"0000004800000000000000490000000000000037000000000000004900000000",
            INIT_1A => X"000000420000000000000042000000000000004e000000000000004100000000",
            INIT_1B => X"0000003f00000000000000360000000000000037000000000000004300000000",
            INIT_1C => X"00000012000000000000001a000000000000002e000000000000002f00000000",
            INIT_1D => X"00000035000000000000002f0000000000000029000000000000002200000000",
            INIT_1E => X"0000003e00000000000000400000000000000044000000000000003d00000000",
            INIT_1F => X"0000003c000000000000003a000000000000002d000000000000003000000000",
            INIT_20 => X"0000005700000000000000540000000000000061000000000000005c00000000",
            INIT_21 => X"0000004b000000000000004c000000000000003f000000000000004900000000",
            INIT_22 => X"0000004b000000000000004b000000000000004a000000000000004a00000000",
            INIT_23 => X"0000003b0000000000000035000000000000003b000000000000004300000000",
            INIT_24 => X"0000001e00000000000000330000000000000034000000000000003b00000000",
            INIT_25 => X"00000027000000000000002e0000000000000029000000000000001f00000000",
            INIT_26 => X"0000003d000000000000003d000000000000003b000000000000002e00000000",
            INIT_27 => X"0000003c000000000000003a0000000000000030000000000000003400000000",
            INIT_28 => X"0000005900000000000000470000000000000066000000000000006500000000",
            INIT_29 => X"0000004c000000000000004c0000000000000046000000000000005100000000",
            INIT_2A => X"00000047000000000000004e0000000000000051000000000000004c00000000",
            INIT_2B => X"0000003100000000000000350000000000000043000000000000004400000000",
            INIT_2C => X"0000003900000000000000480000000000000041000000000000004300000000",
            INIT_2D => X"000000320000000000000042000000000000003e000000000000002b00000000",
            INIT_2E => X"0000003a00000000000000380000000000000036000000000000003800000000",
            INIT_2F => X"00000041000000000000003c000000000000003d000000000000003c00000000",
            INIT_30 => X"0000006300000000000000490000000000000059000000000000007800000000",
            INIT_31 => X"0000004b00000000000000510000000000000050000000000000005300000000",
            INIT_32 => X"0000004200000000000000550000000000000057000000000000005100000000",
            INIT_33 => X"000000350000000000000043000000000000004f000000000000004c00000000",
            INIT_34 => X"0000004d000000000000004a0000000000000040000000000000003c00000000",
            INIT_35 => X"0000002f00000000000000410000000000000040000000000000004100000000",
            INIT_36 => X"00000030000000000000002d0000000000000036000000000000003500000000",
            INIT_37 => X"00000042000000000000003f000000000000003d000000000000003a00000000",
            INIT_38 => X"0000005b000000000000005b000000000000003b000000000000007500000000",
            INIT_39 => X"00000054000000000000004f0000000000000051000000000000005100000000",
            INIT_3A => X"0000004800000000000000560000000000000056000000000000005700000000",
            INIT_3B => X"0000003f000000000000004a000000000000004c000000000000004d00000000",
            INIT_3C => X"00000049000000000000004c0000000000000049000000000000004200000000",
            INIT_3D => X"0000002f0000000000000038000000000000002f000000000000004700000000",
            INIT_3E => X"0000002a00000000000000230000000000000031000000000000002c00000000",
            INIT_3F => X"00000040000000000000003e0000000000000039000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000051000000000000005b0000000000000054000000000000005c00000000",
            INIT_41 => X"000000500000000000000050000000000000004f000000000000005300000000",
            INIT_42 => X"0000004600000000000000490000000000000053000000000000005800000000",
            INIT_43 => X"0000003d00000000000000430000000000000048000000000000005100000000",
            INIT_44 => X"0000004600000000000000460000000000000041000000000000004300000000",
            INIT_45 => X"0000003c000000000000004f0000000000000040000000000000004f00000000",
            INIT_46 => X"0000003b0000000000000034000000000000002d000000000000002c00000000",
            INIT_47 => X"00000040000000000000003d000000000000003d000000000000003a00000000",
            INIT_48 => X"0000005a000000000000004c0000000000000058000000000000006100000000",
            INIT_49 => X"0000004700000000000000530000000000000056000000000000005b00000000",
            INIT_4A => X"0000005300000000000000540000000000000052000000000000004f00000000",
            INIT_4B => X"00000055000000000000004d0000000000000053000000000000005800000000",
            INIT_4C => X"000000460000000000000039000000000000003e000000000000005100000000",
            INIT_4D => X"0000004b00000000000000590000000000000048000000000000005000000000",
            INIT_4E => X"0000003c000000000000003a0000000000000031000000000000002b00000000",
            INIT_4F => X"000000400000000000000039000000000000003f000000000000003a00000000",
            INIT_50 => X"0000006200000000000000560000000000000030000000000000005100000000",
            INIT_51 => X"000000540000000000000052000000000000005b000000000000005900000000",
            INIT_52 => X"0000005000000000000000500000000000000054000000000000005b00000000",
            INIT_53 => X"0000007e00000000000000670000000000000065000000000000005e00000000",
            INIT_54 => X"0000004300000000000000370000000000000049000000000000006b00000000",
            INIT_55 => X"000000440000000000000051000000000000004c000000000000004b00000000",
            INIT_56 => X"0000002d000000000000002f0000000000000031000000000000002000000000",
            INIT_57 => X"00000041000000000000003e000000000000003a000000000000003300000000",
            INIT_58 => X"0000004d0000000000000063000000000000001f000000000000001400000000",
            INIT_59 => X"0000005a000000000000005a0000000000000056000000000000004000000000",
            INIT_5A => X"0000005f00000000000000450000000000000045000000000000005f00000000",
            INIT_5B => X"0000007900000000000000670000000000000088000000000000008f00000000",
            INIT_5C => X"00000050000000000000003f0000000000000052000000000000007600000000",
            INIT_5D => X"000000210000000000000042000000000000004d000000000000005200000000",
            INIT_5E => X"0000002e00000000000000300000000000000030000000000000002100000000",
            INIT_5F => X"0000003f000000000000003b0000000000000036000000000000003000000000",
            INIT_60 => X"0000005c00000000000000700000000000000032000000000000000000000000",
            INIT_61 => X"000000620000000000000069000000000000007a000000000000006e00000000",
            INIT_62 => X"0000007700000000000000540000000000000048000000000000006000000000",
            INIT_63 => X"00000049000000000000005f000000000000007d000000000000009d00000000",
            INIT_64 => X"0000005400000000000000410000000000000047000000000000003400000000",
            INIT_65 => X"0000002a0000000000000041000000000000004f000000000000006000000000",
            INIT_66 => X"0000002900000000000000290000000000000025000000000000002500000000",
            INIT_67 => X"0000003a00000000000000390000000000000038000000000000002d00000000",
            INIT_68 => X"0000005c0000000000000061000000000000003c000000000000001400000000",
            INIT_69 => X"0000006f00000000000000700000000000000078000000000000007d00000000",
            INIT_6A => X"00000080000000000000006e000000000000004c000000000000005900000000",
            INIT_6B => X"0000006c00000000000000620000000000000064000000000000007f00000000",
            INIT_6C => X"0000005b00000000000000620000000000000063000000000000004400000000",
            INIT_6D => X"00000029000000000000003a000000000000004c000000000000006a00000000",
            INIT_6E => X"0000002600000000000000250000000000000023000000000000002100000000",
            INIT_6F => X"0000003500000000000000320000000000000034000000000000002e00000000",
            INIT_70 => X"00000058000000000000003a0000000000000046000000000000003b00000000",
            INIT_71 => X"00000073000000000000006a0000000000000075000000000000007b00000000",
            INIT_72 => X"0000007d00000000000000820000000000000067000000000000006600000000",
            INIT_73 => X"0000008900000000000000660000000000000050000000000000005f00000000",
            INIT_74 => X"00000084000000000000007e000000000000008c000000000000008300000000",
            INIT_75 => X"0000002a0000000000000040000000000000004e000000000000006f00000000",
            INIT_76 => X"00000032000000000000002a0000000000000028000000000000002b00000000",
            INIT_77 => X"00000031000000000000002e0000000000000032000000000000002f00000000",
            INIT_78 => X"0000005e00000000000000320000000000000035000000000000004900000000",
            INIT_79 => X"00000062000000000000006c000000000000007c000000000000007e00000000",
            INIT_7A => X"00000088000000000000008a000000000000007d000000000000007200000000",
            INIT_7B => X"0000008c00000000000000710000000000000062000000000000007b00000000",
            INIT_7C => X"0000008c000000000000008a0000000000000089000000000000008f00000000",
            INIT_7D => X"0000003300000000000000490000000000000069000000000000007500000000",
            INIT_7E => X"0000004d00000000000000320000000000000023000000000000002f00000000",
            INIT_7F => X"00000032000000000000002d000000000000002d000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "sampleifmap_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000056000000000000003a0000000000000041000000000000004800000000",
            INIT_01 => X"0000005300000000000000690000000000000075000000000000007700000000",
            INIT_02 => X"0000008200000000000000930000000000000089000000000000006e00000000",
            INIT_03 => X"00000087000000000000006d000000000000006b000000000000008200000000",
            INIT_04 => X"00000083000000000000007e000000000000007f000000000000008400000000",
            INIT_05 => X"0000002a000000000000003d0000000000000077000000000000008700000000",
            INIT_06 => X"00000055000000000000003c000000000000001b000000000000001a00000000",
            INIT_07 => X"0000003300000000000000240000000000000033000000000000006100000000",
            INIT_08 => X"0000006600000000000000510000000000000048000000000000004700000000",
            INIT_09 => X"00000050000000000000007a000000000000007c000000000000007800000000",
            INIT_0A => X"00000054000000000000006a0000000000000097000000000000006300000000",
            INIT_0B => X"0000005c00000000000000650000000000000079000000000000007c00000000",
            INIT_0C => X"0000006500000000000000680000000000000073000000000000006300000000",
            INIT_0D => X"00000011000000000000001f0000000000000048000000000000005e00000000",
            INIT_0E => X"00000055000000000000003a0000000000000015000000000000000e00000000",
            INIT_0F => X"00000029000000000000001f0000000000000046000000000000006800000000",
            INIT_10 => X"000000640000000000000044000000000000004e000000000000004f00000000",
            INIT_11 => X"0000004b000000000000007d0000000000000088000000000000008600000000",
            INIT_12 => X"00000061000000000000005b0000000000000093000000000000004700000000",
            INIT_13 => X"0000004800000000000000370000000000000071000000000000008e00000000",
            INIT_14 => X"000000320000000000000045000000000000004f000000000000003500000000",
            INIT_15 => X"00000016000000000000000d0000000000000014000000000000002a00000000",
            INIT_16 => X"0000006000000000000000370000000000000023000000000000001400000000",
            INIT_17 => X"00000023000000000000001e000000000000005b000000000000006f00000000",
            INIT_18 => X"0000005800000000000000320000000000000048000000000000005100000000",
            INIT_19 => X"0000005d000000000000008a0000000000000099000000000000008700000000",
            INIT_1A => X"00000071000000000000007f000000000000006f000000000000001f00000000",
            INIT_1B => X"0000008d0000000000000047000000000000005c000000000000007c00000000",
            INIT_1C => X"0000002100000000000000330000000000000041000000000000006700000000",
            INIT_1D => X"0000002c00000000000000240000000000000019000000000000002400000000",
            INIT_1E => X"000000600000000000000036000000000000002b000000000000001a00000000",
            INIT_1F => X"0000001a000000000000001e0000000000000073000000000000008900000000",
            INIT_20 => X"0000005f000000000000004f0000000000000052000000000000005300000000",
            INIT_21 => X"0000006200000000000000860000000000000096000000000000008200000000",
            INIT_22 => X"0000006300000000000000560000000000000017000000000000000a00000000",
            INIT_23 => X"000000740000000000000042000000000000004c000000000000006500000000",
            INIT_24 => X"000000170000000000000027000000000000004e000000000000007a00000000",
            INIT_25 => X"0000002e000000000000002f000000000000002f000000000000002e00000000",
            INIT_26 => X"000000670000000000000034000000000000001b000000000000001400000000",
            INIT_27 => X"00000019000000000000002f0000000000000089000000000000009200000000",
            INIT_28 => X"00000053000000000000004e000000000000005c000000000000005c00000000",
            INIT_29 => X"00000046000000000000006e0000000000000087000000000000007b00000000",
            INIT_2A => X"0000001d00000000000000100000000000000008000000000000000c00000000",
            INIT_2B => X"0000003800000000000000250000000000000034000000000000002f00000000",
            INIT_2C => X"00000012000000000000002b0000000000000039000000000000004600000000",
            INIT_2D => X"0000002c000000000000001d000000000000001c000000000000001900000000",
            INIT_2E => X"0000005e00000000000000310000000000000026000000000000002100000000",
            INIT_2F => X"00000018000000000000003d000000000000008d000000000000008c00000000",
            INIT_30 => X"0000004e0000000000000046000000000000005d000000000000006100000000",
            INIT_31 => X"0000003000000000000000600000000000000076000000000000006b00000000",
            INIT_32 => X"000000130000000000000022000000000000003a000000000000002500000000",
            INIT_33 => X"0000003b0000000000000026000000000000001f000000000000001300000000",
            INIT_34 => X"00000012000000000000001b0000000000000013000000000000002700000000",
            INIT_35 => X"00000018000000000000000a0000000000000011000000000000001100000000",
            INIT_36 => X"000000400000000000000030000000000000002c000000000000002a00000000",
            INIT_37 => X"0000001800000000000000460000000000000080000000000000007800000000",
            INIT_38 => X"000000580000000000000052000000000000004d000000000000005e00000000",
            INIT_39 => X"0000004b000000000000005f000000000000006b000000000000005b00000000",
            INIT_3A => X"0000003900000000000000300000000000000037000000000000004a00000000",
            INIT_3B => X"0000003300000000000000430000000000000035000000000000003a00000000",
            INIT_3C => X"0000000800000000000000030000000000000004000000000000001000000000",
            INIT_3D => X"0000000600000000000000070000000000000013000000000000000e00000000",
            INIT_3E => X"0000002f00000000000000300000000000000017000000000000001100000000",
            INIT_3F => X"0000001b00000000000000570000000000000073000000000000005100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000057000000000000003b000000000000004b00000000",
            INIT_41 => X"0000007e00000000000000750000000000000052000000000000005300000000",
            INIT_42 => X"0000003e00000000000000390000000000000022000000000000005500000000",
            INIT_43 => X"0000002e0000000000000039000000000000003d000000000000004200000000",
            INIT_44 => X"0000000d00000000000000120000000000000017000000000000002400000000",
            INIT_45 => X"0000000e000000000000000c000000000000000e000000000000000f00000000",
            INIT_46 => X"0000001e0000000000000036000000000000001c000000000000000700000000",
            INIT_47 => X"0000003e00000000000000680000000000000055000000000000002800000000",
            INIT_48 => X"000000560000000000000051000000000000004d000000000000004d00000000",
            INIT_49 => X"0000007000000000000000570000000000000045000000000000005500000000",
            INIT_4A => X"0000004f0000000000000064000000000000004f000000000000006f00000000",
            INIT_4B => X"0000003a00000000000000450000000000000043000000000000003b00000000",
            INIT_4C => X"0000001500000000000000200000000000000026000000000000003300000000",
            INIT_4D => X"0000000e0000000000000006000000000000000c000000000000001100000000",
            INIT_4E => X"0000000f00000000000000290000000000000022000000000000000f00000000",
            INIT_4F => X"0000005a000000000000004c000000000000002e000000000000001f00000000",
            INIT_50 => X"0000005500000000000000520000000000000051000000000000004f00000000",
            INIT_51 => X"00000039000000000000004a0000000000000060000000000000006500000000",
            INIT_52 => X"0000003e000000000000003a0000000000000057000000000000006d00000000",
            INIT_53 => X"00000044000000000000005a0000000000000058000000000000003d00000000",
            INIT_54 => X"0000002a000000000000002f0000000000000035000000000000003b00000000",
            INIT_55 => X"0000002300000000000000180000000000000023000000000000002c00000000",
            INIT_56 => X"0000001f000000000000001b000000000000001d000000000000002600000000",
            INIT_57 => X"0000003800000000000000270000000000000052000000000000003900000000",
            INIT_58 => X"0000004a000000000000004a0000000000000057000000000000004c00000000",
            INIT_59 => X"000000390000000000000053000000000000005f000000000000006600000000",
            INIT_5A => X"0000003a00000000000000370000000000000063000000000000004d00000000",
            INIT_5B => X"0000004d00000000000000570000000000000054000000000000003f00000000",
            INIT_5C => X"000000440000000000000043000000000000003c000000000000003900000000",
            INIT_5D => X"0000003f00000000000000310000000000000031000000000000003b00000000",
            INIT_5E => X"0000003300000000000000300000000000000031000000000000003c00000000",
            INIT_5F => X"0000002f000000000000002d0000000000000054000000000000003f00000000",
            INIT_60 => X"000000450000000000000040000000000000005a000000000000005500000000",
            INIT_61 => X"000000440000000000000041000000000000004e000000000000005e00000000",
            INIT_62 => X"0000005a0000000000000042000000000000003c000000000000004c00000000",
            INIT_63 => X"000000510000000000000053000000000000004e000000000000004a00000000",
            INIT_64 => X"00000040000000000000004c0000000000000047000000000000004300000000",
            INIT_65 => X"00000048000000000000003e0000000000000039000000000000003b00000000",
            INIT_66 => X"0000003e00000000000000400000000000000042000000000000004400000000",
            INIT_67 => X"00000053000000000000003d0000000000000029000000000000003200000000",
            INIT_68 => X"0000005c0000000000000049000000000000004b000000000000003d00000000",
            INIT_69 => X"00000050000000000000004e0000000000000051000000000000005700000000",
            INIT_6A => X"000000590000000000000050000000000000004c000000000000005d00000000",
            INIT_6B => X"00000050000000000000004e000000000000004c000000000000004a00000000",
            INIT_6C => X"00000035000000000000003e0000000000000045000000000000004a00000000",
            INIT_6D => X"0000004b00000000000000440000000000000042000000000000004000000000",
            INIT_6E => X"0000004400000000000000480000000000000048000000000000004d00000000",
            INIT_6F => X"00000059000000000000004e0000000000000038000000000000003200000000",
            INIT_70 => X"00000064000000000000005a0000000000000051000000000000004600000000",
            INIT_71 => X"0000005500000000000000570000000000000055000000000000005600000000",
            INIT_72 => X"0000005a000000000000005d0000000000000057000000000000005600000000",
            INIT_73 => X"0000003c000000000000003f0000000000000046000000000000004a00000000",
            INIT_74 => X"0000003e000000000000003e000000000000003c000000000000004200000000",
            INIT_75 => X"0000004c00000000000000470000000000000046000000000000004100000000",
            INIT_76 => X"00000047000000000000004e000000000000004d000000000000005500000000",
            INIT_77 => X"0000004f000000000000004d0000000000000041000000000000003e00000000",
            INIT_78 => X"00000059000000000000005f000000000000005d000000000000004f00000000",
            INIT_79 => X"0000005100000000000000460000000000000039000000000000004600000000",
            INIT_7A => X"0000004700000000000000470000000000000040000000000000005300000000",
            INIT_7B => X"0000002f000000000000003d000000000000004c000000000000004a00000000",
            INIT_7C => X"000000460000000000000048000000000000003f000000000000003800000000",
            INIT_7D => X"00000050000000000000004b000000000000004c000000000000004500000000",
            INIT_7E => X"0000004e0000000000000049000000000000004f000000000000005600000000",
            INIT_7F => X"00000049000000000000004f000000000000004c000000000000004f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "sampleifmap_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d900000000000000d100000000000000b900000000000000a000000000",
            INIT_01 => X"000000f600000000000000f900000000000000f600000000000000e600000000",
            INIT_02 => X"000000dd00000000000000e600000000000000f300000000000000f800000000",
            INIT_03 => X"000000c700000000000000d800000000000000dd00000000000000da00000000",
            INIT_04 => X"000000b400000000000000b800000000000000bb00000000000000bc00000000",
            INIT_05 => X"0000008b0000000000000079000000000000009000000000000000a600000000",
            INIT_06 => X"0000004f00000000000000660000000000000066000000000000006a00000000",
            INIT_07 => X"0000005e000000000000005b0000000000000065000000000000005e00000000",
            INIT_08 => X"000000e600000000000000f200000000000000ef00000000000000e100000000",
            INIT_09 => X"000000eb00000000000000f300000000000000f500000000000000e800000000",
            INIT_0A => X"000000cd00000000000000d800000000000000e600000000000000ed00000000",
            INIT_0B => X"000000ba00000000000000c800000000000000cb00000000000000c900000000",
            INIT_0C => X"0000007f00000000000000a100000000000000ab00000000000000af00000000",
            INIT_0D => X"00000087000000000000007a000000000000008d000000000000008e00000000",
            INIT_0E => X"0000003400000000000000250000000000000052000000000000007600000000",
            INIT_0F => X"000000640000000000000061000000000000006b000000000000005f00000000",
            INIT_10 => X"000000dc00000000000000f100000000000000f900000000000000fc00000000",
            INIT_11 => X"000000d600000000000000df00000000000000e200000000000000d900000000",
            INIT_12 => X"000000b800000000000000c300000000000000cf00000000000000d500000000",
            INIT_13 => X"000000a700000000000000b300000000000000b600000000000000b300000000",
            INIT_14 => X"0000008100000000000000940000000000000098000000000000009f00000000",
            INIT_15 => X"000000720000000000000080000000000000008c000000000000008000000000",
            INIT_16 => X"0000002600000000000000040000000000000028000000000000005700000000",
            INIT_17 => X"0000006900000000000000690000000000000073000000000000006300000000",
            INIT_18 => X"000000d300000000000000de00000000000000e100000000000000e900000000",
            INIT_19 => X"000000c000000000000000c800000000000000cb00000000000000d300000000",
            INIT_1A => X"000000a400000000000000ae00000000000000b700000000000000bb00000000",
            INIT_1B => X"0000009900000000000000a000000000000000a500000000000000a000000000",
            INIT_1C => X"0000008a000000000000008c000000000000008d000000000000009100000000",
            INIT_1D => X"00000069000000000000007f000000000000007d000000000000007d00000000",
            INIT_1E => X"00000037000000000000001a0000000000000025000000000000003b00000000",
            INIT_1F => X"0000006d00000000000000700000000000000078000000000000007000000000",
            INIT_20 => X"000000c900000000000000cf00000000000000c300000000000000cf00000000",
            INIT_21 => X"000000ab00000000000000b300000000000000b400000000000000be00000000",
            INIT_22 => X"000000920000000000000099000000000000009f00000000000000a300000000",
            INIT_23 => X"0000008d00000000000000930000000000000097000000000000009100000000",
            INIT_24 => X"0000008700000000000000830000000000000088000000000000008700000000",
            INIT_25 => X"0000005a0000000000000084000000000000007a000000000000008100000000",
            INIT_26 => X"000000560000000000000030000000000000003d000000000000003a00000000",
            INIT_27 => X"0000006d00000000000000720000000000000078000000000000007500000000",
            INIT_28 => X"000000a200000000000000aa00000000000000ab00000000000000b600000000",
            INIT_29 => X"00000097000000000000009f000000000000009c000000000000009900000000",
            INIT_2A => X"0000008a000000000000008c000000000000008d000000000000009000000000",
            INIT_2B => X"0000008a000000000000008a000000000000008d000000000000008b00000000",
            INIT_2C => X"0000008a0000000000000086000000000000008c000000000000008700000000",
            INIT_2D => X"0000004500000000000000660000000000000089000000000000008c00000000",
            INIT_2E => X"000000740000000000000043000000000000003e000000000000004b00000000",
            INIT_2F => X"0000006e00000000000000700000000000000080000000000000008100000000",
            INIT_30 => X"0000008600000000000000880000000000000088000000000000008d00000000",
            INIT_31 => X"00000085000000000000008c0000000000000086000000000000008800000000",
            INIT_32 => X"0000008d000000000000008b0000000000000089000000000000008700000000",
            INIT_33 => X"00000091000000000000008e0000000000000092000000000000008f00000000",
            INIT_34 => X"0000008f000000000000008a0000000000000091000000000000009100000000",
            INIT_35 => X"00000021000000000000002f000000000000006b000000000000008e00000000",
            INIT_36 => X"0000007f000000000000006c000000000000004b000000000000004800000000",
            INIT_37 => X"00000070000000000000006f0000000000000084000000000000008400000000",
            INIT_38 => X"000000810000000000000080000000000000007d000000000000007600000000",
            INIT_39 => X"00000084000000000000008a0000000000000083000000000000008800000000",
            INIT_3A => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_3B => X"00000099000000000000009a000000000000009e000000000000009600000000",
            INIT_3C => X"0000009400000000000000930000000000000095000000000000009200000000",
            INIT_3D => X"00000011000000000000000d0000000000000042000000000000008000000000",
            INIT_3E => X"0000007a00000000000000800000000000000075000000000000005000000000",
            INIT_3F => X"0000007000000000000000720000000000000080000000000000007b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000850000000000000084000000000000007e000000000000007300000000",
            INIT_41 => X"00000089000000000000008f0000000000000087000000000000008b00000000",
            INIT_42 => X"0000009800000000000000950000000000000091000000000000008b00000000",
            INIT_43 => X"000000aa00000000000000a3000000000000009a000000000000009400000000",
            INIT_44 => X"00000094000000000000009d00000000000000a2000000000000009e00000000",
            INIT_45 => X"0000001e000000000000000e000000000000002c000000000000007300000000",
            INIT_46 => X"0000007e0000000000000088000000000000008b000000000000006900000000",
            INIT_47 => X"0000006f0000000000000074000000000000007a000000000000007700000000",
            INIT_48 => X"0000008800000000000000880000000000000080000000000000007600000000",
            INIT_49 => X"0000008d00000000000000910000000000000088000000000000008d00000000",
            INIT_4A => X"000000a5000000000000009a0000000000000093000000000000008d00000000",
            INIT_4B => X"000000a700000000000000a2000000000000009a000000000000009d00000000",
            INIT_4C => X"0000008a00000000000000910000000000000093000000000000009b00000000",
            INIT_4D => X"00000037000000000000002e0000000000000038000000000000006300000000",
            INIT_4E => X"0000007e000000000000007a000000000000007c000000000000006d00000000",
            INIT_4F => X"0000006e00000000000000750000000000000074000000000000007300000000",
            INIT_50 => X"00000089000000000000008b0000000000000084000000000000007d00000000",
            INIT_51 => X"0000008c00000000000000900000000000000088000000000000008e00000000",
            INIT_52 => X"0000009900000000000000960000000000000090000000000000008b00000000",
            INIT_53 => X"000000980000000000000090000000000000008b000000000000008300000000",
            INIT_54 => X"000000d600000000000000d300000000000000ba00000000000000a600000000",
            INIT_55 => X"0000002a0000000000000045000000000000005c000000000000008000000000",
            INIT_56 => X"000000730000000000000063000000000000005f000000000000005500000000",
            INIT_57 => X"0000006b0000000000000071000000000000006f000000000000007000000000",
            INIT_58 => X"0000008a000000000000008e0000000000000089000000000000008500000000",
            INIT_59 => X"0000008a000000000000008e0000000000000088000000000000008d00000000",
            INIT_5A => X"000000840000000000000088000000000000008f000000000000008900000000",
            INIT_5B => X"000000cb00000000000000c900000000000000b6000000000000008e00000000",
            INIT_5C => X"000000c000000000000000cf00000000000000ce00000000000000d200000000",
            INIT_5D => X"0000002a000000000000009200000000000000bd00000000000000a200000000",
            INIT_5E => X"0000007200000000000000670000000000000028000000000000001b00000000",
            INIT_5F => X"00000068000000000000006c000000000000006a000000000000006d00000000",
            INIT_60 => X"0000008b000000000000008f000000000000008b000000000000008c00000000",
            INIT_61 => X"00000089000000000000008a000000000000008c000000000000008f00000000",
            INIT_62 => X"000000a400000000000000900000000000000085000000000000008700000000",
            INIT_63 => X"00000073000000000000008900000000000000a000000000000000ab00000000",
            INIT_64 => X"0000003b000000000000004b000000000000005d000000000000006a00000000",
            INIT_65 => X"0000005f00000000000000c900000000000000dc000000000000006f00000000",
            INIT_66 => X"00000074000000000000003e0000000000000007000000000000000d00000000",
            INIT_67 => X"0000006400000000000000690000000000000065000000000000006300000000",
            INIT_68 => X"0000008c000000000000008f000000000000008a000000000000009000000000",
            INIT_69 => X"0000008700000000000000820000000000000092000000000000009200000000",
            INIT_6A => X"0000006e000000000000008c0000000000000091000000000000008200000000",
            INIT_6B => X"000000130000000000000031000000000000005c000000000000005e00000000",
            INIT_6C => X"0000001200000000000000190000000000000032000000000000001d00000000",
            INIT_6D => X"0000009d00000000000000d200000000000000d1000000000000007800000000",
            INIT_6E => X"0000004400000000000000130000000000000006000000000000002600000000",
            INIT_6F => X"0000005f00000000000000630000000000000052000000000000004500000000",
            INIT_70 => X"0000008e0000000000000092000000000000008b000000000000009100000000",
            INIT_71 => X"000000800000000000000079000000000000008e000000000000009000000000",
            INIT_72 => X"000000440000000000000054000000000000007f000000000000008500000000",
            INIT_73 => X"00000016000000000000002e0000000000000052000000000000005600000000",
            INIT_74 => X"00000041000000000000001e0000000000000032000000000000001300000000",
            INIT_75 => X"000000cb00000000000000cd00000000000000c900000000000000af00000000",
            INIT_76 => X"0000001600000000000000120000000000000010000000000000006600000000",
            INIT_77 => X"00000058000000000000004f0000000000000038000000000000002300000000",
            INIT_78 => X"000000900000000000000094000000000000008b000000000000008f00000000",
            INIT_79 => X"00000083000000000000008b0000000000000084000000000000008a00000000",
            INIT_7A => X"0000005600000000000000480000000000000042000000000000007500000000",
            INIT_7B => X"000000220000000000000028000000000000004e000000000000006a00000000",
            INIT_7C => X"000000b600000000000000730000000000000046000000000000002400000000",
            INIT_7D => X"000000c300000000000000cd00000000000000c500000000000000cb00000000",
            INIT_7E => X"000000120000000000000025000000000000003d000000000000006c00000000",
            INIT_7F => X"000000530000000000000064000000000000004f000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "sampleifmap_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000900000000000000093000000000000008b000000000000008e00000000",
            INIT_01 => X"0000007900000000000000840000000000000072000000000000008500000000",
            INIT_02 => X"00000045000000000000003c0000000000000059000000000000005100000000",
            INIT_03 => X"0000009b00000000000000530000000000000044000000000000005500000000",
            INIT_04 => X"000000eb00000000000000ed00000000000000db00000000000000c000000000",
            INIT_05 => X"0000007200000000000000d300000000000000d700000000000000d700000000",
            INIT_06 => X"000000140000000000000035000000000000005d000000000000003000000000",
            INIT_07 => X"00000054000000000000008f000000000000008b000000000000004100000000",
            INIT_08 => X"00000089000000000000008e000000000000008d000000000000008f00000000",
            INIT_09 => X"00000043000000000000003a0000000000000045000000000000007400000000",
            INIT_0A => X"0000001c000000000000001d000000000000004b000000000000005100000000",
            INIT_0B => X"000000f2000000000000008c0000000000000019000000000000002400000000",
            INIT_0C => X"000000dc00000000000000e300000000000000eb00000000000000ec00000000",
            INIT_0D => X"0000003a000000000000009500000000000000df00000000000000db00000000",
            INIT_0E => X"0000004e000000000000004e0000000000000054000000000000003900000000",
            INIT_0F => X"0000005b00000000000000a700000000000000a1000000000000008500000000",
            INIT_10 => X"000000860000000000000088000000000000008c000000000000008f00000000",
            INIT_11 => X"00000034000000000000002d0000000000000047000000000000008d00000000",
            INIT_12 => X"0000001600000000000000170000000000000021000000000000004300000000",
            INIT_13 => X"000000d9000000000000009b0000000000000029000000000000002f00000000",
            INIT_14 => X"000000d000000000000000bf00000000000000be00000000000000c700000000",
            INIT_15 => X"0000006700000000000000ad00000000000000df00000000000000dc00000000",
            INIT_16 => X"0000009500000000000000870000000000000073000000000000005d00000000",
            INIT_17 => X"0000005900000000000000a50000000000000094000000000000009800000000",
            INIT_18 => X"000000b5000000000000007e000000000000008c000000000000008f00000000",
            INIT_19 => X"0000002b0000000000000021000000000000004c00000000000000bd00000000",
            INIT_1A => X"0000001700000000000000100000000000000015000000000000003900000000",
            INIT_1B => X"000000c2000000000000009e0000000000000042000000000000003900000000",
            INIT_1C => X"000000c900000000000000c400000000000000b300000000000000b600000000",
            INIT_1D => X"000000b300000000000000de00000000000000ce00000000000000c200000000",
            INIT_1E => X"000000970000000000000095000000000000009c000000000000009700000000",
            INIT_1F => X"0000004200000000000000880000000000000092000000000000009600000000",
            INIT_20 => X"000000ea000000000000009a0000000000000085000000000000008c00000000",
            INIT_21 => X"0000002a0000000000000026000000000000005a00000000000000b500000000",
            INIT_22 => X"0000000b000000000000000b000000000000000b000000000000003400000000",
            INIT_23 => X"000000ba00000000000000a00000000000000031000000000000001400000000",
            INIT_24 => X"0000007300000000000000b900000000000000b900000000000000b000000000",
            INIT_25 => X"000000c400000000000000a1000000000000005a000000000000004500000000",
            INIT_26 => X"0000009900000000000000a000000000000000aa00000000000000b700000000",
            INIT_27 => X"00000026000000000000004d0000000000000088000000000000009300000000",
            INIT_28 => X"000000a300000000000000a30000000000000080000000000000008200000000",
            INIT_29 => X"0000002e000000000000002d000000000000006a000000000000008b00000000",
            INIT_2A => X"0000000f00000000000000090000000000000003000000000000001c00000000",
            INIT_2B => X"000000b400000000000000a20000000000000036000000000000001e00000000",
            INIT_2C => X"00000015000000000000007100000000000000be00000000000000ac00000000",
            INIT_2D => X"0000009500000000000000300000000000000015000000000000001400000000",
            INIT_2E => X"00000085000000000000008e00000000000000ab00000000000000bb00000000",
            INIT_2F => X"0000002700000000000000150000000000000043000000000000008000000000",
            INIT_30 => X"0000001a00000000000000670000000000000084000000000000007c00000000",
            INIT_31 => X"000000300000000000000034000000000000006c000000000000004800000000",
            INIT_32 => X"0000003b000000000000000b0000000000000007000000000000001200000000",
            INIT_33 => X"000000b000000000000000a50000000000000063000000000000005a00000000",
            INIT_34 => X"0000001d000000000000002a00000000000000a900000000000000b100000000",
            INIT_35 => X"00000046000000000000000e0000000000000026000000000000002f00000000",
            INIT_36 => X"0000007500000000000000750000000000000088000000000000009500000000",
            INIT_37 => X"000000300000000000000015000000000000000e000000000000003c00000000",
            INIT_38 => X"0000001e0000000000000049000000000000007c000000000000007900000000",
            INIT_39 => X"0000001f00000000000000440000000000000072000000000000003b00000000",
            INIT_3A => X"000000480000000000000018000000000000000e000000000000000d00000000",
            INIT_3B => X"000000bb00000000000000bb000000000000006c000000000000004f00000000",
            INIT_3C => X"0000002b000000000000001b000000000000008b00000000000000bf00000000",
            INIT_3D => X"0000001b000000000000001c000000000000001b000000000000001e00000000",
            INIT_3E => X"00000059000000000000007b0000000000000084000000000000006c00000000",
            INIT_3F => X"0000003b000000000000002a0000000000000015000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003f00000000000000470000000000000066000000000000006d00000000",
            INIT_41 => X"0000001c000000000000004d0000000000000071000000000000003c00000000",
            INIT_42 => X"000000470000000000000030000000000000001f000000000000001000000000",
            INIT_43 => X"000000b300000000000000bd0000000000000088000000000000004600000000",
            INIT_44 => X"00000036000000000000001f000000000000007400000000000000b400000000",
            INIT_45 => X"0000000e000000000000001b0000000000000029000000000000003500000000",
            INIT_46 => X"0000003c000000000000007c0000000000000085000000000000004800000000",
            INIT_47 => X"0000003b00000000000000320000000000000022000000000000001200000000",
            INIT_48 => X"0000003c000000000000003d0000000000000051000000000000005700000000",
            INIT_49 => X"00000015000000000000004b0000000000000069000000000000003a00000000",
            INIT_4A => X"00000060000000000000004c000000000000002e000000000000001400000000",
            INIT_4B => X"000000a300000000000000a40000000000000091000000000000006100000000",
            INIT_4C => X"000000390000000000000020000000000000007100000000000000aa00000000",
            INIT_4D => X"0000001100000000000000250000000000000031000000000000004700000000",
            INIT_4E => X"000000210000000000000060000000000000006c000000000000002900000000",
            INIT_4F => X"000000320000000000000028000000000000001d000000000000000c00000000",
            INIT_50 => X"0000003c00000000000000400000000000000049000000000000004900000000",
            INIT_51 => X"0000002f0000000000000057000000000000005f000000000000003900000000",
            INIT_52 => X"000000a500000000000000890000000000000062000000000000003d00000000",
            INIT_53 => X"000000b600000000000000b700000000000000b000000000000000a900000000",
            INIT_54 => X"000000360000000000000022000000000000007c00000000000000b600000000",
            INIT_55 => X"0000001b0000000000000033000000000000005c000000000000006000000000",
            INIT_56 => X"0000000c000000000000003b0000000000000046000000000000001100000000",
            INIT_57 => X"00000028000000000000001d0000000000000012000000000000000600000000",
            INIT_58 => X"0000004e00000000000000450000000000000049000000000000004900000000",
            INIT_59 => X"0000002f00000000000000450000000000000059000000000000004100000000",
            INIT_5A => X"00000056000000000000004a000000000000003c000000000000003400000000",
            INIT_5B => X"0000006000000000000000620000000000000060000000000000005b00000000",
            INIT_5C => X"0000003c00000000000000200000000000000053000000000000006200000000",
            INIT_5D => X"00000014000000000000001d000000000000003e000000000000003b00000000",
            INIT_5E => X"00000003000000000000000a0000000000000011000000000000000400000000",
            INIT_5F => X"000000210000000000000011000000000000000a000000000000000700000000",
            INIT_60 => X"0000003600000000000000480000000000000053000000000000004b00000000",
            INIT_61 => X"00000004000000000000000f0000000000000027000000000000002d00000000",
            INIT_62 => X"0000000700000000000000050000000000000002000000000000000300000000",
            INIT_63 => X"0000000b000000000000000a0000000000000008000000000000000700000000",
            INIT_64 => X"000000420000000000000008000000000000000d000000000000000b00000000",
            INIT_65 => X"0000000f0000000000000038000000000000002f000000000000004300000000",
            INIT_66 => X"0000000300000000000000010000000000000002000000000000000200000000",
            INIT_67 => X"00000020000000000000000f000000000000000a000000000000000600000000",
            INIT_68 => X"0000002f00000000000000510000000000000059000000000000005000000000",
            INIT_69 => X"000000190000000000000010000000000000000a000000000000001500000000",
            INIT_6A => X"0000000e000000000000000e000000000000000a000000000000000e00000000",
            INIT_6B => X"0000000c000000000000000e000000000000000e000000000000000e00000000",
            INIT_6C => X"0000001700000000000000060000000000000009000000000000000a00000000",
            INIT_6D => X"00000007000000000000002a0000000000000048000000000000003e00000000",
            INIT_6E => X"0000000500000000000000050000000000000004000000000000000300000000",
            INIT_6F => X"000000210000000000000015000000000000000b000000000000000700000000",
            INIT_70 => X"000000370000000000000049000000000000004f000000000000004900000000",
            INIT_71 => X"0000003a000000000000003b000000000000002f000000000000002e00000000",
            INIT_72 => X"0000001c00000000000000190000000000000011000000000000001a00000000",
            INIT_73 => X"0000001c000000000000001d0000000000000020000000000000001f00000000",
            INIT_74 => X"0000000c00000000000000100000000000000015000000000000001800000000",
            INIT_75 => X"0000000600000000000000080000000000000016000000000000001400000000",
            INIT_76 => X"0000000800000000000000080000000000000007000000000000000800000000",
            INIT_77 => X"0000001f000000000000001b000000000000000f000000000000000b00000000",
            INIT_78 => X"0000004e000000000000004c0000000000000048000000000000004500000000",
            INIT_79 => X"0000003800000000000000480000000000000053000000000000005800000000",
            INIT_7A => X"0000002a000000000000002b0000000000000026000000000000002000000000",
            INIT_7B => X"0000003100000000000000320000000000000033000000000000002f00000000",
            INIT_7C => X"0000001c000000000000001e0000000000000026000000000000002c00000000",
            INIT_7D => X"0000000c00000000000000130000000000000022000000000000002200000000",
            INIT_7E => X"0000000d000000000000000f0000000000000010000000000000000e00000000",
            INIT_7F => X"0000001d000000000000001e000000000000001a000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "sampleifmap_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003a00000000000000390000000000000031000000000000002500000000",
            INIT_01 => X"000000510000000000000050000000000000004e000000000000004200000000",
            INIT_02 => X"0000004200000000000000490000000000000052000000000000005600000000",
            INIT_03 => X"0000003800000000000000430000000000000043000000000000004100000000",
            INIT_04 => X"0000007300000000000000400000000000000032000000000000003200000000",
            INIT_05 => X"0000002700000000000000320000000000000038000000000000003400000000",
            INIT_06 => X"00000024000000000000002e0000000000000022000000000000001600000000",
            INIT_07 => X"0000001300000000000000150000000000000012000000000000001d00000000",
            INIT_08 => X"00000044000000000000004d0000000000000048000000000000004300000000",
            INIT_09 => X"000000420000000000000048000000000000004a000000000000004300000000",
            INIT_0A => X"0000003400000000000000390000000000000040000000000000004400000000",
            INIT_0B => X"0000002e00000000000000370000000000000036000000000000003200000000",
            INIT_0C => X"000000290000000000000027000000000000002a000000000000002900000000",
            INIT_0D => X"00000021000000000000001e0000000000000023000000000000002800000000",
            INIT_0E => X"0000001b000000000000001e000000000000002e000000000000002200000000",
            INIT_0F => X"0000001200000000000000160000000000000015000000000000001c00000000",
            INIT_10 => X"0000003e00000000000000480000000000000044000000000000004800000000",
            INIT_11 => X"000000310000000000000038000000000000003d000000000000003a00000000",
            INIT_12 => X"00000028000000000000002b000000000000002d000000000000003000000000",
            INIT_13 => X"00000026000000000000002b000000000000002a000000000000002600000000",
            INIT_14 => X"0000001c000000000000001e0000000000000023000000000000002200000000",
            INIT_15 => X"00000022000000000000001f0000000000000021000000000000002300000000",
            INIT_16 => X"0000000e000000000000000d0000000000000022000000000000003000000000",
            INIT_17 => X"0000001100000000000000130000000000000014000000000000001500000000",
            INIT_18 => X"0000003c000000000000003d0000000000000036000000000000003800000000",
            INIT_19 => X"00000024000000000000002b0000000000000030000000000000003e00000000",
            INIT_1A => X"0000002000000000000000220000000000000023000000000000002300000000",
            INIT_1B => X"0000002000000000000000220000000000000021000000000000001f00000000",
            INIT_1C => X"0000001d000000000000001b000000000000001e000000000000001d00000000",
            INIT_1D => X"00000025000000000000001d000000000000001c000000000000002000000000",
            INIT_1E => X"0000000f000000000000000b0000000000000012000000000000002a00000000",
            INIT_1F => X"0000001100000000000000100000000000000013000000000000001600000000",
            INIT_20 => X"0000003b00000000000000420000000000000039000000000000003900000000",
            INIT_21 => X"0000001b00000000000000200000000000000024000000000000003400000000",
            INIT_22 => X"0000001a000000000000001c000000000000001d000000000000001c00000000",
            INIT_23 => X"0000001e000000000000001c000000000000001a000000000000001a00000000",
            INIT_24 => X"0000001c000000000000001c000000000000001c000000000000001c00000000",
            INIT_25 => X"0000002a00000000000000430000000000000030000000000000001c00000000",
            INIT_26 => X"00000019000000000000000d0000000000000012000000000000001900000000",
            INIT_27 => X"000000110000000000000013000000000000001f000000000000001b00000000",
            INIT_28 => X"00000021000000000000002f000000000000003a000000000000003b00000000",
            INIT_29 => X"000000160000000000000019000000000000001a000000000000001a00000000",
            INIT_2A => X"00000019000000000000001a0000000000000019000000000000001700000000",
            INIT_2B => X"0000001f000000000000001b0000000000000018000000000000001800000000",
            INIT_2C => X"0000001e0000000000000021000000000000001e000000000000001d00000000",
            INIT_2D => X"0000003c000000000000005e000000000000005d000000000000002100000000",
            INIT_2E => X"0000002c000000000000001e000000000000001b000000000000002900000000",
            INIT_2F => X"000000130000000000000018000000000000002d000000000000002b00000000",
            INIT_30 => X"000000140000000000000017000000000000001c000000000000002200000000",
            INIT_31 => X"0000001500000000000000160000000000000017000000000000001600000000",
            INIT_32 => X"0000001a00000000000000190000000000000016000000000000001600000000",
            INIT_33 => X"00000023000000000000001d0000000000000019000000000000001800000000",
            INIT_34 => X"0000001e0000000000000023000000000000001f000000000000002000000000",
            INIT_35 => X"0000002500000000000000370000000000000059000000000000003300000000",
            INIT_36 => X"0000002d000000000000002b0000000000000028000000000000003800000000",
            INIT_37 => X"000000150000000000000017000000000000001e000000000000002400000000",
            INIT_38 => X"0000001200000000000000100000000000000011000000000000001100000000",
            INIT_39 => X"0000001600000000000000160000000000000017000000000000001600000000",
            INIT_3A => X"0000001b000000000000001a0000000000000017000000000000001800000000",
            INIT_3B => X"00000027000000000000001d000000000000001b000000000000001900000000",
            INIT_3C => X"000000300000000000000033000000000000002d000000000000002800000000",
            INIT_3D => X"0000000b00000000000000120000000000000040000000000000004100000000",
            INIT_3E => X"00000020000000000000001f0000000000000025000000000000002200000000",
            INIT_3F => X"0000001500000000000000160000000000000016000000000000001900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000120000000000000012000000000000001100000000",
            INIT_41 => X"0000001700000000000000170000000000000016000000000000001500000000",
            INIT_42 => X"0000001e000000000000001c0000000000000018000000000000001900000000",
            INIT_43 => X"0000003b00000000000000330000000000000038000000000000002500000000",
            INIT_44 => X"000000360000000000000037000000000000003a000000000000003b00000000",
            INIT_45 => X"0000001000000000000000110000000000000028000000000000003d00000000",
            INIT_46 => X"0000001b00000000000000180000000000000019000000000000001a00000000",
            INIT_47 => X"0000001400000000000000150000000000000017000000000000001a00000000",
            INIT_48 => X"0000001200000000000000120000000000000012000000000000001300000000",
            INIT_49 => X"0000001800000000000000160000000000000014000000000000001500000000",
            INIT_4A => X"0000003100000000000000200000000000000019000000000000001800000000",
            INIT_4B => X"000000340000000000000039000000000000004c000000000000003e00000000",
            INIT_4C => X"0000003a0000000000000032000000000000002e000000000000003100000000",
            INIT_4D => X"0000002c00000000000000300000000000000031000000000000003800000000",
            INIT_4E => X"0000001900000000000000190000000000000023000000000000002900000000",
            INIT_4F => X"0000001400000000000000140000000000000018000000000000001900000000",
            INIT_50 => X"0000001200000000000000130000000000000012000000000000001400000000",
            INIT_51 => X"0000001700000000000000150000000000000015000000000000001500000000",
            INIT_52 => X"0000003500000000000000240000000000000019000000000000001900000000",
            INIT_53 => X"0000004a000000000000003e0000000000000042000000000000003100000000",
            INIT_54 => X"000000b800000000000000a60000000000000089000000000000006800000000",
            INIT_55 => X"00000021000000000000004b0000000000000068000000000000007c00000000",
            INIT_56 => X"000000190000000000000026000000000000003d000000000000003800000000",
            INIT_57 => X"0000001300000000000000120000000000000019000000000000001800000000",
            INIT_58 => X"0000001300000000000000140000000000000012000000000000001500000000",
            INIT_59 => X"0000001800000000000000160000000000000018000000000000001800000000",
            INIT_5A => X"00000030000000000000001f000000000000001d000000000000001900000000",
            INIT_5B => X"000000be00000000000000b20000000000000097000000000000005500000000",
            INIT_5C => X"000000c500000000000000ca00000000000000cd00000000000000cd00000000",
            INIT_5D => X"00000016000000000000009800000000000000d000000000000000b200000000",
            INIT_5E => X"0000002800000000000000460000000000000025000000000000001800000000",
            INIT_5F => X"0000001100000000000000110000000000000016000000000000001500000000",
            INIT_60 => X"0000001500000000000000160000000000000014000000000000001400000000",
            INIT_61 => X"0000001a00000000000000190000000000000018000000000000001800000000",
            INIT_62 => X"0000007000000000000000420000000000000020000000000000001900000000",
            INIT_63 => X"00000075000000000000008c000000000000009b000000000000009000000000",
            INIT_64 => X"0000003d00000000000000470000000000000058000000000000006400000000",
            INIT_65 => X"0000004e00000000000000d500000000000000e8000000000000007500000000",
            INIT_66 => X"000000460000000000000032000000000000000a000000000000000f00000000",
            INIT_67 => X"0000001000000000000000110000000000000015000000000000001a00000000",
            INIT_68 => X"0000001600000000000000190000000000000016000000000000001400000000",
            INIT_69 => X"0000001a00000000000000190000000000000017000000000000001700000000",
            INIT_6A => X"0000005b00000000000000670000000000000048000000000000001a00000000",
            INIT_6B => X"0000001200000000000000340000000000000056000000000000005000000000",
            INIT_6C => X"00000010000000000000000f0000000000000022000000000000001100000000",
            INIT_6D => X"0000009b00000000000000e000000000000000dd000000000000007c00000000",
            INIT_6E => X"0000003b00000000000000160000000000000007000000000000002400000000",
            INIT_6F => X"0000001000000000000000120000000000000013000000000000002100000000",
            INIT_70 => X"00000016000000000000001b0000000000000017000000000000001800000000",
            INIT_71 => X"0000001500000000000000130000000000000019000000000000001800000000",
            INIT_72 => X"00000029000000000000003a0000000000000055000000000000003700000000",
            INIT_73 => X"000000180000000000000032000000000000004e000000000000003d00000000",
            INIT_74 => X"00000049000000000000001e000000000000002b000000000000000b00000000",
            INIT_75 => X"000000cd00000000000000d100000000000000d800000000000000bf00000000",
            INIT_76 => X"000000170000000000000010000000000000000e000000000000006700000000",
            INIT_77 => X"0000001200000000000000140000000000000016000000000000001b00000000",
            INIT_78 => X"00000017000000000000001a0000000000000016000000000000001a00000000",
            INIT_79 => X"00000034000000000000003c0000000000000025000000000000001900000000",
            INIT_7A => X"0000003b00000000000000380000000000000034000000000000004c00000000",
            INIT_7B => X"00000026000000000000002e000000000000004d000000000000005000000000",
            INIT_7C => X"000000c4000000000000007c0000000000000049000000000000002300000000",
            INIT_7D => X"000000d200000000000000d900000000000000d800000000000000df00000000",
            INIT_7E => X"0000000e00000000000000150000000000000039000000000000007600000000",
            INIT_7F => X"00000011000000000000003e0000000000000047000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "sampleifmap_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001700000000000000190000000000000014000000000000001900000000",
            INIT_01 => X"0000005c00000000000000600000000000000035000000000000002100000000",
            INIT_02 => X"00000042000000000000003e000000000000005d000000000000004900000000",
            INIT_03 => X"000000a2000000000000005a0000000000000047000000000000005100000000",
            INIT_04 => X"000000f500000000000000f500000000000000df00000000000000c400000000",
            INIT_05 => X"0000007900000000000000de00000000000000e400000000000000e300000000",
            INIT_06 => X"000000090000000000000011000000000000003b000000000000002500000000",
            INIT_07 => X"000000130000000000000075000000000000008c000000000000004800000000",
            INIT_08 => X"0000001a00000000000000180000000000000015000000000000001900000000",
            INIT_09 => X"000000450000000000000035000000000000002c000000000000002800000000",
            INIT_0A => X"0000002900000000000000250000000000000052000000000000005800000000",
            INIT_0B => X"000000fb00000000000000940000000000000020000000000000003100000000",
            INIT_0C => X"000000e200000000000000e900000000000000f200000000000000f600000000",
            INIT_0D => X"0000001f000000000000008b00000000000000e200000000000000e100000000",
            INIT_0E => X"0000004300000000000000280000000000000019000000000000000b00000000",
            INIT_0F => X"00000022000000000000009700000000000000a2000000000000008500000000",
            INIT_10 => X"0000002600000000000000160000000000000013000000000000001600000000",
            INIT_11 => X"00000036000000000000002e0000000000000046000000000000005d00000000",
            INIT_12 => X"0000001b00000000000000180000000000000026000000000000004b00000000",
            INIT_13 => X"000000e300000000000000a30000000000000031000000000000003800000000",
            INIT_14 => X"000000da00000000000000cb00000000000000cd00000000000000d600000000",
            INIT_15 => X"0000004a00000000000000a300000000000000e400000000000000e500000000",
            INIT_16 => X"000000950000000000000080000000000000005a000000000000003900000000",
            INIT_17 => X"0000003300000000000000a00000000000000096000000000000009700000000",
            INIT_18 => X"0000007c0000000000000026000000000000000f000000000000001300000000",
            INIT_19 => X"0000002a0000000000000024000000000000005a00000000000000af00000000",
            INIT_1A => X"00000015000000000000000b0000000000000017000000000000003f00000000",
            INIT_1B => X"000000d000000000000000aa000000000000004f000000000000004000000000",
            INIT_1C => X"000000d600000000000000d300000000000000c500000000000000c700000000",
            INIT_1D => X"000000b100000000000000e300000000000000d900000000000000ce00000000",
            INIT_1E => X"000000a200000000000000a700000000000000a8000000000000009800000000",
            INIT_1F => X"0000002a00000000000000880000000000000097000000000000009a00000000",
            INIT_20 => X"000000dc0000000000000065000000000000000a000000000000001200000000",
            INIT_21 => X"0000002e000000000000002f000000000000006f00000000000000be00000000",
            INIT_22 => X"0000000e0000000000000009000000000000000a000000000000003900000000",
            INIT_23 => X"000000cc00000000000000b10000000000000042000000000000001f00000000",
            INIT_24 => X"0000007c00000000000000c600000000000000ca00000000000000c200000000",
            INIT_25 => X"000000d300000000000000ac0000000000000066000000000000004f00000000",
            INIT_26 => X"000000a900000000000000b100000000000000b800000000000000c800000000",
            INIT_27 => X"00000011000000000000004a000000000000008c000000000000009c00000000",
            INIT_28 => X"000000a500000000000000840000000000000014000000000000000e00000000",
            INIT_29 => X"0000003400000000000000370000000000000080000000000000009600000000",
            INIT_2A => X"00000016000000000000000a0000000000000003000000000000001e00000000",
            INIT_2B => X"000000c600000000000000b40000000000000048000000000000002d00000000",
            INIT_2C => X"00000019000000000000007b00000000000000cd00000000000000be00000000",
            INIT_2D => X"000000a30000000000000038000000000000001e000000000000001a00000000",
            INIT_2E => X"00000093000000000000009e00000000000000b800000000000000ca00000000",
            INIT_2F => X"00000011000000000000000d0000000000000044000000000000008800000000",
            INIT_30 => X"0000002100000000000000530000000000000023000000000000000a00000000",
            INIT_31 => X"00000035000000000000003e0000000000000082000000000000005300000000",
            INIT_32 => X"0000004800000000000000100000000000000007000000000000001300000000",
            INIT_33 => X"000000c200000000000000b70000000000000075000000000000006c00000000",
            INIT_34 => X"0000001e000000000000002f00000000000000b700000000000000c300000000",
            INIT_35 => X"0000004f0000000000000014000000000000002b000000000000003100000000",
            INIT_36 => X"000000810000000000000084000000000000009400000000000000a100000000",
            INIT_37 => X"000000180000000000000009000000000000000a000000000000004000000000",
            INIT_38 => X"0000002300000000000000370000000000000021000000000000000a00000000",
            INIT_39 => X"00000024000000000000004e0000000000000088000000000000004600000000",
            INIT_3A => X"0000005800000000000000220000000000000011000000000000000f00000000",
            INIT_3B => X"000000cd00000000000000cd000000000000007e000000000000006100000000",
            INIT_3C => X"0000002b0000000000000020000000000000009800000000000000d000000000",
            INIT_3D => X"0000001f0000000000000020000000000000001f000000000000002000000000",
            INIT_3E => X"00000063000000000000008a0000000000000091000000000000007500000000",
            INIT_3F => X"000000210000000000000019000000000000000c000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004100000000000000360000000000000015000000000000000a00000000",
            INIT_41 => X"0000002100000000000000570000000000000088000000000000004700000000",
            INIT_42 => X"00000057000000000000003f0000000000000027000000000000001500000000",
            INIT_43 => X"000000c500000000000000cf000000000000009a000000000000005600000000",
            INIT_44 => X"000000380000000000000025000000000000008100000000000000c600000000",
            INIT_45 => X"0000000f000000000000001c000000000000002c000000000000003700000000",
            INIT_46 => X"00000043000000000000008b0000000000000093000000000000004d00000000",
            INIT_47 => X"0000001f000000000000001c0000000000000014000000000000000e00000000",
            INIT_48 => X"0000003e000000000000002f000000000000000e000000000000000700000000",
            INIT_49 => X"0000001c00000000000000560000000000000080000000000000004500000000",
            INIT_4A => X"0000006f000000000000005e000000000000003c000000000000001e00000000",
            INIT_4B => X"000000b400000000000000b600000000000000a2000000000000006f00000000",
            INIT_4C => X"0000003c0000000000000029000000000000007f00000000000000bc00000000",
            INIT_4D => X"0000000f00000000000000230000000000000035000000000000004b00000000",
            INIT_4E => X"00000026000000000000006f000000000000007a000000000000002c00000000",
            INIT_4F => X"000000160000000000000010000000000000000d000000000000000700000000",
            INIT_50 => X"0000003b00000000000000270000000000000011000000000000000b00000000",
            INIT_51 => X"0000003d00000000000000680000000000000075000000000000004600000000",
            INIT_52 => X"000000b7000000000000009f0000000000000079000000000000005100000000",
            INIT_53 => X"000000c700000000000000c900000000000000c300000000000000b900000000",
            INIT_54 => X"0000003c000000000000002a000000000000008800000000000000c600000000",
            INIT_55 => X"0000001c00000000000000340000000000000062000000000000006600000000",
            INIT_56 => X"000000100000000000000045000000000000004f000000000000001500000000",
            INIT_57 => X"00000016000000000000000c0000000000000007000000000000000300000000",
            INIT_58 => X"00000043000000000000001d0000000000000014000000000000001300000000",
            INIT_59 => X"0000003c00000000000000550000000000000067000000000000004900000000",
            INIT_5A => X"00000064000000000000005b0000000000000050000000000000004500000000",
            INIT_5B => X"0000006d00000000000000710000000000000071000000000000006800000000",
            INIT_5C => X"0000004100000000000000250000000000000059000000000000006d00000000",
            INIT_5D => X"00000017000000000000001f0000000000000042000000000000004000000000",
            INIT_5E => X"00000005000000000000000e0000000000000014000000000000000800000000",
            INIT_5F => X"00000018000000000000000b0000000000000006000000000000000600000000",
            INIT_60 => X"00000025000000000000001d000000000000001c000000000000001700000000",
            INIT_61 => X"000000070000000000000016000000000000002c000000000000002c00000000",
            INIT_62 => X"0000000c000000000000000c000000000000000a000000000000000a00000000",
            INIT_63 => X"0000001000000000000000110000000000000010000000000000000d00000000",
            INIT_64 => X"000000430000000000000009000000000000000f000000000000000f00000000",
            INIT_65 => X"0000001000000000000000380000000000000030000000000000004400000000",
            INIT_66 => X"0000000400000000000000030000000000000003000000000000000400000000",
            INIT_67 => X"00000019000000000000000e0000000000000009000000000000000600000000",
            INIT_68 => X"0000002000000000000000270000000000000025000000000000002100000000",
            INIT_69 => X"0000002000000000000000190000000000000012000000000000001700000000",
            INIT_6A => X"0000001700000000000000170000000000000015000000000000001700000000",
            INIT_6B => X"0000000f00000000000000130000000000000015000000000000001700000000",
            INIT_6C => X"000000180000000000000007000000000000000a000000000000000b00000000",
            INIT_6D => X"0000000800000000000000290000000000000047000000000000003e00000000",
            INIT_6E => X"0000000600000000000000050000000000000005000000000000000400000000",
            INIT_6F => X"0000001d0000000000000018000000000000000e000000000000000900000000",
            INIT_70 => X"0000003200000000000000290000000000000025000000000000002300000000",
            INIT_71 => X"0000004d00000000000000510000000000000043000000000000003c00000000",
            INIT_72 => X"00000030000000000000002d0000000000000024000000000000002c00000000",
            INIT_73 => X"000000230000000000000027000000000000002c000000000000003100000000",
            INIT_74 => X"000000100000000000000015000000000000001b000000000000001d00000000",
            INIT_75 => X"00000009000000000000000a0000000000000019000000000000001700000000",
            INIT_76 => X"0000000b000000000000000a0000000000000009000000000000000b00000000",
            INIT_77 => X"0000001e000000000000001f0000000000000014000000000000000e00000000",
            INIT_78 => X"00000057000000000000003b000000000000002a000000000000002a00000000",
            INIT_79 => X"000000520000000000000066000000000000006f000000000000006d00000000",
            INIT_7A => X"000000470000000000000045000000000000003e000000000000003700000000",
            INIT_7B => X"0000004300000000000000460000000000000048000000000000004a00000000",
            INIT_7C => X"00000029000000000000002b0000000000000033000000000000003b00000000",
            INIT_7D => X"000000120000000000000018000000000000002c000000000000002f00000000",
            INIT_7E => X"0000001300000000000000150000000000000016000000000000001400000000",
            INIT_7F => X"0000001e0000000000000020000000000000001c000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "sampleifmap_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a000000000000000e000000000000000b000000000000000d00000000",
            INIT_01 => X"000000020000000000000005000000000000000a000000000000000900000000",
            INIT_02 => X"0000000200000000000000010000000000000003000000000000000300000000",
            INIT_03 => X"0000000000000000000000050000000000000006000000000000000400000000",
            INIT_04 => X"0000005600000000000000230000000000000000000000000000000100000000",
            INIT_05 => X"00000008000000000000001d0000000000000017000000000000001600000000",
            INIT_06 => X"0000001d0000000000000027000000000000001b000000000000000d00000000",
            INIT_07 => X"0000000500000000000000060000000000000008000000000000001300000000",
            INIT_08 => X"00000004000000000000000a000000000000000c000000000000000d00000000",
            INIT_09 => X"0000000000000000000000030000000000000008000000000000000700000000",
            INIT_0A => X"0000000100000000000000010000000000000002000000000000000400000000",
            INIT_0B => X"0000000100000000000000040000000000000004000000000000000200000000",
            INIT_0C => X"0000001300000000000000100000000000000001000000000000000100000000",
            INIT_0D => X"0000000700000000000000060000000000000006000000000000000700000000",
            INIT_0E => X"000000160000000000000017000000000000002e000000000000002100000000",
            INIT_0F => X"0000000600000000000000040000000000000008000000000000001300000000",
            INIT_10 => X"0000000000000000000000030000000000000004000000000000000700000000",
            INIT_11 => X"0000000000000000000000010000000000000004000000000000000400000000",
            INIT_12 => X"0000000400000000000000040000000000000004000000000000000400000000",
            INIT_13 => X"0000000300000000000000050000000000000006000000000000000400000000",
            INIT_14 => X"00000009000000000000000c0000000000000003000000000000000400000000",
            INIT_15 => X"0000000a00000000000000060000000000000007000000000000000400000000",
            INIT_16 => X"0000000c000000000000000d0000000000000023000000000000002800000000",
            INIT_17 => X"0000000600000000000000030000000000000006000000000000000f00000000",
            INIT_18 => X"0000000b00000000000000080000000000000003000000000000000100000000",
            INIT_19 => X"0000000300000000000000030000000000000004000000000000001200000000",
            INIT_1A => X"0000000700000000000000080000000000000006000000000000000500000000",
            INIT_1B => X"0000000600000000000000060000000000000009000000000000000800000000",
            INIT_1C => X"00000009000000000000000a0000000000000005000000000000000700000000",
            INIT_1D => X"000000170000000000000010000000000000000a000000000000000400000000",
            INIT_1E => X"0000000e00000000000000110000000000000016000000000000001e00000000",
            INIT_1F => X"0000000800000000000000050000000000000006000000000000000f00000000",
            INIT_20 => X"0000001a000000000000001d0000000000000013000000000000000c00000000",
            INIT_21 => X"0000000800000000000000070000000000000006000000000000001700000000",
            INIT_22 => X"0000000800000000000000090000000000000008000000000000000700000000",
            INIT_23 => X"000000080000000000000007000000000000000a000000000000000900000000",
            INIT_24 => X"0000000700000000000000080000000000000007000000000000000900000000",
            INIT_25 => X"0000002700000000000000400000000000000025000000000000000800000000",
            INIT_26 => X"00000015000000000000000e0000000000000010000000000000001000000000",
            INIT_27 => X"00000009000000000000000d000000000000000f000000000000000e00000000",
            INIT_28 => X"0000000c0000000000000016000000000000001e000000000000001800000000",
            INIT_29 => X"0000000800000000000000090000000000000006000000000000000900000000",
            INIT_2A => X"0000000a00000000000000090000000000000005000000000000000500000000",
            INIT_2B => X"000000090000000000000007000000000000000a000000000000000b00000000",
            INIT_2C => X"00000007000000000000000b000000000000000b000000000000000a00000000",
            INIT_2D => X"0000003b000000000000005d0000000000000055000000000000001400000000",
            INIT_2E => X"000000200000000000000013000000000000000e000000000000002200000000",
            INIT_2F => X"000000090000000000000010000000000000001b000000000000001700000000",
            INIT_30 => X"00000007000000000000000a000000000000000b000000000000000c00000000",
            INIT_31 => X"00000007000000000000000a0000000000000008000000000000000800000000",
            INIT_32 => X"0000000e000000000000000a0000000000000005000000000000000600000000",
            INIT_33 => X"0000000c000000000000000a000000000000000c000000000000000d00000000",
            INIT_34 => X"00000007000000000000000e000000000000000e000000000000000900000000",
            INIT_35 => X"00000028000000000000003c0000000000000056000000000000002500000000",
            INIT_36 => X"0000001c000000000000001c000000000000001c000000000000003500000000",
            INIT_37 => X"0000000700000000000000060000000000000010000000000000001400000000",
            INIT_38 => X"0000000700000000000000060000000000000006000000000000000300000000",
            INIT_39 => X"00000009000000000000000c000000000000000a000000000000000b00000000",
            INIT_3A => X"0000000e000000000000000c0000000000000008000000000000000900000000",
            INIT_3B => X"0000001300000000000000100000000000000012000000000000000e00000000",
            INIT_3C => X"00000016000000000000001a0000000000000015000000000000001000000000",
            INIT_3D => X"0000000a0000000000000014000000000000003e000000000000003100000000",
            INIT_3E => X"0000000d0000000000000010000000000000001a000000000000001e00000000",
            INIT_3F => X"0000000700000000000000040000000000000008000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000080000000000000009000000000000000a000000000000000700000000",
            INIT_41 => X"0000000b000000000000000e000000000000000a000000000000000b00000000",
            INIT_42 => X"0000000f000000000000000e000000000000000c000000000000000d00000000",
            INIT_43 => X"0000002800000000000000220000000000000024000000000000001300000000",
            INIT_44 => X"0000002200000000000000220000000000000020000000000000002400000000",
            INIT_45 => X"00000009000000000000000f000000000000002b000000000000003300000000",
            INIT_46 => X"0000000a0000000000000009000000000000000c000000000000001400000000",
            INIT_47 => X"0000000800000000000000080000000000000008000000000000000800000000",
            INIT_48 => X"00000008000000000000000b000000000000000c000000000000000c00000000",
            INIT_49 => X"0000000d000000000000000e000000000000000a000000000000000c00000000",
            INIT_4A => X"000000220000000000000014000000000000000e000000000000000e00000000",
            INIT_4B => X"0000002600000000000000280000000000000031000000000000002700000000",
            INIT_4C => X"000000320000000000000027000000000000001b000000000000002000000000",
            INIT_4D => X"000000260000000000000034000000000000003b000000000000003600000000",
            INIT_4E => X"0000000c000000000000000b0000000000000015000000000000002300000000",
            INIT_4F => X"0000000a000000000000000b0000000000000009000000000000000600000000",
            INIT_50 => X"00000009000000000000000b000000000000000b000000000000000c00000000",
            INIT_51 => X"0000000d000000000000000d000000000000000a000000000000000c00000000",
            INIT_52 => X"00000028000000000000001b0000000000000010000000000000000d00000000",
            INIT_53 => X"0000003f00000000000000320000000000000032000000000000002000000000",
            INIT_54 => X"000000b400000000000000a10000000000000077000000000000005800000000",
            INIT_55 => X"0000002200000000000000540000000000000071000000000000007900000000",
            INIT_56 => X"00000011000000000000001d0000000000000031000000000000003200000000",
            INIT_57 => X"0000000a000000000000000c000000000000000a000000000000000900000000",
            INIT_58 => X"0000000b000000000000000e000000000000000a000000000000000900000000",
            INIT_59 => X"0000000c000000000000000d000000000000000c000000000000000e00000000",
            INIT_5A => X"0000002700000000000000180000000000000012000000000000000c00000000",
            INIT_5B => X"000000ba00000000000000af0000000000000093000000000000004d00000000",
            INIT_5C => X"000000ca00000000000000d200000000000000c800000000000000c800000000",
            INIT_5D => X"0000001c000000000000009e00000000000000d500000000000000b100000000",
            INIT_5E => X"0000002500000000000000460000000000000022000000000000001300000000",
            INIT_5F => X"00000009000000000000000b0000000000000009000000000000000a00000000",
            INIT_60 => X"0000000d000000000000000f000000000000000a000000000000000800000000",
            INIT_61 => X"0000000e000000000000000d000000000000000e000000000000001000000000",
            INIT_62 => X"0000006c000000000000003e0000000000000018000000000000000c00000000",
            INIT_63 => X"0000007d000000000000009300000000000000a2000000000000008e00000000",
            INIT_64 => X"0000004a0000000000000054000000000000005e000000000000006e00000000",
            INIT_65 => X"0000005400000000000000d700000000000000f1000000000000007e00000000",
            INIT_66 => X"0000004900000000000000340000000000000009000000000000000c00000000",
            INIT_67 => X"000000080000000000000009000000000000000d000000000000001900000000",
            INIT_68 => X"0000000e000000000000000f000000000000000b000000000000000b00000000",
            INIT_69 => X"0000000e000000000000000c0000000000000010000000000000001100000000",
            INIT_6A => X"0000005d00000000000000670000000000000044000000000000001400000000",
            INIT_6B => X"00000019000000000000003d000000000000005f000000000000005600000000",
            INIT_6C => X"0000001700000000000000110000000000000023000000000000001600000000",
            INIT_6D => X"000000a700000000000000eb00000000000000eb000000000000008900000000",
            INIT_6E => X"0000004200000000000000170000000000000007000000000000002a00000000",
            INIT_6F => X"0000000700000000000000090000000000000011000000000000002800000000",
            INIT_70 => X"0000000e0000000000000012000000000000000d000000000000000f00000000",
            INIT_71 => X"00000012000000000000000b0000000000000012000000000000001000000000",
            INIT_72 => X"0000002e000000000000003b0000000000000053000000000000003600000000",
            INIT_73 => X"0000001b00000000000000370000000000000053000000000000004400000000",
            INIT_74 => X"0000004c000000000000001c0000000000000027000000000000000c00000000",
            INIT_75 => X"000000e000000000000000e700000000000000e800000000000000c800000000",
            INIT_76 => X"0000001a00000000000000130000000000000016000000000000007300000000",
            INIT_77 => X"00000008000000000000000d0000000000000016000000000000001f00000000",
            INIT_78 => X"0000000e0000000000000013000000000000000d000000000000001000000000",
            INIT_79 => X"000000370000000000000039000000000000001e000000000000000e00000000",
            INIT_7A => X"0000003c00000000000000390000000000000035000000000000004f00000000",
            INIT_7B => X"000000290000000000000032000000000000004e000000000000005200000000",
            INIT_7C => X"000000c8000000000000007c0000000000000047000000000000002300000000",
            INIT_7D => X"000000dd00000000000000ec00000000000000e600000000000000e700000000",
            INIT_7E => X"0000000e000000000000001a0000000000000044000000000000007e00000000",
            INIT_7F => X"00000009000000000000003f0000000000000049000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "sampleifmap_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000110000000000000013000000000000000e000000000000001100000000",
            INIT_01 => X"0000005c000000000000005d000000000000002f000000000000001800000000",
            INIT_02 => X"0000003d000000000000003c0000000000000062000000000000004f00000000",
            INIT_03 => X"000000a6000000000000005e0000000000000047000000000000004c00000000",
            INIT_04 => X"000000fc00000000000000fa00000000000000e200000000000000c600000000",
            INIT_05 => X"0000007c00000000000000e700000000000000f000000000000000ed00000000",
            INIT_06 => X"0000000c000000000000001c000000000000004a000000000000002a00000000",
            INIT_07 => X"00000011000000000000007e0000000000000095000000000000004c00000000",
            INIT_08 => X"0000001500000000000000120000000000000010000000000000001200000000",
            INIT_09 => X"000000480000000000000038000000000000002a000000000000002400000000",
            INIT_0A => X"0000002400000000000000240000000000000058000000000000006000000000",
            INIT_0B => X"00000100000000000000009a0000000000000022000000000000002d00000000",
            INIT_0C => X"000000ed00000000000000f400000000000000f900000000000000fa00000000",
            INIT_0D => X"00000027000000000000009600000000000000ee00000000000000ed00000000",
            INIT_0E => X"0000004d000000000000003b000000000000002e000000000000001500000000",
            INIT_0F => X"0000002600000000000000a300000000000000ae000000000000008e00000000",
            INIT_10 => X"0000002200000000000000100000000000000010000000000000001100000000",
            INIT_11 => X"00000042000000000000003c0000000000000049000000000000005c00000000",
            INIT_12 => X"00000021000000000000001c000000000000002c000000000000005400000000",
            INIT_13 => X"000000f000000000000000ae0000000000000037000000000000003e00000000",
            INIT_14 => X"000000e700000000000000d900000000000000d900000000000000e100000000",
            INIT_15 => X"0000005600000000000000b100000000000000ee00000000000000ef00000000",
            INIT_16 => X"000000a40000000000000092000000000000006a000000000000004500000000",
            INIT_17 => X"0000003700000000000000a900000000000000a100000000000000a400000000",
            INIT_18 => X"0000007d0000000000000020000000000000000a000000000000000d00000000",
            INIT_19 => X"000000380000000000000035000000000000006200000000000000b400000000",
            INIT_1A => X"0000001b000000000000000e000000000000001c000000000000004800000000",
            INIT_1B => X"000000e000000000000000b90000000000000059000000000000004900000000",
            INIT_1C => X"000000e300000000000000e400000000000000d500000000000000d500000000",
            INIT_1D => X"000000c000000000000000f200000000000000e100000000000000d700000000",
            INIT_1E => X"000000b000000000000000b500000000000000b400000000000000a500000000",
            INIT_1F => X"0000002a000000000000008d000000000000009f00000000000000a600000000",
            INIT_20 => X"000000e500000000000000650000000000000007000000000000000c00000000",
            INIT_21 => X"00000039000000000000003e000000000000007b00000000000000c900000000",
            INIT_22 => X"0000000f0000000000000009000000000000000f000000000000004100000000",
            INIT_23 => X"000000da00000000000000bf000000000000004f000000000000002600000000",
            INIT_24 => X"0000008a00000000000000d800000000000000db00000000000000d000000000",
            INIT_25 => X"000000e400000000000000b8000000000000006d000000000000005800000000",
            INIT_26 => X"000000b500000000000000bf00000000000000c900000000000000da00000000",
            INIT_27 => X"0000000e000000000000004d000000000000009300000000000000a600000000",
            INIT_28 => X"000000b3000000000000008b0000000000000018000000000000000d00000000",
            INIT_29 => X"0000003d0000000000000045000000000000008d00000000000000a200000000",
            INIT_2A => X"0000001b000000000000000b0000000000000004000000000000002300000000",
            INIT_2B => X"000000d400000000000000c20000000000000056000000000000003600000000",
            INIT_2C => X"00000024000000000000008800000000000000db00000000000000cc00000000",
            INIT_2D => X"000000b100000000000000400000000000000022000000000000002000000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000cc00000000000000dd00000000",
            INIT_2F => X"0000000d000000000000000f0000000000000049000000000000009000000000",
            INIT_30 => X"00000031000000000000005b0000000000000027000000000000000900000000",
            INIT_31 => X"0000003e000000000000004c000000000000008f000000000000006000000000",
            INIT_32 => X"0000005100000000000000150000000000000007000000000000001500000000",
            INIT_33 => X"000000d000000000000000c50000000000000083000000000000007900000000",
            INIT_34 => X"00000026000000000000003800000000000000c100000000000000d100000000",
            INIT_35 => X"000000590000000000000019000000000000002e000000000000003700000000",
            INIT_36 => X"0000008d000000000000009500000000000000a900000000000000b200000000",
            INIT_37 => X"000000140000000000000008000000000000000e000000000000004800000000",
            INIT_38 => X"00000030000000000000003b0000000000000022000000000000000500000000",
            INIT_39 => X"0000002d000000000000005c0000000000000095000000000000005300000000",
            INIT_3A => X"00000064000000000000002a0000000000000013000000000000000f00000000",
            INIT_3B => X"000000db00000000000000db000000000000008c000000000000006f00000000",
            INIT_3C => X"00000033000000000000002600000000000000a000000000000000de00000000",
            INIT_3D => X"0000002700000000000000240000000000000023000000000000002500000000",
            INIT_3E => X"0000006e000000000000009b00000000000000a4000000000000008200000000",
            INIT_3F => X"0000001e0000000000000016000000000000000c000000000000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d000000000000003a0000000000000017000000000000000700000000",
            INIT_41 => X"0000002a00000000000000650000000000000094000000000000005400000000",
            INIT_42 => X"00000065000000000000004a000000000000002b000000000000001600000000",
            INIT_43 => X"000000d300000000000000dd00000000000000a8000000000000006400000000",
            INIT_44 => X"00000040000000000000002b000000000000008900000000000000d400000000",
            INIT_45 => X"0000001500000000000000230000000000000034000000000000003f00000000",
            INIT_46 => X"0000004e000000000000009a00000000000000a2000000000000005600000000",
            INIT_47 => X"0000001c00000000000000180000000000000012000000000000001300000000",
            INIT_48 => X"0000004c00000000000000370000000000000015000000000000000900000000",
            INIT_49 => X"000000250000000000000065000000000000008c000000000000005200000000",
            INIT_4A => X"0000007f000000000000006c0000000000000043000000000000002100000000",
            INIT_4B => X"000000c200000000000000c300000000000000b0000000000000007e00000000",
            INIT_4C => X"000000460000000000000030000000000000008700000000000000c900000000",
            INIT_4D => X"00000015000000000000002e0000000000000041000000000000005600000000",
            INIT_4E => X"00000031000000000000007b0000000000000083000000000000003200000000",
            INIT_4F => X"00000014000000000000000b000000000000000a000000000000000b00000000",
            INIT_50 => X"0000004900000000000000310000000000000017000000000000000b00000000",
            INIT_51 => X"0000004b00000000000000780000000000000084000000000000005700000000",
            INIT_52 => X"000000c800000000000000b10000000000000086000000000000005d00000000",
            INIT_53 => X"000000d500000000000000d400000000000000cf00000000000000c800000000",
            INIT_54 => X"000000480000000000000035000000000000009400000000000000d600000000",
            INIT_55 => X"000000220000000000000040000000000000006e000000000000007100000000",
            INIT_56 => X"00000016000000000000004c0000000000000055000000000000001800000000",
            INIT_57 => X"00000016000000000000000d0000000000000009000000000000000700000000",
            INIT_58 => X"0000004e00000000000000250000000000000016000000000000000f00000000",
            INIT_59 => X"0000004800000000000000600000000000000073000000000000005700000000",
            INIT_5A => X"000000720000000000000069000000000000005d000000000000005200000000",
            INIT_5B => X"0000007b000000000000007e000000000000007d000000000000007700000000",
            INIT_5C => X"0000004c00000000000000300000000000000066000000000000007c00000000",
            INIT_5D => X"0000001b0000000000000029000000000000004e000000000000004b00000000",
            INIT_5E => X"0000000600000000000000100000000000000018000000000000000900000000",
            INIT_5F => X"00000019000000000000000f000000000000000a000000000000000800000000",
            INIT_60 => X"0000002b0000000000000023000000000000001f000000000000001500000000",
            INIT_61 => X"0000000c00000000000000190000000000000030000000000000003200000000",
            INIT_62 => X"000000110000000000000011000000000000000e000000000000000e00000000",
            INIT_63 => X"00000019000000000000001a0000000000000018000000000000001400000000",
            INIT_64 => X"0000004a000000000000000d0000000000000014000000000000001800000000",
            INIT_65 => X"000000120000000000000041000000000000003b000000000000004e00000000",
            INIT_66 => X"0000000300000000000000040000000000000005000000000000000300000000",
            INIT_67 => X"0000001a000000000000000d0000000000000009000000000000000500000000",
            INIT_68 => X"00000025000000000000002c0000000000000028000000000000002100000000",
            INIT_69 => X"00000025000000000000001e0000000000000017000000000000001e00000000",
            INIT_6A => X"0000001c000000000000001c0000000000000019000000000000001c00000000",
            INIT_6B => X"0000001300000000000000170000000000000018000000000000001b00000000",
            INIT_6C => X"0000001c00000000000000060000000000000009000000000000000f00000000",
            INIT_6D => X"00000008000000000000002f0000000000000053000000000000004700000000",
            INIT_6E => X"0000000400000000000000050000000000000005000000000000000200000000",
            INIT_6F => X"0000001c0000000000000015000000000000000b000000000000000600000000",
            INIT_70 => X"0000003b00000000000000300000000000000029000000000000002500000000",
            INIT_71 => X"00000059000000000000005c000000000000004f000000000000004900000000",
            INIT_72 => X"0000003b0000000000000038000000000000002f000000000000003800000000",
            INIT_73 => X"00000028000000000000002b0000000000000030000000000000003900000000",
            INIT_74 => X"000000150000000000000015000000000000001b000000000000002300000000",
            INIT_75 => X"0000000800000000000000100000000000000025000000000000002100000000",
            INIT_76 => X"0000000a000000000000000a0000000000000009000000000000000800000000",
            INIT_77 => X"0000001c000000000000001d0000000000000012000000000000000d00000000",
            INIT_78 => X"0000006500000000000000460000000000000031000000000000002c00000000",
            INIT_79 => X"0000006300000000000000760000000000000080000000000000008000000000",
            INIT_7A => X"000000550000000000000054000000000000004e000000000000004700000000",
            INIT_7B => X"0000004f00000000000000510000000000000053000000000000005700000000",
            INIT_7C => X"000000310000000000000031000000000000003c000000000000004700000000",
            INIT_7D => X"0000001300000000000000200000000000000038000000000000003a00000000",
            INIT_7E => X"0000001500000000000000180000000000000018000000000000001300000000",
            INIT_7F => X"0000001c0000000000000022000000000000001f000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "sampleifmap_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004d00000000000000510000000000000052000000000000005300000000",
            INIT_01 => X"0000005c000000000000005b0000000000000055000000000000005100000000",
            INIT_02 => X"0000005c0000000000000065000000000000005f000000000000005c00000000",
            INIT_03 => X"0000004c00000000000000500000000000000052000000000000005700000000",
            INIT_04 => X"0000003e000000000000003f0000000000000041000000000000004400000000",
            INIT_05 => X"0000002f00000000000000340000000000000038000000000000003c00000000",
            INIT_06 => X"0000002200000000000000230000000000000025000000000000002a00000000",
            INIT_07 => X"000000150000000000000019000000000000001d000000000000002400000000",
            INIT_08 => X"0000004d00000000000000530000000000000053000000000000005400000000",
            INIT_09 => X"0000005d000000000000005a0000000000000054000000000000005000000000",
            INIT_0A => X"00000061000000000000005f0000000000000058000000000000005a00000000",
            INIT_0B => X"0000004c000000000000004e0000000000000052000000000000005800000000",
            INIT_0C => X"0000004200000000000000400000000000000044000000000000004700000000",
            INIT_0D => X"0000002e00000000000000340000000000000036000000000000003d00000000",
            INIT_0E => X"0000002300000000000000240000000000000026000000000000002a00000000",
            INIT_0F => X"0000001f000000000000001d000000000000001e000000000000002400000000",
            INIT_10 => X"0000004b00000000000000500000000000000051000000000000005200000000",
            INIT_11 => X"0000004c00000000000000580000000000000054000000000000004b00000000",
            INIT_12 => X"0000006300000000000000570000000000000056000000000000005200000000",
            INIT_13 => X"0000004c000000000000004d0000000000000058000000000000006500000000",
            INIT_14 => X"0000004000000000000000400000000000000044000000000000004900000000",
            INIT_15 => X"0000002d00000000000000340000000000000037000000000000003a00000000",
            INIT_16 => X"0000002c00000000000000290000000000000028000000000000002b00000000",
            INIT_17 => X"0000003500000000000000310000000000000030000000000000003100000000",
            INIT_18 => X"0000004e00000000000000500000000000000051000000000000005300000000",
            INIT_19 => X"0000003200000000000000500000000000000057000000000000004a00000000",
            INIT_1A => X"0000005b00000000000000570000000000000061000000000000005500000000",
            INIT_1B => X"0000005000000000000000580000000000000066000000000000006800000000",
            INIT_1C => X"0000003f000000000000003f0000000000000040000000000000004900000000",
            INIT_1D => X"0000003a00000000000000390000000000000038000000000000003b00000000",
            INIT_1E => X"000000470000000000000044000000000000003f000000000000003d00000000",
            INIT_1F => X"0000004500000000000000450000000000000047000000000000004900000000",
            INIT_20 => X"0000004f000000000000004f000000000000004f000000000000004f00000000",
            INIT_21 => X"00000037000000000000004c0000000000000053000000000000004a00000000",
            INIT_22 => X"0000004b000000000000004b0000000000000054000000000000005300000000",
            INIT_23 => X"00000057000000000000005a0000000000000059000000000000004e00000000",
            INIT_24 => X"0000004600000000000000430000000000000042000000000000005300000000",
            INIT_25 => X"0000005700000000000000540000000000000050000000000000004e00000000",
            INIT_26 => X"0000005900000000000000590000000000000056000000000000005700000000",
            INIT_27 => X"00000049000000000000004f0000000000000054000000000000005800000000",
            INIT_28 => X"0000004d000000000000004b000000000000004a000000000000004c00000000",
            INIT_29 => X"0000004600000000000000460000000000000049000000000000004900000000",
            INIT_2A => X"0000004900000000000000470000000000000045000000000000004600000000",
            INIT_2B => X"00000051000000000000004e000000000000004e000000000000004b00000000",
            INIT_2C => X"0000006200000000000000600000000000000059000000000000005a00000000",
            INIT_2D => X"0000006800000000000000660000000000000068000000000000006400000000",
            INIT_2E => X"0000005e0000000000000061000000000000005f000000000000006300000000",
            INIT_2F => X"0000004200000000000000490000000000000050000000000000005700000000",
            INIT_30 => X"0000004900000000000000470000000000000048000000000000004a00000000",
            INIT_31 => X"00000033000000000000002b000000000000003e000000000000004a00000000",
            INIT_32 => X"0000004700000000000000440000000000000040000000000000004400000000",
            INIT_33 => X"0000005e0000000000000051000000000000004a000000000000004b00000000",
            INIT_34 => X"00000072000000000000006e0000000000000062000000000000006000000000",
            INIT_35 => X"0000006d00000000000000680000000000000064000000000000006600000000",
            INIT_36 => X"000000500000000000000055000000000000005b000000000000006300000000",
            INIT_37 => X"0000004300000000000000460000000000000049000000000000004c00000000",
            INIT_38 => X"0000004800000000000000470000000000000048000000000000004700000000",
            INIT_39 => X"00000029000000000000002a000000000000003a000000000000004700000000",
            INIT_3A => X"0000003f000000000000003a0000000000000036000000000000003900000000",
            INIT_3B => X"0000006000000000000000520000000000000047000000000000004100000000",
            INIT_3C => X"00000067000000000000005d000000000000005e000000000000006900000000",
            INIT_3D => X"00000061000000000000006c000000000000006a000000000000006700000000",
            INIT_3E => X"000000500000000000000054000000000000005b000000000000005d00000000",
            INIT_3F => X"0000004d000000000000004f0000000000000050000000000000005000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000052000000000000004b0000000000000049000000000000004900000000",
            INIT_41 => X"0000002e00000000000000570000000000000067000000000000005800000000",
            INIT_42 => X"0000005200000000000000450000000000000038000000000000003800000000",
            INIT_43 => X"00000057000000000000005a0000000000000057000000000000005100000000",
            INIT_44 => X"0000005b000000000000005e0000000000000063000000000000006200000000",
            INIT_45 => X"00000066000000000000006a0000000000000066000000000000006100000000",
            INIT_46 => X"0000005c00000000000000610000000000000063000000000000005e00000000",
            INIT_47 => X"0000005f000000000000005b0000000000000059000000000000005900000000",
            INIT_48 => X"0000007b000000000000006d000000000000005f000000000000005600000000",
            INIT_49 => X"0000003300000000000000680000000000000099000000000000008800000000",
            INIT_4A => X"000000610000000000000049000000000000003b000000000000003c00000000",
            INIT_4B => X"0000005a0000000000000066000000000000006c000000000000006500000000",
            INIT_4C => X"0000005d00000000000000610000000000000061000000000000005f00000000",
            INIT_4D => X"0000006e00000000000000690000000000000063000000000000005d00000000",
            INIT_4E => X"0000006c000000000000006c0000000000000069000000000000006700000000",
            INIT_4F => X"0000006e000000000000006e000000000000006e000000000000006d00000000",
            INIT_50 => X"0000009d0000000000000096000000000000008b000000000000007f00000000",
            INIT_51 => X"00000032000000000000005700000000000000a200000000000000a000000000",
            INIT_52 => X"0000005800000000000000350000000000000038000000000000004300000000",
            INIT_53 => X"0000005a000000000000006b0000000000000070000000000000006500000000",
            INIT_54 => X"00000060000000000000005e0000000000000060000000000000005e00000000",
            INIT_55 => X"000000650000000000000060000000000000005f000000000000006000000000",
            INIT_56 => X"0000007e000000000000007d0000000000000071000000000000006800000000",
            INIT_57 => X"0000007000000000000000740000000000000077000000000000007b00000000",
            INIT_58 => X"000000a2000000000000009f000000000000009d000000000000009800000000",
            INIT_59 => X"0000002c000000000000005a000000000000009f00000000000000a000000000",
            INIT_5A => X"00000056000000000000003a0000000000000045000000000000004800000000",
            INIT_5B => X"0000005c0000000000000061000000000000005a000000000000006700000000",
            INIT_5C => X"0000005e000000000000005f0000000000000060000000000000005a00000000",
            INIT_5D => X"0000005c00000000000000570000000000000062000000000000006300000000",
            INIT_5E => X"0000008300000000000000830000000000000070000000000000006100000000",
            INIT_5F => X"0000006c00000000000000740000000000000079000000000000007f00000000",
            INIT_60 => X"0000009d00000000000000a0000000000000009e000000000000009b00000000",
            INIT_61 => X"0000003000000000000000720000000000000094000000000000009800000000",
            INIT_62 => X"00000067000000000000005e0000000000000058000000000000004400000000",
            INIT_63 => X"0000005d00000000000000580000000000000060000000000000007300000000",
            INIT_64 => X"0000005e00000000000000620000000000000065000000000000005900000000",
            INIT_65 => X"0000005500000000000000540000000000000065000000000000006300000000",
            INIT_66 => X"00000084000000000000007d000000000000006e000000000000006900000000",
            INIT_67 => X"0000005f000000000000006b0000000000000076000000000000007f00000000",
            INIT_68 => X"0000009200000000000000950000000000000094000000000000009400000000",
            INIT_69 => X"000000500000000000000088000000000000008e000000000000009000000000",
            INIT_6A => X"00000068000000000000005e0000000000000048000000000000002f00000000",
            INIT_6B => X"0000005e000000000000005c0000000000000071000000000000007200000000",
            INIT_6C => X"0000005d00000000000000610000000000000067000000000000005d00000000",
            INIT_6D => X"0000005200000000000000550000000000000061000000000000006000000000",
            INIT_6E => X"00000079000000000000006f000000000000006b000000000000006b00000000",
            INIT_6F => X"0000004d00000000000000570000000000000064000000000000007000000000",
            INIT_70 => X"0000008c000000000000008a0000000000000087000000000000008600000000",
            INIT_71 => X"0000008900000000000000970000000000000093000000000000008e00000000",
            INIT_72 => X"0000003e00000000000000320000000000000049000000000000005d00000000",
            INIT_73 => X"00000062000000000000005a000000000000005e000000000000005900000000",
            INIT_74 => X"0000006100000000000000670000000000000069000000000000006600000000",
            INIT_75 => X"000000530000000000000056000000000000005e000000000000005e00000000",
            INIT_76 => X"00000066000000000000005c0000000000000065000000000000005f00000000",
            INIT_77 => X"0000004b000000000000004a0000000000000052000000000000005f00000000",
            INIT_78 => X"00000090000000000000008b0000000000000086000000000000008300000000",
            INIT_79 => X"00000098000000000000009a000000000000009f000000000000009800000000",
            INIT_7A => X"0000003900000000000000350000000000000076000000000000009e00000000",
            INIT_7B => X"00000066000000000000005f0000000000000064000000000000006700000000",
            INIT_7C => X"0000006a000000000000006f0000000000000074000000000000006e00000000",
            INIT_7D => X"000000550000000000000057000000000000005b000000000000006100000000",
            INIT_7E => X"0000005300000000000000550000000000000062000000000000005400000000",
            INIT_7F => X"0000005f000000000000005a0000000000000055000000000000005300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "sampleifmap_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a000000000000000980000000000000090000000000000008700000000",
            INIT_01 => X"00000073000000000000008900000000000000a100000000000000a400000000",
            INIT_02 => X"0000006e00000000000000800000000000000091000000000000009d00000000",
            INIT_03 => X"000000670000000000000068000000000000007a000000000000007b00000000",
            INIT_04 => X"00000068000000000000006c000000000000006d000000000000006900000000",
            INIT_05 => X"000000570000000000000058000000000000005a000000000000006100000000",
            INIT_06 => X"000000550000000000000057000000000000005c000000000000004f00000000",
            INIT_07 => X"0000005e00000000000000690000000000000069000000000000006500000000",
            INIT_08 => X"000000a4000000000000009f000000000000009a000000000000009400000000",
            INIT_09 => X"0000007f00000000000000b000000000000000b300000000000000aa00000000",
            INIT_0A => X"00000098000000000000009d00000000000000c500000000000000b000000000",
            INIT_0B => X"0000006700000000000000800000000000000091000000000000007100000000",
            INIT_0C => X"0000006600000000000000680000000000000065000000000000006700000000",
            INIT_0D => X"00000059000000000000005b000000000000005f000000000000006100000000",
            INIT_0E => X"0000005b000000000000005b0000000000000056000000000000004f00000000",
            INIT_0F => X"0000004600000000000000560000000000000068000000000000006d00000000",
            INIT_10 => X"000000c500000000000000b200000000000000a4000000000000009b00000000",
            INIT_11 => X"000000c400000000000000f800000000000000ee00000000000000dd00000000",
            INIT_12 => X"000000b800000000000000b000000000000000c8000000000000009c00000000",
            INIT_13 => X"0000006a0000000000000089000000000000008e000000000000006c00000000",
            INIT_14 => X"0000006500000000000000640000000000000063000000000000006400000000",
            INIT_15 => X"00000059000000000000005f0000000000000063000000000000006500000000",
            INIT_16 => X"00000053000000000000005c0000000000000051000000000000005000000000",
            INIT_17 => X"0000004700000000000000490000000000000052000000000000005800000000",
            INIT_18 => X"000000f900000000000000eb00000000000000d600000000000000bf00000000",
            INIT_19 => X"000000f400000000000000fb00000000000000f600000000000000fd00000000",
            INIT_1A => X"000000c300000000000000ac000000000000009e00000000000000a000000000",
            INIT_1B => X"0000006e000000000000008b0000000000000072000000000000007100000000",
            INIT_1C => X"0000006300000000000000610000000000000062000000000000006200000000",
            INIT_1D => X"0000005c00000000000000660000000000000068000000000000006700000000",
            INIT_1E => X"000000490000000000000055000000000000004e000000000000005300000000",
            INIT_1F => X"00000048000000000000004a0000000000000050000000000000004b00000000",
            INIT_20 => X"000000fe00000000000000fd00000000000000fc00000000000000f500000000",
            INIT_21 => X"000000c900000000000000ba00000000000000bb00000000000000f300000000",
            INIT_22 => X"0000009c00000000000000970000000000000080000000000000009100000000",
            INIT_23 => X"000000720000000000000080000000000000006a000000000000007400000000",
            INIT_24 => X"0000006700000000000000650000000000000067000000000000006800000000",
            INIT_25 => X"0000005c0000000000000069000000000000006e000000000000006c00000000",
            INIT_26 => X"000000550000000000000054000000000000004c000000000000005200000000",
            INIT_27 => X"00000049000000000000004d0000000000000053000000000000004e00000000",
            INIT_28 => X"0000010000000000000000fc00000000000000fc00000000000000fb00000000",
            INIT_29 => X"00000072000000000000006b000000000000007e00000000000000e900000000",
            INIT_2A => X"0000006e00000000000000780000000000000073000000000000006900000000",
            INIT_2B => X"0000006700000000000000680000000000000063000000000000006300000000",
            INIT_2C => X"0000006b000000000000006b000000000000006e000000000000006d00000000",
            INIT_2D => X"000000560000000000000060000000000000006e000000000000007000000000",
            INIT_2E => X"00000068000000000000005a000000000000004c000000000000004e00000000",
            INIT_2F => X"0000004f00000000000000520000000000000052000000000000005b00000000",
            INIT_30 => X"000000eb00000000000000f600000000000000f800000000000000f800000000",
            INIT_31 => X"000000760000000000000072000000000000007c00000000000000c800000000",
            INIT_32 => X"0000004f00000000000000530000000000000057000000000000005d00000000",
            INIT_33 => X"00000044000000000000004b0000000000000056000000000000005000000000",
            INIT_34 => X"0000006100000000000000620000000000000064000000000000005f00000000",
            INIT_35 => X"0000006100000000000000610000000000000061000000000000006200000000",
            INIT_36 => X"0000006f000000000000005b0000000000000057000000000000005b00000000",
            INIT_37 => X"0000005200000000000000520000000000000055000000000000006e00000000",
            INIT_38 => X"0000009600000000000000b500000000000000d600000000000000eb00000000",
            INIT_39 => X"0000008400000000000000850000000000000088000000000000008a00000000",
            INIT_3A => X"0000003c0000000000000039000000000000003d000000000000006400000000",
            INIT_3B => X"0000003a00000000000000600000000000000059000000000000004300000000",
            INIT_3C => X"0000005000000000000000470000000000000045000000000000003300000000",
            INIT_3D => X"0000006500000000000000680000000000000065000000000000005e00000000",
            INIT_3E => X"0000006d000000000000005e0000000000000057000000000000005d00000000",
            INIT_3F => X"0000005100000000000000510000000000000062000000000000007700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009900000000",
            INIT_41 => X"00000067000000000000006f000000000000007a000000000000007c00000000",
            INIT_42 => X"000000340000000000000039000000000000005a000000000000006a00000000",
            INIT_43 => X"00000053000000000000006a0000000000000066000000000000004500000000",
            INIT_44 => X"00000055000000000000004d0000000000000047000000000000004000000000",
            INIT_45 => X"0000006d00000000000000660000000000000067000000000000006400000000",
            INIT_46 => X"00000063000000000000005d0000000000000057000000000000006a00000000",
            INIT_47 => X"00000050000000000000005c0000000000000073000000000000007100000000",
            INIT_48 => X"0000006d0000000000000072000000000000006f000000000000006d00000000",
            INIT_49 => X"0000006d00000000000000660000000000000061000000000000006500000000",
            INIT_4A => X"0000005500000000000000670000000000000078000000000000007500000000",
            INIT_4B => X"00000059000000000000005f0000000000000065000000000000005d00000000",
            INIT_4C => X"0000005a0000000000000052000000000000004b000000000000004a00000000",
            INIT_4D => X"0000006600000000000000690000000000000077000000000000007200000000",
            INIT_4E => X"00000062000000000000005e000000000000006b000000000000006f00000000",
            INIT_4F => X"0000004f000000000000006b0000000000000075000000000000006500000000",
            INIT_50 => X"0000005b000000000000005d0000000000000062000000000000006900000000",
            INIT_51 => X"00000071000000000000006f000000000000006a000000000000006300000000",
            INIT_52 => X"0000005f00000000000000610000000000000068000000000000007000000000",
            INIT_53 => X"0000005c0000000000000054000000000000004c000000000000005000000000",
            INIT_54 => X"00000059000000000000004f0000000000000048000000000000005100000000",
            INIT_55 => X"0000005e0000000000000069000000000000007b000000000000007500000000",
            INIT_56 => X"0000006500000000000000670000000000000067000000000000006000000000",
            INIT_57 => X"0000005a000000000000006f0000000000000069000000000000006000000000",
            INIT_58 => X"00000065000000000000005e0000000000000057000000000000005700000000",
            INIT_59 => X"00000064000000000000006b000000000000006e000000000000006c00000000",
            INIT_5A => X"0000006800000000000000560000000000000051000000000000005b00000000",
            INIT_5B => X"0000005c000000000000004c0000000000000049000000000000005d00000000",
            INIT_5C => X"0000004f000000000000004f000000000000004d000000000000005800000000",
            INIT_5D => X"00000056000000000000005d0000000000000064000000000000005b00000000",
            INIT_5E => X"000000600000000000000061000000000000005c000000000000005700000000",
            INIT_5F => X"0000006500000000000000660000000000000060000000000000006000000000",
            INIT_60 => X"0000006900000000000000670000000000000060000000000000005a00000000",
            INIT_61 => X"000000500000000000000056000000000000005f000000000000006500000000",
            INIT_62 => X"0000006a00000000000000600000000000000055000000000000005100000000",
            INIT_63 => X"0000005d00000000000000600000000000000055000000000000006200000000",
            INIT_64 => X"0000004c000000000000004f0000000000000051000000000000005800000000",
            INIT_65 => X"0000005b0000000000000054000000000000004c000000000000004700000000",
            INIT_66 => X"0000005a00000000000000530000000000000056000000000000005c00000000",
            INIT_67 => X"00000060000000000000005b0000000000000060000000000000006200000000",
            INIT_68 => X"00000056000000000000005f0000000000000063000000000000006400000000",
            INIT_69 => X"0000004f000000000000004f000000000000004f000000000000005000000000",
            INIT_6A => X"0000006c00000000000000620000000000000053000000000000005200000000",
            INIT_6B => X"0000005900000000000000610000000000000060000000000000006300000000",
            INIT_6C => X"00000051000000000000004f0000000000000054000000000000005c00000000",
            INIT_6D => X"000000590000000000000052000000000000004a000000000000004c00000000",
            INIT_6E => X"0000005600000000000000520000000000000055000000000000005a00000000",
            INIT_6F => X"000000530000000000000053000000000000005c000000000000005d00000000",
            INIT_70 => X"000000470000000000000049000000000000004e000000000000005700000000",
            INIT_71 => X"0000005300000000000000590000000000000057000000000000004d00000000",
            INIT_72 => X"0000006a0000000000000061000000000000004f000000000000005100000000",
            INIT_73 => X"0000005c00000000000000590000000000000067000000000000006400000000",
            INIT_74 => X"0000005900000000000000580000000000000057000000000000006000000000",
            INIT_75 => X"000000530000000000000054000000000000004f000000000000005200000000",
            INIT_76 => X"000000530000000000000056000000000000005a000000000000005600000000",
            INIT_77 => X"00000049000000000000004f0000000000000056000000000000005600000000",
            INIT_78 => X"000000490000000000000046000000000000003f000000000000003e00000000",
            INIT_79 => X"0000005100000000000000530000000000000056000000000000005400000000",
            INIT_7A => X"0000006b000000000000005e000000000000004a000000000000004e00000000",
            INIT_7B => X"00000058000000000000005b0000000000000068000000000000005f00000000",
            INIT_7C => X"0000005900000000000000580000000000000058000000000000005b00000000",
            INIT_7D => X"0000005300000000000000550000000000000050000000000000005500000000",
            INIT_7E => X"0000005000000000000000560000000000000059000000000000005400000000",
            INIT_7F => X"00000048000000000000004c000000000000004d000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "sampleifmap_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000005d000000000000005e000000000000005e00000000",
            INIT_01 => X"000000600000000000000060000000000000005a000000000000005a00000000",
            INIT_02 => X"00000065000000000000006e0000000000000066000000000000006100000000",
            INIT_03 => X"0000005200000000000000550000000000000058000000000000005e00000000",
            INIT_04 => X"000000480000000000000049000000000000004b000000000000004e00000000",
            INIT_05 => X"00000038000000000000003d0000000000000041000000000000004500000000",
            INIT_06 => X"000000270000000000000029000000000000002e000000000000003300000000",
            INIT_07 => X"00000019000000000000001d0000000000000022000000000000002800000000",
            INIT_08 => X"00000059000000000000005f000000000000005f000000000000006000000000",
            INIT_09 => X"00000062000000000000005f0000000000000059000000000000005900000000",
            INIT_0A => X"0000006b000000000000006a0000000000000060000000000000006100000000",
            INIT_0B => X"0000005200000000000000550000000000000059000000000000006000000000",
            INIT_0C => X"000000490000000000000047000000000000004b000000000000004f00000000",
            INIT_0D => X"00000035000000000000003b000000000000003d000000000000004400000000",
            INIT_0E => X"000000250000000000000027000000000000002c000000000000003100000000",
            INIT_0F => X"0000001f000000000000001f0000000000000020000000000000002600000000",
            INIT_10 => X"00000057000000000000005c000000000000005c000000000000005e00000000",
            INIT_11 => X"00000051000000000000005d000000000000005a000000000000005400000000",
            INIT_12 => X"0000006e00000000000000630000000000000060000000000000005900000000",
            INIT_13 => X"0000005400000000000000560000000000000062000000000000007000000000",
            INIT_14 => X"0000004600000000000000440000000000000049000000000000004f00000000",
            INIT_15 => X"000000300000000000000036000000000000003a000000000000003f00000000",
            INIT_16 => X"0000002b0000000000000029000000000000002b000000000000002e00000000",
            INIT_17 => X"000000310000000000000030000000000000002e000000000000002f00000000",
            INIT_18 => X"0000005a000000000000005c000000000000005d000000000000005f00000000",
            INIT_19 => X"000000390000000000000056000000000000005d000000000000005300000000",
            INIT_1A => X"000000680000000000000063000000000000006b000000000000005d00000000",
            INIT_1B => X"0000005a00000000000000650000000000000072000000000000007400000000",
            INIT_1C => X"0000004200000000000000420000000000000043000000000000004e00000000",
            INIT_1D => X"0000003900000000000000380000000000000038000000000000003e00000000",
            INIT_1E => X"000000420000000000000041000000000000003e000000000000003c00000000",
            INIT_1F => X"0000003d000000000000003f0000000000000041000000000000004300000000",
            INIT_20 => X"0000005b000000000000005b000000000000005b000000000000005c00000000",
            INIT_21 => X"0000003e00000000000000520000000000000059000000000000005300000000",
            INIT_22 => X"000000580000000000000058000000000000005f000000000000005c00000000",
            INIT_23 => X"0000006400000000000000690000000000000068000000000000005c00000000",
            INIT_24 => X"0000004800000000000000450000000000000046000000000000005b00000000",
            INIT_25 => X"000000530000000000000050000000000000004d000000000000005000000000",
            INIT_26 => X"0000005000000000000000510000000000000051000000000000005300000000",
            INIT_27 => X"0000003f0000000000000046000000000000004b000000000000004f00000000",
            INIT_28 => X"0000005900000000000000570000000000000056000000000000005800000000",
            INIT_29 => X"0000004d000000000000004c000000000000004f000000000000005200000000",
            INIT_2A => X"0000005700000000000000550000000000000052000000000000005000000000",
            INIT_2B => X"0000005f000000000000005e000000000000005e000000000000005a00000000",
            INIT_2C => X"000000630000000000000062000000000000005e000000000000006300000000",
            INIT_2D => X"0000006200000000000000600000000000000064000000000000006400000000",
            INIT_2E => X"0000005300000000000000580000000000000058000000000000005d00000000",
            INIT_2F => X"00000037000000000000003e0000000000000045000000000000004c00000000",
            INIT_30 => X"0000005400000000000000520000000000000054000000000000005500000000",
            INIT_31 => X"00000037000000000000002a000000000000003d000000000000005100000000",
            INIT_32 => X"0000005900000000000000580000000000000057000000000000005300000000",
            INIT_33 => X"00000065000000000000005d0000000000000057000000000000005b00000000",
            INIT_34 => X"0000007300000000000000700000000000000064000000000000006200000000",
            INIT_35 => X"0000006700000000000000670000000000000067000000000000006900000000",
            INIT_36 => X"0000004a000000000000004e0000000000000050000000000000005b00000000",
            INIT_37 => X"000000360000000000000039000000000000003f000000000000004400000000",
            INIT_38 => X"0000005400000000000000520000000000000053000000000000005200000000",
            INIT_39 => X"0000002c00000000000000260000000000000037000000000000004c00000000",
            INIT_3A => X"0000005100000000000000520000000000000055000000000000004c00000000",
            INIT_3B => X"00000063000000000000005b0000000000000053000000000000005000000000",
            INIT_3C => X"0000006c00000000000000610000000000000060000000000000006700000000",
            INIT_3D => X"0000005e00000000000000710000000000000072000000000000006d00000000",
            INIT_3E => X"0000004b000000000000004d000000000000004d000000000000005200000000",
            INIT_3F => X"0000003b00000000000000400000000000000044000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005b00000000000000540000000000000052000000000000005100000000",
            INIT_41 => X"0000003100000000000000550000000000000068000000000000005e00000000",
            INIT_42 => X"00000063000000000000005b0000000000000054000000000000004900000000",
            INIT_43 => X"0000005e00000000000000650000000000000064000000000000006100000000",
            INIT_44 => X"0000006200000000000000650000000000000068000000000000006500000000",
            INIT_45 => X"000000670000000000000072000000000000006f000000000000006a00000000",
            INIT_46 => X"0000004e00000000000000520000000000000055000000000000005700000000",
            INIT_47 => X"0000004800000000000000470000000000000046000000000000004a00000000",
            INIT_48 => X"0000008000000000000000730000000000000065000000000000005c00000000",
            INIT_49 => X"000000360000000000000068000000000000009d000000000000008e00000000",
            INIT_4A => X"00000071000000000000005d0000000000000054000000000000004b00000000",
            INIT_4B => X"000000650000000000000075000000000000007c000000000000007500000000",
            INIT_4C => X"00000067000000000000006b000000000000006a000000000000006700000000",
            INIT_4D => X"000000760000000000000074000000000000006e000000000000006800000000",
            INIT_4E => X"000000540000000000000055000000000000005a000000000000006400000000",
            INIT_4F => X"0000005200000000000000550000000000000055000000000000005500000000",
            INIT_50 => X"000000a00000000000000099000000000000008e000000000000008200000000",
            INIT_51 => X"00000035000000000000005900000000000000aa00000000000000a600000000",
            INIT_52 => X"000000680000000000000046000000000000004d000000000000005000000000",
            INIT_53 => X"0000006b000000000000007f0000000000000082000000000000007700000000",
            INIT_54 => X"0000006a0000000000000069000000000000006c000000000000006a00000000",
            INIT_55 => X"00000072000000000000006e0000000000000069000000000000006a00000000",
            INIT_56 => X"0000006000000000000000620000000000000062000000000000006900000000",
            INIT_57 => X"000000550000000000000059000000000000005b000000000000005e00000000",
            INIT_58 => X"000000a400000000000000a2000000000000009f000000000000009a00000000",
            INIT_59 => X"0000002e000000000000005d00000000000000a900000000000000a700000000",
            INIT_5A => X"00000067000000000000004a0000000000000056000000000000005100000000",
            INIT_5B => X"00000072000000000000007a0000000000000070000000000000007b00000000",
            INIT_5C => X"00000067000000000000006a000000000000006d000000000000006a00000000",
            INIT_5D => X"0000006e00000000000000670000000000000069000000000000006b00000000",
            INIT_5E => X"0000006300000000000000650000000000000061000000000000006600000000",
            INIT_5F => X"00000055000000000000005a000000000000005e000000000000006000000000",
            INIT_60 => X"0000009e00000000000000a1000000000000009f000000000000009d00000000",
            INIT_61 => X"000000300000000000000075000000000000009f000000000000009e00000000",
            INIT_62 => X"00000078000000000000006c0000000000000065000000000000004900000000",
            INIT_63 => X"0000007500000000000000740000000000000078000000000000008700000000",
            INIT_64 => X"00000066000000000000006c0000000000000073000000000000006b00000000",
            INIT_65 => X"000000690000000000000064000000000000006a000000000000006900000000",
            INIT_66 => X"0000006500000000000000600000000000000060000000000000007000000000",
            INIT_67 => X"0000004c0000000000000055000000000000005d000000000000006200000000",
            INIT_68 => X"0000009300000000000000970000000000000098000000000000009900000000",
            INIT_69 => X"0000004c00000000000000870000000000000093000000000000009300000000",
            INIT_6A => X"0000007500000000000000670000000000000049000000000000002c00000000",
            INIT_6B => X"0000007100000000000000730000000000000085000000000000008300000000",
            INIT_6C => X"0000006b00000000000000710000000000000077000000000000006c00000000",
            INIT_6D => X"000000640000000000000065000000000000006a000000000000006a00000000",
            INIT_6E => X"00000062000000000000005d0000000000000069000000000000007500000000",
            INIT_6F => X"00000040000000000000004a0000000000000055000000000000005d00000000",
            INIT_70 => X"0000008e000000000000008e000000000000008e000000000000008f00000000",
            INIT_71 => X"0000008300000000000000950000000000000094000000000000008f00000000",
            INIT_72 => X"0000004600000000000000350000000000000041000000000000005400000000",
            INIT_73 => X"0000006d0000000000000068000000000000006b000000000000006300000000",
            INIT_74 => X"00000075000000000000007d000000000000007c000000000000007200000000",
            INIT_75 => X"000000620000000000000065000000000000006c000000000000006e00000000",
            INIT_76 => X"0000005a0000000000000058000000000000006f000000000000006c00000000",
            INIT_77 => X"0000003f00000000000000410000000000000048000000000000005500000000",
            INIT_78 => X"00000091000000000000008e000000000000008d000000000000008c00000000",
            INIT_79 => X"00000093000000000000009900000000000000a0000000000000009900000000",
            INIT_7A => X"0000003a0000000000000034000000000000006f000000000000009700000000",
            INIT_7B => X"0000006e00000000000000650000000000000068000000000000006a00000000",
            INIT_7C => X"0000008000000000000000870000000000000089000000000000007b00000000",
            INIT_7D => X"000000650000000000000068000000000000006c000000000000007300000000",
            INIT_7E => X"0000004e0000000000000059000000000000006f000000000000006300000000",
            INIT_7F => X"0000004d000000000000004a0000000000000048000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "sampleifmap_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000000000009b0000000000000095000000000000008f00000000",
            INIT_01 => X"00000072000000000000008800000000000000a000000000000000a400000000",
            INIT_02 => X"00000068000000000000007a000000000000008f000000000000009b00000000",
            INIT_03 => X"0000006c00000000000000660000000000000077000000000000007600000000",
            INIT_04 => X"0000008000000000000000850000000000000084000000000000007800000000",
            INIT_05 => X"0000006a000000000000006b000000000000006d000000000000007500000000",
            INIT_06 => X"000000560000000000000062000000000000006c000000000000006100000000",
            INIT_07 => X"00000044000000000000004f0000000000000054000000000000005a00000000",
            INIT_08 => X"000000a1000000000000009f000000000000009d000000000000009a00000000",
            INIT_09 => X"0000008100000000000000b000000000000000b100000000000000a700000000",
            INIT_0A => X"0000008e000000000000009700000000000000c700000000000000b300000000",
            INIT_0B => X"0000006c000000000000007b0000000000000089000000000000006800000000",
            INIT_0C => X"000000800000000000000083000000000000007e000000000000007900000000",
            INIT_0D => X"0000006e00000000000000700000000000000073000000000000007700000000",
            INIT_0E => X"0000005e000000000000006a0000000000000069000000000000006300000000",
            INIT_0F => X"000000270000000000000034000000000000004a000000000000005c00000000",
            INIT_10 => X"000000c100000000000000b000000000000000a4000000000000009d00000000",
            INIT_11 => X"000000c700000000000000f700000000000000ec00000000000000da00000000",
            INIT_12 => X"000000b100000000000000ad00000000000000ce00000000000000a300000000",
            INIT_13 => X"0000007100000000000000860000000000000088000000000000006500000000",
            INIT_14 => X"000000810000000000000082000000000000007e000000000000007700000000",
            INIT_15 => X"000000710000000000000076000000000000007a000000000000007d00000000",
            INIT_16 => X"00000050000000000000006a0000000000000067000000000000006800000000",
            INIT_17 => X"000000270000000000000025000000000000002c000000000000003e00000000",
            INIT_18 => X"000000f600000000000000e800000000000000d400000000000000c000000000",
            INIT_19 => X"000000f700000000000000fa00000000000000f200000000000000fa00000000",
            INIT_1A => X"000000c100000000000000ae00000000000000aa00000000000000a900000000",
            INIT_1B => X"00000078000000000000008b0000000000000070000000000000006e00000000",
            INIT_1C => X"000000800000000000000080000000000000007e000000000000007600000000",
            INIT_1D => X"00000074000000000000007e000000000000007f000000000000008000000000",
            INIT_1E => X"0000003e00000000000000600000000000000066000000000000006c00000000",
            INIT_1F => X"0000002b00000000000000270000000000000025000000000000002a00000000",
            INIT_20 => X"000000fb00000000000000fa00000000000000fb00000000000000f500000000",
            INIT_21 => X"000000d200000000000000be00000000000000ba00000000000000f100000000",
            INIT_22 => X"000000a0000000000000009c000000000000009200000000000000a100000000",
            INIT_23 => X"0000007a00000000000000870000000000000073000000000000007d00000000",
            INIT_24 => X"000000800000000000000081000000000000007f000000000000007800000000",
            INIT_25 => X"00000074000000000000007d000000000000007f000000000000007f00000000",
            INIT_26 => X"0000004200000000000000570000000000000062000000000000006a00000000",
            INIT_27 => X"000000290000000000000029000000000000002a000000000000002d00000000",
            INIT_28 => X"000000fe00000000000000fb00000000000000fb00000000000000fb00000000",
            INIT_29 => X"000000820000000000000074000000000000008300000000000000ea00000000",
            INIT_2A => X"0000007c0000000000000082000000000000008a000000000000007f00000000",
            INIT_2B => X"0000006b00000000000000720000000000000077000000000000007a00000000",
            INIT_2C => X"0000007f00000000000000820000000000000080000000000000007600000000",
            INIT_2D => X"0000006c000000000000006f0000000000000077000000000000007d00000000",
            INIT_2E => X"000000500000000000000052000000000000005a000000000000006300000000",
            INIT_2F => X"00000029000000000000002c000000000000002f000000000000003d00000000",
            INIT_30 => X"000000ef00000000000000f900000000000000fc00000000000000fc00000000",
            INIT_31 => X"00000083000000000000007b000000000000008000000000000000cb00000000",
            INIT_32 => X"000000670000000000000066000000000000006c000000000000006f00000000",
            INIT_33 => X"0000004400000000000000510000000000000069000000000000006a00000000",
            INIT_34 => X"0000007400000000000000780000000000000075000000000000006600000000",
            INIT_35 => X"000000730000000000000070000000000000006b000000000000006e00000000",
            INIT_36 => X"00000054000000000000004b0000000000000059000000000000006800000000",
            INIT_37 => X"0000002d000000000000002d0000000000000034000000000000005100000000",
            INIT_38 => X"000000a000000000000000bf00000000000000df00000000000000f500000000",
            INIT_39 => X"0000008a00000000000000890000000000000089000000000000009000000000",
            INIT_3A => X"000000570000000000000051000000000000004b000000000000006d00000000",
            INIT_3B => X"0000003a00000000000000630000000000000066000000000000005a00000000",
            INIT_3C => X"00000065000000000000005f0000000000000056000000000000003a00000000",
            INIT_3D => X"00000074000000000000007a0000000000000074000000000000006d00000000",
            INIT_3E => X"000000500000000000000046000000000000004d000000000000006100000000",
            INIT_3F => X"0000002f000000000000002f0000000000000042000000000000005900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000840000000000000086000000000000008d00000000000000a500000000",
            INIT_41 => X"000000690000000000000070000000000000007b000000000000008200000000",
            INIT_42 => X"00000047000000000000004a000000000000005e000000000000006b00000000",
            INIT_43 => X"00000056000000000000006f000000000000006e000000000000005300000000",
            INIT_44 => X"0000006c0000000000000066000000000000005a000000000000004800000000",
            INIT_45 => X"0000007c000000000000007b000000000000007b000000000000007600000000",
            INIT_46 => X"0000004400000000000000420000000000000049000000000000006c00000000",
            INIT_47 => X"00000030000000000000003d0000000000000054000000000000005200000000",
            INIT_48 => X"00000075000000000000007a0000000000000078000000000000007500000000",
            INIT_49 => X"0000006a00000000000000650000000000000061000000000000006a00000000",
            INIT_4A => X"00000057000000000000006a0000000000000073000000000000007000000000",
            INIT_4B => X"0000006100000000000000680000000000000068000000000000005c00000000",
            INIT_4C => X"00000072000000000000006c000000000000005f000000000000005400000000",
            INIT_4D => X"0000007a0000000000000082000000000000008e000000000000008600000000",
            INIT_4E => X"0000004000000000000000450000000000000064000000000000007700000000",
            INIT_4F => X"00000032000000000000004f0000000000000057000000000000004500000000",
            INIT_50 => X"0000005e00000000000000600000000000000066000000000000006c00000000",
            INIT_51 => X"0000006b000000000000006e000000000000006b000000000000006500000000",
            INIT_52 => X"000000510000000000000056000000000000005d000000000000006700000000",
            INIT_53 => X"00000068000000000000005d0000000000000048000000000000004200000000",
            INIT_54 => X"00000071000000000000006b000000000000005f000000000000005e00000000",
            INIT_55 => X"0000007a00000000000000850000000000000094000000000000008900000000",
            INIT_56 => X"000000420000000000000051000000000000006b000000000000007200000000",
            INIT_57 => X"0000003f0000000000000055000000000000004b000000000000004000000000",
            INIT_58 => X"00000063000000000000005d0000000000000057000000000000005800000000",
            INIT_59 => X"000000570000000000000065000000000000006c000000000000006b00000000",
            INIT_5A => X"000000530000000000000041000000000000003c000000000000004900000000",
            INIT_5B => X"0000005e000000000000004e000000000000003f000000000000004a00000000",
            INIT_5C => X"0000005d000000000000005f0000000000000057000000000000005900000000",
            INIT_5D => X"00000072000000000000007a000000000000007b000000000000006900000000",
            INIT_5E => X"0000003b000000000000004e0000000000000068000000000000006d00000000",
            INIT_5F => X"0000004b000000000000004a000000000000003f000000000000003c00000000",
            INIT_60 => X"0000005f0000000000000061000000000000005f000000000000005d00000000",
            INIT_61 => X"0000003800000000000000450000000000000054000000000000005b00000000",
            INIT_62 => X"0000005500000000000000420000000000000031000000000000003200000000",
            INIT_63 => X"0000004800000000000000550000000000000049000000000000005300000000",
            INIT_64 => X"000000440000000000000043000000000000003e000000000000003e00000000",
            INIT_65 => X"0000006800000000000000640000000000000058000000000000004500000000",
            INIT_66 => X"000000330000000000000040000000000000005a000000000000006500000000",
            INIT_67 => X"00000045000000000000003a0000000000000036000000000000003500000000",
            INIT_68 => X"000000440000000000000051000000000000005b000000000000006000000000",
            INIT_69 => X"0000003000000000000000340000000000000037000000000000003b00000000",
            INIT_6A => X"000000520000000000000040000000000000002e000000000000002f00000000",
            INIT_6B => X"00000039000000000000004d000000000000004f000000000000005200000000",
            INIT_6C => X"0000003a00000000000000340000000000000032000000000000003500000000",
            INIT_6D => X"0000004a0000000000000047000000000000003f000000000000003a00000000",
            INIT_6E => X"0000002e00000000000000340000000000000041000000000000004800000000",
            INIT_6F => X"0000003600000000000000300000000000000031000000000000003000000000",
            INIT_70 => X"0000002b0000000000000031000000000000003c000000000000004900000000",
            INIT_71 => X"0000003000000000000000340000000000000030000000000000002c00000000",
            INIT_72 => X"00000049000000000000003a000000000000002c000000000000003000000000",
            INIT_73 => X"00000035000000000000003e000000000000004f000000000000004b00000000",
            INIT_74 => X"000000390000000000000034000000000000002e000000000000003200000000",
            INIT_75 => X"0000002f0000000000000033000000000000002f000000000000003400000000",
            INIT_76 => X"0000002a000000000000002e0000000000000031000000000000002f00000000",
            INIT_77 => X"0000002a000000000000002b000000000000002d000000000000002b00000000",
            INIT_78 => X"0000002500000000000000270000000000000025000000000000002900000000",
            INIT_79 => X"0000002d00000000000000290000000000000029000000000000002a00000000",
            INIT_7A => X"000000470000000000000036000000000000002b000000000000002f00000000",
            INIT_7B => X"0000002e000000000000003b000000000000004c000000000000004300000000",
            INIT_7C => X"00000030000000000000002d000000000000002a000000000000002b00000000",
            INIT_7D => X"0000002d0000000000000031000000000000002d000000000000002f00000000",
            INIT_7E => X"00000027000000000000002a000000000000002d000000000000002b00000000",
            INIT_7F => X"0000002600000000000000280000000000000028000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "sampleifmap_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f00000000000000530000000000000054000000000000005500000000",
            INIT_01 => X"0000005f000000000000005d0000000000000052000000000000005000000000",
            INIT_02 => X"00000048000000000000004f0000000000000055000000000000005a00000000",
            INIT_03 => X"0000004f0000000000000054000000000000004e000000000000004b00000000",
            INIT_04 => X"0000003d000000000000003c000000000000003e000000000000004400000000",
            INIT_05 => X"000000330000000000000038000000000000003b000000000000003c00000000",
            INIT_06 => X"0000002300000000000000250000000000000029000000000000002e00000000",
            INIT_07 => X"000000150000000000000019000000000000001e000000000000002400000000",
            INIT_08 => X"0000004f00000000000000550000000000000055000000000000005600000000",
            INIT_09 => X"0000005d000000000000005a0000000000000050000000000000004e00000000",
            INIT_0A => X"0000004700000000000000460000000000000049000000000000005400000000",
            INIT_0B => X"0000004800000000000000470000000000000045000000000000004400000000",
            INIT_0C => X"0000003e000000000000003e0000000000000043000000000000004600000000",
            INIT_0D => X"0000002e00000000000000340000000000000035000000000000003800000000",
            INIT_0E => X"0000002000000000000000220000000000000025000000000000002900000000",
            INIT_0F => X"0000001b000000000000001a000000000000001b000000000000002100000000",
            INIT_10 => X"0000004e00000000000000520000000000000053000000000000005400000000",
            INIT_11 => X"0000004800000000000000560000000000000050000000000000004900000000",
            INIT_12 => X"0000004300000000000000380000000000000041000000000000004600000000",
            INIT_13 => X"0000003c0000000000000036000000000000003f000000000000004800000000",
            INIT_14 => X"0000003a000000000000003d0000000000000041000000000000004200000000",
            INIT_15 => X"00000026000000000000002d000000000000002f000000000000003000000000",
            INIT_16 => X"0000002500000000000000220000000000000021000000000000002400000000",
            INIT_17 => X"0000002c000000000000002a0000000000000029000000000000002a00000000",
            INIT_18 => X"0000005000000000000000520000000000000053000000000000005500000000",
            INIT_19 => X"0000002b000000000000004d0000000000000052000000000000004800000000",
            INIT_1A => X"0000003400000000000000320000000000000045000000000000004300000000",
            INIT_1B => X"0000002f0000000000000032000000000000003f000000000000004100000000",
            INIT_1C => X"0000003600000000000000390000000000000034000000000000003200000000",
            INIT_1D => X"0000002c000000000000002b000000000000002b000000000000002d00000000",
            INIT_1E => X"0000003b00000000000000380000000000000032000000000000002f00000000",
            INIT_1F => X"000000370000000000000038000000000000003b000000000000003c00000000",
            INIT_20 => X"0000005100000000000000510000000000000051000000000000005200000000",
            INIT_21 => X"0000002c0000000000000046000000000000004c000000000000004800000000",
            INIT_22 => X"0000001d00000000000000220000000000000033000000000000003d00000000",
            INIT_23 => X"0000002300000000000000260000000000000027000000000000001f00000000",
            INIT_24 => X"0000003b0000000000000039000000000000002b000000000000002900000000",
            INIT_25 => X"000000440000000000000041000000000000003d000000000000003d00000000",
            INIT_26 => X"0000004800000000000000470000000000000042000000000000004400000000",
            INIT_27 => X"00000038000000000000003e0000000000000043000000000000004700000000",
            INIT_28 => X"0000004f000000000000004c000000000000004c000000000000004d00000000",
            INIT_29 => X"00000038000000000000003e0000000000000042000000000000004700000000",
            INIT_2A => X"00000017000000000000001a0000000000000021000000000000002c00000000",
            INIT_2B => X"0000000e000000000000000f0000000000000014000000000000001600000000",
            INIT_2C => X"00000054000000000000004f0000000000000035000000000000001f00000000",
            INIT_2D => X"00000050000000000000004e0000000000000052000000000000005300000000",
            INIT_2E => X"0000004b000000000000004d0000000000000048000000000000004c00000000",
            INIT_2F => X"0000002e0000000000000035000000000000003c000000000000004400000000",
            INIT_30 => X"0000004800000000000000460000000000000047000000000000004900000000",
            INIT_31 => X"0000002000000000000000200000000000000037000000000000004700000000",
            INIT_32 => X"0000001300000000000000140000000000000018000000000000002600000000",
            INIT_33 => X"00000015000000000000000e000000000000000b000000000000001200000000",
            INIT_34 => X"0000005900000000000000460000000000000029000000000000001800000000",
            INIT_35 => X"00000052000000000000004f0000000000000050000000000000005600000000",
            INIT_36 => X"0000004300000000000000480000000000000048000000000000004b00000000",
            INIT_37 => X"0000002a000000000000002d0000000000000034000000000000003b00000000",
            INIT_38 => X"0000004500000000000000440000000000000045000000000000004400000000",
            INIT_39 => X"00000011000000000000001c0000000000000033000000000000004300000000",
            INIT_3A => X"0000000b000000000000000a000000000000000c000000000000001700000000",
            INIT_3B => X"000000180000000000000011000000000000000b000000000000000900000000",
            INIT_3C => X"0000003f00000000000000210000000000000016000000000000001c00000000",
            INIT_3D => X"00000040000000000000004d000000000000004f000000000000004d00000000",
            INIT_3E => X"0000004200000000000000480000000000000049000000000000004100000000",
            INIT_3F => X"0000002b000000000000002f0000000000000036000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004e00000000000000470000000000000045000000000000004400000000",
            INIT_41 => X"000000130000000000000046000000000000005d000000000000005200000000",
            INIT_42 => X"000000250000000000000019000000000000000c000000000000001200000000",
            INIT_43 => X"0000001400000000000000210000000000000021000000000000002000000000",
            INIT_44 => X"0000002100000000000000190000000000000018000000000000001600000000",
            INIT_45 => X"0000003b000000000000003c0000000000000038000000000000003100000000",
            INIT_46 => X"0000003f0000000000000049000000000000004b000000000000003b00000000",
            INIT_47 => X"0000003500000000000000340000000000000034000000000000003900000000",
            INIT_48 => X"0000007500000000000000670000000000000059000000000000005000000000",
            INIT_49 => X"000000160000000000000055000000000000008d000000000000008000000000",
            INIT_4A => X"000000380000000000000021000000000000000f000000000000001500000000",
            INIT_4B => X"0000001c0000000000000035000000000000003d000000000000003900000000",
            INIT_4C => X"0000001400000000000000160000000000000016000000000000001500000000",
            INIT_4D => X"0000003a000000000000002d0000000000000023000000000000001800000000",
            INIT_4E => X"0000004100000000000000460000000000000048000000000000003d00000000",
            INIT_4F => X"0000003d000000000000003f0000000000000040000000000000004100000000",
            INIT_50 => X"00000095000000000000008e0000000000000083000000000000007700000000",
            INIT_51 => X"0000001800000000000000470000000000000098000000000000009800000000",
            INIT_52 => X"0000003100000000000000150000000000000011000000000000001e00000000",
            INIT_53 => X"00000021000000000000003f0000000000000044000000000000003c00000000",
            INIT_54 => X"000000110000000000000015000000000000001b000000000000001900000000",
            INIT_55 => X"0000002b000000000000001c0000000000000014000000000000000f00000000",
            INIT_56 => X"0000004a000000000000004d0000000000000046000000000000003700000000",
            INIT_57 => X"0000004100000000000000440000000000000047000000000000004900000000",
            INIT_58 => X"0000009900000000000000960000000000000094000000000000008f00000000",
            INIT_59 => X"00000017000000000000004f0000000000000099000000000000009900000000",
            INIT_5A => X"0000002e00000000000000190000000000000022000000000000002800000000",
            INIT_5B => X"0000002700000000000000370000000000000030000000000000003d00000000",
            INIT_5C => X"00000015000000000000001f0000000000000024000000000000001d00000000",
            INIT_5D => X"0000001f00000000000000120000000000000015000000000000001300000000",
            INIT_5E => X"0000004d000000000000004c000000000000003b000000000000002a00000000",
            INIT_5F => X"00000045000000000000004a000000000000004c000000000000004d00000000",
            INIT_60 => X"0000009400000000000000970000000000000095000000000000009200000000",
            INIT_61 => X"00000020000000000000006b0000000000000092000000000000009200000000",
            INIT_62 => X"0000003b00000000000000340000000000000037000000000000002b00000000",
            INIT_63 => X"00000029000000000000002c0000000000000034000000000000004700000000",
            INIT_64 => X"0000001e000000000000002c0000000000000032000000000000002200000000",
            INIT_65 => X"000000190000000000000012000000000000001c000000000000001a00000000",
            INIT_66 => X"0000005100000000000000450000000000000032000000000000002e00000000",
            INIT_67 => X"000000420000000000000049000000000000004f000000000000005100000000",
            INIT_68 => X"0000008b000000000000008f000000000000008f000000000000009000000000",
            INIT_69 => X"00000040000000000000007e0000000000000089000000000000008a00000000",
            INIT_6A => X"00000041000000000000003d000000000000002e000000000000001a00000000",
            INIT_6B => X"0000002400000000000000280000000000000040000000000000004600000000",
            INIT_6C => X"0000002800000000000000330000000000000036000000000000002400000000",
            INIT_6D => X"000000130000000000000012000000000000001d000000000000002100000000",
            INIT_6E => X"0000004e000000000000003c0000000000000033000000000000002f00000000",
            INIT_6F => X"000000370000000000000040000000000000004a000000000000004f00000000",
            INIT_70 => X"0000008600000000000000860000000000000084000000000000008500000000",
            INIT_71 => X"0000007700000000000000890000000000000088000000000000008600000000",
            INIT_72 => X"00000021000000000000001b0000000000000031000000000000004700000000",
            INIT_73 => X"000000220000000000000020000000000000002a000000000000002e00000000",
            INIT_74 => X"00000032000000000000003d0000000000000039000000000000002800000000",
            INIT_75 => X"000000110000000000000011000000000000001c000000000000002700000000",
            INIT_76 => X"0000004100000000000000300000000000000033000000000000002400000000",
            INIT_77 => X"000000320000000000000036000000000000003e000000000000004600000000",
            INIT_78 => X"000000850000000000000081000000000000007f000000000000007d00000000",
            INIT_79 => X"0000008100000000000000880000000000000091000000000000008c00000000",
            INIT_7A => X"0000001e000000000000001e000000000000005a000000000000008400000000",
            INIT_7B => X"0000002700000000000000270000000000000033000000000000004000000000",
            INIT_7C => X"0000003d00000000000000450000000000000045000000000000003100000000",
            INIT_7D => X"000000130000000000000014000000000000001c000000000000002c00000000",
            INIT_7E => X"0000002d00000000000000290000000000000030000000000000001900000000",
            INIT_7F => X"0000003d000000000000003c0000000000000039000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "sampleifmap_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000091000000000000008b0000000000000084000000000000007d00000000",
            INIT_01 => X"0000005a00000000000000750000000000000091000000000000009500000000",
            INIT_02 => X"0000005000000000000000620000000000000072000000000000008000000000",
            INIT_03 => X"000000280000000000000031000000000000004d000000000000005700000000",
            INIT_04 => X"0000003c0000000000000044000000000000003f000000000000002e00000000",
            INIT_05 => X"000000170000000000000019000000000000001f000000000000002d00000000",
            INIT_06 => X"0000002d000000000000002b000000000000002a000000000000001500000000",
            INIT_07 => X"00000032000000000000003e0000000000000042000000000000004000000000",
            INIT_08 => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_09 => X"00000068000000000000009e00000000000000a4000000000000009a00000000",
            INIT_0A => X"00000077000000000000007a00000000000000a6000000000000009500000000",
            INIT_0B => X"00000029000000000000004b0000000000000067000000000000005000000000",
            INIT_0C => X"0000003c00000000000000410000000000000038000000000000002d00000000",
            INIT_0D => X"0000001b000000000000001f0000000000000028000000000000003000000000",
            INIT_0E => X"00000032000000000000002f0000000000000023000000000000001500000000",
            INIT_0F => X"0000001400000000000000230000000000000039000000000000004100000000",
            INIT_10 => X"000000b600000000000000a40000000000000097000000000000009000000000",
            INIT_11 => X"000000b200000000000000eb00000000000000e600000000000000d200000000",
            INIT_12 => X"00000095000000000000008a00000000000000ab000000000000008500000000",
            INIT_13 => X"0000002d00000000000000550000000000000067000000000000004d00000000",
            INIT_14 => X"0000003c000000000000003f0000000000000038000000000000002b00000000",
            INIT_15 => X"0000001d00000000000000270000000000000030000000000000003500000000",
            INIT_16 => X"00000027000000000000002f000000000000001d000000000000001700000000",
            INIT_17 => X"000000150000000000000016000000000000001f000000000000002700000000",
            INIT_18 => X"000000f000000000000000e100000000000000cd00000000000000b700000000",
            INIT_19 => X"000000e600000000000000f200000000000000f200000000000000f800000000",
            INIT_1A => X"0000009f00000000000000840000000000000084000000000000008d00000000",
            INIT_1B => X"000000310000000000000056000000000000004d000000000000005300000000",
            INIT_1C => X"0000003a000000000000003c0000000000000037000000000000002a00000000",
            INIT_1D => X"00000021000000000000002f0000000000000037000000000000003900000000",
            INIT_1E => X"0000001c0000000000000027000000000000001a000000000000001900000000",
            INIT_1F => X"0000001b000000000000001c000000000000001d000000000000001900000000",
            INIT_20 => X"000000f900000000000000f700000000000000f800000000000000f100000000",
            INIT_21 => X"000000b500000000000000ab00000000000000b000000000000000ec00000000",
            INIT_22 => X"0000007600000000000000720000000000000062000000000000007800000000",
            INIT_23 => X"000000340000000000000047000000000000003c000000000000004d00000000",
            INIT_24 => X"0000003a00000000000000390000000000000036000000000000002e00000000",
            INIT_25 => X"0000002000000000000000300000000000000039000000000000003b00000000",
            INIT_26 => X"0000002500000000000000250000000000000017000000000000001800000000",
            INIT_27 => X"0000001a000000000000001f0000000000000020000000000000001c00000000",
            INIT_28 => X"000000fd00000000000000f900000000000000f900000000000000f800000000",
            INIT_29 => X"000000550000000000000053000000000000006a00000000000000e000000000",
            INIT_2A => X"000000410000000000000051000000000000004e000000000000004700000000",
            INIT_2B => X"000000310000000000000034000000000000002e000000000000003000000000",
            INIT_2C => X"0000003900000000000000360000000000000037000000000000003300000000",
            INIT_2D => X"0000001b00000000000000240000000000000033000000000000003d00000000",
            INIT_2E => X"0000003600000000000000270000000000000016000000000000001500000000",
            INIT_2F => X"0000001c000000000000001f000000000000001f000000000000002800000000",
            INIT_30 => X"000000eb00000000000000f500000000000000f800000000000000f700000000",
            INIT_31 => X"0000005e0000000000000060000000000000006d00000000000000c200000000",
            INIT_32 => X"0000001900000000000000230000000000000035000000000000004100000000",
            INIT_33 => X"00000020000000000000002d000000000000002b000000000000001c00000000",
            INIT_34 => X"0000002f000000000000002f0000000000000033000000000000002e00000000",
            INIT_35 => X"00000029000000000000002b000000000000002d000000000000003000000000",
            INIT_36 => X"0000003a0000000000000024000000000000001e000000000000002200000000",
            INIT_37 => X"0000001e000000000000001d0000000000000021000000000000003900000000",
            INIT_38 => X"0000009800000000000000b600000000000000d700000000000000ec00000000",
            INIT_39 => X"00000074000000000000007a0000000000000081000000000000008800000000",
            INIT_3A => X"00000009000000000000000d0000000000000023000000000000005100000000",
            INIT_3B => X"0000002200000000000000490000000000000034000000000000001400000000",
            INIT_3C => X"00000020000000000000001a000000000000001c000000000000001100000000",
            INIT_3D => X"00000031000000000000003b000000000000003b000000000000002f00000000",
            INIT_3E => X"000000340000000000000022000000000000001a000000000000002300000000",
            INIT_3F => X"0000001d000000000000001c000000000000002c000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009a00000000",
            INIT_41 => X"0000005c00000000000000680000000000000076000000000000007b00000000",
            INIT_42 => X"00000012000000000000001f0000000000000046000000000000005a00000000",
            INIT_43 => X"000000340000000000000045000000000000003d000000000000001d00000000",
            INIT_44 => X"0000002800000000000000240000000000000024000000000000002200000000",
            INIT_45 => X"0000003d00000000000000410000000000000047000000000000003a00000000",
            INIT_46 => X"00000028000000000000001f0000000000000017000000000000003000000000",
            INIT_47 => X"0000001c0000000000000027000000000000003c000000000000003800000000",
            INIT_48 => X"00000068000000000000006d000000000000006b000000000000006900000000",
            INIT_49 => X"0000005d000000000000005b0000000000000058000000000000005f00000000",
            INIT_4A => X"0000003e00000000000000560000000000000062000000000000006000000000",
            INIT_4B => X"00000031000000000000002f0000000000000038000000000000003800000000",
            INIT_4C => X"00000030000000000000002a0000000000000025000000000000002800000000",
            INIT_4D => X"000000390000000000000048000000000000005b000000000000004c00000000",
            INIT_4E => X"00000023000000000000001d000000000000002c000000000000003600000000",
            INIT_4F => X"0000001d0000000000000037000000000000003d000000000000002a00000000",
            INIT_50 => X"0000005100000000000000530000000000000059000000000000005f00000000",
            INIT_51 => X"00000058000000000000005b0000000000000058000000000000005600000000",
            INIT_52 => X"0000003e00000000000000440000000000000049000000000000005300000000",
            INIT_53 => X"00000034000000000000002c0000000000000023000000000000002800000000",
            INIT_54 => X"000000310000000000000027000000000000001e000000000000002800000000",
            INIT_55 => X"000000320000000000000047000000000000005f000000000000005100000000",
            INIT_56 => X"000000230000000000000025000000000000002a000000000000002900000000",
            INIT_57 => X"00000028000000000000003a0000000000000030000000000000002200000000",
            INIT_58 => X"00000055000000000000004f0000000000000049000000000000004b00000000",
            INIT_59 => X"00000040000000000000004c0000000000000053000000000000005700000000",
            INIT_5A => X"0000003b000000000000002a0000000000000027000000000000003300000000",
            INIT_5B => X"0000003100000000000000290000000000000022000000000000003200000000",
            INIT_5C => X"000000270000000000000024000000000000001e000000000000002600000000",
            INIT_5D => X"0000002d000000000000003c0000000000000045000000000000003700000000",
            INIT_5E => X"0000001d00000000000000220000000000000026000000000000002600000000",
            INIT_5F => X"0000003300000000000000300000000000000024000000000000002000000000",
            INIT_60 => X"0000004d000000000000004f000000000000004e000000000000004c00000000",
            INIT_61 => X"00000021000000000000002c0000000000000039000000000000004400000000",
            INIT_62 => X"0000003d000000000000002e000000000000001e000000000000001d00000000",
            INIT_63 => X"0000002600000000000000320000000000000029000000000000003700000000",
            INIT_64 => X"0000001e000000000000001d000000000000001a000000000000001d00000000",
            INIT_65 => X"00000030000000000000002e0000000000000025000000000000001d00000000",
            INIT_66 => X"0000001800000000000000190000000000000025000000000000002e00000000",
            INIT_67 => X"0000002f00000000000000240000000000000020000000000000001e00000000",
            INIT_68 => X"000000320000000000000040000000000000004a000000000000005000000000",
            INIT_69 => X"0000001b000000000000001e0000000000000020000000000000002600000000",
            INIT_6A => X"0000003c000000000000002d000000000000001b000000000000001b00000000",
            INIT_6B => X"0000001d000000000000002c000000000000002f000000000000003500000000",
            INIT_6C => X"0000001c00000000000000170000000000000017000000000000001c00000000",
            INIT_6D => X"0000002500000000000000200000000000000018000000000000001900000000",
            INIT_6E => X"000000150000000000000015000000000000001d000000000000002300000000",
            INIT_6F => X"00000022000000000000001c000000000000001e000000000000001a00000000",
            INIT_70 => X"0000001a0000000000000021000000000000002d000000000000003a00000000",
            INIT_71 => X"0000001c0000000000000021000000000000001d000000000000001a00000000",
            INIT_72 => X"0000003300000000000000270000000000000018000000000000001b00000000",
            INIT_73 => X"0000001c00000000000000210000000000000032000000000000003100000000",
            INIT_74 => X"0000001d00000000000000190000000000000015000000000000001b00000000",
            INIT_75 => X"0000001700000000000000190000000000000015000000000000001800000000",
            INIT_76 => X"000000120000000000000016000000000000001a000000000000001700000000",
            INIT_77 => X"000000170000000000000019000000000000001a000000000000001500000000",
            INIT_78 => X"0000001500000000000000180000000000000017000000000000001b00000000",
            INIT_79 => X"0000001900000000000000180000000000000019000000000000001a00000000",
            INIT_7A => X"0000003000000000000000210000000000000016000000000000001a00000000",
            INIT_7B => X"0000001800000000000000230000000000000033000000000000002a00000000",
            INIT_7C => X"0000001800000000000000150000000000000014000000000000001500000000",
            INIT_7D => X"00000019000000000000001d0000000000000017000000000000001700000000",
            INIT_7E => X"000000120000000000000016000000000000001b000000000000001800000000",
            INIT_7F => X"0000001600000000000000180000000000000016000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "sampleifmap_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004100000000000000150000000000000013000000000000001700000000",
            INIT_01 => X"000000b200000000000000b700000000000000bc00000000000000a400000000",
            INIT_02 => X"000000ba00000000000000ba00000000000000ac00000000000000aa00000000",
            INIT_03 => X"000000b700000000000000b600000000000000b700000000000000b800000000",
            INIT_04 => X"0000005c000000000000007f00000000000000a400000000000000b400000000",
            INIT_05 => X"000000c20000000000000099000000000000006e000000000000006b00000000",
            INIT_06 => X"000000c600000000000000c500000000000000c900000000000000c300000000",
            INIT_07 => X"000000c500000000000000c700000000000000c800000000000000c900000000",
            INIT_08 => X"0000002e00000000000000150000000000000013000000000000001700000000",
            INIT_09 => X"000000b200000000000000bf00000000000000ca000000000000009900000000",
            INIT_0A => X"000000b700000000000000a9000000000000009e00000000000000a400000000",
            INIT_0B => X"000000b200000000000000b400000000000000b800000000000000ba00000000",
            INIT_0C => X"00000056000000000000008a00000000000000ad00000000000000b400000000",
            INIT_0D => X"000000ce00000000000000b4000000000000006a000000000000004a00000000",
            INIT_0E => X"000000ce00000000000000d000000000000000d500000000000000cf00000000",
            INIT_0F => X"000000ca00000000000000cc00000000000000cd00000000000000cf00000000",
            INIT_10 => X"0000001f00000000000000170000000000000014000000000000001700000000",
            INIT_11 => X"000000a800000000000000b900000000000000c8000000000000007f00000000",
            INIT_12 => X"000000a2000000000000009a000000000000009e000000000000009f00000000",
            INIT_13 => X"000000b200000000000000b300000000000000b200000000000000b200000000",
            INIT_14 => X"0000007d00000000000000b600000000000000be00000000000000b500000000",
            INIT_15 => X"000000d100000000000000c50000000000000072000000000000004700000000",
            INIT_16 => X"000000d300000000000000d500000000000000d800000000000000d500000000",
            INIT_17 => X"000000ce00000000000000d000000000000000d300000000000000d400000000",
            INIT_18 => X"0000001700000000000000180000000000000015000000000000001700000000",
            INIT_19 => X"000000a000000000000000af00000000000000bd000000000000006300000000",
            INIT_1A => X"0000009500000000000000a600000000000000a800000000000000a800000000",
            INIT_1B => X"000000c300000000000000bf00000000000000ba00000000000000aa00000000",
            INIT_1C => X"0000008d00000000000000bc00000000000000c800000000000000c300000000",
            INIT_1D => X"000000d600000000000000d20000000000000092000000000000006300000000",
            INIT_1E => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1F => X"000000d600000000000000d700000000000000d900000000000000d900000000",
            INIT_20 => X"0000001500000000000000170000000000000017000000000000001900000000",
            INIT_21 => X"0000009700000000000000a500000000000000aa000000000000004800000000",
            INIT_22 => X"0000009b00000000000000b900000000000000b700000000000000af00000000",
            INIT_23 => X"000000bc00000000000000a9000000000000009d000000000000009200000000",
            INIT_24 => X"0000008d00000000000000b200000000000000c400000000000000c500000000",
            INIT_25 => X"000000db00000000000000d300000000000000ac000000000000007900000000",
            INIT_26 => X"000000d900000000000000d900000000000000d900000000000000dd00000000",
            INIT_27 => X"000000ce00000000000000d100000000000000d400000000000000d600000000",
            INIT_28 => X"00000017000000000000001a000000000000001b000000000000001a00000000",
            INIT_29 => X"0000009a00000000000000a4000000000000008f000000000000003100000000",
            INIT_2A => X"000000a600000000000000c800000000000000c200000000000000a900000000",
            INIT_2B => X"000000970000000000000080000000000000007d000000000000008200000000",
            INIT_2C => X"0000008f000000000000009400000000000000a500000000000000a500000000",
            INIT_2D => X"000000c900000000000000bc00000000000000b6000000000000009300000000",
            INIT_2E => X"000000db00000000000000d500000000000000d900000000000000d400000000",
            INIT_2F => X"000000d300000000000000d700000000000000d700000000000000dc00000000",
            INIT_30 => X"00000019000000000000001b000000000000001a000000000000001e00000000",
            INIT_31 => X"000000ab00000000000000b4000000000000007d000000000000002500000000",
            INIT_32 => X"000000b300000000000000ca00000000000000c500000000000000a900000000",
            INIT_33 => X"00000082000000000000007a0000000000000071000000000000008b00000000",
            INIT_34 => X"0000008c000000000000007a0000000000000085000000000000007700000000",
            INIT_35 => X"000000c900000000000000bf00000000000000cb00000000000000b900000000",
            INIT_36 => X"000000db00000000000000d700000000000000da00000000000000d700000000",
            INIT_37 => X"000000e000000000000000dc00000000000000da00000000000000dc00000000",
            INIT_38 => X"00000024000000000000001f0000000000000030000000000000005e00000000",
            INIT_39 => X"000000a800000000000000c100000000000000af000000000000006400000000",
            INIT_3A => X"000000c300000000000000c600000000000000c000000000000000a300000000",
            INIT_3B => X"00000084000000000000008e000000000000009100000000000000ae00000000",
            INIT_3C => X"0000008b000000000000007a0000000000000079000000000000006a00000000",
            INIT_3D => X"000000d500000000000000bd00000000000000d100000000000000c000000000",
            INIT_3E => X"000000e800000000000000ef00000000000000ed00000000000000f200000000",
            INIT_3F => X"000000e500000000000000de00000000000000d500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007a0000000000000072000000000000009e00000000000000b400000000",
            INIT_41 => X"000000a000000000000000be00000000000000be00000000000000b100000000",
            INIT_42 => X"000000c800000000000000c500000000000000ad000000000000008500000000",
            INIT_43 => X"0000009200000000000000a700000000000000b900000000000000c200000000",
            INIT_44 => X"0000008d00000000000000850000000000000081000000000000008100000000",
            INIT_45 => X"000000dc00000000000000bd00000000000000c900000000000000b100000000",
            INIT_46 => X"000000d500000000000000e800000000000000eb00000000000000f100000000",
            INIT_47 => X"000000ea00000000000000e100000000000000c700000000000000bd00000000",
            INIT_48 => X"000000ba00000000000000b200000000000000c000000000000000c500000000",
            INIT_49 => X"0000009d00000000000000c500000000000000c300000000000000c100000000",
            INIT_4A => X"000000bf00000000000000b900000000000000a3000000000000008000000000",
            INIT_4B => X"0000009700000000000000b200000000000000c300000000000000c100000000",
            INIT_4C => X"0000008600000000000000830000000000000081000000000000007200000000",
            INIT_4D => X"000000ea00000000000000d000000000000000c200000000000000aa00000000",
            INIT_4E => X"000000c900000000000000eb00000000000000f000000000000000ec00000000",
            INIT_4F => X"000000eb00000000000000d000000000000000bb00000000000000b900000000",
            INIT_50 => X"000000c000000000000000bb00000000000000c400000000000000ca00000000",
            INIT_51 => X"0000009700000000000000c500000000000000cd00000000000000c800000000",
            INIT_52 => X"000000bd00000000000000b800000000000000af000000000000009500000000",
            INIT_53 => X"0000008800000000000000a800000000000000bb00000000000000c100000000",
            INIT_54 => X"0000008100000000000000800000000000000080000000000000007500000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b500000000000000a700000000",
            INIT_56 => X"000000ce00000000000000ee00000000000000f300000000000000f300000000",
            INIT_57 => X"000000dd00000000000000c100000000000000bb00000000000000ba00000000",
            INIT_58 => X"000000c000000000000000c500000000000000cd00000000000000cd00000000",
            INIT_59 => X"000000a000000000000000c200000000000000d000000000000000cb00000000",
            INIT_5A => X"000000bf00000000000000c100000000000000bf00000000000000a800000000",
            INIT_5B => X"00000077000000000000009200000000000000ac00000000000000c100000000",
            INIT_5C => X"000000870000000000000085000000000000008e000000000000007c00000000",
            INIT_5D => X"000000ea00000000000000bf00000000000000b000000000000000a700000000",
            INIT_5E => X"000000d700000000000000ec00000000000000f100000000000000f300000000",
            INIT_5F => X"000000c400000000000000b900000000000000b800000000000000ba00000000",
            INIT_60 => X"000000c100000000000000c800000000000000cc00000000000000ce00000000",
            INIT_61 => X"000000b400000000000000bf00000000000000c700000000000000c500000000",
            INIT_62 => X"000000ad00000000000000b700000000000000b300000000000000ac00000000",
            INIT_63 => X"00000083000000000000009800000000000000ae00000000000000ae00000000",
            INIT_64 => X"0000009a000000000000008e00000000000000a6000000000000008d00000000",
            INIT_65 => X"000000e600000000000000bf00000000000000ac00000000000000a900000000",
            INIT_66 => X"000000e400000000000000ef00000000000000f100000000000000f000000000",
            INIT_67 => X"000000c000000000000000b800000000000000ba00000000000000c800000000",
            INIT_68 => X"000000bf00000000000000c600000000000000ca00000000000000d200000000",
            INIT_69 => X"000000ca00000000000000b100000000000000b400000000000000c900000000",
            INIT_6A => X"0000008e000000000000008e000000000000009a00000000000000ab00000000",
            INIT_6B => X"0000009c000000000000009300000000000000a800000000000000a800000000",
            INIT_6C => X"000000a4000000000000009600000000000000a900000000000000af00000000",
            INIT_6D => X"000000e600000000000000c500000000000000a0000000000000009e00000000",
            INIT_6E => X"000000f200000000000000f400000000000000f100000000000000f100000000",
            INIT_6F => X"000000d700000000000000c300000000000000bf00000000000000e200000000",
            INIT_70 => X"000000c000000000000000c700000000000000c900000000000000d300000000",
            INIT_71 => X"000000d700000000000000a100000000000000aa00000000000000cf00000000",
            INIT_72 => X"000000ac00000000000000ad00000000000000ba00000000000000bd00000000",
            INIT_73 => X"0000007f000000000000008900000000000000b100000000000000be00000000",
            INIT_74 => X"000000a0000000000000009600000000000000ae00000000000000b400000000",
            INIT_75 => X"000000ec00000000000000c100000000000000b000000000000000af00000000",
            INIT_76 => X"000000fb00000000000000f300000000000000f200000000000000f500000000",
            INIT_77 => X"000000e100000000000000d400000000000000c900000000000000ef00000000",
            INIT_78 => X"000000c100000000000000c500000000000000c400000000000000d300000000",
            INIT_79 => X"000000d9000000000000009a00000000000000b500000000000000d100000000",
            INIT_7A => X"000000b900000000000000c300000000000000c500000000000000ce00000000",
            INIT_7B => X"0000009800000000000000a600000000000000ad00000000000000aa00000000",
            INIT_7C => X"0000009800000000000000a600000000000000b800000000000000a300000000",
            INIT_7D => X"000000cc00000000000000af00000000000000b500000000000000c000000000",
            INIT_7E => X"000000f700000000000000f400000000000000f300000000000000ee00000000",
            INIT_7F => X"000000e200000000000000e200000000000000d500000000000000df00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "sampleifmap_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b500000000000000b400000000000000c200000000000000d600000000",
            INIT_01 => X"000000c6000000000000009b00000000000000c400000000000000c500000000",
            INIT_02 => X"000000b700000000000000ae00000000000000c000000000000000d600000000",
            INIT_03 => X"000000b200000000000000ae00000000000000a100000000000000ad00000000",
            INIT_04 => X"0000009300000000000000bd00000000000000a4000000000000008000000000",
            INIT_05 => X"00000076000000000000009c00000000000000b400000000000000a700000000",
            INIT_06 => X"000000eb00000000000000ef00000000000000d7000000000000009d00000000",
            INIT_07 => X"000000e400000000000000ea00000000000000d600000000000000ce00000000",
            INIT_08 => X"000000a300000000000000a600000000000000c600000000000000d700000000",
            INIT_09 => X"000000b900000000000000be00000000000000ca00000000000000b400000000",
            INIT_0A => X"000000d600000000000000cd00000000000000d200000000000000cf00000000",
            INIT_0B => X"000000ad00000000000000b000000000000000ae00000000000000c100000000",
            INIT_0C => X"0000009900000000000000bf0000000000000089000000000000008100000000",
            INIT_0D => X"0000008700000000000000ab00000000000000c800000000000000a300000000",
            INIT_0E => X"000000c100000000000000b80000000000000090000000000000007400000000",
            INIT_0F => X"000000eb00000000000000ef00000000000000d200000000000000bb00000000",
            INIT_10 => X"000000a400000000000000ae00000000000000cd00000000000000d800000000",
            INIT_11 => X"000000c200000000000000d200000000000000cb00000000000000b900000000",
            INIT_12 => X"000000e200000000000000da00000000000000d300000000000000bf00000000",
            INIT_13 => X"000000b300000000000000be00000000000000cb00000000000000e100000000",
            INIT_14 => X"0000009e00000000000000a80000000000000079000000000000009700000000",
            INIT_15 => X"000000ac00000000000000aa00000000000000c200000000000000a700000000",
            INIT_16 => X"000000a900000000000000990000000000000083000000000000009a00000000",
            INIT_17 => X"000000ec00000000000000de00000000000000b800000000000000a200000000",
            INIT_18 => X"000000b400000000000000c000000000000000d000000000000000d800000000",
            INIT_19 => X"000000d200000000000000d100000000000000ca00000000000000c500000000",
            INIT_1A => X"000000cc00000000000000c500000000000000bd00000000000000ba00000000",
            INIT_1B => X"000000b500000000000000cf00000000000000d500000000000000d100000000",
            INIT_1C => X"000000af0000000000000092000000000000009500000000000000b200000000",
            INIT_1D => X"000000ab000000000000009c00000000000000ae00000000000000b700000000",
            INIT_1E => X"000000b400000000000000a9000000000000009400000000000000a300000000",
            INIT_1F => X"000000cc00000000000000ac00000000000000a000000000000000a600000000",
            INIT_20 => X"000000b600000000000000ca00000000000000d500000000000000da00000000",
            INIT_21 => X"000000ca00000000000000c900000000000000cb00000000000000bf00000000",
            INIT_22 => X"000000c000000000000000c100000000000000c300000000000000ca00000000",
            INIT_23 => X"000000c700000000000000cf00000000000000c600000000000000b200000000",
            INIT_24 => X"000000bb00000000000000a600000000000000cb00000000000000d300000000",
            INIT_25 => X"000000a60000000000000093000000000000009b00000000000000b100000000",
            INIT_26 => X"000000af00000000000000b600000000000000ab00000000000000a700000000",
            INIT_27 => X"000000a7000000000000009f000000000000009c000000000000009c00000000",
            INIT_28 => X"000000ba00000000000000d100000000000000d700000000000000d900000000",
            INIT_29 => X"000000c800000000000000d000000000000000c800000000000000b300000000",
            INIT_2A => X"000000ba00000000000000d200000000000000d700000000000000d100000000",
            INIT_2B => X"000000c200000000000000c400000000000000b600000000000000a100000000",
            INIT_2C => X"000000b900000000000000be00000000000000cf00000000000000cb00000000",
            INIT_2D => X"000000a6000000000000009b000000000000008e000000000000009b00000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000b300000000000000ac00000000",
            INIT_2F => X"0000008f000000000000009e000000000000009e000000000000009600000000",
            INIT_30 => X"000000c000000000000000d600000000000000d500000000000000d600000000",
            INIT_31 => X"000000d900000000000000da00000000000000c500000000000000a900000000",
            INIT_32 => X"000000c300000000000000d400000000000000d900000000000000d700000000",
            INIT_33 => X"000000bf00000000000000c300000000000000b300000000000000aa00000000",
            INIT_34 => X"000000aa00000000000000c000000000000000c000000000000000be00000000",
            INIT_35 => X"000000aa00000000000000a7000000000000008e000000000000008400000000",
            INIT_36 => X"0000009d00000000000000ad00000000000000b300000000000000aa00000000",
            INIT_37 => X"0000007d00000000000000860000000000000093000000000000009d00000000",
            INIT_38 => X"000000ca00000000000000d300000000000000d100000000000000d500000000",
            INIT_39 => X"000000de00000000000000d800000000000000c100000000000000a800000000",
            INIT_3A => X"000000cd00000000000000d300000000000000de00000000000000df00000000",
            INIT_3B => X"000000c600000000000000c900000000000000c200000000000000c200000000",
            INIT_3C => X"0000009900000000000000bc00000000000000c400000000000000c600000000",
            INIT_3D => X"000000a700000000000000ab000000000000009b000000000000008600000000",
            INIT_3E => X"000000a500000000000000b200000000000000bd00000000000000a600000000",
            INIT_3F => X"000000890000000000000085000000000000008e00000000000000a300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ca00000000000000ce00000000000000ce00000000000000d300000000",
            INIT_41 => X"000000d500000000000000d300000000000000bf00000000000000af00000000",
            INIT_42 => X"000000ab00000000000000c600000000000000d800000000000000d600000000",
            INIT_43 => X"000000c900000000000000c900000000000000ce00000000000000c200000000",
            INIT_44 => X"0000009600000000000000b100000000000000c500000000000000c800000000",
            INIT_45 => X"0000009d00000000000000a7000000000000009e000000000000009000000000",
            INIT_46 => X"000000a800000000000000b000000000000000b5000000000000009f00000000",
            INIT_47 => X"0000009000000000000000950000000000000096000000000000009800000000",
            INIT_48 => X"000000c100000000000000c900000000000000cc00000000000000d200000000",
            INIT_49 => X"000000d200000000000000d000000000000000bc00000000000000b500000000",
            INIT_4A => X"0000007a00000000000000a000000000000000ce00000000000000cd00000000",
            INIT_4B => X"000000c200000000000000c600000000000000d000000000000000b100000000",
            INIT_4C => X"0000009600000000000000a600000000000000b800000000000000c100000000",
            INIT_4D => X"0000009900000000000000a0000000000000009c000000000000008b00000000",
            INIT_4E => X"0000009b000000000000009f00000000000000a0000000000000009b00000000",
            INIT_4F => X"00000083000000000000008c0000000000000098000000000000009800000000",
            INIT_50 => X"000000bb00000000000000c600000000000000ca00000000000000d200000000",
            INIT_51 => X"000000d600000000000000cd00000000000000b200000000000000ae00000000",
            INIT_52 => X"0000008300000000000000a400000000000000cb00000000000000d100000000",
            INIT_53 => X"000000b600000000000000bb00000000000000ca00000000000000b400000000",
            INIT_54 => X"0000008b000000000000009d00000000000000a900000000000000b600000000",
            INIT_55 => X"00000090000000000000009a0000000000000099000000000000008600000000",
            INIT_56 => X"0000008d0000000000000083000000000000008d000000000000009700000000",
            INIT_57 => X"000000930000000000000096000000000000009b000000000000009d00000000",
            INIT_58 => X"000000b500000000000000c200000000000000c800000000000000d200000000",
            INIT_59 => X"000000d700000000000000c400000000000000a800000000000000a800000000",
            INIT_5A => X"000000b800000000000000bd00000000000000c700000000000000d400000000",
            INIT_5B => X"000000ac00000000000000ad00000000000000b900000000000000cb00000000",
            INIT_5C => X"000000760000000000000093000000000000009b00000000000000a300000000",
            INIT_5D => X"0000008d00000000000000910000000000000094000000000000008300000000",
            INIT_5E => X"00000085000000000000007f0000000000000084000000000000009000000000",
            INIT_5F => X"0000009c00000000000000a200000000000000a3000000000000009500000000",
            INIT_60 => X"000000b400000000000000bd00000000000000c200000000000000d000000000",
            INIT_61 => X"000000d300000000000000bd000000000000009e00000000000000a200000000",
            INIT_62 => X"000000c700000000000000c200000000000000c500000000000000d300000000",
            INIT_63 => X"000000a400000000000000a300000000000000ac00000000000000bf00000000",
            INIT_64 => X"0000006d00000000000000820000000000000093000000000000009e00000000",
            INIT_65 => X"0000009100000000000000900000000000000090000000000000008900000000",
            INIT_66 => X"00000086000000000000007c0000000000000084000000000000009000000000",
            INIT_67 => X"00000093000000000000009f00000000000000a2000000000000009700000000",
            INIT_68 => X"000000b500000000000000b000000000000000b100000000000000c200000000",
            INIT_69 => X"000000cd00000000000000b3000000000000008f000000000000009f00000000",
            INIT_6A => X"000000be00000000000000c200000000000000c700000000000000d000000000",
            INIT_6B => X"000000a1000000000000009c00000000000000a500000000000000b500000000",
            INIT_6C => X"0000007200000000000000700000000000000088000000000000009500000000",
            INIT_6D => X"00000092000000000000008a0000000000000085000000000000008900000000",
            INIT_6E => X"0000009000000000000000830000000000000083000000000000009200000000",
            INIT_6F => X"0000008d00000000000000940000000000000095000000000000009600000000",
            INIT_70 => X"000000b200000000000000a5000000000000009d00000000000000ac00000000",
            INIT_71 => X"000000c7000000000000009c000000000000008500000000000000a700000000",
            INIT_72 => X"000000c200000000000000c700000000000000c700000000000000ce00000000",
            INIT_73 => X"0000008b0000000000000084000000000000008500000000000000a000000000",
            INIT_74 => X"0000007e000000000000006b000000000000007e000000000000008c00000000",
            INIT_75 => X"00000095000000000000008a0000000000000081000000000000008200000000",
            INIT_76 => X"0000008e0000000000000091000000000000008c000000000000008d00000000",
            INIT_77 => X"000000980000000000000095000000000000008c000000000000008800000000",
            INIT_78 => X"0000009b00000000000000900000000000000086000000000000009700000000",
            INIT_79 => X"000000b70000000000000082000000000000007d000000000000009e00000000",
            INIT_7A => X"000000a500000000000000b700000000000000bf00000000000000c500000000",
            INIT_7B => X"00000069000000000000005e0000000000000067000000000000008000000000",
            INIT_7C => X"0000007c00000000000000750000000000000070000000000000007700000000",
            INIT_7D => X"0000008f000000000000008b000000000000007d000000000000007900000000",
            INIT_7E => X"0000007d0000000000000081000000000000008c000000000000008b00000000",
            INIT_7F => X"00000096000000000000009b0000000000000095000000000000008400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "sampleifmap_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000100000000000000015000000000000001300000000",
            INIT_01 => X"0000008e00000000000000930000000000000093000000000000008300000000",
            INIT_02 => X"0000008e00000000000000900000000000000089000000000000008700000000",
            INIT_03 => X"0000008f000000000000008c000000000000008c000000000000008d00000000",
            INIT_04 => X"000000490000000000000060000000000000007e000000000000008c00000000",
            INIT_05 => X"000000a40000000000000082000000000000005d000000000000005f00000000",
            INIT_06 => X"0000009d000000000000009b000000000000009c000000000000009b00000000",
            INIT_07 => X"000000970000000000000098000000000000009b000000000000009e00000000",
            INIT_08 => X"0000001f00000000000000110000000000000014000000000000001400000000",
            INIT_09 => X"00000092000000000000009b00000000000000a1000000000000007a00000000",
            INIT_0A => X"00000095000000000000008b0000000000000088000000000000008a00000000",
            INIT_0B => X"0000009700000000000000920000000000000096000000000000009800000000",
            INIT_0C => X"0000004900000000000000750000000000000096000000000000009f00000000",
            INIT_0D => X"000000af000000000000009c0000000000000058000000000000004100000000",
            INIT_0E => X"000000ad00000000000000ab00000000000000a900000000000000a800000000",
            INIT_0F => X"000000a300000000000000a400000000000000a800000000000000ac00000000",
            INIT_10 => X"0000001500000000000000140000000000000014000000000000001400000000",
            INIT_11 => X"0000008c000000000000009700000000000000a2000000000000006600000000",
            INIT_12 => X"0000008b00000000000000880000000000000095000000000000008d00000000",
            INIT_13 => X"0000009f00000000000000980000000000000099000000000000009a00000000",
            INIT_14 => X"0000006d00000000000000a100000000000000ab00000000000000a600000000",
            INIT_15 => X"000000b700000000000000b10000000000000061000000000000003a00000000",
            INIT_16 => X"000000b200000000000000b100000000000000b200000000000000b300000000",
            INIT_17 => X"000000a600000000000000a900000000000000ad00000000000000b100000000",
            INIT_18 => X"0000001100000000000000150000000000000014000000000000001400000000",
            INIT_19 => X"00000082000000000000008c0000000000000099000000000000004f00000000",
            INIT_1A => X"00000087000000000000009d00000000000000a4000000000000009700000000",
            INIT_1B => X"000000b000000000000000a900000000000000a6000000000000009900000000",
            INIT_1C => X"0000007600000000000000a100000000000000af00000000000000b000000000",
            INIT_1D => X"000000c300000000000000c40000000000000085000000000000005200000000",
            INIT_1E => X"000000b300000000000000b400000000000000b700000000000000bd00000000",
            INIT_1F => X"000000ab00000000000000ad00000000000000b100000000000000b300000000",
            INIT_20 => X"0000001300000000000000150000000000000014000000000000001500000000",
            INIT_21 => X"0000007700000000000000820000000000000089000000000000003800000000",
            INIT_22 => X"0000009200000000000000b300000000000000b2000000000000009c00000000",
            INIT_23 => X"000000a70000000000000094000000000000008b000000000000008400000000",
            INIT_24 => X"00000078000000000000009800000000000000a900000000000000af00000000",
            INIT_25 => X"000000d200000000000000ce00000000000000a7000000000000006d00000000",
            INIT_26 => X"000000bf00000000000000c300000000000000c900000000000000d100000000",
            INIT_27 => X"000000ac00000000000000b100000000000000b600000000000000ba00000000",
            INIT_28 => X"0000001600000000000000170000000000000016000000000000001600000000",
            INIT_29 => X"0000007800000000000000820000000000000073000000000000002600000000",
            INIT_2A => X"0000009e00000000000000c300000000000000b9000000000000009200000000",
            INIT_2B => X"00000084000000000000006b000000000000006c000000000000007600000000",
            INIT_2C => X"000000840000000000000081000000000000008f000000000000009200000000",
            INIT_2D => X"000000c700000000000000be00000000000000b7000000000000008f00000000",
            INIT_2E => X"000000d100000000000000cc00000000000000d100000000000000cf00000000",
            INIT_2F => X"000000c200000000000000c700000000000000ca00000000000000d100000000",
            INIT_30 => X"0000001400000000000000150000000000000013000000000000001800000000",
            INIT_31 => X"0000009400000000000000a10000000000000071000000000000001e00000000",
            INIT_32 => X"000000aa00000000000000c200000000000000ba000000000000009700000000",
            INIT_33 => X"0000007100000000000000690000000000000062000000000000008000000000",
            INIT_34 => X"00000080000000000000006b0000000000000074000000000000006800000000",
            INIT_35 => X"000000c500000000000000c000000000000000ca00000000000000b200000000",
            INIT_36 => X"000000d700000000000000d100000000000000cf00000000000000ce00000000",
            INIT_37 => X"000000da00000000000000d700000000000000d600000000000000d800000000",
            INIT_38 => X"0000001d00000000000000180000000000000029000000000000005800000000",
            INIT_39 => X"0000009c00000000000000ba00000000000000ae000000000000006000000000",
            INIT_3A => X"000000ba00000000000000bd00000000000000b5000000000000009500000000",
            INIT_3B => X"000000760000000000000081000000000000008400000000000000a400000000",
            INIT_3C => X"0000007c000000000000006c000000000000006b000000000000005c00000000",
            INIT_3D => X"000000ce00000000000000bb00000000000000cc00000000000000b400000000",
            INIT_3E => X"000000e400000000000000e700000000000000e000000000000000e600000000",
            INIT_3F => X"000000e200000000000000dc00000000000000d300000000000000cd00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000075000000000000006d000000000000009900000000000000b100000000",
            INIT_41 => X"0000009300000000000000b700000000000000bd00000000000000af00000000",
            INIT_42 => X"000000c000000000000000bc00000000000000a1000000000000007800000000",
            INIT_43 => X"00000083000000000000009a00000000000000ad00000000000000b800000000",
            INIT_44 => X"0000007f00000000000000770000000000000073000000000000007300000000",
            INIT_45 => X"000000d800000000000000bc00000000000000c500000000000000a600000000",
            INIT_46 => X"000000d300000000000000e300000000000000e200000000000000e900000000",
            INIT_47 => X"000000e800000000000000e000000000000000c600000000000000bc00000000",
            INIT_48 => X"000000b600000000000000af00000000000000bc00000000000000c200000000",
            INIT_49 => X"0000009000000000000000be00000000000000c200000000000000bf00000000",
            INIT_4A => X"000000b600000000000000b10000000000000098000000000000007300000000",
            INIT_4B => X"0000008a00000000000000a400000000000000b600000000000000b700000000",
            INIT_4C => X"0000007b00000000000000770000000000000076000000000000006600000000",
            INIT_4D => X"000000e900000000000000d000000000000000bd00000000000000a000000000",
            INIT_4E => X"000000cb00000000000000ea00000000000000eb00000000000000e800000000",
            INIT_4F => X"000000eb00000000000000d100000000000000bd00000000000000bb00000000",
            INIT_50 => X"000000bb00000000000000b700000000000000c000000000000000c700000000",
            INIT_51 => X"0000008a00000000000000bf00000000000000cd00000000000000c600000000",
            INIT_52 => X"000000b500000000000000b000000000000000a5000000000000008800000000",
            INIT_53 => X"0000007c000000000000009a00000000000000af00000000000000b800000000",
            INIT_54 => X"0000007800000000000000770000000000000076000000000000006b00000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b0000000000000009e00000000",
            INIT_56 => X"000000d400000000000000f200000000000000f400000000000000f300000000",
            INIT_57 => X"000000e000000000000000c600000000000000c000000000000000c000000000",
            INIT_58 => X"000000bb00000000000000c100000000000000c900000000000000c900000000",
            INIT_59 => X"0000009200000000000000bc00000000000000d100000000000000c900000000",
            INIT_5A => X"000000b700000000000000b900000000000000b6000000000000009b00000000",
            INIT_5B => X"0000006b0000000000000084000000000000009f00000000000000b700000000",
            INIT_5C => X"0000007e000000000000007c0000000000000085000000000000007300000000",
            INIT_5D => X"000000eb00000000000000bd00000000000000aa000000000000009e00000000",
            INIT_5E => X"000000de00000000000000f200000000000000f600000000000000f600000000",
            INIT_5F => X"000000ca00000000000000c000000000000000c000000000000000c200000000",
            INIT_60 => X"000000bd00000000000000c500000000000000c900000000000000cb00000000",
            INIT_61 => X"000000a500000000000000b700000000000000c600000000000000c400000000",
            INIT_62 => X"000000a500000000000000b000000000000000aa000000000000009f00000000",
            INIT_63 => X"00000078000000000000008a00000000000000a200000000000000a400000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008500000000",
            INIT_65 => X"000000e700000000000000bd00000000000000a500000000000000a100000000",
            INIT_66 => X"000000ea00000000000000f700000000000000f800000000000000f400000000",
            INIT_67 => X"000000c700000000000000c100000000000000c300000000000000d000000000",
            INIT_68 => X"000000b900000000000000c400000000000000ca00000000000000d000000000",
            INIT_69 => X"000000b9000000000000009c00000000000000a700000000000000c100000000",
            INIT_6A => X"000000870000000000000087000000000000009100000000000000a100000000",
            INIT_6B => X"0000008f0000000000000089000000000000009e00000000000000a100000000",
            INIT_6C => X"000000a2000000000000009500000000000000a400000000000000a400000000",
            INIT_6D => X"000000e400000000000000c3000000000000009d000000000000009900000000",
            INIT_6E => X"000000f500000000000000f900000000000000f700000000000000f200000000",
            INIT_6F => X"000000de00000000000000cc00000000000000c700000000000000e800000000",
            INIT_70 => X"000000b600000000000000c500000000000000cc00000000000000d200000000",
            INIT_71 => X"000000c1000000000000007d000000000000008e00000000000000bf00000000",
            INIT_72 => X"000000a700000000000000a600000000000000b100000000000000b500000000",
            INIT_73 => X"00000072000000000000008200000000000000aa00000000000000b800000000",
            INIT_74 => X"0000009e000000000000009800000000000000aa00000000000000a500000000",
            INIT_75 => X"000000e700000000000000bd00000000000000ae00000000000000ab00000000",
            INIT_76 => X"000000fb00000000000000f500000000000000f400000000000000f200000000",
            INIT_77 => X"000000e900000000000000dd00000000000000cf00000000000000f200000000",
            INIT_78 => X"000000b900000000000000c500000000000000c800000000000000d400000000",
            INIT_79 => X"000000c00000000000000070000000000000009100000000000000bd00000000",
            INIT_7A => X"000000b400000000000000bd00000000000000be00000000000000c700000000",
            INIT_7B => X"0000008900000000000000a000000000000000a700000000000000a400000000",
            INIT_7C => X"0000009100000000000000a200000000000000b0000000000000009200000000",
            INIT_7D => X"000000c300000000000000a800000000000000b100000000000000b800000000",
            INIT_7E => X"000000f900000000000000f500000000000000f100000000000000e800000000",
            INIT_7F => X"000000eb00000000000000ec00000000000000dd00000000000000e400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "sampleifmap_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ae00000000000000b600000000000000c700000000000000d800000000",
            INIT_01 => X"000000ad000000000000006e000000000000009b00000000000000b000000000",
            INIT_02 => X"000000b200000000000000a800000000000000ba00000000000000d000000000",
            INIT_03 => X"000000a400000000000000a7000000000000009b00000000000000a800000000",
            INIT_04 => X"0000008600000000000000b10000000000000096000000000000006e00000000",
            INIT_05 => X"00000068000000000000009000000000000000ab000000000000009a00000000",
            INIT_06 => X"000000ed00000000000000ee00000000000000d1000000000000009100000000",
            INIT_07 => X"000000ed00000000000000f300000000000000dd00000000000000d200000000",
            INIT_08 => X"0000009e00000000000000a900000000000000ce00000000000000db00000000",
            INIT_09 => X"000000a2000000000000009500000000000000a700000000000000a300000000",
            INIT_0A => X"000000d100000000000000c800000000000000cd00000000000000ca00000000",
            INIT_0B => X"000000a100000000000000aa00000000000000a800000000000000bc00000000",
            INIT_0C => X"0000008700000000000000ad0000000000000078000000000000007000000000",
            INIT_0D => X"00000073000000000000009b00000000000000ba000000000000009300000000",
            INIT_0E => X"000000bc00000000000000b20000000000000084000000000000006200000000",
            INIT_0F => X"000000ef00000000000000f300000000000000d400000000000000b900000000",
            INIT_10 => X"000000a100000000000000b300000000000000d600000000000000dd00000000",
            INIT_11 => X"000000b100000000000000b300000000000000b500000000000000af00000000",
            INIT_12 => X"000000dd00000000000000d400000000000000cf00000000000000bd00000000",
            INIT_13 => X"000000ab00000000000000b800000000000000c500000000000000dc00000000",
            INIT_14 => X"0000008c00000000000000950000000000000067000000000000008b00000000",
            INIT_15 => X"00000093000000000000009400000000000000b1000000000000009700000000",
            INIT_16 => X"0000009c000000000000008a0000000000000070000000000000008300000000",
            INIT_17 => X"000000ea00000000000000d900000000000000b1000000000000009700000000",
            INIT_18 => X"000000b200000000000000c600000000000000da00000000000000df00000000",
            INIT_19 => X"000000c800000000000000be00000000000000c200000000000000c200000000",
            INIT_1A => X"000000c700000000000000bf00000000000000b800000000000000ba00000000",
            INIT_1B => X"000000b100000000000000c800000000000000d000000000000000cb00000000",
            INIT_1C => X"0000009e000000000000007f000000000000008700000000000000ab00000000",
            INIT_1D => X"0000008f0000000000000083000000000000009b00000000000000a800000000",
            INIT_1E => X"0000009f0000000000000094000000000000007e000000000000008900000000",
            INIT_1F => X"000000c5000000000000009e0000000000000090000000000000009300000000",
            INIT_20 => X"000000b700000000000000d000000000000000dd00000000000000e100000000",
            INIT_21 => X"000000c200000000000000be00000000000000c700000000000000bf00000000",
            INIT_22 => X"000000ba00000000000000be00000000000000bc00000000000000c600000000",
            INIT_23 => X"000000bf00000000000000c600000000000000c100000000000000ab00000000",
            INIT_24 => X"000000a9000000000000009400000000000000bf00000000000000cf00000000",
            INIT_25 => X"0000008d000000000000007b000000000000008700000000000000a000000000",
            INIT_26 => X"00000098000000000000009f0000000000000095000000000000008e00000000",
            INIT_27 => X"0000009a000000000000008c0000000000000088000000000000008700000000",
            INIT_28 => X"000000be00000000000000d600000000000000dd00000000000000de00000000",
            INIT_29 => X"000000be00000000000000c800000000000000c300000000000000b300000000",
            INIT_2A => X"000000b200000000000000d100000000000000cd00000000000000c600000000",
            INIT_2B => X"000000b500000000000000b600000000000000b3000000000000009700000000",
            INIT_2C => X"000000a500000000000000ae00000000000000c400000000000000c500000000",
            INIT_2D => X"000000930000000000000089000000000000007c000000000000008600000000",
            INIT_2E => X"0000008b000000000000009900000000000000a1000000000000009900000000",
            INIT_2F => X"0000007d000000000000008b000000000000008b000000000000008300000000",
            INIT_30 => X"000000c600000000000000db00000000000000da00000000000000db00000000",
            INIT_31 => X"000000cf00000000000000d200000000000000bf00000000000000aa00000000",
            INIT_32 => X"000000b400000000000000cf00000000000000ce00000000000000cb00000000",
            INIT_33 => X"000000b000000000000000b400000000000000ae000000000000009c00000000",
            INIT_34 => X"0000009600000000000000b000000000000000b500000000000000b600000000",
            INIT_35 => X"000000980000000000000096000000000000007d000000000000006f00000000",
            INIT_36 => X"0000008a000000000000009a00000000000000a1000000000000009800000000",
            INIT_37 => X"0000006a00000000000000730000000000000080000000000000008a00000000",
            INIT_38 => X"000000cf00000000000000d900000000000000d600000000000000da00000000",
            INIT_39 => X"000000d500000000000000d200000000000000bc00000000000000aa00000000",
            INIT_3A => X"000000b600000000000000c700000000000000d300000000000000d400000000",
            INIT_3B => X"000000b500000000000000ba00000000000000ba00000000000000ae00000000",
            INIT_3C => X"0000008500000000000000ab00000000000000b600000000000000ba00000000",
            INIT_3D => X"00000095000000000000009a0000000000000089000000000000007200000000",
            INIT_3E => X"00000092000000000000009f00000000000000ab000000000000009400000000",
            INIT_3F => X"000000760000000000000073000000000000007b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000d400000000000000d400000000000000d800000000",
            INIT_41 => X"000000cd00000000000000cf00000000000000bd00000000000000b300000000",
            INIT_42 => X"0000008a00000000000000b100000000000000cd00000000000000cd00000000",
            INIT_43 => X"000000b600000000000000bb00000000000000c300000000000000a700000000",
            INIT_44 => X"00000082000000000000009e00000000000000b500000000000000b900000000",
            INIT_45 => X"0000008c0000000000000096000000000000008d000000000000007d00000000",
            INIT_46 => X"00000095000000000000009d00000000000000a3000000000000008d00000000",
            INIT_47 => X"0000007c00000000000000820000000000000083000000000000008500000000",
            INIT_48 => X"000000c800000000000000d000000000000000d200000000000000d700000000",
            INIT_49 => X"000000cc00000000000000ce00000000000000be00000000000000bb00000000",
            INIT_4A => X"00000050000000000000008300000000000000c400000000000000c600000000",
            INIT_4B => X"000000ae00000000000000b800000000000000c2000000000000009100000000",
            INIT_4C => X"00000083000000000000009300000000000000a500000000000000ae00000000",
            INIT_4D => X"00000088000000000000008f000000000000008b000000000000007800000000",
            INIT_4E => X"00000088000000000000008c000000000000008e000000000000008900000000",
            INIT_4F => X"0000007000000000000000790000000000000085000000000000008500000000",
            INIT_50 => X"000000c200000000000000cd00000000000000d000000000000000d700000000",
            INIT_51 => X"000000d100000000000000cd00000000000000b700000000000000b500000000",
            INIT_52 => X"00000051000000000000008100000000000000c200000000000000cc00000000",
            INIT_53 => X"000000a100000000000000ab00000000000000ba000000000000008e00000000",
            INIT_54 => X"000000780000000000000089000000000000009500000000000000a100000000",
            INIT_55 => X"0000007e00000000000000890000000000000087000000000000007300000000",
            INIT_56 => X"0000007a0000000000000070000000000000007b000000000000008500000000",
            INIT_57 => X"0000008000000000000000830000000000000088000000000000008a00000000",
            INIT_58 => X"000000bc00000000000000c800000000000000cd00000000000000d600000000",
            INIT_59 => X"000000d400000000000000c600000000000000af00000000000000b000000000",
            INIT_5A => X"0000008e00000000000000a000000000000000c000000000000000d000000000",
            INIT_5B => X"00000095000000000000009b00000000000000a800000000000000aa00000000",
            INIT_5C => X"00000064000000000000007f0000000000000085000000000000008d00000000",
            INIT_5D => X"0000007b00000000000000800000000000000083000000000000007100000000",
            INIT_5E => X"00000072000000000000006c0000000000000072000000000000007e00000000",
            INIT_5F => X"0000008900000000000000900000000000000090000000000000008200000000",
            INIT_60 => X"000000b700000000000000c000000000000000c400000000000000d200000000",
            INIT_61 => X"000000d200000000000000c000000000000000a600000000000000a900000000",
            INIT_62 => X"000000b400000000000000b600000000000000c000000000000000d100000000",
            INIT_63 => X"0000008c000000000000008d000000000000009900000000000000ab00000000",
            INIT_64 => X"0000005c000000000000006f000000000000007d000000000000008600000000",
            INIT_65 => X"0000007f000000000000007e000000000000007e000000000000007800000000",
            INIT_66 => X"0000007400000000000000690000000000000072000000000000007e00000000",
            INIT_67 => X"00000081000000000000008d0000000000000090000000000000008500000000",
            INIT_68 => X"000000b900000000000000b300000000000000b300000000000000c400000000",
            INIT_69 => X"000000cc00000000000000b5000000000000009700000000000000a600000000",
            INIT_6A => X"000000b300000000000000ba00000000000000c200000000000000cd00000000",
            INIT_6B => X"000000880000000000000085000000000000009200000000000000a600000000",
            INIT_6C => X"00000061000000000000005d0000000000000072000000000000007e00000000",
            INIT_6D => X"0000008000000000000000780000000000000073000000000000007800000000",
            INIT_6E => X"0000007e00000000000000710000000000000071000000000000008000000000",
            INIT_6F => X"0000007b00000000000000820000000000000083000000000000008400000000",
            INIT_70 => X"000000b800000000000000aa00000000000000a100000000000000b100000000",
            INIT_71 => X"000000c3000000000000009c000000000000008c00000000000000ae00000000",
            INIT_72 => X"000000b600000000000000bf00000000000000c100000000000000c900000000",
            INIT_73 => X"00000073000000000000006c0000000000000071000000000000009100000000",
            INIT_74 => X"0000006e0000000000000059000000000000006a000000000000007600000000",
            INIT_75 => X"0000008300000000000000780000000000000070000000000000007200000000",
            INIT_76 => X"0000007c000000000000007f000000000000007a000000000000007b00000000",
            INIT_77 => X"000000860000000000000082000000000000007a000000000000007500000000",
            INIT_78 => X"000000a10000000000000097000000000000008c000000000000009d00000000",
            INIT_79 => X"000000b10000000000000080000000000000008200000000000000a600000000",
            INIT_7A => X"0000009a00000000000000af00000000000000b700000000000000bf00000000",
            INIT_7B => X"0000005300000000000000470000000000000053000000000000007000000000",
            INIT_7C => X"0000006e0000000000000065000000000000005e000000000000006300000000",
            INIT_7D => X"0000007e0000000000000079000000000000006c000000000000006c00000000",
            INIT_7E => X"0000006b000000000000006f000000000000007a000000000000007900000000",
            INIT_7F => X"0000008400000000000000890000000000000084000000000000007300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "sampleifmap_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000280000000000000013000000000000001c000000000000001700000000",
            INIT_01 => X"00000074000000000000006d0000000000000073000000000000007100000000",
            INIT_02 => X"00000069000000000000006a0000000000000067000000000000007100000000",
            INIT_03 => X"0000006b00000000000000690000000000000069000000000000006900000000",
            INIT_04 => X"0000003a000000000000004c0000000000000063000000000000006a00000000",
            INIT_05 => X"0000008900000000000000720000000000000056000000000000005400000000",
            INIT_06 => X"0000007d000000000000007c000000000000007d000000000000007c00000000",
            INIT_07 => X"00000078000000000000007a000000000000007d000000000000007f00000000",
            INIT_08 => X"0000001a0000000000000014000000000000001b000000000000001800000000",
            INIT_09 => X"0000007c00000000000000760000000000000082000000000000006a00000000",
            INIT_0A => X"00000075000000000000006d0000000000000072000000000000007d00000000",
            INIT_0B => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_0C => X"00000044000000000000006a0000000000000083000000000000008500000000",
            INIT_0D => X"00000096000000000000008c0000000000000051000000000000003e00000000",
            INIT_0E => X"000000880000000000000089000000000000008c000000000000008a00000000",
            INIT_0F => X"0000008000000000000000810000000000000085000000000000008800000000",
            INIT_10 => X"000000120000000000000017000000000000001a000000000000001800000000",
            INIT_11 => X"0000007b00000000000000740000000000000083000000000000005800000000",
            INIT_12 => X"000000740000000000000074000000000000008d000000000000008b00000000",
            INIT_13 => X"00000084000000000000007d000000000000007f000000000000008100000000",
            INIT_14 => X"000000690000000000000098000000000000009a000000000000008e00000000",
            INIT_15 => X"0000009e000000000000009f0000000000000059000000000000003700000000",
            INIT_16 => X"0000008e00000000000000920000000000000097000000000000009700000000",
            INIT_17 => X"000000840000000000000088000000000000008b000000000000008e00000000",
            INIT_18 => X"0000001200000000000000190000000000000019000000000000001800000000",
            INIT_19 => X"00000073000000000000006a000000000000007c000000000000004500000000",
            INIT_1A => X"00000078000000000000009200000000000000a6000000000000009c00000000",
            INIT_1B => X"0000009700000000000000950000000000000094000000000000008900000000",
            INIT_1C => X"0000006d0000000000000094000000000000009c000000000000009600000000",
            INIT_1D => X"000000a900000000000000b1000000000000007a000000000000004a00000000",
            INIT_1E => X"000000950000000000000098000000000000009d00000000000000a100000000",
            INIT_1F => X"0000008e00000000000000910000000000000094000000000000009600000000",
            INIT_20 => X"0000001700000000000000190000000000000018000000000000001900000000",
            INIT_21 => X"000000680000000000000060000000000000006d000000000000003300000000",
            INIT_22 => X"0000008d00000000000000b200000000000000b800000000000000a100000000",
            INIT_23 => X"0000009300000000000000860000000000000080000000000000007c00000000",
            INIT_24 => X"0000006c00000000000000890000000000000096000000000000009700000000",
            INIT_25 => X"000000b500000000000000b70000000000000098000000000000006000000000",
            INIT_26 => X"000000a400000000000000a800000000000000ae00000000000000b300000000",
            INIT_27 => X"000000930000000000000098000000000000009c00000000000000a000000000",
            INIT_28 => X"0000001c000000000000001b000000000000001a000000000000001a00000000",
            INIT_29 => X"00000066000000000000005f0000000000000059000000000000002300000000",
            INIT_2A => X"0000009f00000000000000c700000000000000c1000000000000009600000000",
            INIT_2B => X"0000007600000000000000620000000000000066000000000000007400000000",
            INIT_2C => X"0000007a00000000000000770000000000000083000000000000008200000000",
            INIT_2D => X"000000aa00000000000000a600000000000000a7000000000000008400000000",
            INIT_2E => X"000000b700000000000000b300000000000000b700000000000000b200000000",
            INIT_2F => X"000000a900000000000000af00000000000000b100000000000000b700000000",
            INIT_30 => X"0000001a00000000000000190000000000000016000000000000001a00000000",
            INIT_31 => X"0000007b0000000000000080000000000000005c000000000000001d00000000",
            INIT_32 => X"000000ab00000000000000c700000000000000c3000000000000009300000000",
            INIT_33 => X"0000006a0000000000000063000000000000005e000000000000007e00000000",
            INIT_34 => X"0000007a0000000000000065000000000000006d000000000000006000000000",
            INIT_35 => X"000000b000000000000000aa00000000000000c000000000000000ac00000000",
            INIT_36 => X"000000ca00000000000000c500000000000000c400000000000000c300000000",
            INIT_37 => X"000000c200000000000000bf00000000000000bf00000000000000c500000000",
            INIT_38 => X"0000001900000000000000110000000000000021000000000000004d00000000",
            INIT_39 => X"0000007e000000000000009b000000000000009a000000000000005800000000",
            INIT_3A => X"000000b900000000000000c100000000000000be000000000000008c00000000",
            INIT_3B => X"00000071000000000000007b000000000000008100000000000000a300000000",
            INIT_3C => X"0000007900000000000000680000000000000067000000000000005800000000",
            INIT_3D => X"000000bd00000000000000a500000000000000c600000000000000b100000000",
            INIT_3E => X"000000da00000000000000e000000000000000db00000000000000e400000000",
            INIT_3F => X"000000cd00000000000000c400000000000000bb00000000000000ba00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006000000000000000560000000000000080000000000000009500000000",
            INIT_41 => X"00000077000000000000009900000000000000a7000000000000009b00000000",
            INIT_42 => X"000000bf00000000000000bf00000000000000a8000000000000006f00000000",
            INIT_43 => X"0000007f000000000000009400000000000000aa00000000000000b700000000",
            INIT_44 => X"0000007c00000000000000740000000000000070000000000000007000000000",
            INIT_45 => X"000000c100000000000000a200000000000000bb00000000000000a300000000",
            INIT_46 => X"000000bb00000000000000cf00000000000000d500000000000000df00000000",
            INIT_47 => X"000000d200000000000000c400000000000000a6000000000000009d00000000",
            INIT_48 => X"0000009b0000000000000092000000000000009e00000000000000a100000000",
            INIT_49 => X"00000075000000000000009f00000000000000a900000000000000a700000000",
            INIT_4A => X"000000b500000000000000b3000000000000009b000000000000006800000000",
            INIT_4B => X"00000087000000000000009f00000000000000b400000000000000b600000000",
            INIT_4C => X"0000007900000000000000750000000000000074000000000000006400000000",
            INIT_4D => X"000000cc00000000000000b200000000000000b2000000000000009e00000000",
            INIT_4E => X"000000a700000000000000cb00000000000000d600000000000000d800000000",
            INIT_4F => X"000000cf00000000000000b00000000000000096000000000000009300000000",
            INIT_50 => X"000000a5000000000000009e00000000000000a500000000000000aa00000000",
            INIT_51 => X"0000007000000000000000a000000000000000b000000000000000af00000000",
            INIT_52 => X"000000b400000000000000b100000000000000a4000000000000007b00000000",
            INIT_53 => X"00000079000000000000009500000000000000ac00000000000000b600000000",
            INIT_54 => X"0000007600000000000000750000000000000074000000000000006a00000000",
            INIT_55 => X"000000d100000000000000af00000000000000a6000000000000009c00000000",
            INIT_56 => X"000000a900000000000000cd00000000000000d800000000000000de00000000",
            INIT_57 => X"000000ba000000000000009f0000000000000093000000000000009100000000",
            INIT_58 => X"000000a600000000000000a900000000000000ae00000000000000ac00000000",
            INIT_59 => X"0000007a000000000000009d00000000000000b000000000000000b000000000",
            INIT_5A => X"000000b600000000000000b900000000000000b1000000000000008d00000000",
            INIT_5B => X"00000068000000000000007f000000000000009d00000000000000b600000000",
            INIT_5C => X"0000007d000000000000007b0000000000000084000000000000007300000000",
            INIT_5D => X"000000ce00000000000000a300000000000000a4000000000000009f00000000",
            INIT_5E => X"000000b500000000000000cd00000000000000d900000000000000e000000000",
            INIT_5F => X"0000009c0000000000000093000000000000008e000000000000009200000000",
            INIT_60 => X"000000a000000000000000a500000000000000a700000000000000a700000000",
            INIT_61 => X"0000008f000000000000009900000000000000a400000000000000a500000000",
            INIT_62 => X"000000a400000000000000ae00000000000000a3000000000000009100000000",
            INIT_63 => X"000000760000000000000085000000000000009f00000000000000a300000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008600000000",
            INIT_65 => X"000000cd00000000000000a800000000000000a300000000000000a300000000",
            INIT_66 => X"000000c700000000000000d600000000000000dc00000000000000df00000000",
            INIT_67 => X"000000980000000000000090000000000000009000000000000000a300000000",
            INIT_68 => X"0000009b00000000000000a000000000000000a200000000000000a900000000",
            INIT_69 => X"000000a40000000000000083000000000000008800000000000000a300000000",
            INIT_6A => X"0000008500000000000000840000000000000088000000000000009200000000",
            INIT_6B => X"000000920000000000000087000000000000009e000000000000009f00000000",
            INIT_6C => X"0000009e000000000000009000000000000000a200000000000000a700000000",
            INIT_6D => X"000000cb00000000000000b00000000000000098000000000000009800000000",
            INIT_6E => X"000000da00000000000000dd00000000000000d800000000000000d700000000",
            INIT_6F => X"000000b600000000000000a2000000000000009f00000000000000c500000000",
            INIT_70 => X"0000009d00000000000000a200000000000000a400000000000000ae00000000",
            INIT_71 => X"000000b2000000000000006d000000000000007800000000000000a800000000",
            INIT_72 => X"000000a300000000000000a100000000000000a700000000000000a600000000",
            INIT_73 => X"00000078000000000000008400000000000000ab00000000000000b600000000",
            INIT_74 => X"00000095000000000000008c00000000000000a300000000000000a900000000",
            INIT_75 => X"000000cc00000000000000aa00000000000000a400000000000000a600000000",
            INIT_76 => X"000000e400000000000000da00000000000000d500000000000000d300000000",
            INIT_77 => X"000000c700000000000000bb00000000000000b000000000000000d600000000",
            INIT_78 => X"0000009f00000000000000a100000000000000a000000000000000af00000000",
            INIT_79 => X"000000b70000000000000068000000000000008400000000000000aa00000000",
            INIT_7A => X"000000b000000000000000b800000000000000b600000000000000bc00000000",
            INIT_7B => X"0000008d00000000000000a300000000000000a800000000000000a200000000",
            INIT_7C => X"00000085000000000000009200000000000000a5000000000000009100000000",
            INIT_7D => X"000000a9000000000000009600000000000000a500000000000000af00000000",
            INIT_7E => X"000000dd00000000000000d900000000000000d400000000000000ca00000000",
            INIT_7F => X"000000c700000000000000c700000000000000ba00000000000000c400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "sampleifmap_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000940000000000000092000000000000009f00000000000000b300000000",
            INIT_01 => X"000000a8000000000000006d000000000000009700000000000000a100000000",
            INIT_02 => X"000000ae00000000000000a400000000000000b500000000000000c700000000",
            INIT_03 => X"000000a600000000000000aa000000000000009c00000000000000a500000000",
            INIT_04 => X"00000077000000000000009f0000000000000088000000000000006900000000",
            INIT_05 => X"00000050000000000000007e000000000000009e000000000000008f00000000",
            INIT_06 => X"000000cd00000000000000d100000000000000b7000000000000007600000000",
            INIT_07 => X"000000c500000000000000c900000000000000b700000000000000af00000000",
            INIT_08 => X"00000083000000000000008500000000000000a400000000000000b500000000",
            INIT_09 => X"0000009f000000000000009700000000000000a5000000000000009500000000",
            INIT_0A => X"000000cd00000000000000c400000000000000c700000000000000c200000000",
            INIT_0B => X"000000a200000000000000ac00000000000000a800000000000000b900000000",
            INIT_0C => X"00000077000000000000009b0000000000000069000000000000006800000000",
            INIT_0D => X"0000005c000000000000008800000000000000ad000000000000008600000000",
            INIT_0E => X"0000009e0000000000000098000000000000006f000000000000004b00000000",
            INIT_0F => X"000000c800000000000000cb00000000000000b0000000000000009800000000",
            INIT_10 => X"00000085000000000000008e00000000000000ac00000000000000b700000000",
            INIT_11 => X"000000aa00000000000000b100000000000000b0000000000000009f00000000",
            INIT_12 => X"000000d900000000000000cf00000000000000c500000000000000b100000000",
            INIT_13 => X"000000aa00000000000000bb00000000000000c600000000000000d900000000",
            INIT_14 => X"0000007e0000000000000085000000000000005a000000000000008300000000",
            INIT_15 => X"0000007e000000000000008200000000000000a2000000000000008b00000000",
            INIT_16 => X"0000008400000000000000760000000000000060000000000000006f00000000",
            INIT_17 => X"000000c700000000000000b80000000000000092000000000000007c00000000",
            INIT_18 => X"0000009500000000000000a100000000000000b000000000000000b900000000",
            INIT_19 => X"000000bc00000000000000b600000000000000b700000000000000af00000000",
            INIT_1A => X"000000c200000000000000b900000000000000aa00000000000000aa00000000",
            INIT_1B => X"000000af00000000000000ca00000000000000d000000000000000c900000000",
            INIT_1C => X"000000910000000000000071000000000000007b00000000000000a400000000",
            INIT_1D => X"0000007b0000000000000071000000000000008c000000000000009d00000000",
            INIT_1E => X"0000008e00000000000000860000000000000070000000000000007700000000",
            INIT_1F => X"000000a600000000000000840000000000000079000000000000007f00000000",
            INIT_20 => X"0000009b00000000000000ad00000000000000b700000000000000bd00000000",
            INIT_21 => X"000000b200000000000000b100000000000000ba00000000000000ab00000000",
            INIT_22 => X"000000b100000000000000b200000000000000ac00000000000000b400000000",
            INIT_23 => X"000000bd00000000000000c300000000000000bc00000000000000a400000000",
            INIT_24 => X"0000009d000000000000008800000000000000b600000000000000c900000000",
            INIT_25 => X"0000007c000000000000006a0000000000000078000000000000009300000000",
            INIT_26 => X"0000008a0000000000000094000000000000008a000000000000008000000000",
            INIT_27 => X"00000082000000000000007a0000000000000077000000000000007800000000",
            INIT_28 => X"000000a100000000000000b700000000000000bc00000000000000bd00000000",
            INIT_29 => X"000000b000000000000000bb00000000000000b7000000000000009e00000000",
            INIT_2A => X"000000a400000000000000c000000000000000bf00000000000000b800000000",
            INIT_2B => X"000000b100000000000000ad00000000000000a6000000000000008b00000000",
            INIT_2C => X"0000009600000000000000a200000000000000bc00000000000000c000000000",
            INIT_2D => X"000000850000000000000079000000000000006b000000000000007600000000",
            INIT_2E => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_2F => X"0000006c000000000000007d000000000000007c000000000000007500000000",
            INIT_30 => X"000000a600000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_31 => X"000000c500000000000000c700000000000000b4000000000000009400000000",
            INIT_32 => X"000000a800000000000000c000000000000000c300000000000000c100000000",
            INIT_33 => X"000000aa00000000000000a9000000000000009f000000000000009100000000",
            INIT_34 => X"0000008600000000000000a300000000000000ac00000000000000af00000000",
            INIT_35 => X"0000008b0000000000000086000000000000006c000000000000005d00000000",
            INIT_36 => X"0000007c000000000000008e0000000000000097000000000000008d00000000",
            INIT_37 => X"0000005b00000000000000650000000000000072000000000000007c00000000",
            INIT_38 => X"000000ac00000000000000b700000000000000b500000000000000ba00000000",
            INIT_39 => X"000000cf00000000000000c900000000000000b0000000000000008f00000000",
            INIT_3A => X"000000af00000000000000bd00000000000000cb00000000000000ce00000000",
            INIT_3B => X"000000ac00000000000000ae00000000000000ab00000000000000a500000000",
            INIT_3C => X"00000075000000000000009e00000000000000ab00000000000000b200000000",
            INIT_3D => X"00000088000000000000008a0000000000000078000000000000006100000000",
            INIT_3E => X"00000084000000000000009200000000000000a1000000000000008a00000000",
            INIT_3F => X"000000680000000000000064000000000000006d000000000000008200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a900000000000000af00000000000000b200000000000000b800000000",
            INIT_41 => X"000000ca00000000000000c600000000000000aa000000000000009200000000",
            INIT_42 => X"0000008800000000000000ab00000000000000c500000000000000c800000000",
            INIT_43 => X"000000aa00000000000000ab00000000000000b400000000000000a100000000",
            INIT_44 => X"00000073000000000000009000000000000000a800000000000000ad00000000",
            INIT_45 => X"0000007e0000000000000086000000000000007c000000000000006c00000000",
            INIT_46 => X"0000008700000000000000910000000000000099000000000000008200000000",
            INIT_47 => X"0000006f00000000000000740000000000000075000000000000007700000000",
            INIT_48 => X"0000009d00000000000000a800000000000000b000000000000000b800000000",
            INIT_49 => X"000000c800000000000000c000000000000000a2000000000000009300000000",
            INIT_4A => X"00000052000000000000008100000000000000b900000000000000bf00000000",
            INIT_4B => X"0000009f00000000000000a600000000000000b3000000000000008d00000000",
            INIT_4C => X"0000007400000000000000840000000000000096000000000000009f00000000",
            INIT_4D => X"0000007a000000000000007f000000000000007a000000000000006900000000",
            INIT_4E => X"0000007a00000000000000800000000000000084000000000000007f00000000",
            INIT_4F => X"00000062000000000000006b0000000000000077000000000000007700000000",
            INIT_50 => X"0000009400000000000000a300000000000000ac00000000000000b800000000",
            INIT_51 => X"000000ca00000000000000ba0000000000000092000000000000008600000000",
            INIT_52 => X"00000058000000000000008200000000000000b200000000000000c000000000",
            INIT_53 => X"00000090000000000000009800000000000000ac000000000000008c00000000",
            INIT_54 => X"00000069000000000000007a0000000000000084000000000000009100000000",
            INIT_55 => X"0000007000000000000000790000000000000077000000000000006400000000",
            INIT_56 => X"0000006c00000000000000640000000000000071000000000000007a00000000",
            INIT_57 => X"000000720000000000000075000000000000007a000000000000007c00000000",
            INIT_58 => X"0000008e000000000000009e00000000000000a900000000000000b700000000",
            INIT_59 => X"000000cc00000000000000b20000000000000084000000000000007e00000000",
            INIT_5A => X"00000090000000000000009d00000000000000af00000000000000c300000000",
            INIT_5B => X"000000830000000000000087000000000000009800000000000000a400000000",
            INIT_5C => X"00000054000000000000006f0000000000000074000000000000007c00000000",
            INIT_5D => X"0000006d00000000000000710000000000000073000000000000006100000000",
            INIT_5E => X"00000064000000000000005f0000000000000066000000000000007200000000",
            INIT_5F => X"0000007b00000000000000820000000000000082000000000000007400000000",
            INIT_60 => X"0000008e000000000000009900000000000000a100000000000000b100000000",
            INIT_61 => X"000000cc00000000000000b2000000000000007a000000000000007700000000",
            INIT_62 => X"000000a800000000000000aa00000000000000b400000000000000c500000000",
            INIT_63 => X"0000007b000000000000007a0000000000000087000000000000009d00000000",
            INIT_64 => X"0000004b000000000000005e000000000000006d000000000000007700000000",
            INIT_65 => X"000000710000000000000070000000000000006f000000000000006800000000",
            INIT_66 => X"00000066000000000000005c0000000000000064000000000000007000000000",
            INIT_67 => X"00000073000000000000007e0000000000000082000000000000007700000000",
            INIT_68 => X"00000091000000000000008d000000000000009000000000000000a300000000",
            INIT_69 => X"000000c800000000000000a9000000000000006b000000000000007400000000",
            INIT_6A => X"000000a300000000000000ac00000000000000b700000000000000c200000000",
            INIT_6B => X"0000007900000000000000730000000000000081000000000000009600000000",
            INIT_6C => X"00000051000000000000004e0000000000000064000000000000007000000000",
            INIT_6D => X"00000072000000000000006a0000000000000065000000000000006800000000",
            INIT_6E => X"0000007000000000000000630000000000000063000000000000007200000000",
            INIT_6F => X"0000006e00000000000000740000000000000075000000000000007600000000",
            INIT_70 => X"0000008f0000000000000083000000000000007e000000000000008e00000000",
            INIT_71 => X"000000c00000000000000091000000000000005f000000000000007c00000000",
            INIT_72 => X"000000a800000000000000b200000000000000b700000000000000be00000000",
            INIT_73 => X"00000065000000000000005c0000000000000062000000000000008200000000",
            INIT_74 => X"0000005f000000000000004b000000000000005c000000000000006800000000",
            INIT_75 => X"00000074000000000000006a0000000000000061000000000000006300000000",
            INIT_76 => X"0000006e0000000000000071000000000000006c000000000000006d00000000",
            INIT_77 => X"000000770000000000000074000000000000006c000000000000006700000000",
            INIT_78 => X"0000007800000000000000700000000000000068000000000000007b00000000",
            INIT_79 => X"000000ae00000000000000760000000000000057000000000000007400000000",
            INIT_7A => X"0000008d00000000000000a400000000000000ae00000000000000b500000000",
            INIT_7B => X"0000004600000000000000390000000000000045000000000000006300000000",
            INIT_7C => X"0000006000000000000000580000000000000051000000000000005700000000",
            INIT_7D => X"00000070000000000000006b000000000000005e000000000000005d00000000",
            INIT_7E => X"0000005d0000000000000061000000000000006c000000000000006b00000000",
            INIT_7F => X"00000076000000000000007b0000000000000076000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "sampleifmap_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c700000000000000cd00000000000000d200000000000000d900000000",
            INIT_01 => X"000000bd00000000000000cf00000000000000d600000000000000da00000000",
            INIT_02 => X"000000a900000000000000a600000000000000ae00000000000000bb00000000",
            INIT_03 => X"0000008f000000000000008c000000000000009a000000000000009600000000",
            INIT_04 => X"000000df00000000000000db00000000000000bf00000000000000a700000000",
            INIT_05 => X"000000e100000000000000e200000000000000d700000000000000db00000000",
            INIT_06 => X"000000bb00000000000000af00000000000000be00000000000000db00000000",
            INIT_07 => X"000000a200000000000000a100000000000000aa00000000000000c800000000",
            INIT_08 => X"000000d700000000000000dc00000000000000dd00000000000000de00000000",
            INIT_09 => X"000000b300000000000000d300000000000000e100000000000000d800000000",
            INIT_0A => X"000000bc00000000000000be00000000000000c000000000000000b400000000",
            INIT_0B => X"000000db00000000000000d100000000000000ce00000000000000c700000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000eb00000000000000e500000000",
            INIT_0D => X"000000e500000000000000e100000000000000e200000000000000e900000000",
            INIT_0E => X"000000cd00000000000000d000000000000000d400000000000000e700000000",
            INIT_0F => X"000000c800000000000000ba00000000000000b700000000000000d800000000",
            INIT_10 => X"000000e800000000000000e700000000000000e900000000000000ea00000000",
            INIT_11 => X"000000ad00000000000000d900000000000000ef00000000000000e900000000",
            INIT_12 => X"000000b700000000000000ad00000000000000b400000000000000a400000000",
            INIT_13 => X"000000e000000000000000d400000000000000bc00000000000000be00000000",
            INIT_14 => X"000000e100000000000000e300000000000000eb00000000000000da00000000",
            INIT_15 => X"000000e100000000000000d600000000000000df00000000000000e500000000",
            INIT_16 => X"000000d800000000000000e600000000000000e800000000000000ea00000000",
            INIT_17 => X"000000d300000000000000d000000000000000ca00000000000000d100000000",
            INIT_18 => X"000000f200000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009e00000000000000e400000000000000f300000000000000f400000000",
            INIT_1A => X"0000009f0000000000000083000000000000009d000000000000009200000000",
            INIT_1B => X"0000009f00000000000000a20000000000000088000000000000009100000000",
            INIT_1C => X"000000d300000000000000c300000000000000cb00000000000000a900000000",
            INIT_1D => X"000000e200000000000000d000000000000000cb00000000000000d100000000",
            INIT_1E => X"000000d500000000000000e400000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e000000000000000db00000000000000c700000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000007500000000000000cf00000000000000f100000000000000f500000000",
            INIT_22 => X"0000006b0000000000000059000000000000006c000000000000006300000000",
            INIT_23 => X"0000005c0000000000000064000000000000005b000000000000006400000000",
            INIT_24 => X"00000095000000000000007c000000000000007c000000000000006600000000",
            INIT_25 => X"000000e900000000000000ca00000000000000b900000000000000b600000000",
            INIT_26 => X"000000cd00000000000000e300000000000000e200000000000000e100000000",
            INIT_27 => X"000000de00000000000000e200000000000000d500000000000000c200000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007e00000000000000d800000000000000ed00000000000000f500000000",
            INIT_2A => X"00000066000000000000005b000000000000005a000000000000004800000000",
            INIT_2B => X"00000063000000000000006b0000000000000067000000000000006500000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005900000000",
            INIT_2D => X"000000eb00000000000000d800000000000000be000000000000007e00000000",
            INIT_2E => X"000000c400000000000000d800000000000000df00000000000000e700000000",
            INIT_2F => X"000000ec00000000000000d900000000000000bd00000000000000ae00000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009e00000000000000d900000000000000db00000000000000f100000000",
            INIT_32 => X"0000009700000000000000840000000000000072000000000000005000000000",
            INIT_33 => X"0000008a000000000000008f0000000000000084000000000000008c00000000",
            INIT_34 => X"000000780000000000000072000000000000007a000000000000008200000000",
            INIT_35 => X"000000e900000000000000dd000000000000009b000000000000006e00000000",
            INIT_36 => X"000000c000000000000000c600000000000000e000000000000000eb00000000",
            INIT_37 => X"000000eb00000000000000cc00000000000000ab00000000000000a700000000",
            INIT_38 => X"000000f600000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009900000000000000d700000000000000c700000000000000e300000000",
            INIT_3A => X"000000ca00000000000000bb0000000000000092000000000000005100000000",
            INIT_3B => X"000000830000000000000083000000000000009e00000000000000cf00000000",
            INIT_3C => X"000000840000000000000083000000000000008d000000000000008100000000",
            INIT_3D => X"000000d7000000000000009f0000000000000084000000000000009f00000000",
            INIT_3E => X"000000d100000000000000d400000000000000d700000000000000e500000000",
            INIT_3F => X"000000dd00000000000000b200000000000000ab00000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000008200000000000000da00000000000000ce00000000000000e300000000",
            INIT_42 => X"0000008100000000000000800000000000000082000000000000005100000000",
            INIT_43 => X"0000007d0000000000000074000000000000009100000000000000b800000000",
            INIT_44 => X"0000007d000000000000008e0000000000000089000000000000007c00000000",
            INIT_45 => X"000000c600000000000000900000000000000093000000000000009900000000",
            INIT_46 => X"000000dc00000000000000e900000000000000db00000000000000d600000000",
            INIT_47 => X"000000c900000000000000a900000000000000a400000000000000b800000000",
            INIT_48 => X"000000f200000000000000f400000000000000f300000000000000f300000000",
            INIT_49 => X"0000006e00000000000000a800000000000000be00000000000000e400000000",
            INIT_4A => X"0000006e00000000000000770000000000000086000000000000005300000000",
            INIT_4B => X"0000007800000000000000730000000000000080000000000000008f00000000",
            INIT_4C => X"0000007d00000000000000920000000000000083000000000000007d00000000",
            INIT_4D => X"000000c4000000000000008c000000000000009b000000000000009500000000",
            INIT_4E => X"000000e900000000000000f000000000000000f000000000000000e900000000",
            INIT_4F => X"000000dc00000000000000d700000000000000c800000000000000c800000000",
            INIT_50 => X"000000f500000000000000f400000000000000f100000000000000ef00000000",
            INIT_51 => X"0000005f0000000000000082000000000000008500000000000000dc00000000",
            INIT_52 => X"0000006c00000000000000740000000000000074000000000000004e00000000",
            INIT_53 => X"0000006c000000000000006d000000000000006b000000000000006d00000000",
            INIT_54 => X"0000007300000000000000780000000000000078000000000000007300000000",
            INIT_55 => X"000000a7000000000000008f0000000000000096000000000000008800000000",
            INIT_56 => X"000000f300000000000000f500000000000000e400000000000000d000000000",
            INIT_57 => X"000000f400000000000000f500000000000000f500000000000000f400000000",
            INIT_58 => X"000000f400000000000000f200000000000000e900000000000000de00000000",
            INIT_59 => X"0000005900000000000000a500000000000000a900000000000000d800000000",
            INIT_5A => X"00000064000000000000005b0000000000000043000000000000003d00000000",
            INIT_5B => X"000000600000000000000062000000000000005f000000000000005f00000000",
            INIT_5C => X"00000061000000000000005a000000000000005f000000000000006000000000",
            INIT_5D => X"0000007e00000000000000810000000000000079000000000000006900000000",
            INIT_5E => X"000000f300000000000000f800000000000000d8000000000000009b00000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e300000000000000ec00000000000000df00000000000000d000000000",
            INIT_61 => X"0000006400000000000000b500000000000000b700000000000000bf00000000",
            INIT_62 => X"0000006500000000000000580000000000000038000000000000003700000000",
            INIT_63 => X"0000005400000000000000560000000000000063000000000000006f00000000",
            INIT_64 => X"00000071000000000000005d0000000000000054000000000000005200000000",
            INIT_65 => X"0000008100000000000000700000000000000062000000000000006d00000000",
            INIT_66 => X"000000f400000000000000f500000000000000e200000000000000ae00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c300000000000000db00000000000000cc00000000000000c800000000",
            INIT_69 => X"00000066000000000000009c000000000000009a00000000000000aa00000000",
            INIT_6A => X"00000066000000000000006c0000000000000063000000000000006800000000",
            INIT_6B => X"00000055000000000000005e0000000000000075000000000000007300000000",
            INIT_6C => X"0000008c000000000000007a000000000000006a000000000000005a00000000",
            INIT_6D => X"0000007c000000000000006c0000000000000068000000000000008000000000",
            INIT_6E => X"000000d400000000000000c300000000000000b3000000000000009600000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a900000000000000cf00000000000000d200000000000000c800000000",
            INIT_71 => X"0000008a0000000000000093000000000000009400000000000000a400000000",
            INIT_72 => X"0000005d000000000000006a000000000000005c000000000000008100000000",
            INIT_73 => X"0000004d0000000000000054000000000000005d000000000000005900000000",
            INIT_74 => X"0000005100000000000000510000000000000051000000000000004c00000000",
            INIT_75 => X"00000052000000000000004b000000000000004a000000000000004f00000000",
            INIT_76 => X"0000008f000000000000008c000000000000007b000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bf00000000",
            INIT_78 => X"0000007700000000000000c400000000000000e200000000000000d200000000",
            INIT_79 => X"000000c000000000000000ba0000000000000096000000000000007000000000",
            INIT_7A => X"00000037000000000000004d000000000000004d000000000000006c00000000",
            INIT_7B => X"0000003f000000000000003c000000000000002f000000000000002d00000000",
            INIT_7C => X"00000036000000000000003b000000000000003f000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000032000000000000003100000000",
            INIT_7E => X"00000067000000000000005b000000000000004b000000000000004700000000",
            INIT_7F => X"000000f400000000000000f600000000000000e1000000000000008700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "sampleifmap_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006000000000000000b400000000000000c100000000000000c700000000",
            INIT_01 => X"000000a100000000000000c00000000000000091000000000000005d00000000",
            INIT_02 => X"00000062000000000000005c0000000000000049000000000000005600000000",
            INIT_03 => X"00000047000000000000004f000000000000004f000000000000006800000000",
            INIT_04 => X"0000001b000000000000001e000000000000001c000000000000002500000000",
            INIT_05 => X"0000001c00000000000000160000000000000032000000000000003400000000",
            INIT_06 => X"00000068000000000000005b0000000000000035000000000000001800000000",
            INIT_07 => X"000000f300000000000000f700000000000000ce000000000000008000000000",
            INIT_08 => X"0000007100000000000000c200000000000000c700000000000000d300000000",
            INIT_09 => X"00000047000000000000009f000000000000009d000000000000007800000000",
            INIT_0A => X"0000007c0000000000000074000000000000005a000000000000004400000000",
            INIT_0B => X"0000006600000000000000800000000000000079000000000000009500000000",
            INIT_0C => X"0000006400000000000000700000000000000062000000000000004e00000000",
            INIT_0D => X"00000063000000000000005c0000000000000093000000000000009400000000",
            INIT_0E => X"0000008e0000000000000087000000000000006c000000000000005e00000000",
            INIT_0F => X"000000f500000000000000f200000000000000b7000000000000009c00000000",
            INIT_10 => X"0000006600000000000000b700000000000000ca00000000000000dc00000000",
            INIT_11 => X"0000001e000000000000008400000000000000a5000000000000006e00000000",
            INIT_12 => X"00000053000000000000006b0000000000000062000000000000003900000000",
            INIT_13 => X"0000006400000000000000810000000000000065000000000000005200000000",
            INIT_14 => X"0000009f000000000000009e00000000000000ae000000000000009900000000",
            INIT_15 => X"000000a300000000000000a200000000000000a800000000000000ac00000000",
            INIT_16 => X"00000077000000000000009c00000000000000af00000000000000a000000000",
            INIT_17 => X"000000f700000000000000e40000000000000087000000000000007200000000",
            INIT_18 => X"0000006200000000000000bc00000000000000cf00000000000000db00000000",
            INIT_19 => X"0000002a000000000000006f000000000000008d000000000000005300000000",
            INIT_1A => X"0000003e000000000000004c0000000000000048000000000000003a00000000",
            INIT_1B => X"0000005d00000000000000400000000000000038000000000000003500000000",
            INIT_1C => X"00000065000000000000005b000000000000007c00000000000000a000000000",
            INIT_1D => X"000000670000000000000067000000000000006b000000000000007400000000",
            INIT_1E => X"00000043000000000000007e000000000000009b000000000000006300000000",
            INIT_1F => X"000000f800000000000000d90000000000000076000000000000005100000000",
            INIT_20 => X"0000006500000000000000c700000000000000d200000000000000d900000000",
            INIT_21 => X"0000003c000000000000005d0000000000000058000000000000003800000000",
            INIT_22 => X"00000046000000000000003f000000000000002e000000000000003800000000",
            INIT_23 => X"0000004100000000000000400000000000000036000000000000003c00000000",
            INIT_24 => X"0000006700000000000000690000000000000072000000000000006300000000",
            INIT_25 => X"00000061000000000000005d0000000000000060000000000000006400000000",
            INIT_26 => X"000000490000000000000064000000000000006f000000000000006600000000",
            INIT_27 => X"000000f900000000000000d40000000000000072000000000000005200000000",
            INIT_28 => X"0000007500000000000000ca00000000000000cd00000000000000d100000000",
            INIT_29 => X"0000004400000000000000510000000000000046000000000000005300000000",
            INIT_2A => X"00000033000000000000002b0000000000000023000000000000003200000000",
            INIT_2B => X"0000003f0000000000000057000000000000004d000000000000004400000000",
            INIT_2C => X"0000004800000000000000520000000000000047000000000000003400000000",
            INIT_2D => X"0000005d000000000000003e0000000000000043000000000000004000000000",
            INIT_2E => X"0000006c0000000000000053000000000000003c000000000000005800000000",
            INIT_2F => X"000000fa00000000000000cc000000000000006c000000000000007000000000",
            INIT_30 => X"0000006800000000000000c500000000000000ca00000000000000cd00000000",
            INIT_31 => X"000000490000000000000047000000000000006f000000000000005d00000000",
            INIT_32 => X"0000002200000000000000260000000000000029000000000000003f00000000",
            INIT_33 => X"0000004f000000000000008e0000000000000063000000000000004b00000000",
            INIT_34 => X"0000007600000000000000930000000000000056000000000000001e00000000",
            INIT_35 => X"0000009900000000000000660000000000000072000000000000006300000000",
            INIT_36 => X"0000008d000000000000004a000000000000003f00000000000000b200000000",
            INIT_37 => X"000000f600000000000000c3000000000000005a000000000000007700000000",
            INIT_38 => X"0000005700000000000000b900000000000000c200000000000000c600000000",
            INIT_39 => X"000000630000000000000061000000000000006c000000000000003100000000",
            INIT_3A => X"0000002400000000000000270000000000000033000000000000005f00000000",
            INIT_3B => X"0000003700000000000000570000000000000032000000000000002800000000",
            INIT_3C => X"0000007f0000000000000097000000000000004f000000000000002000000000",
            INIT_3D => X"0000009c00000000000000740000000000000088000000000000007a00000000",
            INIT_3E => X"0000004a00000000000000350000000000000037000000000000009f00000000",
            INIT_3F => X"000000f000000000000000c2000000000000004e000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d00000000000000a900000000000000b400000000000000b600000000",
            INIT_41 => X"00000090000000000000006c000000000000003b000000000000002500000000",
            INIT_42 => X"00000020000000000000002b000000000000003c000000000000006a00000000",
            INIT_43 => X"00000021000000000000001e000000000000001c000000000000001d00000000",
            INIT_44 => X"00000058000000000000003a000000000000002a000000000000002700000000",
            INIT_45 => X"00000075000000000000007a0000000000000079000000000000006a00000000",
            INIT_46 => X"000000320000000000000033000000000000002f000000000000004300000000",
            INIT_47 => X"000000e100000000000000ba0000000000000050000000000000003300000000",
            INIT_48 => X"0000007d00000000000000a400000000000000a500000000000000a800000000",
            INIT_49 => X"0000008d000000000000006f0000000000000060000000000000005b00000000",
            INIT_4A => X"000000240000000000000037000000000000004a000000000000006000000000",
            INIT_4B => X"0000001f000000000000001d000000000000001e000000000000001e00000000",
            INIT_4C => X"000000ae00000000000000400000000000000018000000000000002300000000",
            INIT_4D => X"000000b500000000000000b300000000000000cb00000000000000cd00000000",
            INIT_4E => X"00000030000000000000002b0000000000000026000000000000005700000000",
            INIT_4F => X"000000d300000000000000ae000000000000005b000000000000004200000000",
            INIT_50 => X"000000b400000000000000af00000000000000a300000000000000a200000000",
            INIT_51 => X"0000008d000000000000006c0000000000000076000000000000009800000000",
            INIT_52 => X"00000030000000000000004e0000000000000053000000000000005b00000000",
            INIT_53 => X"0000001d00000000000000190000000000000018000000000000001900000000",
            INIT_54 => X"000000a400000000000000470000000000000026000000000000002700000000",
            INIT_55 => X"000000a600000000000000a900000000000000b100000000000000b800000000",
            INIT_56 => X"00000031000000000000001e000000000000001e000000000000005100000000",
            INIT_57 => X"000000ce00000000000000a9000000000000005f000000000000004e00000000",
            INIT_58 => X"000000a600000000000000b300000000000000ac000000000000009a00000000",
            INIT_59 => X"0000009200000000000000670000000000000075000000000000009200000000",
            INIT_5A => X"0000003600000000000000520000000000000055000000000000005700000000",
            INIT_5B => X"000000250000000000000021000000000000001e000000000000002000000000",
            INIT_5C => X"000000650000000000000056000000000000004d000000000000003600000000",
            INIT_5D => X"00000089000000000000008e0000000000000079000000000000006b00000000",
            INIT_5E => X"000000360000000000000021000000000000001e000000000000003c00000000",
            INIT_5F => X"000000c700000000000000a5000000000000005b000000000000004e00000000",
            INIT_60 => X"00000094000000000000009e00000000000000a900000000000000a600000000",
            INIT_61 => X"0000007100000000000000670000000000000085000000000000008f00000000",
            INIT_62 => X"0000003c000000000000004b0000000000000051000000000000004f00000000",
            INIT_63 => X"0000002c000000000000002a0000000000000027000000000000002a00000000",
            INIT_64 => X"0000004d00000000000000410000000000000036000000000000003000000000",
            INIT_65 => X"0000008b0000000000000083000000000000006e000000000000005a00000000",
            INIT_66 => X"000000360000000000000026000000000000001d000000000000003500000000",
            INIT_67 => X"000000c400000000000000a9000000000000005b000000000000004600000000",
            INIT_68 => X"0000008d0000000000000093000000000000009700000000000000a200000000",
            INIT_69 => X"0000004e000000000000006b0000000000000085000000000000008900000000",
            INIT_6A => X"0000003c0000000000000046000000000000004e000000000000004800000000",
            INIT_6B => X"00000030000000000000002e000000000000002a000000000000003200000000",
            INIT_6C => X"00000042000000000000003b0000000000000033000000000000003100000000",
            INIT_6D => X"0000007100000000000000650000000000000059000000000000004c00000000",
            INIT_6E => X"000000340000000000000023000000000000001d000000000000004500000000",
            INIT_6F => X"000000ba00000000000000ae0000000000000062000000000000003f00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009400000000",
            INIT_71 => X"0000003c000000000000006a000000000000008c000000000000008f00000000",
            INIT_72 => X"000000370000000000000042000000000000004a000000000000004200000000",
            INIT_73 => X"0000003a00000000000000360000000000000034000000000000003900000000",
            INIT_74 => X"000000460000000000000041000000000000003a000000000000003a00000000",
            INIT_75 => X"0000005d00000000000000570000000000000050000000000000004900000000",
            INIT_76 => X"0000003700000000000000260000000000000025000000000000004d00000000",
            INIT_77 => X"000000b400000000000000b30000000000000083000000000000004a00000000",
            INIT_78 => X"000000a200000000000000a00000000000000095000000000000009000000000",
            INIT_79 => X"0000003d000000000000007e0000000000000092000000000000009e00000000",
            INIT_7A => X"00000043000000000000003a0000000000000039000000000000003900000000",
            INIT_7B => X"0000004800000000000000490000000000000045000000000000004600000000",
            INIT_7C => X"0000006200000000000000590000000000000049000000000000004400000000",
            INIT_7D => X"0000006100000000000000630000000000000061000000000000005e00000000",
            INIT_7E => X"0000004700000000000000400000000000000045000000000000005200000000",
            INIT_7F => X"000000ba00000000000000b600000000000000a4000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "sampleifmap_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ca00000000000000d000000000000000d000000000000000d700000000",
            INIT_01 => X"000000b900000000000000ca00000000000000d100000000000000d700000000",
            INIT_02 => X"000000a0000000000000009800000000000000a800000000000000b800000000",
            INIT_03 => X"0000009d000000000000009a00000000000000a7000000000000009d00000000",
            INIT_04 => X"000000e100000000000000e100000000000000cb00000000000000b500000000",
            INIT_05 => X"000000e400000000000000e500000000000000db00000000000000de00000000",
            INIT_06 => X"000000c400000000000000b800000000000000c500000000000000dd00000000",
            INIT_07 => X"000000a500000000000000b000000000000000b800000000000000d000000000",
            INIT_08 => X"000000d900000000000000e100000000000000e000000000000000e200000000",
            INIT_09 => X"000000ab00000000000000cc00000000000000dd00000000000000d500000000",
            INIT_0A => X"000000b100000000000000b200000000000000bd00000000000000b400000000",
            INIT_0B => X"000000e000000000000000d000000000000000cd00000000000000c400000000",
            INIT_0C => X"000000f300000000000000f200000000000000f000000000000000ec00000000",
            INIT_0D => X"000000e700000000000000e400000000000000e500000000000000ee00000000",
            INIT_0E => X"000000d200000000000000d400000000000000d600000000000000e700000000",
            INIT_0F => X"000000c500000000000000bf00000000000000be00000000000000de00000000",
            INIT_10 => X"000000eb00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_11 => X"000000a600000000000000d600000000000000ef00000000000000ea00000000",
            INIT_12 => X"000000b100000000000000a800000000000000b100000000000000a600000000",
            INIT_13 => X"000000df00000000000000ce00000000000000b700000000000000b800000000",
            INIT_14 => X"000000e800000000000000e300000000000000ec00000000000000dc00000000",
            INIT_15 => X"000000e000000000000000d900000000000000e400000000000000eb00000000",
            INIT_16 => X"000000dd00000000000000e600000000000000e900000000000000e900000000",
            INIT_17 => X"000000d200000000000000d100000000000000ce00000000000000d900000000",
            INIT_18 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009900000000000000e300000000000000f400000000000000f400000000",
            INIT_1A => X"0000009f0000000000000082000000000000009b000000000000009200000000",
            INIT_1B => X"000000a000000000000000a2000000000000008a000000000000009000000000",
            INIT_1C => X"000000dc00000000000000c200000000000000cd00000000000000ac00000000",
            INIT_1D => X"000000e000000000000000d300000000000000d300000000000000de00000000",
            INIT_1E => X"000000db00000000000000e500000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e200000000000000df00000000000000cf00000000",
            INIT_20 => X"000000f400000000000000f400000000000000f400000000000000f500000000",
            INIT_21 => X"0000007000000000000000cd00000000000000f000000000000000f500000000",
            INIT_22 => X"0000006d000000000000005b000000000000006d000000000000006200000000",
            INIT_23 => X"0000005c0000000000000064000000000000005c000000000000006500000000",
            INIT_24 => X"0000009a000000000000007c000000000000007d000000000000006800000000",
            INIT_25 => X"000000e300000000000000c900000000000000c200000000000000c200000000",
            INIT_26 => X"000000d300000000000000e300000000000000de00000000000000dc00000000",
            INIT_27 => X"000000e100000000000000e800000000000000dc00000000000000cb00000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007b00000000000000d400000000000000eb00000000000000f600000000",
            INIT_2A => X"00000069000000000000005f000000000000005d000000000000004700000000",
            INIT_2B => X"00000066000000000000006e000000000000006a000000000000006700000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005b00000000",
            INIT_2D => X"000000e600000000000000d900000000000000c5000000000000008100000000",
            INIT_2E => X"000000c600000000000000d600000000000000da00000000000000dd00000000",
            INIT_2F => X"000000ed00000000000000e200000000000000c500000000000000b400000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009c00000000000000d500000000000000d600000000000000f000000000",
            INIT_32 => X"0000009a00000000000000890000000000000077000000000000004f00000000",
            INIT_33 => X"00000096000000000000009b000000000000008b000000000000009000000000",
            INIT_34 => X"0000007e00000000000000790000000000000080000000000000008e00000000",
            INIT_35 => X"000000e900000000000000e100000000000000a0000000000000007200000000",
            INIT_36 => X"000000ba00000000000000c000000000000000da00000000000000e900000000",
            INIT_37 => X"000000ec00000000000000d400000000000000b000000000000000a500000000",
            INIT_38 => X"000000f700000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009600000000000000d300000000000000c100000000000000e200000000",
            INIT_3A => X"000000c800000000000000bc0000000000000098000000000000005100000000",
            INIT_3B => X"00000090000000000000008d00000000000000a500000000000000cd00000000",
            INIT_3C => X"0000008f000000000000008d0000000000000096000000000000008e00000000",
            INIT_3D => X"000000d600000000000000a3000000000000008c00000000000000a700000000",
            INIT_3E => X"000000d200000000000000d300000000000000d100000000000000e000000000",
            INIT_3F => X"000000dc00000000000000af00000000000000ae00000000000000c700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000007f00000000000000d800000000000000ca00000000000000e100000000",
            INIT_42 => X"0000008700000000000000840000000000000086000000000000005100000000",
            INIT_43 => X"00000087000000000000007c000000000000009700000000000000b900000000",
            INIT_44 => X"0000008800000000000000960000000000000091000000000000008600000000",
            INIT_45 => X"000000c0000000000000008e000000000000009e00000000000000a400000000",
            INIT_46 => X"000000d700000000000000e700000000000000d800000000000000cf00000000",
            INIT_47 => X"000000c4000000000000009c000000000000009e00000000000000b100000000",
            INIT_48 => X"000000f200000000000000f400000000000000f200000000000000f200000000",
            INIT_49 => X"0000006e00000000000000a800000000000000bd00000000000000e300000000",
            INIT_4A => X"000000760000000000000080000000000000008c000000000000005300000000",
            INIT_4B => X"00000081000000000000007c0000000000000087000000000000009300000000",
            INIT_4C => X"000000860000000000000097000000000000008b000000000000008500000000",
            INIT_4D => X"000000c1000000000000009100000000000000a4000000000000009e00000000",
            INIT_4E => X"000000e600000000000000ef00000000000000ef00000000000000e500000000",
            INIT_4F => X"000000d700000000000000cc00000000000000be00000000000000c100000000",
            INIT_50 => X"000000f400000000000000f300000000000000ef00000000000000e800000000",
            INIT_51 => X"0000005e0000000000000080000000000000008100000000000000da00000000",
            INIT_52 => X"00000070000000000000007a000000000000007a000000000000004f00000000",
            INIT_53 => X"0000007300000000000000730000000000000070000000000000007100000000",
            INIT_54 => X"0000007e000000000000007f0000000000000080000000000000007c00000000",
            INIT_55 => X"000000aa0000000000000099000000000000009e000000000000009000000000",
            INIT_56 => X"000000f400000000000000f600000000000000e300000000000000ce00000000",
            INIT_57 => X"000000f400000000000000f500000000000000f300000000000000f300000000",
            INIT_58 => X"000000f200000000000000f200000000000000e300000000000000cd00000000",
            INIT_59 => X"00000058000000000000009f00000000000000a100000000000000d300000000",
            INIT_5A => X"00000066000000000000005e0000000000000045000000000000003c00000000",
            INIT_5B => X"0000006600000000000000670000000000000061000000000000006200000000",
            INIT_5C => X"00000067000000000000005f0000000000000064000000000000006800000000",
            INIT_5D => X"000000800000000000000089000000000000007f000000000000007100000000",
            INIT_5E => X"000000f300000000000000f800000000000000d7000000000000009900000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000dc00000000000000e400000000000000d500000000000000bc00000000",
            INIT_61 => X"0000006300000000000000ad00000000000000aa00000000000000b400000000",
            INIT_62 => X"00000066000000000000005a0000000000000039000000000000003700000000",
            INIT_63 => X"0000005500000000000000580000000000000067000000000000007200000000",
            INIT_64 => X"00000073000000000000005d0000000000000055000000000000005500000000",
            INIT_65 => X"0000008600000000000000760000000000000065000000000000007000000000",
            INIT_66 => X"000000f400000000000000f500000000000000e100000000000000b000000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000b500000000000000ca00000000000000bc00000000000000b800000000",
            INIT_69 => X"00000063000000000000008d0000000000000086000000000000009800000000",
            INIT_6A => X"00000067000000000000006f0000000000000066000000000000006700000000",
            INIT_6B => X"0000005600000000000000600000000000000078000000000000007600000000",
            INIT_6C => X"00000092000000000000007d000000000000006b000000000000005c00000000",
            INIT_6D => X"0000007f000000000000006e000000000000006a000000000000008400000000",
            INIT_6E => X"000000d200000000000000c300000000000000b3000000000000009800000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ee00000000",
            INIT_70 => X"0000009800000000000000bd00000000000000c200000000000000b600000000",
            INIT_71 => X"0000007e000000000000007f000000000000007b000000000000009200000000",
            INIT_72 => X"0000005e0000000000000069000000000000005d000000000000007c00000000",
            INIT_73 => X"0000004f0000000000000055000000000000005d000000000000005a00000000",
            INIT_74 => X"0000005500000000000000540000000000000053000000000000004e00000000",
            INIT_75 => X"00000053000000000000004c000000000000004b000000000000005100000000",
            INIT_76 => X"0000008a000000000000008a000000000000007a000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bc00000000",
            INIT_78 => X"0000006500000000000000a700000000000000cc00000000000000bd00000000",
            INIT_79 => X"000000ae00000000000000a9000000000000007d000000000000006500000000",
            INIT_7A => X"00000036000000000000004f000000000000004d000000000000006700000000",
            INIT_7B => X"0000003e000000000000003b000000000000002f000000000000002b00000000",
            INIT_7C => X"000000340000000000000039000000000000003e000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000030000000000000002f00000000",
            INIT_7E => X"00000061000000000000005a000000000000004a000000000000004600000000",
            INIT_7F => X"000000f400000000000000f600000000000000df000000000000008000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "sampleifmap_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000054000000000000009700000000000000a400000000000000ae00000000",
            INIT_01 => X"0000009200000000000000ac000000000000007c000000000000005200000000",
            INIT_02 => X"0000005a00000000000000570000000000000049000000000000005300000000",
            INIT_03 => X"00000044000000000000004c000000000000004b000000000000006400000000",
            INIT_04 => X"00000017000000000000001a0000000000000017000000000000002100000000",
            INIT_05 => X"000000190000000000000014000000000000002f000000000000003000000000",
            INIT_06 => X"0000006400000000000000560000000000000032000000000000001500000000",
            INIT_07 => X"000000f300000000000000f700000000000000ca000000000000007800000000",
            INIT_08 => X"0000006800000000000000b300000000000000b400000000000000c000000000",
            INIT_09 => X"00000040000000000000008e0000000000000087000000000000006800000000",
            INIT_0A => X"00000078000000000000006c0000000000000057000000000000004100000000",
            INIT_0B => X"00000062000000000000007d0000000000000076000000000000009500000000",
            INIT_0C => X"00000060000000000000006a0000000000000059000000000000004600000000",
            INIT_0D => X"0000006000000000000000590000000000000090000000000000009000000000",
            INIT_0E => X"0000008b00000000000000820000000000000067000000000000005a00000000",
            INIT_0F => X"000000f400000000000000f100000000000000b2000000000000009700000000",
            INIT_10 => X"0000005e00000000000000ab00000000000000bd00000000000000d100000000",
            INIT_11 => X"0000001c00000000000000760000000000000092000000000000006200000000",
            INIT_12 => X"0000004f0000000000000067000000000000005f000000000000003600000000",
            INIT_13 => X"0000005f00000000000000800000000000000064000000000000005300000000",
            INIT_14 => X"0000009e000000000000009b00000000000000aa000000000000009200000000",
            INIT_15 => X"000000a100000000000000a000000000000000a800000000000000ab00000000",
            INIT_16 => X"00000077000000000000009b00000000000000ac000000000000009e00000000",
            INIT_17 => X"000000f700000000000000e20000000000000080000000000000006f00000000",
            INIT_18 => X"0000005b00000000000000b000000000000000c100000000000000d000000000",
            INIT_19 => X"000000280000000000000064000000000000007f000000000000004c00000000",
            INIT_1A => X"0000003900000000000000490000000000000044000000000000003500000000",
            INIT_1B => X"00000059000000000000003d0000000000000035000000000000003200000000",
            INIT_1C => X"0000006200000000000000570000000000000077000000000000009c00000000",
            INIT_1D => X"0000006400000000000000630000000000000068000000000000007100000000",
            INIT_1E => X"0000003f000000000000007a0000000000000098000000000000006000000000",
            INIT_1F => X"000000f800000000000000d60000000000000070000000000000004d00000000",
            INIT_20 => X"0000005f00000000000000be00000000000000c300000000000000ca00000000",
            INIT_21 => X"000000380000000000000053000000000000004e000000000000003300000000",
            INIT_22 => X"00000044000000000000003c0000000000000027000000000000003300000000",
            INIT_23 => X"0000003d000000000000003b0000000000000033000000000000003900000000",
            INIT_24 => X"000000650000000000000066000000000000006e000000000000005f00000000",
            INIT_25 => X"00000060000000000000005c000000000000005f000000000000006300000000",
            INIT_26 => X"000000460000000000000060000000000000006c000000000000006400000000",
            INIT_27 => X"000000f900000000000000d0000000000000006c000000000000004f00000000",
            INIT_28 => X"0000006e00000000000000c000000000000000c000000000000000c200000000",
            INIT_29 => X"0000003f0000000000000049000000000000003e000000000000004c00000000",
            INIT_2A => X"000000300000000000000028000000000000001d000000000000002e00000000",
            INIT_2B => X"0000003b00000000000000530000000000000048000000000000004100000000",
            INIT_2C => X"00000043000000000000004d0000000000000043000000000000003000000000",
            INIT_2D => X"00000058000000000000003b0000000000000040000000000000003c00000000",
            INIT_2E => X"00000069000000000000004e0000000000000036000000000000005200000000",
            INIT_2F => X"000000f900000000000000c90000000000000065000000000000006b00000000",
            INIT_30 => X"0000006100000000000000bb00000000000000be00000000000000c300000000",
            INIT_31 => X"0000004300000000000000410000000000000063000000000000005500000000",
            INIT_32 => X"0000002000000000000000230000000000000026000000000000003a00000000",
            INIT_33 => X"0000004c000000000000008d0000000000000060000000000000004800000000",
            INIT_34 => X"00000071000000000000008c000000000000004f000000000000001900000000",
            INIT_35 => X"000000920000000000000061000000000000006d000000000000005e00000000",
            INIT_36 => X"0000008a0000000000000045000000000000003a00000000000000ab00000000",
            INIT_37 => X"000000f400000000000000c00000000000000053000000000000007400000000",
            INIT_38 => X"0000005200000000000000b000000000000000b700000000000000bd00000000",
            INIT_39 => X"0000005e00000000000000590000000000000063000000000000002c00000000",
            INIT_3A => X"0000002100000000000000240000000000000030000000000000005a00000000",
            INIT_3B => X"000000340000000000000055000000000000002f000000000000002600000000",
            INIT_3C => X"0000007b0000000000000091000000000000004a000000000000001c00000000",
            INIT_3D => X"0000009700000000000000710000000000000086000000000000007700000000",
            INIT_3E => X"0000004700000000000000320000000000000033000000000000009c00000000",
            INIT_3F => X"000000ee00000000000000c00000000000000047000000000000003b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004800000000000000a300000000000000ad00000000000000ae00000000",
            INIT_41 => X"0000008b00000000000000650000000000000036000000000000002200000000",
            INIT_42 => X"0000001e0000000000000028000000000000003a000000000000006600000000",
            INIT_43 => X"0000001e000000000000001a0000000000000019000000000000001a00000000",
            INIT_44 => X"0000005600000000000000350000000000000026000000000000002500000000",
            INIT_45 => X"0000007200000000000000760000000000000075000000000000006800000000",
            INIT_46 => X"0000002e0000000000000030000000000000002b000000000000003e00000000",
            INIT_47 => X"000000df00000000000000b8000000000000004b000000000000002f00000000",
            INIT_48 => X"00000078000000000000009e00000000000000a000000000000000a200000000",
            INIT_49 => X"0000008800000000000000670000000000000059000000000000005700000000",
            INIT_4A => X"0000002200000000000000340000000000000048000000000000005c00000000",
            INIT_4B => X"0000001d000000000000001b000000000000001b000000000000001c00000000",
            INIT_4C => X"000000af000000000000003d0000000000000015000000000000002000000000",
            INIT_4D => X"000000b400000000000000b100000000000000ca00000000000000cf00000000",
            INIT_4E => X"0000002c00000000000000280000000000000022000000000000005400000000",
            INIT_4F => X"000000d100000000000000ab0000000000000057000000000000003e00000000",
            INIT_50 => X"000000b000000000000000a8000000000000009c000000000000009c00000000",
            INIT_51 => X"0000008800000000000000660000000000000070000000000000009300000000",
            INIT_52 => X"0000002d000000000000004b0000000000000051000000000000005600000000",
            INIT_53 => X"0000001a00000000000000170000000000000016000000000000001600000000",
            INIT_54 => X"000000a400000000000000450000000000000022000000000000002300000000",
            INIT_55 => X"000000a500000000000000a900000000000000b100000000000000b900000000",
            INIT_56 => X"0000002d000000000000001a0000000000000019000000000000004e00000000",
            INIT_57 => X"000000cc00000000000000a7000000000000005c000000000000004b00000000",
            INIT_58 => X"000000a100000000000000ad00000000000000a7000000000000009500000000",
            INIT_59 => X"0000008e00000000000000630000000000000071000000000000008d00000000",
            INIT_5A => X"00000033000000000000004f0000000000000053000000000000005300000000",
            INIT_5B => X"00000022000000000000001f000000000000001c000000000000001d00000000",
            INIT_5C => X"0000006100000000000000510000000000000048000000000000003200000000",
            INIT_5D => X"00000085000000000000008a0000000000000074000000000000006600000000",
            INIT_5E => X"00000032000000000000001d000000000000001b000000000000003700000000",
            INIT_5F => X"000000c600000000000000a40000000000000059000000000000004c00000000",
            INIT_60 => X"00000090000000000000009b00000000000000a600000000000000a400000000",
            INIT_61 => X"0000006c00000000000000630000000000000082000000000000008b00000000",
            INIT_62 => X"0000003800000000000000480000000000000050000000000000004c00000000",
            INIT_63 => X"0000002900000000000000270000000000000024000000000000002600000000",
            INIT_64 => X"00000048000000000000003d0000000000000033000000000000002d00000000",
            INIT_65 => X"00000083000000000000007c0000000000000067000000000000005400000000",
            INIT_66 => X"000000320000000000000021000000000000001a000000000000003100000000",
            INIT_67 => X"000000c300000000000000a90000000000000059000000000000004500000000",
            INIT_68 => X"0000008d0000000000000092000000000000009400000000000000a000000000",
            INIT_69 => X"0000004900000000000000660000000000000082000000000000008700000000",
            INIT_6A => X"000000380000000000000042000000000000004d000000000000004500000000",
            INIT_6B => X"0000002d000000000000002b0000000000000028000000000000002f00000000",
            INIT_6C => X"0000003d00000000000000360000000000000030000000000000002e00000000",
            INIT_6D => X"0000006a000000000000005e0000000000000054000000000000004600000000",
            INIT_6E => X"00000030000000000000001f000000000000001a000000000000004000000000",
            INIT_6F => X"000000ba00000000000000af0000000000000062000000000000003d00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009300000000",
            INIT_71 => X"000000390000000000000068000000000000008b000000000000008f00000000",
            INIT_72 => X"00000034000000000000003f000000000000004a000000000000004000000000",
            INIT_73 => X"0000003600000000000000330000000000000031000000000000003700000000",
            INIT_74 => X"00000042000000000000003d0000000000000036000000000000003600000000",
            INIT_75 => X"000000570000000000000051000000000000004a000000000000004400000000",
            INIT_76 => X"0000003400000000000000230000000000000021000000000000004800000000",
            INIT_77 => X"000000b500000000000000b60000000000000084000000000000004800000000",
            INIT_78 => X"000000a300000000000000a10000000000000096000000000000009200000000",
            INIT_79 => X"0000003a000000000000007c0000000000000091000000000000009d00000000",
            INIT_7A => X"0000004100000000000000390000000000000038000000000000003700000000",
            INIT_7B => X"0000004500000000000000460000000000000042000000000000004300000000",
            INIT_7C => X"0000005f00000000000000570000000000000048000000000000004300000000",
            INIT_7D => X"0000005e0000000000000060000000000000005f000000000000005c00000000",
            INIT_7E => X"00000046000000000000003e0000000000000044000000000000005100000000",
            INIT_7F => X"000000b900000000000000b600000000000000a3000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "sampleifmap_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000bf00000000000000ca00000000000000d100000000",
            INIT_01 => X"000000af00000000000000c600000000000000d100000000000000d100000000",
            INIT_02 => X"000000a0000000000000009d00000000000000a500000000000000ab00000000",
            INIT_03 => X"0000008f000000000000008d000000000000009a000000000000009500000000",
            INIT_04 => X"000000db00000000000000d600000000000000bc00000000000000a400000000",
            INIT_05 => X"000000d600000000000000d900000000000000ca00000000000000d100000000",
            INIT_06 => X"000000ad00000000000000a100000000000000b100000000000000d000000000",
            INIT_07 => X"000000950000000000000095000000000000009d00000000000000b700000000",
            INIT_08 => X"000000cd00000000000000d200000000000000d400000000000000d400000000",
            INIT_09 => X"000000a300000000000000c800000000000000db00000000000000cf00000000",
            INIT_0A => X"000000b600000000000000b800000000000000b600000000000000a500000000",
            INIT_0B => X"000000d700000000000000cd00000000000000c900000000000000c200000000",
            INIT_0C => X"000000e400000000000000e300000000000000e300000000000000df00000000",
            INIT_0D => X"000000d700000000000000d300000000000000d400000000000000dd00000000",
            INIT_0E => X"000000bb00000000000000c300000000000000cd00000000000000df00000000",
            INIT_0F => X"000000ba00000000000000ad00000000000000aa00000000000000c600000000",
            INIT_10 => X"000000e200000000000000e300000000000000e500000000000000e600000000",
            INIT_11 => X"000000a400000000000000d300000000000000ec00000000000000e300000000",
            INIT_12 => X"000000b800000000000000b700000000000000ad000000000000009f00000000",
            INIT_13 => X"000000e000000000000000cf00000000000000bf00000000000000bc00000000",
            INIT_14 => X"000000d600000000000000e000000000000000e500000000000000db00000000",
            INIT_15 => X"000000d300000000000000c800000000000000d000000000000000d600000000",
            INIT_16 => X"000000c500000000000000db00000000000000e000000000000000de00000000",
            INIT_17 => X"000000c600000000000000c500000000000000bc00000000000000b900000000",
            INIT_18 => X"000000f100000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"000000af00000000000000e300000000000000f100000000000000f200000000",
            INIT_1A => X"000000bb00000000000000a100000000000000b000000000000000a800000000",
            INIT_1B => X"000000b600000000000000b800000000000000a000000000000000ae00000000",
            INIT_1C => X"000000ca00000000000000d000000000000000d500000000000000b900000000",
            INIT_1D => X"000000d400000000000000c400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000bb00000000000000d500000000000000dc00000000000000d700000000",
            INIT_1F => X"000000c800000000000000d400000000000000c500000000000000a900000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000008400000000000000cd00000000000000f100000000000000f500000000",
            INIT_22 => X"000000a7000000000000008a00000000000000a1000000000000008b00000000",
            INIT_23 => X"0000008d000000000000009b000000000000008b000000000000009f00000000",
            INIT_24 => X"000000a4000000000000009900000000000000a6000000000000008e00000000",
            INIT_25 => X"000000e000000000000000c400000000000000a900000000000000a900000000",
            INIT_26 => X"000000b100000000000000d400000000000000d100000000000000d100000000",
            INIT_27 => X"000000d200000000000000cc00000000000000b800000000000000a000000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000008100000000000000d700000000000000ee00000000000000f600000000",
            INIT_2A => X"000000aa00000000000000a0000000000000009c000000000000007100000000",
            INIT_2B => X"000000a700000000000000b100000000000000aa00000000000000aa00000000",
            INIT_2C => X"0000008f0000000000000098000000000000009d000000000000009d00000000",
            INIT_2D => X"000000e400000000000000cd00000000000000b3000000000000009400000000",
            INIT_2E => X"000000aa00000000000000c100000000000000ce00000000000000da00000000",
            INIT_2F => X"000000df00000000000000c000000000000000a0000000000000009300000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"000000b400000000000000dd00000000000000dd00000000000000f100000000",
            INIT_32 => X"000000cf00000000000000c400000000000000b4000000000000008300000000",
            INIT_33 => X"000000d300000000000000d900000000000000cb00000000000000c800000000",
            INIT_34 => X"000000bf00000000000000c000000000000000c300000000000000cc00000000",
            INIT_35 => X"000000e100000000000000cd00000000000000a600000000000000a300000000",
            INIT_36 => X"000000a900000000000000b100000000000000d500000000000000e300000000",
            INIT_37 => X"000000da00000000000000b20000000000000092000000000000009100000000",
            INIT_38 => X"000000f700000000000000f200000000000000f200000000000000f400000000",
            INIT_39 => X"000000c000000000000000d900000000000000ca00000000000000e600000000",
            INIT_3A => X"000000e800000000000000e000000000000000c2000000000000008600000000",
            INIT_3B => X"000000d100000000000000ce00000000000000d700000000000000ea00000000",
            INIT_3C => X"000000cf00000000000000ca00000000000000d000000000000000cf00000000",
            INIT_3D => X"000000cc000000000000009a00000000000000b400000000000000e000000000",
            INIT_3E => X"000000bc00000000000000c400000000000000c900000000000000dc00000000",
            INIT_3F => X"000000c7000000000000009a000000000000009200000000000000ab00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f300000000000000f300000000000000f500000000",
            INIT_41 => X"000000ae00000000000000df00000000000000d100000000000000e300000000",
            INIT_42 => X"000000c100000000000000c100000000000000ba000000000000008700000000",
            INIT_43 => X"000000c900000000000000c100000000000000cc00000000000000dd00000000",
            INIT_44 => X"000000c600000000000000cd00000000000000cd00000000000000ca00000000",
            INIT_45 => X"000000bc00000000000000a300000000000000d000000000000000dc00000000",
            INIT_46 => X"000000cb00000000000000df00000000000000d100000000000000cb00000000",
            INIT_47 => X"000000b20000000000000094000000000000008b00000000000000a100000000",
            INIT_48 => X"000000f200000000000000f300000000000000f100000000000000f200000000",
            INIT_49 => X"000000a400000000000000c200000000000000cd00000000000000e500000000",
            INIT_4A => X"000000b800000000000000bd00000000000000c1000000000000008c00000000",
            INIT_4B => X"000000c400000000000000c000000000000000c400000000000000ca00000000",
            INIT_4C => X"000000c600000000000000d000000000000000ca00000000000000c700000000",
            INIT_4D => X"000000c800000000000000bc00000000000000e000000000000000d700000000",
            INIT_4E => X"000000e300000000000000ed00000000000000ee00000000000000e600000000",
            INIT_4F => X"000000d300000000000000ca00000000000000ba00000000000000bc00000000",
            INIT_50 => X"000000f400000000000000f300000000000000ee00000000000000ea00000000",
            INIT_51 => X"0000009c00000000000000a900000000000000a000000000000000df00000000",
            INIT_52 => X"000000ac00000000000000b300000000000000b1000000000000008600000000",
            INIT_53 => X"000000b700000000000000b400000000000000ae00000000000000ae00000000",
            INIT_54 => X"000000be00000000000000bc00000000000000be00000000000000bb00000000",
            INIT_55 => X"000000c400000000000000d000000000000000dc00000000000000cd00000000",
            INIT_56 => X"000000f400000000000000f600000000000000e600000000000000d900000000",
            INIT_57 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_58 => X"000000f200000000000000f200000000000000e600000000000000d300000000",
            INIT_59 => X"0000009700000000000000be00000000000000b600000000000000d800000000",
            INIT_5A => X"000000a00000000000000093000000000000006e000000000000006a00000000",
            INIT_5B => X"000000aa00000000000000a6000000000000009f000000000000009e00000000",
            INIT_5C => X"000000a6000000000000009e00000000000000a300000000000000a900000000",
            INIT_5D => X"000000af00000000000000c600000000000000bd00000000000000ad00000000",
            INIT_5E => X"000000f300000000000000f800000000000000e000000000000000b700000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e100000000000000e900000000000000da00000000000000c400000000",
            INIT_61 => X"0000009f00000000000000c300000000000000b400000000000000bd00000000",
            INIT_62 => X"000000a0000000000000008d000000000000005c000000000000005d00000000",
            INIT_63 => X"0000008c000000000000008f00000000000000a800000000000000ba00000000",
            INIT_64 => X"000000a700000000000000920000000000000089000000000000008b00000000",
            INIT_65 => X"00000096000000000000008f0000000000000083000000000000009800000000",
            INIT_66 => X"000000f400000000000000f300000000000000e300000000000000bc00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c100000000000000d300000000000000c700000000000000c300000000",
            INIT_69 => X"0000008900000000000000a2000000000000009500000000000000a400000000",
            INIT_6A => X"000000a600000000000000b200000000000000aa000000000000009600000000",
            INIT_6B => X"0000009200000000000000a600000000000000cd00000000000000bd00000000",
            INIT_6C => X"000000d300000000000000c000000000000000ac000000000000009900000000",
            INIT_6D => X"0000008a0000000000000080000000000000008000000000000000af00000000",
            INIT_6E => X"000000d300000000000000bf00000000000000b100000000000000a000000000",
            INIT_6F => X"000000f300000000000000f300000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a200000000000000c800000000000000cf00000000000000c200000000",
            INIT_71 => X"00000089000000000000008e0000000000000088000000000000009c00000000",
            INIT_72 => X"0000009f00000000000000b100000000000000b200000000000000a200000000",
            INIT_73 => X"0000008b000000000000009500000000000000a3000000000000009600000000",
            INIT_74 => X"0000009300000000000000920000000000000092000000000000008d00000000",
            INIT_75 => X"00000085000000000000007f000000000000007c000000000000008600000000",
            INIT_76 => X"000000a600000000000000ad00000000000000a3000000000000009500000000",
            INIT_77 => X"000000f400000000000000f300000000000000f500000000000000cc00000000",
            INIT_78 => X"0000006e00000000000000ad00000000000000d000000000000000c300000000",
            INIT_79 => X"000000b900000000000000b4000000000000008b000000000000007100000000",
            INIT_7A => X"00000057000000000000007f000000000000009a000000000000008500000000",
            INIT_7B => X"0000005f0000000000000059000000000000004c000000000000004900000000",
            INIT_7C => X"00000058000000000000005e0000000000000060000000000000005c00000000",
            INIT_7D => X"0000006700000000000000630000000000000056000000000000005600000000",
            INIT_7E => X"0000009b000000000000008f0000000000000074000000000000006d00000000",
            INIT_7F => X"000000f500000000000000f500000000000000e800000000000000af00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "sampleifmap_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006500000000000000a100000000000000aa00000000000000b700000000",
            INIT_01 => X"000000a100000000000000b50000000000000088000000000000006000000000",
            INIT_02 => X"0000008700000000000000810000000000000084000000000000008000000000",
            INIT_03 => X"0000006a000000000000007d000000000000007d000000000000008c00000000",
            INIT_04 => X"00000027000000000000002c000000000000002b000000000000003500000000",
            INIT_05 => X"0000002800000000000000230000000000000047000000000000004d00000000",
            INIT_06 => X"0000009700000000000000910000000000000050000000000000002000000000",
            INIT_07 => X"000000f300000000000000f600000000000000db00000000000000a700000000",
            INIT_08 => X"0000007c00000000000000c200000000000000c100000000000000ca00000000",
            INIT_09 => X"0000004900000000000000990000000000000092000000000000007800000000",
            INIT_0A => X"0000009400000000000000830000000000000087000000000000006900000000",
            INIT_0B => X"0000008300000000000000a9000000000000009f00000000000000b800000000",
            INIT_0C => X"0000007a00000000000000840000000000000076000000000000006600000000",
            INIT_0D => X"00000073000000000000006f00000000000000aa00000000000000af00000000",
            INIT_0E => X"000000b500000000000000b20000000000000091000000000000006f00000000",
            INIT_0F => X"000000f400000000000000f200000000000000c500000000000000bb00000000",
            INIT_10 => X"0000007200000000000000b800000000000000c800000000000000d800000000",
            INIT_11 => X"000000240000000000000082000000000000009d000000000000007300000000",
            INIT_12 => X"0000006300000000000000810000000000000095000000000000004f00000000",
            INIT_13 => X"00000084000000000000009d0000000000000081000000000000006f00000000",
            INIT_14 => X"000000b900000000000000b700000000000000c100000000000000b100000000",
            INIT_15 => X"000000bd00000000000000ba00000000000000c100000000000000c800000000",
            INIT_16 => X"0000009700000000000000b600000000000000c700000000000000b500000000",
            INIT_17 => X"000000f600000000000000e800000000000000a2000000000000009400000000",
            INIT_18 => X"0000007100000000000000bb00000000000000cc00000000000000d900000000",
            INIT_19 => X"0000003d0000000000000071000000000000008b000000000000006000000000",
            INIT_1A => X"0000005d00000000000000730000000000000070000000000000004e00000000",
            INIT_1B => X"0000007d000000000000005e0000000000000053000000000000005500000000",
            INIT_1C => X"0000008a000000000000007f000000000000009f00000000000000bf00000000",
            INIT_1D => X"0000008f000000000000008c000000000000009500000000000000a000000000",
            INIT_1E => X"00000063000000000000009f00000000000000bd000000000000008a00000000",
            INIT_1F => X"000000f700000000000000e2000000000000009a000000000000007300000000",
            INIT_20 => X"0000007500000000000000c700000000000000d000000000000000d500000000",
            INIT_21 => X"000000540000000000000063000000000000005c000000000000004900000000",
            INIT_22 => X"0000006900000000000000610000000000000041000000000000004b00000000",
            INIT_23 => X"0000005f00000000000000670000000000000057000000000000005f00000000",
            INIT_24 => X"00000097000000000000009900000000000000a2000000000000008600000000",
            INIT_25 => X"0000008f00000000000000890000000000000090000000000000009600000000",
            INIT_26 => X"0000006f000000000000008f0000000000000099000000000000009300000000",
            INIT_27 => X"000000f700000000000000de0000000000000092000000000000007300000000",
            INIT_28 => X"0000008300000000000000cc00000000000000ce00000000000000cc00000000",
            INIT_29 => X"0000005a000000000000005c0000000000000051000000000000006500000000",
            INIT_2A => X"000000450000000000000039000000000000002d000000000000004600000000",
            INIT_2B => X"00000057000000000000007d000000000000006f000000000000006200000000",
            INIT_2C => X"0000006700000000000000700000000000000066000000000000004a00000000",
            INIT_2D => X"0000007d000000000000005e0000000000000065000000000000006200000000",
            INIT_2E => X"0000009500000000000000710000000000000052000000000000007300000000",
            INIT_2F => X"000000f800000000000000d40000000000000089000000000000009a00000000",
            INIT_30 => X"0000007500000000000000ce00000000000000d000000000000000d100000000",
            INIT_31 => X"0000005e0000000000000056000000000000007a000000000000006900000000",
            INIT_32 => X"0000002f00000000000000330000000000000036000000000000005600000000",
            INIT_33 => X"0000006300000000000000ad0000000000000083000000000000006600000000",
            INIT_34 => X"00000082000000000000009e0000000000000064000000000000002d00000000",
            INIT_35 => X"000000ab000000000000007c000000000000008a000000000000007900000000",
            INIT_36 => X"000000ab000000000000005f000000000000004b00000000000000bb00000000",
            INIT_37 => X"000000fa00000000000000cf0000000000000075000000000000009800000000",
            INIT_38 => X"0000006800000000000000cc00000000000000d600000000000000dd00000000",
            INIT_39 => X"0000008000000000000000720000000000000074000000000000003b00000000",
            INIT_3A => X"0000003000000000000000340000000000000041000000000000007c00000000",
            INIT_3B => X"0000004b000000000000006c0000000000000046000000000000003800000000",
            INIT_3C => X"0000008f00000000000000a6000000000000005f000000000000003000000000",
            INIT_3D => X"000000af000000000000008f00000000000000a7000000000000009100000000",
            INIT_3E => X"000000620000000000000048000000000000004a00000000000000af00000000",
            INIT_3F => X"000000fb00000000000000d60000000000000068000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006300000000000000c900000000000000d400000000000000d700000000",
            INIT_41 => X"000000b000000000000000800000000000000044000000000000002f00000000",
            INIT_42 => X"0000002d00000000000000380000000000000050000000000000008700000000",
            INIT_43 => X"0000002f000000000000002b0000000000000027000000000000002800000000",
            INIT_44 => X"0000006e0000000000000050000000000000003c000000000000003700000000",
            INIT_45 => X"0000008b00000000000000900000000000000093000000000000007d00000000",
            INIT_46 => X"0000004300000000000000460000000000000043000000000000005c00000000",
            INIT_47 => X"000000fb00000000000000d9000000000000006d000000000000004500000000",
            INIT_48 => X"0000009d00000000000000cb00000000000000cf00000000000000cf00000000",
            INIT_49 => X"000000aa00000000000000850000000000000075000000000000007300000000",
            INIT_4A => X"0000003000000000000000480000000000000065000000000000007e00000000",
            INIT_4B => X"0000002d00000000000000290000000000000029000000000000002800000000",
            INIT_4C => X"000000c000000000000000530000000000000027000000000000003200000000",
            INIT_4D => X"000000c900000000000000c700000000000000dc00000000000000da00000000",
            INIT_4E => X"0000003f00000000000000380000000000000034000000000000006b00000000",
            INIT_4F => X"000000f700000000000000d2000000000000007e000000000000005a00000000",
            INIT_50 => X"000000d800000000000000ce00000000000000c000000000000000bc00000000",
            INIT_51 => X"000000a10000000000000086000000000000009a00000000000000bf00000000",
            INIT_52 => X"0000003e00000000000000680000000000000073000000000000007900000000",
            INIT_53 => X"0000002900000000000000230000000000000022000000000000002100000000",
            INIT_54 => X"000000b300000000000000550000000000000031000000000000003300000000",
            INIT_55 => X"000000bb00000000000000be00000000000000c000000000000000c700000000",
            INIT_56 => X"0000004200000000000000260000000000000027000000000000006000000000",
            INIT_57 => X"000000f500000000000000d10000000000000085000000000000006f00000000",
            INIT_58 => X"000000c600000000000000cd00000000000000c600000000000000bf00000000",
            INIT_59 => X"000000a00000000000000084000000000000009e00000000000000b500000000",
            INIT_5A => X"00000046000000000000006f0000000000000076000000000000007200000000",
            INIT_5B => X"00000031000000000000002c0000000000000026000000000000002700000000",
            INIT_5C => X"0000007e0000000000000069000000000000005d000000000000004400000000",
            INIT_5D => X"000000a600000000000000ad0000000000000096000000000000008700000000",
            INIT_5E => X"00000047000000000000002a0000000000000028000000000000004800000000",
            INIT_5F => X"000000f200000000000000cf0000000000000082000000000000007100000000",
            INIT_60 => X"000000b800000000000000c600000000000000d100000000000000ce00000000",
            INIT_61 => X"00000085000000000000008200000000000000a300000000000000ab00000000",
            INIT_62 => X"0000004d0000000000000068000000000000006f000000000000006b00000000",
            INIT_63 => X"000000390000000000000035000000000000002f000000000000003200000000",
            INIT_64 => X"0000006800000000000000570000000000000048000000000000003f00000000",
            INIT_65 => X"000000b000000000000000a80000000000000091000000000000007800000000",
            INIT_66 => X"0000004700000000000000300000000000000028000000000000004500000000",
            INIT_67 => X"000000ee00000000000000d4000000000000007e000000000000006600000000",
            INIT_68 => X"000000bd00000000000000c200000000000000c200000000000000c700000000",
            INIT_69 => X"00000065000000000000008600000000000000a600000000000000b200000000",
            INIT_6A => X"0000004f00000000000000600000000000000069000000000000006300000000",
            INIT_6B => X"0000003e000000000000003b0000000000000036000000000000003e00000000",
            INIT_6C => X"00000057000000000000004e0000000000000045000000000000004100000000",
            INIT_6D => X"0000008f00000000000000810000000000000074000000000000006400000000",
            INIT_6E => X"00000047000000000000002c0000000000000027000000000000005700000000",
            INIT_6F => X"000000e800000000000000df0000000000000085000000000000005900000000",
            INIT_70 => X"000000bc00000000000000be00000000000000bc00000000000000c100000000",
            INIT_71 => X"00000050000000000000009000000000000000bc00000000000000bd00000000",
            INIT_72 => X"0000004600000000000000580000000000000063000000000000005a00000000",
            INIT_73 => X"0000004e000000000000004a0000000000000045000000000000004900000000",
            INIT_74 => X"0000005d0000000000000056000000000000004e000000000000004e00000000",
            INIT_75 => X"00000072000000000000006d0000000000000066000000000000006100000000",
            INIT_76 => X"0000004a00000000000000300000000000000030000000000000005e00000000",
            INIT_77 => X"000000e700000000000000e800000000000000ad000000000000006400000000",
            INIT_78 => X"000000cd00000000000000d000000000000000c700000000000000c400000000",
            INIT_79 => X"0000005500000000000000a500000000000000bb00000000000000c800000000",
            INIT_7A => X"00000054000000000000004e000000000000004c000000000000004c00000000",
            INIT_7B => X"0000006300000000000000620000000000000059000000000000005400000000",
            INIT_7C => X"0000007c00000000000000720000000000000063000000000000005e00000000",
            INIT_7D => X"0000007f00000000000000800000000000000081000000000000007d00000000",
            INIT_7E => X"000000600000000000000054000000000000005b000000000000007000000000",
            INIT_7F => X"000000df00000000000000e100000000000000cc000000000000009400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "samplegold_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000d00000000000000000000000000000000000000000000000a00000000",
            INIT_0A => X"0000000000000000000000140000000000000017000000000000002400000000",
            INIT_0B => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002b00000000000000100000000000000016000000000000001200000000",
            INIT_0E => X"00000000000000000000000b000000000000001b000000000000001c00000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000002300000000",
            INIT_10 => X"0000001d0000000000000025000000000000001a000000000000000000000000",
            INIT_11 => X"0000001a00000000000000130000000000000006000000000000001b00000000",
            INIT_12 => X"000000470000000000000000000000000000000a000000000000000b00000000",
            INIT_13 => X"0000003300000000000000220000000000000008000000000000003000000000",
            INIT_14 => X"000000120000000000000011000000000000002e000000000000003c00000000",
            INIT_15 => X"0000000d00000000000000280000000000000040000000000000000000000000",
            INIT_16 => X"00000047000000000000003f0000000000000007000000000000001100000000",
            INIT_17 => X"0000001e00000000000000090000000000000000000000000000000300000000",
            INIT_18 => X"000000150000000000000016000000000000002c000000000000002d00000000",
            INIT_19 => X"0000000f0000000000000014000000000000001d000000000000003a00000000",
            INIT_1A => X"000000130000000000000033000000000000004b000000000000001400000000",
            INIT_1B => X"00000050000000000000001e0000000000000000000000000000000000000000",
            INIT_1C => X"00000039000000000000001c000000000000001a000000000000003200000000",
            INIT_1D => X"0000000b000000000000001f0000000000000011000000000000002000000000",
            INIT_1E => X"00000018000000000000004b0000000000000042000000000000005400000000",
            INIT_1F => X"000000130000000000000019000000000000002d000000000000001c00000000",
            INIT_20 => X"00000028000000000000000f0000000000000017000000000000000200000000",
            INIT_21 => X"0000004e00000000000000000000000000000003000000000000001200000000",
            INIT_22 => X"0000001b00000000000000210000000000000042000000000000004b00000000",
            INIT_23 => X"00000023000000000000001a0000000000000011000000000000002200000000",
            INIT_24 => X"0000000000000000000000030000000000000024000000000000002000000000",
            INIT_25 => X"0000004300000000000000340000000000000000000000000000000000000000",
            INIT_26 => X"0000001400000000000000440000000000000011000000000000004300000000",
            INIT_27 => X"000000170000000000000038000000000000004d000000000000003a00000000",
            INIT_28 => X"0000001400000000000000210000000000000013000000000000000400000000",
            INIT_29 => X"00000034000000000000004f0000000000000042000000000000001400000000",
            INIT_2A => X"00000042000000000000005a0000000000000083000000000000003c00000000",
            INIT_2B => X"0000003700000000000000300000000000000038000000000000003f00000000",
            INIT_2C => X"0000004500000000000000460000000000000041000000000000003d00000000",
            INIT_2D => X"00000065000000000000003c0000000000000045000000000000005000000000",
            INIT_2E => X"0000003a000000000000003d000000000000003b000000000000005900000000",
            INIT_2F => X"0000003e000000000000003b0000000000000037000000000000003700000000",
            INIT_30 => X"000000520000000000000043000000000000004a000000000000004a00000000",
            INIT_31 => X"00000041000000000000006b0000000000000042000000000000004400000000",
            INIT_32 => X"0000003c0000000000000039000000000000003f000000000000003b00000000",
            INIT_33 => X"0000004e000000000000004d000000000000004b000000000000004000000000",
            INIT_34 => X"0000004c000000000000005a000000000000006a000000000000004600000000",
            INIT_35 => X"0000003f000000000000003d0000000000000034000000000000005400000000",
            INIT_36 => X"00000042000000000000003d000000000000003f000000000000004300000000",
            INIT_37 => X"00000056000000000000003c0000000000000042000000000000004700000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000003000000000000000200000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_43 => X"0000003d00000000000000000000000000000001000000000000000a00000000",
            INIT_44 => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_45 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"00000000000000000000002e0000000000000000000000000000002600000000",
            INIT_48 => X"00000000000000000000000c0000000000000000000000000000003d00000000",
            INIT_49 => X"0000000000000000000000410000000000000000000000000000000000000000",
            INIT_4A => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000007d000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4F => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_53 => X"0000002a000000000000002c0000000000000000000000000000000700000000",
            INIT_54 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_58 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_59 => X"00000010000000000000000f0000000000000000000000000000000000000000",
            INIT_5A => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5D => X"0000000d0000000000000000000000000000001c000000000000002000000000",
            INIT_5E => X"0000000000000000000000750000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000019000000000000001100000000",
            INIT_60 => X"000000140000000000000013000000000000000e000000000000000000000000",
            INIT_61 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000046000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000002d000000000000001d0000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000900000000000000000000000000000000000000000000000700000000",
            INIT_69 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000060000000000000005c0000000000000000000000000000000000000000",
            INIT_71 => X"0000005a00000000000000610000000000000061000000000000006000000000",
            INIT_72 => X"0000004d00000000000000680000000000000071000000000000006400000000",
            INIT_73 => X"00000050000000000000004a0000000000000043000000000000003d00000000",
            INIT_74 => X"000000630000000000000069000000000000005e000000000000005400000000",
            INIT_75 => X"0000004d00000000000000500000000000000061000000000000006400000000",
            INIT_76 => X"0000000000000000000000180000000000000039000000000000005500000000",
            INIT_77 => X"0000004d000000000000003b000000000000001d000000000000000200000000",
            INIT_78 => X"0000006b000000000000006a000000000000004a000000000000003c00000000",
            INIT_79 => X"0000001b00000000000000370000000000000054000000000000006900000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"00000000000000000000003a0000000000000006000000000000000000000000",
            INIT_7C => X"0000005700000000000000680000000000000058000000000000000a00000000",
            INIT_7D => X"0000000000000000000000000000000000000005000000000000003500000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000001a000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "samplegold_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000038000000000000003b00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000d000000000000004e00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000056000000000000001f0000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000006000000000000000d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000006000000000000001c0000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_0F => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_10 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000c00000000000000000000000000000000000000000000000500000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000004300000000000000260000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000ba00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000bf00000000000000c200000000000000bd00000000000000c100000000",
            INIT_2A => X"000000bb00000000000000c200000000000000c600000000000000bc00000000",
            INIT_2B => X"000000a7000000000000009f00000000000000a500000000000000b500000000",
            INIT_2C => X"000000bd00000000000000b5000000000000009e00000000000000aa00000000",
            INIT_2D => X"000000e300000000000000bf00000000000000c900000000000000c200000000",
            INIT_2E => X"0000008600000000000000ac00000000000000c100000000000000e300000000",
            INIT_2F => X"0000008b000000000000007e000000000000008f00000000000000a100000000",
            INIT_30 => X"000000c0000000000000008800000000000000b600000000000000a300000000",
            INIT_31 => X"000000bf00000000000000ea00000000000000c200000000000000c300000000",
            INIT_32 => X"000000de00000000000000a20000000000000061000000000000007e00000000",
            INIT_33 => X"0000008e000000000000006900000000000000a700000000000000ae00000000",
            INIT_34 => X"000000bf00000000000000c8000000000000006800000000000000c800000000",
            INIT_35 => X"000000a300000000000000d5000000000000009e00000000000000d000000000",
            INIT_36 => X"000000ad00000000000000ef00000000000000a0000000000000009200000000",
            INIT_37 => X"00000103000000000000005e0000000000000062000000000000008e00000000",
            INIT_38 => X"0000014400000000000000b000000000000000f200000000000000ed00000000",
            INIT_39 => X"0000008a00000000000000b50000000000000115000000000000012f00000000",
            INIT_3A => X"0000008c00000000000000ce00000000000000f7000000000000006200000000",
            INIT_3B => X"00000118000000000000011e0000000000000056000000000000007d00000000",
            INIT_3C => X"0000011500000000000000f000000000000000db000000000000010300000000",
            INIT_3D => X"0000007a00000000000000a800000000000000d2000000000000012b00000000",
            INIT_3E => X"00000097000000000000009000000000000000c7000000000000014600000000",
            INIT_3F => X"000000c000000000000001450000000000000113000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000015000000000000000ed00000000000000ac00000000000000c600000000",
            INIT_41 => X"0000012700000000000000be00000000000000cc000000000000010300000000",
            INIT_42 => X"000000a70000000000000096000000000000008c00000000000000ba00000000",
            INIT_43 => X"000000d000000000000000de0000000000000139000000000000013900000000",
            INIT_44 => X"000000de0000000000000146000000000000012400000000000000ac00000000",
            INIT_45 => X"000000c0000000000000010600000000000000cd00000000000000b000000000",
            INIT_46 => X"0000016200000000000000a000000000000000b8000000000000008500000000",
            INIT_47 => X"000000e200000000000000c40000000000000114000000000000014600000000",
            INIT_48 => X"0000009900000000000000bd00000000000000c600000000000000cc00000000",
            INIT_49 => X"00000061000000000000009e00000000000000a800000000000000ec00000000",
            INIT_4A => X"00000149000000000000014900000000000000b7000000000000008400000000",
            INIT_4B => X"000000a800000000000000f500000000000000ca000000000000012a00000000",
            INIT_4C => X"000000b600000000000000d5000000000000011700000000000000b300000000",
            INIT_4D => X"000000b200000000000000610000000000000043000000000000009b00000000",
            INIT_4E => X"0000012e0000000000000146000000000000010900000000000000c800000000",
            INIT_4F => X"0000010f0000000000000109000000000000018d00000000000000d400000000",
            INIT_50 => X"00000058000000000000009100000000000000e9000000000000013700000000",
            INIT_51 => X"000000aa00000000000000ad0000000000000091000000000000006f00000000",
            INIT_52 => X"000001790000000000000128000000000000010e00000000000000cc00000000",
            INIT_53 => X"0000009c00000000000000a300000000000000c700000000000001c800000000",
            INIT_54 => X"00000093000000000000008a0000000000000083000000000000008900000000",
            INIT_55 => X"000000b200000000000000a600000000000000ab000000000000009a00000000",
            INIT_56 => X"000000ff00000000000001c000000000000000e500000000000000b500000000",
            INIT_57 => X"00000087000000000000008c0000000000000097000000000000009500000000",
            INIT_58 => X"000000b400000000000000a1000000000000008f000000000000008500000000",
            INIT_59 => X"0000009500000000000000ae00000000000000b000000000000000aa00000000",
            INIT_5A => X"0000009a00000000000000ac000000000000016a00000000000000bb00000000",
            INIT_5B => X"00000096000000000000008b000000000000008f000000000000009f00000000",
            INIT_5C => X"0000009e000000000000009e00000000000000a300000000000000a200000000",
            INIT_5D => X"000000a3000000000000009500000000000000c100000000000000db00000000",
            INIT_5E => X"0000008f000000000000007c000000000000008b00000000000000ae00000000",
            INIT_5F => X"000000aa00000000000000ad000000000000009d000000000000009200000000",
            INIT_60 => X"000000af00000000000000f300000000000000a7000000000000009000000000",
            INIT_61 => X"0000007b0000000000000078000000000000007e000000000000007600000000",
            INIT_62 => X"0000008500000000000000820000000000000074000000000000007700000000",
            INIT_63 => X"0000006200000000000000620000000000000070000000000000007b00000000",
            INIT_64 => X"000000750000000000000067000000000000006a000000000000006200000000",
            INIT_65 => X"000000770000000000000080000000000000007e000000000000007d00000000",
            INIT_66 => X"0000005f00000000000000790000000000000079000000000000006f00000000",
            INIT_67 => X"0000003f000000000000002e0000000000000026000000000000003400000000",
            INIT_68 => X"00000063000000000000006e0000000000000065000000000000005b00000000",
            INIT_69 => X"00000084000000000000007d0000000000000081000000000000007d00000000",
            INIT_6A => X"00000016000000000000001f0000000000000037000000000000006200000000",
            INIT_6B => X"0000002f00000000000000250000000000000021000000000000003200000000",
            INIT_6C => X"0000007c000000000000001c0000000000000040000000000000005900000000",
            INIT_6D => X"0000004500000000000000420000000000000077000000000000007c00000000",
            INIT_6E => X"0000004100000000000000260000000000000018000000000000002100000000",
            INIT_6F => X"0000003a000000000000001d0000000000000023000000000000003000000000",
            INIT_70 => X"0000005000000000000000740000000000000034000000000000003200000000",
            INIT_71 => X"0000002e000000000000004f0000000000000031000000000000006200000000",
            INIT_72 => X"0000003100000000000000400000000000000000000000000000002100000000",
            INIT_73 => X"000000270000000000000015000000000000001b000000000000001d00000000",
            INIT_74 => X"0000006f000000000000004e0000000000000077000000000000004e00000000",
            INIT_75 => X"000000270000000000000039000000000000005d000000000000005600000000",
            INIT_76 => X"0000002200000000000000360000000000000051000000000000000300000000",
            INIT_77 => X"00000054000000000000001f000000000000000d000000000000001900000000",
            INIT_78 => X"00000040000000000000003d0000000000000075000000000000006900000000",
            INIT_79 => X"0000001300000000000000400000000000000039000000000000007200000000",
            INIT_7A => X"0000001a00000000000000130000000000000029000000000000004f00000000",
            INIT_7B => X"0000002c0000000000000049000000000000002d000000000000002900000000",
            INIT_7C => X"000000500000000000000060000000000000002e000000000000005700000000",
            INIT_7D => X"000000490000000000000031000000000000003c000000000000004300000000",
            INIT_7E => X"00000042000000000000002f000000000000001b000000000000003300000000",
            INIT_7F => X"0000003d000000000000002d0000000000000040000000000000003c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "samplegold_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003200000000000000450000000000000039000000000000003000000000",
            INIT_01 => X"0000003100000000000000550000000000000036000000000000002800000000",
            INIT_02 => X"0000004b000000000000005f000000000000003c000000000000001100000000",
            INIT_03 => X"00000054000000000000000c0000000000000046000000000000003f00000000",
            INIT_04 => X"000000240000000000000042000000000000001c000000000000001500000000",
            INIT_05 => X"00000017000000000000000a0000000000000029000000000000005000000000",
            INIT_06 => X"000000400000000000000039000000000000006c000000000000004e00000000",
            INIT_07 => X"00000024000000000000003e000000000000000e000000000000004600000000",
            INIT_08 => X"000000010000000000000033000000000000004c000000000000002100000000",
            INIT_09 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000003c0000000000000028000000000000000b000000000000001400000000",
            INIT_0B => X"00000000000000000000001b0000000000000073000000000000003b00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000006e000000000000000f0000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000005000000000000000500000000",
            INIT_1B => X"0000000300000000000000050000000000000008000000000000000400000000",
            INIT_1C => X"0000000c00000000000000060000000000000000000000000000000000000000",
            INIT_1D => X"0000000600000000000000000000000000000000000000000000000100000000",
            INIT_1E => X"00000009000000000000001a0000000000000000000000000000000000000000",
            INIT_1F => X"00000008000000000000000b0000000000000000000000000000000a00000000",
            INIT_20 => X"0000001a00000000000000060000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000012000000000000002b000000000000000000000000",
            INIT_23 => X"0000001f00000000000000110000000000000017000000000000000000000000",
            INIT_24 => X"00000000000000000000005a0000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000016000000000000000e00000000",
            INIT_27 => X"0000001600000000000000220000000000000002000000000000003500000000",
            INIT_28 => X"0000001e00000000000000000000000000000048000000000000000000000000",
            INIT_29 => X"0000003400000000000000060000000000000005000000000000000000000000",
            INIT_2A => X"0000000d0000000000000000000000000000001b000000000000003000000000",
            INIT_2B => X"0000000000000000000000270000000000000004000000000000003300000000",
            INIT_2C => X"00000005000000000000002c0000000000000000000000000000003200000000",
            INIT_2D => X"0000002400000000000000320000000000000006000000000000000000000000",
            INIT_2E => X"00000040000000000000003c0000000000000000000000000000004200000000",
            INIT_2F => X"0000003100000000000000140000000000000018000000000000000000000000",
            INIT_30 => X"00000000000000000000003a0000000000000000000000000000001e00000000",
            INIT_31 => X"000000420000000000000027000000000000000c000000000000000000000000",
            INIT_32 => X"00000000000000000000002d0000000000000045000000000000000000000000",
            INIT_33 => X"0000002200000000000000230000000000000019000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_35 => X"000000000000000000000027000000000000000b000000000000005400000000",
            INIT_36 => X"0000000000000000000000000000000000000036000000000000002900000000",
            INIT_37 => X"0000005d0000000000000000000000000000002d000000000000001200000000",
            INIT_38 => X"0000001800000000000000000000000000000016000000000000000000000000",
            INIT_39 => X"0000000000000000000000120000000000000000000000000000001000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_3B => X"0000000000000000000000650000000000000000000000000000000e00000000",
            INIT_3C => X"0000001500000000000000000000000000000006000000000000002800000000",
            INIT_3D => X"000000000000000000000033000000000000000d000000000000000f00000000",
            INIT_3E => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_3F => X"000000560000000000000000000000000000005a000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003e000000000000000e0000000000000000000000000000001300000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003900000000000000610000000000000000000000000000001300000000",
            INIT_44 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000000b000000000000000500000000",
            INIT_47 => X"000000010000000000000000000000000000007f000000000000000c00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000005100000000000000000000000000000000000000000000001600000000",
            INIT_4B => X"00000000000000000000000b0000000000000000000000000000002100000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000002000000000000000080000000000000000000000000000000100000000",
            INIT_4E => X"0000000b00000000000000010000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000002c000000000000001200000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001e00000000000000040000000000000004000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_5C => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_72 => X"0000000000000000000000070000000000000003000000000000003400000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_75 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_7A => X"0000001900000000000000060000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001c0000000000000031000000000000002a000000000000003f00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7E => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000002d0000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "samplegold_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_06 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000050000000000000011000000000000000900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000004000000000000000200000000",
            INIT_0B => X"0000000200000000000000000000000000000000000000000000000700000000",
            INIT_0C => X"00000007000000000000000b0000000000000003000000000000000000000000",
            INIT_0D => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_0E => X"0000001f00000000000000070000000000000000000000000000000400000000",
            INIT_0F => X"0000001f00000000000000000000000000000001000000000000000000000000",
            INIT_10 => X"0000000f000000000000000b0000000000000000000000000000000000000000",
            INIT_11 => X"0000000100000000000000260000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_13 => X"00000000000000000000002a000000000000000b000000000000000000000000",
            INIT_14 => X"0000001500000000000000040000000000000000000000000000000000000000",
            INIT_15 => X"0000000a00000000000000000000000000000039000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_18 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000003a0000000000000000000000000000000f00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000100000000000000000000000000000000000000000000004b00000000",
            INIT_1C => X"0000000c00000000000000000000000000000009000000000000000000000000",
            INIT_1D => X"0000000000000000000000490000000000000000000000000000000000000000",
            INIT_1E => X"0000008100000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000002f000000000000003a000000000000000000000000",
            INIT_22 => X"0000000000000000000000600000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000c0000000000000003000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000002b000000000000001b00000000",
            INIT_26 => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_28 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_29 => X"0000001800000000000000000000000000000000000000000000000100000000",
            INIT_2A => X"000000110000000000000000000000000000000b000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2C => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_2E => X"0000001400000000000000220000000000000004000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_30 => X"0000001a00000000000000000000000000000000000000000000007200000000",
            INIT_31 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000d0000000000000010000000000000000d00000000",
            INIT_33 => X"0000003a00000000000000000000000000000021000000000000001f00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000045000000000000001a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000050000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_42 => X"0000004600000000000000440000000000000045000000000000003f00000000",
            INIT_43 => X"0000004b00000000000000470000000000000041000000000000004300000000",
            INIT_44 => X"0000002d000000000000002a0000000000000034000000000000004300000000",
            INIT_45 => X"00000043000000000000003b000000000000003d000000000000003500000000",
            INIT_46 => X"0000004400000000000000480000000000000049000000000000004800000000",
            INIT_47 => X"0000002200000000000000380000000000000041000000000000004500000000",
            INIT_48 => X"00000015000000000000000e000000000000000e000000000000001100000000",
            INIT_49 => X"00000025000000000000002b0000000000000038000000000000002700000000",
            INIT_4A => X"0000003100000000000000470000000000000049000000000000004400000000",
            INIT_4B => X"0000000d000000000000000d000000000000000e000000000000002000000000",
            INIT_4C => X"00000010000000000000000f0000000000000011000000000000001500000000",
            INIT_4D => X"0000003c0000000000000019000000000000001c000000000000002900000000",
            INIT_4E => X"00000023000000000000001e000000000000003a000000000000004300000000",
            INIT_4F => X"00000019000000000000000c000000000000000b000000000000001500000000",
            INIT_50 => X"00000019000000000000000c000000000000000a000000000000001100000000",
            INIT_51 => X"0000002e000000000000003a0000000000000022000000000000001600000000",
            INIT_52 => X"000000150000000000000020000000000000002c000000000000003b00000000",
            INIT_53 => X"0000001a000000000000001d0000000000000004000000000000000a00000000",
            INIT_54 => X"00000009000000000000000e000000000000000f000000000000000f00000000",
            INIT_55 => X"00000011000000000000002a000000000000003c000000000000001600000000",
            INIT_56 => X"00000014000000000000001d0000000000000026000000000000001e00000000",
            INIT_57 => X"0000000d000000000000000f000000000000001b000000000000000b00000000",
            INIT_58 => X"00000011000000000000000e0000000000000010000000000000000c00000000",
            INIT_59 => X"0000001b000000000000001b0000000000000036000000000000002300000000",
            INIT_5A => X"0000000700000000000000180000000000000017000000000000001f00000000",
            INIT_5B => X"0000000b00000000000000080000000000000010000000000000001400000000",
            INIT_5C => X"0000001600000000000000110000000000000011000000000000001900000000",
            INIT_5D => X"00000016000000000000001f000000000000001c000000000000002300000000",
            INIT_5E => X"0000001700000000000000170000000000000018000000000000000d00000000",
            INIT_5F => X"0000002700000000000000140000000000000008000000000000000f00000000",
            INIT_60 => X"0000000f000000000000000c000000000000000a000000000000000f00000000",
            INIT_61 => X"0000001200000000000000150000000000000009000000000000001700000000",
            INIT_62 => X"0000000800000000000000120000000000000014000000000000001100000000",
            INIT_63 => X"0000000f000000000000003a0000000000000020000000000000000800000000",
            INIT_64 => X"0000001700000000000000000000000000000011000000000000000e00000000",
            INIT_65 => X"00000015000000000000001b000000000000000c000000000000000f00000000",
            INIT_66 => X"0000001400000000000000000000000000000004000000000000001200000000",
            INIT_67 => X"0000000c00000000000000000000000000000035000000000000002d00000000",
            INIT_68 => X"000000190000000000000023000000000000000c000000000000000e00000000",
            INIT_69 => X"0000000000000000000000060000000000000000000000000000000500000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "samplegold_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000150000000000000010000000000000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000003000000000000000600000000",
            INIT_27 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_28 => X"0000000400000000000000020000000000000000000000000000000000000000",
            INIT_29 => X"00000009000000000000000a0000000000000006000000000000000400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2B => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_2C => X"0000000600000000000000030000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000030000000000000006000000000000000700000000",
            INIT_2E => X"0000000500000000000000000000000000000003000000000000000300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_30 => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000002000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000004000000000000001c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000003000000000000000a0000000000000004000000000000000000000000",
            INIT_75 => X"000000000000000000000000000000000000000a000000000000000b00000000",
            INIT_76 => X"000000000000000000000000000000000000001a000000000000002500000000",
            INIT_77 => X"0000000a000000000000001e0000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000005f00000000000000000000000000000000000000000000003800000000",
            INIT_7B => X"0000000000000000000000070000000000000001000000000000003600000000",
            INIT_7C => X"0000000a0000000000000016000000000000001e000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000d000000000000001d0000000000000018000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "samplegold_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000e000000000000002200000000",
            INIT_02 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_04 => X"00000010000000000000000c0000000000000000000000000000000900000000",
            INIT_05 => X"0000001200000000000000180000000000000013000000000000000900000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0A => X"0000000600000000000000070000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0D => X"0000000000000000000000020000000000000002000000000000000a00000000",
            INIT_0E => X"0000000000000000000000000000000000000035000000000000000200000000",
            INIT_0F => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000005c0000000000000080000000000000002e00000000",
            INIT_12 => X"00000029000000000000000d0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000013000000000000003400000000",
            INIT_14 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"0000000a00000000000000040000000000000005000000000000000a00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000500000000000000010000000000000002000000000000000500000000",
            INIT_1A => X"0000000000000000000000190000000000000013000000000000000c00000000",
            INIT_1B => X"0000000300000000000000070000000000000023000000000000000000000000",
            INIT_1C => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000700000000000000010000000000000006000000000000001100000000",
            INIT_1E => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000030000000000000009000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000a000000000000001b0000000000000014000000000000000000000000",
            INIT_22 => X"0000000e0000000000000023000000000000002c000000000000000600000000",
            INIT_23 => X"0000003400000000000000340000000000000032000000000000003300000000",
            INIT_24 => X"0000003900000000000000350000000000000030000000000000003700000000",
            INIT_25 => X"000000280000000000000025000000000000002c000000000000003600000000",
            INIT_26 => X"00000037000000000000002f000000000000002d000000000000002900000000",
            INIT_27 => X"0000003700000000000000340000000000000038000000000000003400000000",
            INIT_28 => X"00000020000000000000002a0000000000000029000000000000003400000000",
            INIT_29 => X"0000002100000000000000170000000000000013000000000000001f00000000",
            INIT_2A => X"00000035000000000000001e000000000000002d000000000000002b00000000",
            INIT_2B => X"0000003800000000000000390000000000000037000000000000003600000000",
            INIT_2C => X"000000210000000000000013000000000000001a000000000000001600000000",
            INIT_2D => X"00000021000000000000000f000000000000000a000000000000000100000000",
            INIT_2E => X"00000032000000000000003d0000000000000000000000000000002d00000000",
            INIT_2F => X"000000130000000000000028000000000000002b000000000000003a00000000",
            INIT_30 => X"000000000000000000000023000000000000000f000000000000000600000000",
            INIT_31 => X"00000037000000000000000e0000000000000004000000000000000c00000000",
            INIT_32 => X"0000003e00000000000000210000000000000025000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000a000000000000000f00000000",
            INIT_34 => X"00000000000000000000000b000000000000002b000000000000000900000000",
            INIT_35 => X"0000000000000000000000250000000000000009000000000000001100000000",
            INIT_36 => X"00000018000000000000001d0000000000000012000000000000000e00000000",
            INIT_37 => X"0000000300000000000000070000000000000000000000000000000000000000",
            INIT_38 => X"0000001400000000000000000000000000000000000000000000003b00000000",
            INIT_39 => X"000000040000000000000000000000000000000c000000000000000900000000",
            INIT_3A => X"0000001700000000000000340000000000000018000000000000001900000000",
            INIT_3B => X"0000003900000000000000000000000000000000000000000000000400000000",
            INIT_3C => X"0000001100000000000000130000000000000000000000000000000000000000",
            INIT_3D => X"0000000d00000000000000000000000000000000000000000000000700000000",
            INIT_3E => X"000000000000000000000017000000000000002d000000000000001500000000",
            INIT_3F => X"0000000000000000000000310000000000000000000000000000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000000c0000000000000014000000000000000000000000",
            INIT_41 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000f000000000000000a0000000000000013000000000000000300000000",
            INIT_43 => X"00000000000000000000000e0000000000000020000000000000001b00000000",
            INIT_44 => X"0000000000000000000000300000000000000026000000000000001400000000",
            INIT_45 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_46 => X"0000000500000000000000050000000000000019000000000000000800000000",
            INIT_47 => X"00000020000000000000000e0000000000000002000000000000000400000000",
            INIT_48 => X"0000000000000000000000110000000000000029000000000000003300000000",
            INIT_49 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_4A => X"0000000400000000000000000000000000000000000000000000000700000000",
            INIT_4B => X"00000015000000000000000b0000000000000004000000000000000700000000",
            INIT_4C => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"00000000000000000000000b0000000000000008000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000f0000000000000003000000000000000e000000000000000000000000",
            INIT_66 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_69 => X"0000000600000000000000070000000000000008000000000000000700000000",
            INIT_6A => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_6B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_6D => X"0000000000000000000000050000000000000000000000000000000200000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000002000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_70 => X"0000000c00000000000000180000000000000000000000000000000c00000000",
            INIT_71 => X"0000000900000000000000000000000000000005000000000000000200000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_73 => X"0000000f00000000000000000000000000000015000000000000000000000000",
            INIT_74 => X"0000000200000000000000050000000000000017000000000000000000000000",
            INIT_75 => X"0000001800000000000000110000000000000000000000000000000000000000",
            INIT_76 => X"0000000400000000000000000000000000000000000000000000000300000000",
            INIT_77 => X"0000000000000000000000000000000000000015000000000000002500000000",
            INIT_78 => X"000000080000000000000004000000000000000c000000000000000e00000000",
            INIT_79 => X"0000002200000000000000230000000000000023000000000000000000000000",
            INIT_7A => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000001000000000000001700000000",
            INIT_7D => X"0000001000000000000000290000000000000021000000000000001900000000",
            INIT_7E => X"0000000200000000000000000000000000000000000000000000001100000000",
            INIT_7F => X"0000000700000000000000200000000000000007000000000000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "samplegold_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000f0000000000000000000000000000002c000000000000001600000000",
            INIT_02 => X"0000002f000000000000003c0000000000000029000000000000000b00000000",
            INIT_03 => X"00000034000000000000001f0000000000000011000000000000001800000000",
            INIT_04 => X"000000320000000000000067000000000000002a000000000000003100000000",
            INIT_05 => X"0000005000000000000000710000000000000010000000000000001100000000",
            INIT_06 => X"0000004500000000000000460000000000000048000000000000004d00000000",
            INIT_07 => X"0000005700000000000000510000000000000053000000000000004f00000000",
            INIT_08 => X"0000000a0000000000000059000000000000006f000000000000005400000000",
            INIT_09 => X"0000004f0000000000000048000000000000004d000000000000004500000000",
            INIT_0A => X"00000052000000000000004a0000000000000049000000000000004900000000",
            INIT_0B => X"0000005400000000000000600000000000000061000000000000005300000000",
            INIT_0C => X"0000006600000000000000440000000000000062000000000000006f00000000",
            INIT_0D => X"0000004b000000000000004b000000000000004a000000000000004100000000",
            INIT_0E => X"0000006700000000000000610000000000000052000000000000004d00000000",
            INIT_0F => X"0000006f000000000000008a000000000000005d000000000000006500000000",
            INIT_10 => X"00000051000000000000005a0000000000000063000000000000006700000000",
            INIT_11 => X"00000048000000000000004b0000000000000056000000000000005300000000",
            INIT_12 => X"000000450000000000000054000000000000005b000000000000004e00000000",
            INIT_13 => X"0000003900000000000000380000000000000071000000000000006d00000000",
            INIT_14 => X"0000003600000000000000340000000000000036000000000000003900000000",
            INIT_15 => X"0000002d0000000000000034000000000000003f000000000000003e00000000",
            INIT_16 => X"00000030000000000000002f0000000000000030000000000000002c00000000",
            INIT_17 => X"0000003b000000000000003b0000000000000036000000000000002c00000000",
            INIT_18 => X"00000029000000000000001c0000000000000036000000000000003900000000",
            INIT_19 => X"00000000000000000000000b000000000000002b000000000000003300000000",
            INIT_1A => X"0000002d0000000000000030000000000000001d000000000000000300000000",
            INIT_1B => X"0000003b000000000000003c0000000000000043000000000000002700000000",
            INIT_1C => X"0000000900000000000000160000000000000028000000000000003c00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1E => X"00000000000000000000002e000000000000001c000000000000000000000000",
            INIT_1F => X"0000002600000000000000370000000000000036000000000000001c00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_22 => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000029000000000000002100000000",
            INIT_24 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001f00000000000000000000000000000000000000000000001700000000",
            INIT_27 => X"00000000000000000000000a000000000000001d000000000000002900000000",
            INIT_28 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000019000000000000002a0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000007000000000000001700000000",
            INIT_2C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000f00000000000000090000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_31 => X"000000000000000000000000000000000000000d000000000000000300000000",
            INIT_32 => X"0000000700000000000000020000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_34 => X"0000001200000000000000080000000000000000000000000000001100000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_38 => X"0000001f000000000000001c0000000000000009000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"00000048000000000000004b000000000000004b000000000000004400000000",
            INIT_4D => X"000000470000000000000051000000000000004e000000000000004200000000",
            INIT_4E => X"000000390000000000000033000000000000002e000000000000003700000000",
            INIT_4F => X"000000480000000000000049000000000000003f000000000000004000000000",
            INIT_50 => X"0000001e000000000000004e000000000000004b000000000000004d00000000",
            INIT_51 => X"0000001500000000000000260000000000000034000000000000004c00000000",
            INIT_52 => X"000000350000000000000018000000000000000c000000000000000700000000",
            INIT_53 => X"0000004e0000000000000035000000000000001a000000000000003d00000000",
            INIT_54 => X"000000240000000000000019000000000000004e000000000000004c00000000",
            INIT_55 => X"0000001000000000000000000000000000000023000000000000001800000000",
            INIT_56 => X"0000002a00000000000000220000000000000002000000000000001000000000",
            INIT_57 => X"00000048000000000000004c0000000000000014000000000000000600000000",
            INIT_58 => X"0000001f0000000000000012000000000000002e000000000000002d00000000",
            INIT_59 => X"0000001200000000000000090000000000000019000000000000000800000000",
            INIT_5A => X"0000001f0000000000000020000000000000000f000000000000000a00000000",
            INIT_5B => X"000000110000000000000059000000000000004f000000000000000000000000",
            INIT_5C => X"0000000000000000000000120000000000000010000000000000002c00000000",
            INIT_5D => X"00000006000000000000001a0000000000000015000000000000001f00000000",
            INIT_5E => X"0000000000000000000000330000000000000019000000000000000700000000",
            INIT_5F => X"0000003900000000000000000000000000000033000000000000005600000000",
            INIT_60 => X"0000000e0000000000000000000000000000001a000000000000000400000000",
            INIT_61 => X"0000000b000000000000000c000000000000001a000000000000001400000000",
            INIT_62 => X"0000004100000000000000000000000000000047000000000000001200000000",
            INIT_63 => X"00000003000000000000001b0000000000000000000000000000003100000000",
            INIT_64 => X"0000001700000000000000000000000000000008000000000000001700000000",
            INIT_65 => X"0000001b000000000000000e0000000000000007000000000000001200000000",
            INIT_66 => X"00000020000000000000002f0000000000000000000000000000003100000000",
            INIT_67 => X"00000009000000000000000e000000000000000c000000000000002d00000000",
            INIT_68 => X"0000000e000000000000000f0000000000000002000000000000001c00000000",
            INIT_69 => X"0000001100000000000000350000000000000011000000000000000d00000000",
            INIT_6A => X"0000002c0000000000000001000000000000001c000000000000000000000000",
            INIT_6B => X"0000001e0000000000000000000000000000001b000000000000001100000000",
            INIT_6C => X"0000000a000000000000000a0000000000000019000000000000000000000000",
            INIT_6D => X"000000070000000000000004000000000000003c000000000000002200000000",
            INIT_6E => X"0000002200000000000000250000000000000000000000000000000200000000",
            INIT_6F => X"0000001c000000000000001b0000000000000000000000000000001a00000000",
            INIT_70 => X"0000002300000000000000080000000000000009000000000000000000000000",
            INIT_71 => X"00000000000000000000000d0000000000000000000000000000003900000000",
            INIT_72 => X"00000000000000000000001f0000000000000003000000000000000e00000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000080000000000000000000000000000001c000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "samplegold_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000005c000000000000005c000000000000005c000000000000005d00000000",
            INIT_05 => X"0000005c000000000000005c000000000000005c000000000000005c00000000",
            INIT_06 => X"0000005c000000000000005e000000000000005d000000000000005c00000000",
            INIT_07 => X"0000005e000000000000005c000000000000005c000000000000005b00000000",
            INIT_08 => X"0000005c000000000000005d000000000000005c000000000000005c00000000",
            INIT_09 => X"0000005c000000000000005c000000000000005c000000000000005c00000000",
            INIT_0A => X"0000005c0000000000000057000000000000005b000000000000006c00000000",
            INIT_0B => X"0000005e000000000000005f000000000000005c000000000000005c00000000",
            INIT_0C => X"0000005e000000000000005c000000000000005c000000000000005d00000000",
            INIT_0D => X"0000005600000000000000640000000000000067000000000000005d00000000",
            INIT_0E => X"0000005d000000000000005e000000000000005c000000000000005200000000",
            INIT_0F => X"0000005c000000000000005d0000000000000058000000000000005d00000000",
            INIT_10 => X"000000560000000000000067000000000000005f000000000000005c00000000",
            INIT_11 => X"000000420000000000000048000000000000004c000000000000005900000000",
            INIT_12 => X"0000005d000000000000005d000000000000005e000000000000004500000000",
            INIT_13 => X"0000005d0000000000000056000000000000005a000000000000006600000000",
            INIT_14 => X"0000005600000000000000500000000000000053000000000000005e00000000",
            INIT_15 => X"0000007500000000000000730000000000000064000000000000005b00000000",
            INIT_16 => X"00000038000000000000005e0000000000000055000000000000006c00000000",
            INIT_17 => X"00000062000000000000005e0000000000000054000000000000004000000000",
            INIT_18 => X"00000069000000000000006f0000000000000072000000000000006e00000000",
            INIT_19 => X"00000041000000000000003a0000000000000043000000000000006100000000",
            INIT_1A => X"00000062000000000000006b000000000000005b000000000000003f00000000",
            INIT_1B => X"0000004a00000000000000560000000000000048000000000000005300000000",
            INIT_1C => X"000000620000000000000031000000000000001f000000000000002900000000",
            INIT_1D => X"0000007000000000000000640000000000000075000000000000007000000000",
            INIT_1E => X"00000040000000000000002d000000000000001d000000000000006000000000",
            INIT_1F => X"0000003500000000000000350000000000000047000000000000004400000000",
            INIT_20 => X"0000004000000000000000530000000000000064000000000000006500000000",
            INIT_21 => X"00000041000000000000002a000000000000002a000000000000002c00000000",
            INIT_22 => X"000000400000000000000035000000000000003d000000000000000000000000",
            INIT_23 => X"0000005900000000000000650000000000000069000000000000005b00000000",
            INIT_24 => X"00000064000000000000005d000000000000005b000000000000004d00000000",
            INIT_25 => X"0000005700000000000000590000000000000069000000000000006800000000",
            INIT_26 => X"0000006f0000000000000070000000000000006f000000000000006f00000000",
            INIT_27 => X"0000005200000000000000530000000000000060000000000000006400000000",
            INIT_28 => X"0000003b00000000000000480000000000000050000000000000005100000000",
            INIT_29 => X"00000032000000000000002d000000000000003f000000000000003d00000000",
            INIT_2A => X"00000053000000000000004b0000000000000047000000000000004000000000",
            INIT_2B => X"00000053000000000000005a000000000000005f000000000000005e00000000",
            INIT_2C => X"0000002d0000000000000034000000000000003d000000000000004600000000",
            INIT_2D => X"000000120000000000000000000000000000000b000000000000003300000000",
            INIT_2E => X"0000000400000000000000000000000000000000000000000000000800000000",
            INIT_2F => X"0000000f00000000000000110000000000000010000000000000001000000000",
            INIT_30 => X"000000250000000000000034000000000000003d000000000000001800000000",
            INIT_31 => X"0000000300000000000000050000000000000002000000000000000000000000",
            INIT_32 => X"0000004700000000000000060000000000000000000000000000000000000000",
            INIT_33 => X"0000002c00000000000000480000000000000041000000000000003c00000000",
            INIT_34 => X"0000000d000000000000002c0000000000000020000000000000001200000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000001b00000000000000140000000000000000000000000000000000000000",
            INIT_37 => X"00000020000000000000000d0000000000000000000000000000000300000000",
            INIT_38 => X"0000000000000000000000090000000000000036000000000000002600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000002a000000000000001f000000000000001d000000000000001a00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_4A => X"000000000000000000000000000000000000002b000000000000000a00000000",
            INIT_4B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_4F => X"000000000000000000000001000000000000001a000000000000000f00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_53 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_54 => X"00000047000000000000002e000000000000000c000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000002400000000000000260000000000000000000000000000000000000000",
            INIT_57 => X"000000030000000000000000000000000000001b000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_59 => X"0000001600000000000000140000000000000003000000000000000000000000",
            INIT_5A => X"0000000e000000000000000000000000000000a2000000000000001900000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000280000000000000000000000000000000f000000000000000d00000000",
            INIT_66 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"00000020000000000000001c0000000000000019000000000000003300000000",
            INIT_68 => X"000000000000000000000006000000000000002f000000000000003000000000",
            INIT_69 => X"0000000000000000000000060000000000000000000000000000001900000000",
            INIT_6A => X"0000005e00000000000000010000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000001a00000000000000120000000000000010000000000000000000000000",
            INIT_6D => X"0000000000000000000000050000000000000002000000000000000000000000",
            INIT_6E => X"0000000500000000000000420000000000000002000000000000000200000000",
            INIT_6F => X"0000001e00000000000000230000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000000f000000000000000e000000000000000000000000",
            INIT_71 => X"0000000700000000000000050000000000000006000000000000000100000000",
            INIT_72 => X"00000022000000000000000b0000000000000023000000000000000a00000000",
            INIT_73 => X"0000000700000000000000000000000000000004000000000000003200000000",
            INIT_74 => X"000000000000000000000000000000000000000e000000000000000b00000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "samplegold_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000010000000000000002000000000000000c000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000006000000000000000200000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000050000000000000033000000000000005f000000000000006c00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2C => X"000001b900000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"000001b600000000000001b600000000000001b600000000000001b600000000",
            INIT_2E => X"000001b400000000000001b800000000000001b700000000000001b700000000",
            INIT_2F => X"000001b600000000000001b600000000000001b300000000000001b700000000",
            INIT_30 => X"000001b700000000000001ba00000000000001b600000000000001b600000000",
            INIT_31 => X"000001b600000000000001b600000000000001b700000000000001b700000000",
            INIT_32 => X"000001af00000000000001b600000000000001b700000000000001b600000000",
            INIT_33 => X"000001b600000000000001b8000000000000019c000000000000017200000000",
            INIT_34 => X"000001b700000000000001b500000000000001b500000000000001b700000000",
            INIT_35 => X"000001b100000000000001bb00000000000001b800000000000001b900000000",
            INIT_36 => X"0000014d0000000000000158000000000000018300000000000001ba00000000",
            INIT_37 => X"000001ba00000000000001b800000000000001b9000000000000017e00000000",
            INIT_38 => X"000001ba00000000000001b600000000000001b200000000000001a300000000",
            INIT_39 => X"000001a8000000000000018700000000000001c100000000000001bc00000000",
            INIT_3A => X"0000017c000000000000015d0000000000000172000000000000017100000000",
            INIT_3B => X"0000011d00000000000001bb00000000000001b700000000000001b800000000",
            INIT_3C => X"000001b700000000000001b3000000000000016e000000000000011d00000000",
            INIT_3D => X"000001ac00000000000001b000000000000001a400000000000001b000000000",
            INIT_3E => X"000001550000000000000175000000000000019f00000000000001b000000000",
            INIT_3F => X"0000016b000000000000015700000000000001b3000000000000014400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000001800000000000000188000000000000018a00000000000001aa00000000",
            INIT_41 => X"000001a3000000000000017c0000000000000166000000000000015700000000",
            INIT_42 => X"000001560000000000000165000000000000016b000000000000017300000000",
            INIT_43 => X"0000012c00000000000000f000000000000000f300000000000001b000000000",
            INIT_44 => X"000000a80000000000000103000000000000019b000000000000014a00000000",
            INIT_45 => X"0000019800000000000001ac000000000000013a00000000000000d200000000",
            INIT_46 => X"0000014d000000000000016d0000000000000154000000000000017600000000",
            INIT_47 => X"00000118000000000000010200000000000000e7000000000000004c00000000",
            INIT_48 => X"0000019f00000000000001630000000000000150000000000000015900000000",
            INIT_49 => X"000000ed00000000000001090000000000000128000000000000014d00000000",
            INIT_4A => X"000000450000000000000148000000000000011900000000000000fe00000000",
            INIT_4B => X"0000019c000000000000017a0000000000000153000000000000017c00000000",
            INIT_4C => X"0000014e000000000000016c000000000000019200000000000001a900000000",
            INIT_4D => X"0000012e000000000000014e0000000000000145000000000000015200000000",
            INIT_4E => X"0000011300000000000001020000000000000114000000000000012900000000",
            INIT_4F => X"00000122000000000000011f000000000000011c000000000000011900000000",
            INIT_50 => X"000000ec00000000000001030000000000000104000000000000012600000000",
            INIT_51 => X"000000c700000000000000b900000000000000c800000000000000e600000000",
            INIT_52 => X"00000058000000000000003a000000000000004500000000000000dd00000000",
            INIT_53 => X"0000007e00000000000000620000000000000052000000000000004a00000000",
            INIT_54 => X"00000078000000000000008a0000000000000096000000000000008900000000",
            INIT_55 => X"000000d800000000000000bd0000000000000090000000000000007c00000000",
            INIT_56 => X"0000003800000000000000590000000000000011000000000000001c00000000",
            INIT_57 => X"0000009000000000000000270000000000000000000000000000000500000000",
            INIT_58 => X"000000b2000000000000007e0000000000000065000000000000006800000000",
            INIT_59 => X"0000003400000000000000de00000000000000cf00000000000000dd00000000",
            INIT_5A => X"00000000000000000000000e0000000000000011000000000000000000000000",
            INIT_5B => X"000000fc00000000000000fa0000000000000042000000000000000000000000",
            INIT_5C => X"0000009f000000000000009600000000000000cd00000000000000ee00000000",
            INIT_5D => X"000000000000000000000072000000000000010a00000000000000d800000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000004700000000000000750000000000000080000000000000000700000000",
            INIT_60 => X"000000e800000000000000d900000000000000b4000000000000006200000000",
            INIT_61 => X"00000000000000000000000d0000000000000070000000000000012500000000",
            INIT_62 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000d60000000000000091000000000000003f000000000000002b00000000",
            INIT_64 => X"00000135000000000000010300000000000000de00000000000000d200000000",
            INIT_65 => X"0000005e000000000000005e000000000000005e000000000000005f00000000",
            INIT_66 => X"00000060000000000000005e000000000000005e000000000000005e00000000",
            INIT_67 => X"0000005e000000000000005c000000000000005d000000000000005f00000000",
            INIT_68 => X"0000005f000000000000005e000000000000005e000000000000005e00000000",
            INIT_69 => X"0000005e000000000000005e000000000000005e000000000000005e00000000",
            INIT_6A => X"00000060000000000000005f000000000000005e000000000000005e00000000",
            INIT_6B => X"0000005e000000000000005b0000000000000050000000000000006400000000",
            INIT_6C => X"0000005f000000000000005f000000000000005e000000000000005e00000000",
            INIT_6D => X"00000062000000000000005e000000000000005f000000000000005e00000000",
            INIT_6E => X"0000004d00000000000000550000000000000063000000000000005b00000000",
            INIT_6F => X"0000005e0000000000000060000000000000004a000000000000003d00000000",
            INIT_70 => X"0000005d00000000000000560000000000000053000000000000005f00000000",
            INIT_71 => X"00000054000000000000006a0000000000000061000000000000006000000000",
            INIT_72 => X"0000001d000000000000002a0000000000000033000000000000005a00000000",
            INIT_73 => X"0000005d000000000000005b000000000000005b000000000000003300000000",
            INIT_74 => X"0000005f00000000000000570000000000000044000000000000003d00000000",
            INIT_75 => X"0000005d000000000000004e0000000000000063000000000000006100000000",
            INIT_76 => X"0000004e00000000000000560000000000000056000000000000004d00000000",
            INIT_77 => X"0000001d000000000000005a0000000000000044000000000000005200000000",
            INIT_78 => X"0000006200000000000000600000000000000046000000000000001c00000000",
            INIT_79 => X"0000004e000000000000005e000000000000005e000000000000006d00000000",
            INIT_7A => X"0000002500000000000000280000000000000036000000000000004e00000000",
            INIT_7B => X"0000002f00000000000000350000000000000054000000000000002100000000",
            INIT_7C => X"00000012000000000000004d000000000000003a000000000000005400000000",
            INIT_7D => X"0000005e00000000000000280000000000000000000000000000000000000000",
            INIT_7E => X"0000004f000000000000005e000000000000005d000000000000006100000000",
            INIT_7F => X"0000001c00000000000000090000000000000000000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "samplegold_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c000000000000002d0000000000000047000000000000003200000000",
            INIT_01 => X"0000002200000000000000360000000000000042000000000000004000000000",
            INIT_02 => X"00000023000000000000001a000000000000000e000000000000001700000000",
            INIT_03 => X"00000037000000000000002c0000000000000043000000000000000000000000",
            INIT_04 => X"00000054000000000000005c0000000000000056000000000000004500000000",
            INIT_05 => X"0000003800000000000000320000000000000033000000000000002b00000000",
            INIT_06 => X"0000000c00000000000000300000000000000030000000000000003300000000",
            INIT_07 => X"00000028000000000000002e000000000000002b000000000000003200000000",
            INIT_08 => X"0000001b00000000000000140000000000000020000000000000002a00000000",
            INIT_09 => X"00000003000000000000000e000000000000000e000000000000000f00000000",
            INIT_0A => X"0000000000000000000000000000000000000011000000000000000a00000000",
            INIT_0B => X"0000000c000000000000000d0000000000000006000000000000000300000000",
            INIT_0C => X"00000005000000000000000b000000000000000c000000000000000e00000000",
            INIT_0D => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000500000000000000000000000000000000000000000000001700000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000200000000000000020000000000000001c000000000000000600000000",
            INIT_12 => X"0000000a000000000000000b0000000000000000000000000000000000000000",
            INIT_13 => X"0000006a00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000003300000000000000480000000000000058000000000000005c00000000",
            INIT_15 => X"0000001a0000000000000027000000000000001f000000000000002b00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000007900000000000000850000000000000005000000000000000000000000",
            INIT_18 => X"00000028000000000000001f0000000000000024000000000000003f00000000",
            INIT_19 => X"000000000000000000000020000000000000002e000000000000002500000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000190000000000000021000000000000002c000000000000000000000000",
            INIT_1C => X"00000028000000000000002a000000000000002b000000000000002f00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000001e000000000000000100000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000a00000000000000130000000000000000000000000000000100000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000e00000000000000020000000000000024000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_2E => X"0000000b000000000000000c0000000000000000000000000000000300000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_32 => X"00000005000000000000000f000000000000000f000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_34 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000006200000000",
            INIT_36 => X"00000000000000000000000a0000000000000007000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001900000000000000000000000000000000000000000000000a00000000",
            INIT_39 => X"0000000d00000000000000010000000000000011000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_3E => X"0000000200000000000000000000000000000000000000000000000900000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000005000000000000000b0000000000000000000000000000000000000000",
            INIT_41 => X"0000001100000000000000000000000000000017000000000000000000000000",
            INIT_42 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_44 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_46 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_47 => X"00000000000000000000000f0000000000000022000000000000001600000000",
            INIT_48 => X"000000000000000000000004000000000000001d000000000000000000000000",
            INIT_49 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000000c000000000000001800000000",
            INIT_4C => X"000000120000000000000023000000000000001e000000000000001a00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_4E => X"0000000700000000000000000000000000000004000000000000006000000000",
            INIT_4F => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_51 => X"0000005500000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000200000000000000040000000000000005000000000000000d00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000004100000000000000400000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000001400000000000000150000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"000000000000000000000029000000000000003c000000000000003500000000",
            INIT_6D => X"0000000e00000000000000100000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001100000000000000060000000000000000000000000000000000000000",
            INIT_70 => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_71 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000000b0000000000000019000000000000002000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000001900000000000000140000000000000000000000000000001600000000",
            INIT_78 => X"0000000d000000000000001d000000000000001a000000000000002000000000",
            INIT_79 => X"000000080000000000000008000000000000000e000000000000001300000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_7B => X"000000480000000000000041000000000000003e000000000000003f00000000",
            INIT_7C => X"00000032000000000000003d0000000000000047000000000000004900000000",
            INIT_7D => X"0000001100000000000000230000000000000025000000000000002700000000",
            INIT_7E => X"0000000500000000000000000000000000000000000000000000000600000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "samplegold_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"00000005000000000000000f0000000000000020000000000000002400000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_05 => X"000000000000000000000008000000000000001f000000000000000000000000",
            INIT_06 => X"0000000600000000000000050000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000070000000000000008000000000000000c00000000",
            INIT_08 => X"0000000000000000000000180000000000000006000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0B => X"0000000900000000000000000000000000000001000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000002000000000000001100000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_1B => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000027000000000000001400000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000110000000000000008000000000000000700000000",
            INIT_23 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000e000000000000001f0000000000000000000000000000000000000000",
            INIT_25 => X"0000000800000000000000000000000000000000000000000000001800000000",
            INIT_26 => X"0000000000000000000000000000000000000021000000000000001e00000000",
            INIT_27 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002800000000000000000000000000000017000000000000003800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000009500000000000000000000000000000003000000000000000200000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000030000000000000001000000000000000300000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000150000000000000000000000000000000a00000000",
            INIT_34 => X"0000000d000000000000000f0000000000000006000000000000000000000000",
            INIT_35 => X"0000000300000000000000000000000000000002000000000000000800000000",
            INIT_36 => X"0000000800000000000000000000000000000012000000000000000700000000",
            INIT_37 => X"0000000000000000000000000000000000000026000000000000000000000000",
            INIT_38 => X"00000000000000000000004f000000000000000c000000000000000000000000",
            INIT_39 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000160000000000000002000000000000000000000000",
            INIT_3B => X"000000000000000000000000000000000000000b000000000000000c00000000",
            INIT_3C => X"0000000000000000000000000000000000000059000000000000000400000000",
            INIT_3D => X"0000001100000000000000130000000000000000000000000000000000000000",
            INIT_3E => X"0000000200000000000000000000000000000018000000000000000e00000000",
            INIT_3F => X"0000000500000000000000040000000000000002000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002900000000000000160000000000000023000000000000003400000000",
            INIT_41 => X"0000000f0000000000000001000000000000000e000000000000002000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_43 => X"0000001800000000000000040000000000000002000000000000000000000000",
            INIT_44 => X"000000000000000000000018000000000000001e000000000000001e00000000",
            INIT_45 => X"0000000f000000000000000a0000000000000007000000000000000000000000",
            INIT_46 => X"0000001400000000000000140000000000000014000000000000001400000000",
            INIT_47 => X"0000001500000000000000130000000000000014000000000000001400000000",
            INIT_48 => X"0000001300000000000000120000000000000012000000000000001500000000",
            INIT_49 => X"0000001300000000000000140000000000000014000000000000001400000000",
            INIT_4A => X"0000001300000000000000130000000000000013000000000000001300000000",
            INIT_4B => X"0000001100000000000000130000000000000013000000000000001300000000",
            INIT_4C => X"00000014000000000000000e0000000000000001000000000000000a00000000",
            INIT_4D => X"0000001300000000000000130000000000000013000000000000001300000000",
            INIT_4E => X"0000001400000000000000140000000000000014000000000000001300000000",
            INIT_4F => X"000000000000000000000000000000000000000d000000000000001000000000",
            INIT_50 => X"0000001300000000000000130000000000000004000000000000000000000000",
            INIT_51 => X"00000011000000000000000c0000000000000009000000000000001300000000",
            INIT_52 => X"0000000c00000000000000140000000000000014000000000000001300000000",
            INIT_53 => X"00000009000000000000000a000000000000000c000000000000001100000000",
            INIT_54 => X"00000010000000000000000e000000000000000c000000000000000800000000",
            INIT_55 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_56 => X"0000001300000000000000120000000000000013000000000000001300000000",
            INIT_57 => X"000000000000000000000005000000000000000f000000000000001100000000",
            INIT_58 => X"00000016000000000000000c0000000000000000000000000000000000000000",
            INIT_59 => X"00000009000000000000000b0000000000000011000000000000001700000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5B => X"000000130000000000000012000000000000000c000000000000000600000000",
            INIT_5C => X"000000000000000000000000000000000000000b000000000000000c00000000",
            INIT_5D => X"00000000000000000000000b0000000000000006000000000000000000000000",
            INIT_5E => X"00000010000000000000000c0000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000020000000000000001000000000000000900000000",
            INIT_60 => X"00000002000000000000000a0000000000000000000000000000000000000000",
            INIT_61 => X"0000001e000000000000001a0000000000000007000000000000000200000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_63 => X"0000000800000000000000050000000000000000000000000000000000000000",
            INIT_64 => X"0000001400000000000000130000000000000010000000000000000000000000",
            INIT_65 => X"0000000400000000000000000000000000000004000000000000000a00000000",
            INIT_66 => X"0000000000000000000000000000000000000001000000000000000400000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000c00000000000000000000000000000001000000000000000700000000",
            INIT_70 => X"0000000000000000000000000000000000000004000000000000000c00000000",
            INIT_71 => X"0000000900000000000000000000000000000000000000000000000500000000",
            INIT_72 => X"0000000d000000000000000a0000000000000014000000000000001800000000",
            INIT_73 => X"0000000500000000000000000000000000000000000000000000000d00000000",
            INIT_74 => X"00000041000000000000000a0000000000000001000000000000000300000000",
            INIT_75 => X"0000000d00000000000000220000000000000041000000000000004d00000000",
            INIT_76 => X"0000000e000000000000000a000000000000000d000000000000001300000000",
            INIT_77 => X"0000000300000000000000030000000000000001000000000000000400000000",
            INIT_78 => X"0000003e000000000000004a0000000000000010000000000000000300000000",
            INIT_79 => X"0000000d0000000000000018000000000000001a000000000000001b00000000",
            INIT_7A => X"0000000b000000000000000b0000000000000007000000000000000900000000",
            INIT_7B => X"0000000500000000000000060000000000000005000000000000000700000000",
            INIT_7C => X"00000020000000000000001e000000000000000d000000000000000000000000",
            INIT_7D => X"0000000a000000000000000c000000000000000b000000000000001a00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "samplegold_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000013000000000000001f0000000000000000000000000000000000000000",
            INIT_28 => X"0000002f00000000000000300000000000000029000000000000001600000000",
            INIT_29 => X"0000001a000000000000001c0000000000000021000000000000001d00000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_2B => X"0000001000000000000000230000000000000026000000000000000000000000",
            INIT_2C => X"00000000000000000000002f000000000000002c000000000000001c00000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000002d000000000000002e000000000000002f000000000000001500000000",
            INIT_30 => X"0000000000000000000000100000000000000031000000000000003000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000002c000000000000002a0000000000000029000000000000002500000000",
            INIT_34 => X"000000010000000000000000000000000000001c000000000000002c00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001200000000000000410000000000000032000000000000001c00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "samplegold_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000005500000000000000580000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000260000000000000053000000000000004f000000000000003100000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000800000000000000050000000000000002000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000002a000000000000003900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000046000000000000000000000000",
            INIT_0A => X"00000000000000000000006f0000000000000066000000000000000000000000",
            INIT_0B => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"00000053000000000000001a0000000000000040000000000000002c00000000",
            INIT_0D => X"0000000000000000000000270000000000000048000000000000001a00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_18 => X"0000001d00000000000000130000000000000000000000000000000000000000",
            INIT_19 => X"0000008f00000000000000550000000000000000000000000000000500000000",
            INIT_1A => X"000000540000000000000065000000000000005f000000000000006000000000",
            INIT_1B => X"0000001b000000000000000e0000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000200000000000000170000000000000007000000000000000a00000000",
            INIT_20 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000020000000000000003900000000",
            INIT_23 => X"00000018000000000000001d0000000000000006000000000000000000000000",
            INIT_24 => X"0000000100000000000000180000000000000016000000000000001300000000",
            INIT_25 => X"00000002000000000000002d0000000000000044000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_36 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000100000000000000000000000000000000000000000000000f00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000000000000000000000a0000000000000015000000000000000f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000003000000000000000a0000000000000015000000000000000000000000",
            INIT_42 => X"0000000100000000000000000000000000000000000000000000001400000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000010000000000000008000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000900000000000000010000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"00000001000000000000001d0000000000000007000000000000000800000000",
            INIT_51 => X"0000001f0000000000000010000000000000000d000000000000000700000000",
            INIT_52 => X"0000000700000000000000030000000000000004000000000000000000000000",
            INIT_53 => X"0000001000000000000000050000000000000000000000000000000000000000",
            INIT_54 => X"0000000a0000000000000014000000000000001a000000000000000b00000000",
            INIT_55 => X"0000000000000000000000300000000000000016000000000000001200000000",
            INIT_56 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000140000000000000013000000000000000a00000000",
            INIT_58 => X"0000001700000000000000140000000000000018000000000000001800000000",
            INIT_59 => X"0000000000000000000000000000000000000025000000000000001800000000",
            INIT_5A => X"00000011000000000000001a0000000000000017000000000000000c00000000",
            INIT_5B => X"0000001c00000000000000000000000000000011000000000000001200000000",
            INIT_5C => X"0000001c000000000000001b000000000000001c000000000000001c00000000",
            INIT_5D => X"000000240000000000000016000000000000001e000000000000002200000000",
            INIT_5E => X"0000001100000000000000130000000000000011000000000000001500000000",
            INIT_5F => X"0000002200000000000000220000000000000022000000000000000f00000000",
            INIT_60 => X"0000002200000000000000220000000000000022000000000000002200000000",
            INIT_61 => X"000000250000000000000024000000000000001f000000000000002200000000",
            INIT_62 => X"0000002200000000000000220000000000000022000000000000002200000000",
            INIT_63 => X"0000002300000000000000220000000000000022000000000000002300000000",
            INIT_64 => X"0000002200000000000000220000000000000022000000000000002200000000",
            INIT_65 => X"0000001f000000000000002c0000000000000041000000000000002500000000",
            INIT_66 => X"0000002400000000000000220000000000000022000000000000002200000000",
            INIT_67 => X"0000002100000000000000220000000000000021000000000000002300000000",
            INIT_68 => X"0000004100000000000000360000000000000025000000000000002400000000",
            INIT_69 => X"0000002200000000000000290000000000000038000000000000003c00000000",
            INIT_6A => X"0000002800000000000000270000000000000023000000000000002200000000",
            INIT_6B => X"0000003100000000000000220000000000000021000000000000002400000000",
            INIT_6C => X"00000024000000000000001e0000000000000025000000000000001c00000000",
            INIT_6D => X"000000260000000000000029000000000000001c000000000000001b00000000",
            INIT_6E => X"00000024000000000000003e0000000000000050000000000000002400000000",
            INIT_6F => X"0000001d00000000000000230000000000000023000000000000002200000000",
            INIT_70 => X"0000005000000000000000310000000000000023000000000000002100000000",
            INIT_71 => X"00000028000000000000002a000000000000004f000000000000005500000000",
            INIT_72 => X"0000003000000000000000340000000000000015000000000000001700000000",
            INIT_73 => X"0000004d00000000000000550000000000000057000000000000002f00000000",
            INIT_74 => X"0000001300000000000000190000000000000032000000000000003d00000000",
            INIT_75 => X"0000005d000000000000002c0000000000000011000000000000001d00000000",
            INIT_76 => X"0000003d00000000000000150000000000000034000000000000004b00000000",
            INIT_77 => X"0000000500000000000000020000000000000021000000000000003000000000",
            INIT_78 => X"00000042000000000000004f0000000000000049000000000000003700000000",
            INIT_79 => X"0000000d00000000000000170000000000000037000000000000005200000000",
            INIT_7A => X"00000001000000000000001b0000000000000019000000000000002700000000",
            INIT_7B => X"0000003200000000000000440000000000000048000000000000000700000000",
            INIT_7C => X"0000000d00000000000000110000000000000014000000000000002400000000",
            INIT_7D => X"0000001200000000000000300000000000000000000000000000002200000000",
            INIT_7E => X"0000004400000000000000410000000000000035000000000000001e00000000",
            INIT_7F => X"00000049000000000000004e0000000000000035000000000000003d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "samplegold_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004000000000000000580000000000000059000000000000005700000000",
            INIT_01 => X"0000006600000000000000670000000000000062000000000000005d00000000",
            INIT_02 => X"0000004800000000000000580000000000000057000000000000006000000000",
            INIT_03 => X"0000004400000000000000500000000000000041000000000000004a00000000",
            INIT_04 => X"00000030000000000000002d0000000000000035000000000000003a00000000",
            INIT_05 => X"0000004b0000000000000047000000000000003f000000000000002e00000000",
            INIT_06 => X"0000005e00000000000000620000000000000066000000000000005300000000",
            INIT_07 => X"0000002a000000000000003e000000000000004a000000000000005800000000",
            INIT_08 => X"00000005000000000000000c000000000000001b000000000000001e00000000",
            INIT_09 => X"000000050000000000000008000000000000000c000000000000000d00000000",
            INIT_0A => X"0000000e0000000000000015000000000000000e000000000000000000000000",
            INIT_0B => X"0000001400000000000000250000000000000006000000000000000000000000",
            INIT_0C => X"0000000800000000000000070000000000000001000000000000000300000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0E => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000b00000000000000050000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000800000000000000160000000000000008000000000000000700000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000500000000000000080000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000016000000000000000c00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000200000000000000020000000000000005000000000000000f00000000",
            INIT_46 => X"00000022000000000000002f0000000000000035000000000000003f00000000",
            INIT_47 => X"0000000000000000000000000000000000000004000000000000001b00000000",
            INIT_48 => X"0000000600000000000000010000000000000000000000000000000000000000",
            INIT_49 => X"0000004500000000000000010000000000000003000000000000000400000000",
            INIT_4A => X"00000008000000000000002d000000000000005a000000000000006e00000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000002800000000000000140000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000005000000000000001700000000",
            INIT_4F => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000b000000000000000a000000000000000a000000000000000a00000000",
            INIT_51 => X"0000000c000000000000000b000000000000000b000000000000000a00000000",
            INIT_52 => X"0000000a000000000000000b0000000000000006000000000000000900000000",
            INIT_53 => X"0000000a000000000000000c000000000000000a000000000000000a00000000",
            INIT_54 => X"0000000a000000000000000a000000000000000a000000000000000a00000000",
            INIT_55 => X"000000000000000000000006000000000000000a000000000000000b00000000",
            INIT_56 => X"0000000a000000000000000a000000000000000a000000000000000000000000",
            INIT_57 => X"0000000a000000000000000b000000000000000b000000000000000a00000000",
            INIT_58 => X"0000000a0000000000000008000000000000000b000000000000000a00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000a000000000000000b000000000000000c000000000000000000000000",
            INIT_5B => X"0000000c00000000000000090000000000000004000000000000000400000000",
            INIT_5C => X"00000006000000000000000b0000000000000000000000000000000a00000000",
            INIT_5D => X"0000000200000000000000000000000000000001000000000000000a00000000",
            INIT_5E => X"0000000000000000000000090000000000000007000000000000000700000000",
            INIT_5F => X"0000000a000000000000000c0000000000000000000000000000000400000000",
            INIT_60 => X"00000007000000000000000a0000000000000005000000000000000400000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_62 => X"00000006000000000000000c0000000000000005000000000000000c00000000",
            INIT_63 => X"0000000f00000000000000000000000000000010000000000000000000000000",
            INIT_64 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_65 => X"000000010000000000000000000000000000000d000000000000000c00000000",
            INIT_66 => X"0000000400000000000000000000000000000000000000000000000400000000",
            INIT_67 => X"00000000000000000000000d0000000000000000000000000000000d00000000",
            INIT_68 => X"0000000400000000000000040000000000000012000000000000000000000000",
            INIT_69 => X"0000000400000000000000000000000000000005000000000000000100000000",
            INIT_6A => X"0000000000000000000000040000000000000000000000000000000600000000",
            INIT_6B => X"00000000000000000000000d000000000000001b000000000000000500000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000e00000000000000040000000000000001000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_6F => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000000000000000000002000000000000000c000000000000000a00000000",
            INIT_7A => X"0000000000000000000000000000000000000005000000000000000200000000",
            INIT_7B => X"0000000c00000000000000030000000000000000000000000000000000000000",
            INIT_7C => X"0000000d000000000000000b0000000000000000000000000000000200000000",
            INIT_7D => X"0000000800000000000000080000000000000000000000000000000300000000",
            INIT_7E => X"000000320000000000000039000000000000000f000000000000000300000000",
            INIT_7F => X"0000001700000000000000050000000000000006000000000000002200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "samplegold_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000006000000000000000c0000000000000005000000000000000700000000",
            INIT_01 => X"0000000400000000000000050000000000000004000000000000000100000000",
            INIT_02 => X"0000000700000000000000100000000000000014000000000000001800000000",
            INIT_03 => X"0000000d0000000000000008000000000000000d000000000000001800000000",
            INIT_04 => X"00000009000000000000000d0000000000000019000000000000000400000000",
            INIT_05 => X"0000000100000000000000070000000000000008000000000000000700000000",
            INIT_06 => X"0000000e0000000000000018000000000000001e000000000000000000000000",
            INIT_07 => X"00000005000000000000000b000000000000000f000000000000000e00000000",
            INIT_08 => X"0000006900000000000000630000000000000058000000000000006300000000",
            INIT_09 => X"0000006300000000000000640000000000000066000000000000006a00000000",
            INIT_0A => X"0000006000000000000000670000000000000065000000000000005e00000000",
            INIT_0B => X"00000060000000000000005e0000000000000062000000000000006200000000",
            INIT_0C => X"000000610000000000000064000000000000005d000000000000005400000000",
            INIT_0D => X"0000005d000000000000005f0000000000000062000000000000006200000000",
            INIT_0E => X"00000064000000000000005c0000000000000050000000000000007100000000",
            INIT_0F => X"0000004e000000000000005b0000000000000061000000000000006200000000",
            INIT_10 => X"0000005700000000000000560000000000000059000000000000005500000000",
            INIT_11 => X"0000006c00000000000000580000000000000058000000000000005a00000000",
            INIT_12 => X"0000005b00000000000000660000000000000062000000000000004000000000",
            INIT_13 => X"00000058000000000000004b0000000000000059000000000000005b00000000",
            INIT_14 => X"0000004b00000000000000500000000000000052000000000000005700000000",
            INIT_15 => X"00000042000000000000003f0000000000000064000000000000005200000000",
            INIT_16 => X"0000005500000000000000560000000000000041000000000000004900000000",
            INIT_17 => X"00000042000000000000003e0000000000000048000000000000004700000000",
            INIT_18 => X"00000049000000000000004b000000000000004a000000000000004700000000",
            INIT_19 => X"0000001a0000000000000039000000000000003c000000000000003d00000000",
            INIT_1A => X"0000001c00000000000000390000000000000042000000000000003000000000",
            INIT_1B => X"0000002400000000000000200000000000000033000000000000001d00000000",
            INIT_1C => X"000000380000000000000041000000000000003d000000000000002500000000",
            INIT_1D => X"00000042000000000000002a000000000000001d000000000000002e00000000",
            INIT_1E => X"000000390000000000000034000000000000002e000000000000001a00000000",
            INIT_1F => X"00000044000000000000003b0000000000000035000000000000002e00000000",
            INIT_20 => X"0000002f000000000000002f0000000000000038000000000000003e00000000",
            INIT_21 => X"000000310000000000000037000000000000004b000000000000003700000000",
            INIT_22 => X"0000002c00000000000000300000000000000036000000000000004600000000",
            INIT_23 => X"000000560000000000000054000000000000004d000000000000003f00000000",
            INIT_24 => X"00000041000000000000005d0000000000000059000000000000005f00000000",
            INIT_25 => X"000000030000000000000035000000000000003c000000000000003800000000",
            INIT_26 => X"0000005a000000000000004b0000000000000059000000000000005000000000",
            INIT_27 => X"00000049000000000000005e0000000000000068000000000000006500000000",
            INIT_28 => X"0000003a00000000000000290000000000000036000000000000003d00000000",
            INIT_29 => X"0000003c0000000000000038000000000000003e000000000000004100000000",
            INIT_2A => X"0000004e000000000000005c0000000000000050000000000000003000000000",
            INIT_2B => X"0000004f0000000000000055000000000000004c000000000000004600000000",
            INIT_2C => X"0000004e000000000000004b0000000000000046000000000000004600000000",
            INIT_2D => X"00000050000000000000004e0000000000000030000000000000004200000000",
            INIT_2E => X"0000005300000000000000580000000000000056000000000000005300000000",
            INIT_2F => X"00000045000000000000002a000000000000003d000000000000005600000000",
            INIT_30 => X"0000002100000000000000300000000000000040000000000000005200000000",
            INIT_31 => X"00000054000000000000004f000000000000003d000000000000002500000000",
            INIT_32 => X"0000004a0000000000000038000000000000002d000000000000003900000000",
            INIT_33 => X"0000002f000000000000002f0000000000000037000000000000003e00000000",
            INIT_34 => X"0000000f000000000000001d000000000000001c000000000000002a00000000",
            INIT_35 => X"0000004300000000000000480000000000000050000000000000003900000000",
            INIT_36 => X"0000002800000000000000280000000000000036000000000000004300000000",
            INIT_37 => X"0000001c000000000000001b000000000000002b000000000000002f00000000",
            INIT_38 => X"0000002a000000000000000b0000000000000010000000000000001e00000000",
            INIT_39 => X"00000020000000000000001b000000000000001e000000000000002400000000",
            INIT_3A => X"0000000c000000000000001d0000000000000021000000000000002200000000",
            INIT_3B => X"0000001000000000000000160000000000000017000000000000002100000000",
            INIT_3C => X"00000009000000000000000c000000000000000e000000000000000c00000000",
            INIT_3D => X"00000010000000000000000b000000000000000c000000000000000b00000000",
            INIT_3E => X"0000002000000000000000160000000000000018000000000000001700000000",
            INIT_3F => X"0000000c000000000000000d000000000000000f000000000000001200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000300000000000000100000000000000000000000000000001200000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000000000000000000004000000000000000b000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000005000000000000000800000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_4B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000016000000000000001900000000",
            INIT_53 => X"0000000d00000000000000000000000000000019000000000000000e00000000",
            INIT_54 => X"000000000000000000000000000000000000000b000000000000000800000000",
            INIT_55 => X"0000002000000000000000310000000000000000000000000000000000000000",
            INIT_56 => X"0000000400000000000000000000000000000006000000000000000000000000",
            INIT_57 => X"0000000a00000000000000130000000000000000000000000000000000000000",
            INIT_58 => X"0000000e00000000000000020000000000000002000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000027000000000000000c00000000",
            INIT_5A => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000090000000000000019000000000000001900000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000a00000000000000000000000000000000000000000000001600000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000001c00000000000000000000000000000009000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000020000000000000023000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_6A => X"0000001b00000000000000030000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000400000000000000020000000000000001000000000000000100000000",
            INIT_76 => X"0000001700000000000000000000000000000000000000000000000200000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "samplegold_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000016b00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"000001a40000000000000198000000000000017d000000000000013900000000",
            INIT_32 => X"000001ab00000000000001bc00000000000001b400000000000001a400000000",
            INIT_33 => X"000001c100000000000001be00000000000001be00000000000001c100000000",
            INIT_34 => X"0000013e000000000000017500000000000001b700000000000001c600000000",
            INIT_35 => X"000001a100000000000001a4000000000000019c000000000000018200000000",
            INIT_36 => X"000001c200000000000001ac00000000000001ab00000000000001a800000000",
            INIT_37 => X"000001c500000000000001c400000000000001b4000000000000014f00000000",
            INIT_38 => X"0000017a0000000000000139000000000000017a00000000000001b500000000",
            INIT_39 => X"0000019d000000000000019300000000000001a4000000000000019700000000",
            INIT_3A => X"000001070000000000000198000000000000017a000000000000017900000000",
            INIT_3B => X"000001a700000000000001a900000000000001b3000000000000018d00000000",
            INIT_3C => X"00000171000000000000016b0000000000000122000000000000016600000000",
            INIT_3D => X"0000016a0000000000000185000000000000017e000000000000019000000000",
            INIT_3E => X"000000cd00000000000000c400000000000000d4000000000000013b00000000",
            INIT_3F => X"000000cd0000000000000168000000000000017300000000000000f300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000fa00000000000000e200000000000000d400000000000000c600000000",
            INIT_41 => X"000000d10000000000000118000000000000010a000000000000010500000000",
            INIT_42 => X"000000f400000000000000a600000000000000b200000000000000ca00000000",
            INIT_43 => X"000000a4000000000000008700000000000000e2000000000000012700000000",
            INIT_44 => X"000000d700000000000000d700000000000000a100000000000000d200000000",
            INIT_45 => X"000000c100000000000000c400000000000000e000000000000000ea00000000",
            INIT_46 => X"000000fb0000000000000146000000000000012700000000000000b500000000",
            INIT_47 => X"000000a800000000000000b300000000000000b700000000000000ef00000000",
            INIT_48 => X"000000fd00000000000000fe00000000000000e600000000000000ac00000000",
            INIT_49 => X"0000010f00000000000000fb00000000000000f400000000000000f100000000",
            INIT_4A => X"000000be00000000000001160000000000000144000000000000015600000000",
            INIT_4B => X"0000011500000000000000e700000000000000df00000000000000d600000000",
            INIT_4C => X"0000014400000000000001460000000000000142000000000000013100000000",
            INIT_4D => X"0000011700000000000000ec0000000000000132000000000000013100000000",
            INIT_4E => X"000000e900000000000000b000000000000000fe000000000000013100000000",
            INIT_4F => X"00000141000000000000012200000000000000df00000000000000ea00000000",
            INIT_50 => X"0000011200000000000001160000000000000127000000000000013600000000",
            INIT_51 => X"00000126000000000000012d000000000000010a000000000000011b00000000",
            INIT_52 => X"000000cc00000000000000ca0000000000000117000000000000011400000000",
            INIT_53 => X"000001170000000000000103000000000000011e000000000000011300000000",
            INIT_54 => X"000001210000000000000105000000000000012d000000000000012b00000000",
            INIT_55 => X"000000d6000000000000010a000000000000012d000000000000012c00000000",
            INIT_56 => X"00000108000000000000010500000000000000d900000000000000a200000000",
            INIT_57 => X"0000012200000000000000fa00000000000000f500000000000000ff00000000",
            INIT_58 => X"000000fc00000000000000fd000000000000009c00000000000000c000000000",
            INIT_59 => X"0000007b000000000000007e00000000000000a400000000000000d000000000",
            INIT_5A => X"000000a900000000000000fb00000000000000f100000000000000ba00000000",
            INIT_5B => X"000000ba00000000000000f500000000000000d500000000000000a400000000",
            INIT_5C => X"0000008500000000000000a100000000000000af00000000000000ae00000000",
            INIT_5D => X"000000a60000000000000040000000000000005b000000000000006f00000000",
            INIT_5E => X"0000009e00000000000000a000000000000000bc00000000000000ce00000000",
            INIT_5F => X"0000008c000000000000008b0000000000000083000000000000009100000000",
            INIT_60 => X"0000006000000000000000620000000000000066000000000000007c00000000",
            INIT_61 => X"0000004700000000000000540000000000000037000000000000003a00000000",
            INIT_62 => X"000000650000000000000063000000000000004e000000000000004b00000000",
            INIT_63 => X"00000088000000000000004f0000000000000062000000000000006200000000",
            INIT_64 => X"00000037000000000000003a0000000000000049000000000000004f00000000",
            INIT_65 => X"0000003a000000000000002f0000000000000032000000000000003c00000000",
            INIT_66 => X"0000005800000000000000510000000000000046000000000000004000000000",
            INIT_67 => X"0000003f000000000000006f000000000000004b000000000000005400000000",
            INIT_68 => X"0000004100000000000000360000000000000033000000000000003500000000",
            INIT_69 => X"00000037000000000000002a000000000000000c000000000000002a00000000",
            INIT_6A => X"0000005c00000000000000530000000000000046000000000000004300000000",
            INIT_6B => X"0000005c000000000000005c000000000000005d000000000000005000000000",
            INIT_6C => X"000000380000000000000056000000000000005e000000000000005900000000",
            INIT_6D => X"000000530000000000000049000000000000003a000000000000001c00000000",
            INIT_6E => X"00000055000000000000005f000000000000005e000000000000005200000000",
            INIT_6F => X"0000005f000000000000005d0000000000000044000000000000006800000000",
            INIT_70 => X"0000002500000000000000470000000000000058000000000000006700000000",
            INIT_71 => X"0000005700000000000000620000000000000055000000000000004500000000",
            INIT_72 => X"0000006300000000000000550000000000000059000000000000006500000000",
            INIT_73 => X"0000006a00000000000000640000000000000057000000000000003000000000",
            INIT_74 => X"0000005b000000000000002e0000000000000053000000000000005d00000000",
            INIT_75 => X"00000066000000000000005e000000000000006e000000000000006100000000",
            INIT_76 => X"0000000600000000000000340000000000000039000000000000005300000000",
            INIT_77 => X"00000060000000000000006c000000000000005a000000000000002b00000000",
            INIT_78 => X"00000042000000000000003b0000000000000027000000000000003900000000",
            INIT_79 => X"000000440000000000000044000000000000004f000000000000005300000000",
            INIT_7A => X"0000000f0000000000000002000000000000000d000000000000001900000000",
            INIT_7B => X"00000000000000000000003d000000000000004a000000000000001600000000",
            INIT_7C => X"0000000d00000000000000000000000000000013000000000000000100000000",
            INIT_7D => X"000000060000000000000012000000000000000a000000000000000c00000000",
            INIT_7E => X"0000003700000000000000230000000000000000000000000000000700000000",
            INIT_7F => X"0000000300000000000000000000000000000026000000000000005400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "samplegold_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000006000000000000000b0000000000000000000000000000000900000000",
            INIT_01 => X"0000000700000000000000000000000000000000000000000000000200000000",
            INIT_02 => X"0000004500000000000000620000000000000048000000000000001800000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_04 => X"000000190000000000000012000000000000000c000000000000000000000000",
            INIT_05 => X"0000002e00000000000000380000000000000027000000000000001d00000000",
            INIT_06 => X"0000001200000000000000250000000000000045000000000000004700000000",
            INIT_07 => X"000000160000000000000004000000000000000c000000000000001000000000",
            INIT_08 => X"0000001d000000000000001b000000000000001e000000000000001f00000000",
            INIT_09 => X"00000031000000000000001b000000000000002d000000000000002000000000",
            INIT_0A => X"000000000000000000000046000000000000003d000000000000003600000000",
            INIT_0B => X"0000000d00000000000000100000000000000003000000000000000000000000",
            INIT_0C => X"00000022000000000000002f000000000000001f000000000000001300000000",
            INIT_0D => X"0000003a00000000000000420000000000000030000000000000002e00000000",
            INIT_0E => X"0000000300000000000000000000000000000020000000000000003600000000",
            INIT_0F => X"000000150000000000000019000000000000001b000000000000001000000000",
            INIT_10 => X"0000003100000000000000000000000000000011000000000000002800000000",
            INIT_11 => X"0000000e000000000000001e000000000000002c000000000000003000000000",
            INIT_12 => X"0000001100000000000000080000000000000000000000000000001200000000",
            INIT_13 => X"00000031000000000000000d0000000000000000000000000000000000000000",
            INIT_14 => X"0000001700000000000000170000000000000003000000000000000e00000000",
            INIT_15 => X"0000000100000000000000000000000000000009000000000000000200000000",
            INIT_16 => X"00000005000000000000001b0000000000000013000000000000000100000000",
            INIT_17 => X"00000007000000000000000c000000000000000b000000000000000300000000",
            INIT_18 => X"0000000000000000000000050000000000000004000000000000000700000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000600000000000000000000000000000001000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000016000000000000000600000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_24 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_28 => X"0000001a00000000000000000000000000000000000000000000000700000000",
            INIT_29 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_2B => X"0000000d00000000000000000000000000000000000000000000006300000000",
            INIT_2C => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_2E => X"00000029000000000000001a0000000000000014000000000000001000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000090000000000000014000000000000001900000000",
            INIT_33 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_35 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_37 => X"0000000000000000000000340000000000000000000000000000003d00000000",
            INIT_38 => X"000000000000000000000000000000000000000e000000000000000400000000",
            INIT_39 => X"0000000000000000000000050000000000000000000000000000000500000000",
            INIT_3A => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000052000000000000000500000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000002600000000000000000000000000000008000000000000000000000000",
            INIT_3E => X"0000004b00000000000000040000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000200000000000000000000000000000000400000000",
            INIT_42 => X"00000000000000000000000f0000000000000001000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_44 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000002000000000000001e000000000000000e00000000",
            INIT_47 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000200000000000000022000000000000000000000000",
            INIT_49 => X"00000012000000000000001b0000000000000008000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000007000000000000000e00000000",
            INIT_4B => X"0000000000000000000000000000000000000009000000000000002000000000",
            INIT_4C => X"000000050000000000000000000000000000000c000000000000001e00000000",
            INIT_4D => X"000000070000000000000010000000000000000a000000000000000c00000000",
            INIT_4E => X"0000001200000000000000000000000000000000000000000000001200000000",
            INIT_4F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000e00000000000000050000000000000001000000000000000000000000",
            INIT_51 => X"0000000500000000000000040000000000000017000000000000000000000000",
            INIT_52 => X"0000000000000000000000010000000000000001000000000000000100000000",
            INIT_53 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000400000000000000050000000000000017000000000000000000000000",
            INIT_55 => X"0000000400000000000000050000000000000000000000000000000800000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000050000000000000000000000000000002f00000000",
            INIT_59 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000004300000000000000550000000000000018000000000000004f00000000",
            INIT_68 => X"0000001000000000000000270000000000000000000000000000000000000000",
            INIT_69 => X"0000001a0000000000000023000000000000001f000000000000002800000000",
            INIT_6A => X"0000000000000000000000000000000000000011000000000000001900000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000015000000000000000d0000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "samplegold_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001600000000000000000000000000000000000000000000001700000000",
            INIT_02 => X"0000000000000000000000000000000000000009000000000000000c00000000",
            INIT_03 => X"0000000500000000000000150000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000001100000000000000020000000000000005000000000000000f00000000",
            INIT_06 => X"0000000000000000000000000000000000000010000000000000000200000000",
            INIT_07 => X"0000002100000000000000030000000000000000000000000000000700000000",
            INIT_08 => X"0000000c00000000000000000000000000000000000000000000001900000000",
            INIT_09 => X"0000000700000000000000030000000000000000000000000000001100000000",
            INIT_0A => X"0000001500000000000000270000000000000019000000000000000000000000",
            INIT_0B => X"0000000b00000000000000000000000000000000000000000000000a00000000",
            INIT_0C => X"0000000600000000000000000000000000000006000000000000001100000000",
            INIT_0D => X"0000000000000000000000000000000000000008000000000000000400000000",
            INIT_0E => X"0000000400000000000000030000000000000002000000000000000200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_10 => X"0000000800000000000000000000000000000006000000000000000400000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_12 => X"0000000000000000000000000000000000000001000000000000000100000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000003000000000000001a00000000",
            INIT_19 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000003800000000000000000000000000000007000000000000000000000000",
            INIT_1C => X"0000000200000000000000000000000000000000000000000000000d00000000",
            INIT_1D => X"0000000700000000000000000000000000000004000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_20 => X"0000000300000000000000060000000000000000000000000000003e00000000",
            INIT_21 => X"00000007000000000000000f0000000000000001000000000000000500000000",
            INIT_22 => X"0000000000000000000000000000000000000009000000000000000b00000000",
            INIT_23 => X"00000004000000000000000a0000000000000000000000000000000000000000",
            INIT_24 => X"0000000200000000000000140000000000000006000000000000000000000000",
            INIT_25 => X"000000000000000000000004000000000000000e000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000001800000000000000000000000000000008000000000000001b00000000",
            INIT_28 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000000b000000000000001a00000000",
            INIT_2A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000100000000000000070000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000c00000000000000110000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000080000000000000018000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_33 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_38 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_3C => X"000000000000000000000000000000000000000f000000000000000100000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_44 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000002000000000000000200000000",
            INIT_48 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_49 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_4A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000010000000000000000d000000000000000a000000000000000600000000",
            INIT_4C => X"0000001200000000000000110000000000000011000000000000000d00000000",
            INIT_4D => X"0000000000000000000000110000000000000012000000000000001200000000",
            INIT_4E => X"0000000d000000000000000b0000000000000004000000000000000000000000",
            INIT_4F => X"0000000f000000000000000f0000000000000010000000000000000f00000000",
            INIT_50 => X"0000001400000000000000110000000000000000000000000000000b00000000",
            INIT_51 => X"0000000500000000000000080000000000000012000000000000001300000000",
            INIT_52 => X"0000001200000000000000150000000000000013000000000000000b00000000",
            INIT_53 => X"00000009000000000000000a000000000000000a000000000000001300000000",
            INIT_54 => X"0000001400000000000000120000000000000008000000000000000000000000",
            INIT_55 => X"00000015000000000000000d000000000000000d000000000000001500000000",
            INIT_56 => X"000000170000000000000019000000000000001c000000000000001700000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_58 => X"0000001300000000000000110000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000000000000000000001000000000000000c000000000000000c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001b00000000000000180000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000010000000000000001300000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001400000000000000180000000000000010000000000000000900000000",
            INIT_64 => X"0000000100000000000000000000000000000000000000000000000300000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"00000013000000000000000d000000000000000e000000000000000b00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000a000000000000000d000000000000000b000000000000000000000000",
            INIT_6B => X"00000000000000000000000b000000000000000e000000000000000700000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000080000000000000004000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "samplegold_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000001800000000000000130000000000000007000000000000000300000000",
            INIT_33 => X"0000000400000000000000030000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000f00000000000000090000000000000006000000000000000400000000",
            INIT_36 => X"0000001600000000000000170000000000000017000000000000001400000000",
            INIT_37 => X"0000000f00000000000000100000000000000013000000000000001600000000",
            INIT_38 => X"000000000000000000000009000000000000000b000000000000000f00000000",
            INIT_39 => X"0000001800000000000000170000000000000014000000000000000600000000",
            INIT_3A => X"0000000000000000000000000000000000000017000000000000001600000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "samplegold_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_05 => X"0000001300000000000000100000000000000000000000000000000000000000",
            INIT_06 => X"0000001c0000000000000029000000000000000a000000000000000300000000",
            INIT_07 => X"0000000a00000000000000000000000000000000000000000000000200000000",
            INIT_08 => X"0000000000000000000000260000000000000046000000000000002c00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0A => X"0000002400000000000000150000000000000000000000000000000000000000",
            INIT_0B => X"000000140000000000000038000000000000004b000000000000003a00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"00000040000000000000004b0000000000000038000000000000002400000000",
            INIT_0E => X"00000000000000000000000c0000000000000014000000000000002100000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000006b0000000000000021000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000026000000000000002200000000",
            INIT_14 => X"0000002e000000000000001c0000000000000000000000000000000000000000",
            INIT_15 => X"0000001200000000000000000000000000000000000000000000000600000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000003000000000000000a0000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000060000000000000007000000000000000200000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000000000000000000000000000000000c000000000000000400000000",
            INIT_3A => X"0000000700000000000000010000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000b00000000000000070000000000000004000000000000001200000000",
            INIT_3E => X"00000007000000000000000c0000000000000000000000000000000400000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000b000000000000000b000000000000000000000000",
            INIT_41 => X"0000000000000000000000020000000000000000000000000000001800000000",
            INIT_42 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000004000000000000000a00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000d00000000000000000000000000000000000000000000000700000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_53 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000a000000000000000500000000",
            INIT_55 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000010000000000000005000000000000000000000000",
            INIT_57 => X"0000000700000000000000070000000000000002000000000000000700000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_59 => X"0000000200000000000000000000000000000003000000000000000000000000",
            INIT_5A => X"0000000a00000000000000030000000000000006000000000000000300000000",
            INIT_5B => X"00000006000000000000000c000000000000000a000000000000000200000000",
            INIT_5C => X"0000000900000000000000090000000000000008000000000000000600000000",
            INIT_5D => X"0000000f0000000000000008000000000000000a000000000000000a00000000",
            INIT_5E => X"0000000900000000000000080000000000000009000000000000000200000000",
            INIT_5F => X"00000011000000000000000d000000000000000a000000000000000d00000000",
            INIT_60 => X"0000000c000000000000000e0000000000000010000000000000001100000000",
            INIT_61 => X"0000000000000000000000180000000000000008000000000000000c00000000",
            INIT_62 => X"0000000e000000000000000c0000000000000009000000000000000b00000000",
            INIT_63 => X"000000400000000000000037000000000000004d000000000000000700000000",
            INIT_64 => X"0000002e0000000000000032000000000000003b000000000000004000000000",
            INIT_65 => X"0000002c000000000000002c000000000000002a000000000000003000000000",
            INIT_66 => X"00000021000000000000002b0000000000000027000000000000002400000000",
            INIT_67 => X"000000320000000000000032000000000000002b000000000000004300000000",
            INIT_68 => X"0000002b000000000000002b0000000000000029000000000000002e00000000",
            INIT_69 => X"0000002000000000000000190000000000000049000000000000002600000000",
            INIT_6A => X"00000038000000000000001f0000000000000029000000000000002500000000",
            INIT_6B => X"0000002200000000000000200000000000000024000000000000002300000000",
            INIT_6C => X"00000023000000000000002e000000000000002b000000000000002000000000",
            INIT_6D => X"00000028000000000000002e000000000000001c000000000000004c00000000",
            INIT_6E => X"000000140000000000000032000000000000001e000000000000002100000000",
            INIT_6F => X"0000001500000000000000180000000000000016000000000000002200000000",
            INIT_70 => X"00000037000000000000004f0000000000000028000000000000001e00000000",
            INIT_71 => X"0000002900000000000000200000000000000036000000000000003800000000",
            INIT_72 => X"0000003000000000000000300000000000000036000000000000001800000000",
            INIT_73 => X"0000002d000000000000002c000000000000002a000000000000002f00000000",
            INIT_74 => X"0000003500000000000000390000000000000030000000000000004000000000",
            INIT_75 => X"0000001d000000000000001d0000000000000017000000000000000300000000",
            INIT_76 => X"00000016000000000000002f0000000000000017000000000000001e00000000",
            INIT_77 => X"0000004100000000000000390000000000000021000000000000001d00000000",
            INIT_78 => X"0000000600000000000000060000000000000028000000000000003300000000",
            INIT_79 => X"00000038000000000000001e0000000000000007000000000000001a00000000",
            INIT_7A => X"00000030000000000000002c000000000000002f000000000000002d00000000",
            INIT_7B => X"00000024000000000000002c0000000000000035000000000000003300000000",
            INIT_7C => X"00000013000000000000001d0000000000000015000000000000002300000000",
            INIT_7D => X"000000240000000000000033000000000000001e000000000000001e00000000",
            INIT_7E => X"00000041000000000000003d0000000000000033000000000000002000000000",
            INIT_7F => X"0000004a00000000000000440000000000000049000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "samplegold_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001100000000000000140000000000000010000000000000002300000000",
            INIT_01 => X"0000003a0000000000000055000000000000004d000000000000000000000000",
            INIT_02 => X"0000004e00000000000000580000000000000056000000000000004700000000",
            INIT_03 => X"00000010000000000000001f0000000000000026000000000000003600000000",
            INIT_04 => X"00000024000000000000001a0000000000000021000000000000001c00000000",
            INIT_05 => X"00000050000000000000004a000000000000002c000000000000003700000000",
            INIT_06 => X"0000004600000000000000390000000000000035000000000000003c00000000",
            INIT_07 => X"0000002f0000000000000028000000000000002d000000000000003900000000",
            INIT_08 => X"0000004700000000000000210000000000000033000000000000003a00000000",
            INIT_09 => X"00000051000000000000004f000000000000004a000000000000004b00000000",
            INIT_0A => X"000000170000000000000034000000000000004d000000000000004100000000",
            INIT_0B => X"0000002c00000000000000370000000000000043000000000000003a00000000",
            INIT_0C => X"00000045000000000000003e0000000000000028000000000000002300000000",
            INIT_0D => X"00000033000000000000002b0000000000000036000000000000005200000000",
            INIT_0E => X"0000002a000000000000002e0000000000000035000000000000004700000000",
            INIT_0F => X"00000022000000000000001f000000000000002e000000000000003100000000",
            INIT_10 => X"0000004b000000000000004e000000000000003d000000000000001600000000",
            INIT_11 => X"000000250000000000000034000000000000003f000000000000004200000000",
            INIT_12 => X"0000001d000000000000002d0000000000000035000000000000002900000000",
            INIT_13 => X"0000001600000000000000180000000000000025000000000000002100000000",
            INIT_14 => X"0000002100000000000000240000000000000026000000000000002c00000000",
            INIT_15 => X"0000002100000000000000260000000000000028000000000000002700000000",
            INIT_16 => X"0000001b000000000000001e000000000000002a000000000000000d00000000",
            INIT_17 => X"0000001200000000000000140000000000000015000000000000001800000000",
            INIT_18 => X"0000001400000000000000130000000000000013000000000000000f00000000",
            INIT_19 => X"0000001400000000000000200000000000000020000000000000001800000000",
            INIT_1A => X"000000160000000000000015000000000000001a000000000000002500000000",
            INIT_1B => X"000000000000000000000000000000000000001d000000000000001500000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000100000000000000030000000000000004000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_55 => X"0000000200000000000000000000000000000003000000000000000700000000",
            INIT_56 => X"00000010000000000000000a0000000000000011000000000000000500000000",
            INIT_57 => X"0000001100000000000000000000000000000012000000000000000000000000",
            INIT_58 => X"0000000c00000000000000000000000000000009000000000000000000000000",
            INIT_59 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000130000000000000009000000000000001d00000000",
            INIT_5B => X"0000000900000000000000200000000000000000000000000000001200000000",
            INIT_5C => X"00000000000000000000000d0000000000000003000000000000001200000000",
            INIT_5D => X"0000001000000000000000000000000000000012000000000000000500000000",
            INIT_5E => X"0000000f0000000000000006000000000000000c000000000000000900000000",
            INIT_5F => X"00000013000000000000000a0000000000000026000000000000000100000000",
            INIT_60 => X"00000000000000000000000c0000000000000012000000000000001000000000",
            INIT_61 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000210000000000000003000000000000000d00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"00000009000000000000001a0000000000000000000000000000000000000000",
            INIT_66 => X"0000001000000000000000000000000000000009000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000006000000000000001400000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000170000000000000015000000000000000e000000000000000800000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"000000000000000000000006000000000000000f000000000000000c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000300000000000000010000000000000003000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "samplegold_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000004900000000000000550000000000000055000000000000003f00000000",
            INIT_0D => X"00000045000000000000004b000000000000004f000000000000004900000000",
            INIT_0E => X"00000049000000000000004a0000000000000048000000000000004900000000",
            INIT_0F => X"000000490000000000000055000000000000004d000000000000004300000000",
            INIT_10 => X"0000004b000000000000005d000000000000005c000000000000005f00000000",
            INIT_11 => X"0000005c0000000000000059000000000000005b000000000000005b00000000",
            INIT_12 => X"000000590000000000000055000000000000005e000000000000005900000000",
            INIT_13 => X"0000005e000000000000004b000000000000005d000000000000005c00000000",
            INIT_14 => X"000000290000000000000035000000000000004d000000000000005d00000000",
            INIT_15 => X"00000030000000000000002e0000000000000025000000000000003100000000",
            INIT_16 => X"0000005e000000000000005c000000000000003c000000000000002e00000000",
            INIT_17 => X"0000005f000000000000005b000000000000004c000000000000006000000000",
            INIT_18 => X"000000390000000000000040000000000000003c000000000000003d00000000",
            INIT_19 => X"00000041000000000000004a000000000000004a000000000000004200000000",
            INIT_1A => X"0000005f000000000000005e0000000000000041000000000000004300000000",
            INIT_1B => X"000000580000000000000055000000000000005b000000000000005300000000",
            INIT_1C => X"0000004c000000000000004d0000000000000050000000000000004f00000000",
            INIT_1D => X"00000042000000000000004a000000000000004e000000000000005300000000",
            INIT_1E => X"000000500000000000000061000000000000005c000000000000005a00000000",
            INIT_1F => X"0000004c00000000000000530000000000000064000000000000005d00000000",
            INIT_20 => X"000000520000000000000051000000000000004e000000000000004d00000000",
            INIT_21 => X"0000005e000000000000005c000000000000004c000000000000004e00000000",
            INIT_22 => X"0000005a000000000000004f000000000000005d000000000000005b00000000",
            INIT_23 => X"00000065000000000000005d0000000000000048000000000000004900000000",
            INIT_24 => X"00000060000000000000005f0000000000000061000000000000006000000000",
            INIT_25 => X"0000006200000000000000600000000000000060000000000000005f00000000",
            INIT_26 => X"0000004200000000000000600000000000000050000000000000006200000000",
            INIT_27 => X"0000006000000000000000470000000000000033000000000000003700000000",
            INIT_28 => X"0000005b000000000000005e0000000000000061000000000000006400000000",
            INIT_29 => X"0000005f000000000000005d000000000000005d000000000000005d00000000",
            INIT_2A => X"0000004f000000000000005f000000000000005e000000000000005100000000",
            INIT_2B => X"0000004c0000000000000039000000000000001e000000000000004b00000000",
            INIT_2C => X"0000005e000000000000005f0000000000000068000000000000006100000000",
            INIT_2D => X"0000004f0000000000000061000000000000005f000000000000005f00000000",
            INIT_2E => X"000000540000000000000066000000000000005d000000000000005c00000000",
            INIT_2F => X"0000002600000000000000170000000000000011000000000000001000000000",
            INIT_30 => X"00000063000000000000005e0000000000000049000000000000003a00000000",
            INIT_31 => X"0000005e000000000000004d0000000000000061000000000000006300000000",
            INIT_32 => X"0000001a00000000000000110000000000000055000000000000005e00000000",
            INIT_33 => X"0000000600000000000000170000000000000000000000000000000000000000",
            INIT_34 => X"0000004000000000000000070000000000000005000000000000000600000000",
            INIT_35 => X"0000006f00000000000000710000000000000059000000000000005300000000",
            INIT_36 => X"00000053000000000000005b0000000000000070000000000000006e00000000",
            INIT_37 => X"0000005b000000000000005d0000000000000065000000000000006300000000",
            INIT_38 => X"0000006500000000000000650000000000000063000000000000005700000000",
            INIT_39 => X"0000002d00000000000000300000000000000033000000000000002a00000000",
            INIT_3A => X"0000003c000000000000002f000000000000002b000000000000002c00000000",
            INIT_3B => X"0000004c000000000000004a0000000000000046000000000000004700000000",
            INIT_3C => X"0000002300000000000000540000000000000054000000000000005000000000",
            INIT_3D => X"00000017000000000000001d0000000000000026000000000000002800000000",
            INIT_3E => X"0000001000000000000000160000000000000016000000000000001500000000",
            INIT_3F => X"0000000b000000000000000b000000000000000b000000000000000f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d000000000000000f0000000000000000000000000000000700000000",
            INIT_41 => X"0000000400000000000000080000000000000009000000000000000a00000000",
            INIT_42 => X"0000000200000000000000040000000000000003000000000000000700000000",
            INIT_43 => X"0000000000000000000000000000000000000006000000000000000400000000",
            INIT_44 => X"000000000000000000000000000000000000000a000000000000003000000000",
            INIT_45 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000800000000000000110000000000000000000000000000000c00000000",
            INIT_4E => X"0000000800000000000000020000000000000002000000000000000300000000",
            INIT_4F => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_52 => X"00000000000000000000001a0000000000000000000000000000000200000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000100000000000000020000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000f000000000000005e0000000000000022000000000000000000000000",
            INIT_6C => X"000000510000000000000017000000000000001f000000000000000d00000000",
            INIT_6D => X"0000000000000000000000000000000000000003000000000000001200000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000210000000000000002000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000090000000000000002000000000000000600000000",
            INIT_7B => X"0000000e00000000000000000000000000000000000000000000000400000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "samplegold_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000012c00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000014100000000000001440000000000000161000000000000016300000000",
            INIT_36 => X"00000156000000000000014c0000000000000159000000000000015800000000",
            INIT_37 => X"000001580000000000000159000000000000015b000000000000015500000000",
            INIT_38 => X"00000162000000000000012f0000000000000182000000000000017b00000000",
            INIT_39 => X"00000146000000000000012e000000000000015c000000000000016f00000000",
            INIT_3A => X"0000015400000000000001540000000000000140000000000000014a00000000",
            INIT_3B => X"0000018300000000000001740000000000000146000000000000015200000000",
            INIT_3C => X"00000174000000000000015b000000000000012a000000000000018900000000",
            INIT_3D => X"0000012a00000000000001200000000000000138000000000000014200000000",
            INIT_3E => X"0000013d00000000000001460000000000000139000000000000012200000000",
            INIT_3F => X"0000018900000000000001840000000000000168000000000000014800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000011d00000000000001680000000000000155000000000000013300000000",
            INIT_41 => X"0000012700000000000001290000000000000127000000000000012500000000",
            INIT_42 => X"0000013b00000000000001260000000000000137000000000000013200000000",
            INIT_43 => X"0000014c00000000000001800000000000000179000000000000013400000000",
            INIT_44 => X"0000013500000000000001650000000000000160000000000000015600000000",
            INIT_45 => X"00000146000000000000013f0000000000000133000000000000013600000000",
            INIT_46 => X"000001760000000000000141000000000000013a000000000000013e00000000",
            INIT_47 => X"0000016b000000000000015f000000000000017d000000000000017d00000000",
            INIT_48 => X"0000015f0000000000000166000000000000014d000000000000015700000000",
            INIT_49 => X"00000168000000000000016b0000000000000170000000000000016600000000",
            INIT_4A => X"0000017b00000000000001780000000000000173000000000000016700000000",
            INIT_4B => X"0000013100000000000001680000000000000167000000000000017d00000000",
            INIT_4C => X"0000017a000000000000015b000000000000010300000000000000f500000000",
            INIT_4D => X"0000017a00000000000001830000000000000184000000000000018500000000",
            INIT_4E => X"0000017d000000000000017e000000000000017c000000000000017d00000000",
            INIT_4F => X"0000015000000000000001770000000000000188000000000000016c00000000",
            INIT_50 => X"0000017d000000000000013000000000000000d000000000000000ec00000000",
            INIT_51 => X"000001790000000000000177000000000000017d000000000000018800000000",
            INIT_52 => X"0000017200000000000001780000000000000179000000000000017a00000000",
            INIT_53 => X"00000139000000000000018a0000000000000197000000000000019100000000",
            INIT_54 => X"0000011500000000000000db00000000000000af000000000000008900000000",
            INIT_55 => X"0000017f00000000000001820000000000000162000000000000015000000000",
            INIT_56 => X"0000019000000000000001720000000000000179000000000000017a00000000",
            INIT_57 => X"00000060000000000000011d000000000000019a000000000000019400000000",
            INIT_58 => X"000000a600000000000000a00000000000000086000000000000006900000000",
            INIT_59 => X"00000153000000000000011a00000000000000e5000000000000009d00000000",
            INIT_5A => X"0000018e000000000000018b0000000000000168000000000000017400000000",
            INIT_5B => X"0000009600000000000001030000000000000110000000000000018500000000",
            INIT_5C => X"000000cc00000000000000df000000000000011e000000000000009f00000000",
            INIT_5D => X"00000160000000000000014a00000000000000d300000000000000c900000000",
            INIT_5E => X"00000131000000000000013c0000000000000145000000000000012a00000000",
            INIT_5F => X"0000011b00000000000001010000000000000112000000000000012a00000000",
            INIT_60 => X"000001210000000000000128000000000000011b000000000000013100000000",
            INIT_61 => X"000000c900000000000001310000000000000130000000000000013800000000",
            INIT_62 => X"000000b900000000000000c000000000000000ca00000000000000cc00000000",
            INIT_63 => X"000000c000000000000000b900000000000000ad00000000000000af00000000",
            INIT_64 => X"000000b300000000000000ae00000000000000b200000000000000b100000000",
            INIT_65 => X"0000007f000000000000008900000000000000a900000000000000b700000000",
            INIT_66 => X"0000006700000000000000750000000000000071000000000000007a00000000",
            INIT_67 => X"0000006100000000000000690000000000000066000000000000006400000000",
            INIT_68 => X"00000057000000000000005d000000000000005e000000000000005800000000",
            INIT_69 => X"000000600000000000000063000000000000006f000000000000005e00000000",
            INIT_6A => X"0000006d000000000000005d000000000000005f000000000000006100000000",
            INIT_6B => X"00000069000000000000006b0000000000000073000000000000006900000000",
            INIT_6C => X"000000c600000000000000890000000000000054000000000000005f00000000",
            INIT_6D => X"00000039000000000000002f0000000000000031000000000000002700000000",
            INIT_6E => X"00000038000000000000003c0000000000000039000000000000003300000000",
            INIT_6F => X"0000003c000000000000003c0000000000000037000000000000003600000000",
            INIT_70 => X"0000002000000000000000460000000000000045000000000000003a00000000",
            INIT_71 => X"0000005b000000000000004f000000000000003a000000000000002b00000000",
            INIT_72 => X"00000064000000000000005d0000000000000061000000000000005f00000000",
            INIT_73 => X"00000044000000000000004f0000000000000061000000000000006300000000",
            INIT_74 => X"0000002600000000000000220000000000000046000000000000004800000000",
            INIT_75 => X"0000005a00000000000000600000000000000063000000000000003d00000000",
            INIT_76 => X"0000005f00000000000000590000000000000059000000000000005d00000000",
            INIT_77 => X"00000044000000000000004a000000000000004e000000000000005800000000",
            INIT_78 => X"0000004800000000000000250000000000000021000000000000004300000000",
            INIT_79 => X"0000004b00000000000000440000000000000049000000000000004c00000000",
            INIT_7A => X"0000005200000000000000550000000000000046000000000000004700000000",
            INIT_7B => X"0000003d0000000000000040000000000000003b000000000000005300000000",
            INIT_7C => X"0000003e00000000000000340000000000000026000000000000002a00000000",
            INIT_7D => X"0000003600000000000000310000000000000033000000000000003400000000",
            INIT_7E => X"000000380000000000000037000000000000003a000000000000003c00000000",
            INIT_7F => X"00000038000000000000003a000000000000003d000000000000003b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "samplegold_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d00000000000000330000000000000037000000000000003a00000000",
            INIT_01 => X"000000330000000000000034000000000000002e000000000000002c00000000",
            INIT_02 => X"0000003d000000000000002e0000000000000031000000000000003100000000",
            INIT_03 => X"0000002a000000000000003a0000000000000039000000000000003c00000000",
            INIT_04 => X"000000340000000000000044000000000000003e000000000000002800000000",
            INIT_05 => X"00000040000000000000003f000000000000003e000000000000003a00000000",
            INIT_06 => X"00000040000000000000003d000000000000003f000000000000003e00000000",
            INIT_07 => X"0000004d000000000000003e000000000000003c000000000000003f00000000",
            INIT_08 => X"0000004300000000000000350000000000000017000000000000002f00000000",
            INIT_09 => X"0000003f00000000000000440000000000000045000000000000004200000000",
            INIT_0A => X"00000037000000000000003a000000000000003c000000000000003e00000000",
            INIT_0B => X"00000053000000000000004a0000000000000048000000000000004300000000",
            INIT_0C => X"0000004d000000000000001b0000000000000017000000000000004600000000",
            INIT_0D => X"0000003e00000000000000380000000000000048000000000000005600000000",
            INIT_0E => X"000000480000000000000038000000000000003d000000000000003f00000000",
            INIT_0F => X"00000052000000000000005f000000000000004b000000000000004b00000000",
            INIT_10 => X"00000015000000000000001b0000000000000019000000000000001700000000",
            INIT_11 => X"0000004f000000000000005b0000000000000033000000000000002400000000",
            INIT_12 => X"000000480000000000000041000000000000003a000000000000004100000000",
            INIT_13 => X"000000000000000000000029000000000000004c000000000000004a00000000",
            INIT_14 => X"0000000300000000000000170000000000000004000000000000000000000000",
            INIT_15 => X"0000001f000000000000000c0000000000000000000000000000000000000000",
            INIT_16 => X"0000005a0000000000000059000000000000004d000000000000003b00000000",
            INIT_17 => X"0000003c000000000000005e0000000000000057000000000000005a00000000",
            INIT_18 => X"00000034000000000000003d0000000000000045000000000000002e00000000",
            INIT_19 => X"0000003b00000000000000350000000000000028000000000000003800000000",
            INIT_1A => X"0000001f000000000000001f000000000000001f000000000000001b00000000",
            INIT_1B => X"000000170000000000000016000000000000001c000000000000002000000000",
            INIT_1C => X"0000002400000000000000230000000000000024000000000000002500000000",
            INIT_1D => X"0000001b0000000000000027000000000000002a000000000000002700000000",
            INIT_1E => X"0000001e000000000000001b0000000000000021000000000000001e00000000",
            INIT_1F => X"0000001a00000000000000150000000000000015000000000000001500000000",
            INIT_20 => X"0000001000000000000000120000000000000011000000000000001200000000",
            INIT_21 => X"0000001000000000000000160000000000000000000000000000000a00000000",
            INIT_22 => X"0000000700000000000000110000000000000010000000000000001200000000",
            INIT_23 => X"0000000d000000000000000e000000000000000d000000000000000f00000000",
            INIT_24 => X"0000000b00000000000000000000000000000013000000000000001100000000",
            INIT_25 => X"0000001a00000000000000000000000000000000000000000000001200000000",
            INIT_26 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000002c00000000000000080000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000160000000000000003000000000000000000000000",
            INIT_2B => X"0000000000000000000000040000000000000009000000000000000c00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000d000000000000000d0000000000000005000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000007000000000000001c00000000",
            INIT_32 => X"0000001400000000000000030000000000000000000000000000000400000000",
            INIT_33 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_36 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000030000000000000002200000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000012000000000000004b000000000000001600000000",
            INIT_41 => X"0000000200000000000000010000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000095000000000000001000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000009c00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002a000000000000002c0000000000000000000000000000000000000000",
            INIT_4C => X"0000000d00000000000000000000000000000000000000000000004d00000000",
            INIT_4D => X"0000000000000000000000100000000000000000000000000000002b00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000200000000000000010000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000900000000000000020000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000070000000000000003000000000000000500000000",
            INIT_54 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_55 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000060000000000000000000000000000001000000000",
            INIT_57 => X"0000000000000000000000000000000000000002000000000000000700000000",
            INIT_58 => X"0000000000000000000000000000000000000006000000000000000400000000",
            INIT_59 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000300000000000000000000000000000002000000000000000300000000",
            INIT_5B => X"0000000700000000000000000000000000000004000000000000000000000000",
            INIT_5C => X"0000000000000000000000050000000000000005000000000000000500000000",
            INIT_5D => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000000f0000000000000042000000000000000c00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "samplegold_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000000000140000000000000000000000000000000000000000",
            INIT_01 => X"0000005900000000000000300000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000003b00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000700000000000000040000000000000000000000000000000000000000",
            INIT_08 => X"0000000900000000000000000000000000000000000000000000001000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000008000000000000000800000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000100000000000000040000000000000003000000000000000000000000",
            INIT_0E => X"0000002200000000000000200000000000000015000000000000000f00000000",
            INIT_0F => X"0000001200000000000000140000000000000015000000000000001a00000000",
            INIT_10 => X"000000060000000000000002000000000000000c000000000000000d00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_1C => X"00000000000000000000000e0000000000000005000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_1E => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_1F => X"0000000500000000000000000000000000000005000000000000001500000000",
            INIT_20 => X"0000000000000000000000000000000000000012000000000000000300000000",
            INIT_21 => X"0000000000000000000000000000000000000001000000000000001000000000",
            INIT_22 => X"0000000800000000000000000000000000000003000000000000000a00000000",
            INIT_23 => X"00000004000000000000000e0000000000000000000000000000000600000000",
            INIT_24 => X"0000000300000000000000000000000000000000000000000000001c00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_2D => X"00000000000000000000000f000000000000002b000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_31 => X"00000000000000000000002a000000000000002b000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000001b00000000000000190000000000000010000000000000000700000000",
            INIT_36 => X"000000000000000000000000000000000000000b000000000000000a00000000",
            INIT_37 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000009000000000000001100000000",
            INIT_3A => X"0000000f000000000000001f0000000000000017000000000000001e00000000",
            INIT_3B => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_3E => X"0000000000000000000000000000000000000030000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000001300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001400000000000000020000000000000000000000000000000000000000",
            INIT_41 => X"0000000200000000000000010000000000000000000000000000000000000000",
            INIT_42 => X"0000000300000000000000030000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_4B => X"0000000000000000000000080000000000000000000000000000000100000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_4D => X"00000000000000000000000b0000000000000015000000000000000000000000",
            INIT_4E => X"0000000800000000000000030000000000000000000000000000000100000000",
            INIT_4F => X"0000000700000000000000070000000000000004000000000000000500000000",
            INIT_50 => X"0000000800000000000000080000000000000007000000000000000800000000",
            INIT_51 => X"00000000000000000000000a000000000000000d000000000000000900000000",
            INIT_52 => X"0000002e000000000000001a0000000000000003000000000000000000000000",
            INIT_53 => X"0000002a00000000000000270000000000000029000000000000002c00000000",
            INIT_54 => X"0000001100000000000000180000000000000024000000000000002a00000000",
            INIT_55 => X"000000000000000000000000000000000000000b000000000000000b00000000",
            INIT_56 => X"000000250000000000000022000000000000001f000000000000000600000000",
            INIT_57 => X"00000021000000000000001e0000000000000024000000000000002700000000",
            INIT_58 => X"0000000900000000000000100000000000000021000000000000002500000000",
            INIT_59 => X"0000000500000000000000000000000000000002000000000000000800000000",
            INIT_5A => X"00000019000000000000001a000000000000001d000000000000002600000000",
            INIT_5B => X"0000001d000000000000001e000000000000001e000000000000001f00000000",
            INIT_5C => X"0000000300000000000000080000000000000016000000000000001f00000000",
            INIT_5D => X"0000000300000000000000000000000000000000000000000000000600000000",
            INIT_5E => X"0000000200000000000000000000000000000000000000000000000100000000",
            INIT_5F => X"0000000000000000000000030000000000000001000000000000000300000000",
            INIT_60 => X"0000000900000000000000040000000000000004000000000000000a00000000",
            INIT_61 => X"0000000800000000000000000000000000000000000000000000000500000000",
            INIT_62 => X"0000000b000000000000000a0000000000000009000000000000000700000000",
            INIT_63 => X"0000000300000000000000050000000000000009000000000000000900000000",
            INIT_64 => X"0000000400000000000000080000000000000006000000000000000400000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_66 => X"0000000900000000000000090000000000000007000000000000000600000000",
            INIT_67 => X"0000000400000000000000040000000000000007000000000000000700000000",
            INIT_68 => X"0000001100000000000000070000000000000009000000000000000300000000",
            INIT_69 => X"000000000000000000000000000000000000000c000000000000001c00000000",
            INIT_6A => X"0000000700000000000000070000000000000008000000000000000700000000",
            INIT_6B => X"0000000200000000000000040000000000000006000000000000000700000000",
            INIT_6C => X"00000010000000000000000b000000000000000b000000000000000d00000000",
            INIT_6D => X"0000000000000000000000000000000000000006000000000000001900000000",
            INIT_6E => X"0000000800000000000000030000000000000005000000000000000000000000",
            INIT_6F => X"0000000e00000000000000030000000000000005000000000000000700000000",
            INIT_70 => X"0000000d0000000000000010000000000000000a000000000000000c00000000",
            INIT_71 => X"00000003000000000000000c0000000000000006000000000000000400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"00000009000000000000000a0000000000000005000000000000000300000000",
            INIT_74 => X"0000001d000000000000001d000000000000000c000000000000000b00000000",
            INIT_75 => X"00000016000000000000001e0000000000000013000000000000000900000000",
            INIT_76 => X"0000000b000000000000000d000000000000000f000000000000001600000000",
            INIT_77 => X"0000000000000000000000000000000000000001000000000000000700000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000a00000000000000090000000000000007000000000000000900000000",
            INIT_7C => X"000000030000000000000008000000000000000a000000000000000c00000000",
            INIT_7D => X"0000000000000000000000000000000000000002000000000000000200000000",
            INIT_7E => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000400000000000000030000000000000002000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "samplegold_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000000000050000000000000003000000000000000200000000",
            INIT_01 => X"0000000600000000000000080000000000000006000000000000000600000000",
            INIT_02 => X"00000007000000000000000e0000000000000001000000000000000200000000",
            INIT_03 => X"0000000900000000000000080000000000000007000000000000000700000000",
            INIT_04 => X"0000000d000000000000000d000000000000000c000000000000000d00000000",
            INIT_05 => X"000000070000000000000002000000000000000a000000000000000d00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_78 => X"0000000700000000000000020000000000000001000000000000000000000000",
            INIT_79 => X"0000000700000000000000000000000000000001000000000000000300000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000700000000000000190000000000000007000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "samplegold_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000018000000000000001b000000000000001d000000000000001100000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_02 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"00000004000000000000000d0000000000000006000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000400000000000000000000000000000000000000000000000200000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000001e00000000000000230000000000000000000000000000000000000000",
            INIT_0B => X"00000018000000000000001c0000000000000019000000000000001c00000000",
            INIT_0C => X"0000000000000000000000000000000000000002000000000000001500000000",
            INIT_0D => X"0000001800000000000000170000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000006d00000000000000200000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000002000000000000000010000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000006e00000000000000a70000000000000088000000000000000900000000",
            INIT_1E => X"0000008f00000000000000840000000000000089000000000000007700000000",
            INIT_1F => X"0000000000000000000000200000000000000051000000000000007a00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_2C => X"00000013000000000000000d0000000000000000000000000000000000000000",
            INIT_2D => X"0000000700000000000000150000000000000012000000000000001000000000",
            INIT_2E => X"00000000000000000000002c0000000000000013000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000020000000000000013000000000000000f000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"00000011000000000000000d000000000000000f000000000000001000000000",
            INIT_53 => X"0000000000000000000000000000000000000006000000000000000800000000",
            INIT_54 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"000000000000000000000004000000000000001b000000000000001500000000",
            INIT_57 => X"000000000000000000000019000000000000000e000000000000000e00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000e000000000000000e0000000000000007000000000000000700000000",
            INIT_61 => X"00000010000000000000000f000000000000000c000000000000000d00000000",
            INIT_62 => X"0000001400000000000000140000000000000013000000000000001100000000",
            INIT_63 => X"00000012000000000000000a0000000000000020000000000000001900000000",
            INIT_64 => X"0000001400000000000000120000000000000013000000000000001100000000",
            INIT_65 => X"0000001400000000000000150000000000000017000000000000001100000000",
            INIT_66 => X"0000001700000000000000220000000000000016000000000000001300000000",
            INIT_67 => X"0000003300000000000000360000000000000029000000000000001500000000",
            INIT_68 => X"0000002400000000000000250000000000000027000000000000002100000000",
            INIT_69 => X"000000220000000000000020000000000000001f000000000000001f00000000",
            INIT_6A => X"0000002800000000000000230000000000000019000000000000002100000000",
            INIT_6B => X"00000014000000000000003b0000000000000043000000000000003100000000",
            INIT_6C => X"0000000900000000000000120000000000000013000000000000000000000000",
            INIT_6D => X"0000000e00000000000000160000000000000016000000000000001300000000",
            INIT_6E => X"000000310000000000000029000000000000002e000000000000002e00000000",
            INIT_6F => X"00000011000000000000000b0000000000000043000000000000004100000000",
            INIT_70 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"00000028000000000000000e000000000000000b000000000000000d00000000",
            INIT_72 => X"0000003e0000000000000032000000000000002d000000000000003100000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_75 => X"0000002f00000000000000000000000000000005000000000000000000000000",
            INIT_76 => X"0000003a000000000000003e0000000000000034000000000000003500000000",
            INIT_77 => X"0000002c00000000000000330000000000000030000000000000004100000000",
            INIT_78 => X"0000002900000000000000310000000000000032000000000000002e00000000",
            INIT_79 => X"000000360000000000000037000000000000002d000000000000002800000000",
            INIT_7A => X"0000003100000000000000490000000000000042000000000000003000000000",
            INIT_7B => X"0000002d000000000000002b000000000000002b000000000000002f00000000",
            INIT_7C => X"00000034000000000000002b000000000000002d000000000000002b00000000",
            INIT_7D => X"0000002b00000000000000300000000000000033000000000000003800000000",
            INIT_7E => X"0000003900000000000000350000000000000025000000000000003200000000",
            INIT_7F => X"0000003200000000000000350000000000000033000000000000003a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "samplegold_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003800000000000000370000000000000034000000000000003500000000",
            INIT_01 => X"00000035000000000000002b0000000000000037000000000000003800000000",
            INIT_02 => X"0000002f0000000000000023000000000000000f000000000000002000000000",
            INIT_03 => X"0000003300000000000000340000000000000032000000000000003600000000",
            INIT_04 => X"0000003500000000000000340000000000000032000000000000003000000000",
            INIT_05 => X"0000002f000000000000002f000000000000002a000000000000003600000000",
            INIT_06 => X"00000021000000000000000d000000000000002b000000000000002600000000",
            INIT_07 => X"00000031000000000000003c000000000000003a000000000000003300000000",
            INIT_08 => X"0000003600000000000000360000000000000034000000000000003100000000",
            INIT_09 => X"0000003a000000000000002e000000000000002b000000000000002800000000",
            INIT_0A => X"0000000200000000000000040000000000000010000000000000003a00000000",
            INIT_0B => X"000000420000000000000037000000000000002d000000000000001300000000",
            INIT_0C => X"0000002800000000000000330000000000000038000000000000003d00000000",
            INIT_0D => X"00000000000000000000002e000000000000002e000000000000002d00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000005200000000000000460000000000000027000000000000001900000000",
            INIT_11 => X"0000004800000000000000540000000000000052000000000000005200000000",
            INIT_12 => X"0000004400000000000000500000000000000049000000000000004400000000",
            INIT_13 => X"0000005000000000000000510000000000000042000000000000004a00000000",
            INIT_14 => X"0000001d000000000000001d0000000000000019000000000000004a00000000",
            INIT_15 => X"00000020000000000000001b0000000000000019000000000000001c00000000",
            INIT_16 => X"0000003700000000000000340000000000000033000000000000002c00000000",
            INIT_17 => X"00000038000000000000003f000000000000003b000000000000003800000000",
            INIT_18 => X"0000000d00000000000000160000000000000018000000000000001400000000",
            INIT_19 => X"00000009000000000000000c000000000000000c000000000000000c00000000",
            INIT_1A => X"0000000300000000000000020000000000000006000000000000000700000000",
            INIT_1B => X"0000000000000000000000000000000000000001000000000000000400000000",
            INIT_1C => X"0000000000000000000000020000000000000004000000000000000400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000008000000000000000f0000000000000012000000000000000000000000",
            INIT_25 => X"00000008000000000000000f0000000000000010000000000000001000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000001b000000000000001b0000000000000016000000000000000900000000",
            INIT_29 => X"0000000f000000000000000f0000000000000012000000000000001000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000000000000000000004000000000000000f000000000000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_43 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_5A => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000003000000000000000200000000",
            INIT_5C => X"0000001800000000000000170000000000000016000000000000000000000000",
            INIT_5D => X"00000016000000000000001d000000000000001f000000000000001800000000",
            INIT_5E => X"0000000000000000000000000000000000000023000000000000001700000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_60 => X"0000001700000000000000040000000000000000000000000000003200000000",
            INIT_61 => X"0000000300000000000000050000000000000005000000000000000b00000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_63 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000010000000000000006000000000000000400000000",
            INIT_65 => X"0000000000000000000000020000000000000000000000000000000400000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000003000000000000000600000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000001000000000000000a0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000001400000000000000030000000000000000000000000000000000000000",
            INIT_77 => X"0000000700000000000000070000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000009000000000000000b0000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000008000000000000000700000000",
            INIT_7C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_7F => X"0000000000000000000000180000000000000000000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "samplegold_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000006000000000000000400000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000700000000000000050000000000000002000000000000000100000000",
            INIT_06 => X"0000000000000000000000000000000000000002000000000000000700000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_09 => X"0000000400000000000000080000000000000007000000000000000000000000",
            INIT_0A => X"0000000800000000000000070000000000000007000000000000000500000000",
            INIT_0B => X"0000000600000000000000080000000000000009000000000000000a00000000",
            INIT_0C => X"0000000700000000000000080000000000000015000000000000000a00000000",
            INIT_0D => X"0000000b0000000000000007000000000000000b000000000000000800000000",
            INIT_0E => X"00000011000000000000000f000000000000000d000000000000000e00000000",
            INIT_0F => X"00000000000000000000000b0000000000000006000000000000000d00000000",
            INIT_10 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_12 => X"00000000000000000000000d000000000000000a000000000000000700000000",
            INIT_13 => X"0000000800000000000000000000000000000000000000000000001600000000",
            INIT_14 => X"0000000500000000000000080000000000000003000000000000000000000000",
            INIT_15 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000700000000000000000000000000000008000000000000000400000000",
            INIT_17 => X"00000017000000000000001f0000000000000010000000000000000000000000",
            INIT_18 => X"0000000000000000000000060000000000000010000000000000000700000000",
            INIT_19 => X"00000014000000000000000a0000000000000009000000000000000000000000",
            INIT_1A => X"0000000d000000000000001a0000000000000000000000000000000000000000",
            INIT_1B => X"0000000900000000000000000000000000000001000000000000000900000000",
            INIT_1C => X"0000000800000000000000000000000000000000000000000000001200000000",
            INIT_1D => X"0000000000000000000000070000000000000000000000000000000700000000",
            INIT_1E => X"0000002800000000000000180000000000000022000000000000000b00000000",
            INIT_1F => X"00000000000000000000001c0000000000000002000000000000000b00000000",
            INIT_20 => X"0000000000000000000000070000000000000004000000000000000100000000",
            INIT_21 => X"00000004000000000000000e0000000000000000000000000000000000000000",
            INIT_22 => X"000000160000000000000024000000000000001e000000000000001800000000",
            INIT_23 => X"00000000000000000000000e0000000000000018000000000000000900000000",
            INIT_24 => X"0000000e000000000000000e0000000000000004000000000000000d00000000",
            INIT_25 => X"0000001d00000000000000010000000000000003000000000000000e00000000",
            INIT_26 => X"00000005000000000000000b000000000000001a000000000000002100000000",
            INIT_27 => X"0000000f0000000000000017000000000000001e000000000000001800000000",
            INIT_28 => X"0000001400000000000000140000000000000014000000000000000c00000000",
            INIT_29 => X"0000001500000000000000130000000000000019000000000000001400000000",
            INIT_2A => X"0000001b00000000000000080000000000000015000000000000001000000000",
            INIT_2B => X"00000012000000000000000c000000000000001b000000000000001d00000000",
            INIT_2C => X"00000015000000000000000a0000000000000014000000000000000c00000000",
            INIT_2D => X"00000022000000000000001b000000000000002a000000000000001c00000000",
            INIT_2E => X"0000001a0000000000000020000000000000000f000000000000000500000000",
            INIT_2F => X"0000001b0000000000000013000000000000002e000000000000001800000000",
            INIT_30 => X"0000002a00000000000000140000000000000021000000000000002200000000",
            INIT_31 => X"0000001c00000000000000150000000000000027000000000000002200000000",
            INIT_32 => X"000000220000000000000016000000000000001d000000000000002500000000",
            INIT_33 => X"0000001d0000000000000027000000000000002a000000000000000b00000000",
            INIT_34 => X"00000023000000000000001e0000000000000020000000000000002c00000000",
            INIT_35 => X"00000006000000000000002a0000000000000000000000000000000c00000000",
            INIT_36 => X"0000002400000000000000080000000000000000000000000000000b00000000",
            INIT_37 => X"0000002600000000000000330000000000000030000000000000000800000000",
            INIT_38 => X"000000080000000000000016000000000000001a000000000000002900000000",
            INIT_39 => X"0000000600000000000000030000000000000000000000000000001c00000000",
            INIT_3A => X"000000280000000000000004000000000000001a000000000000000800000000",
            INIT_3B => X"0000001e0000000000000026000000000000002b000000000000002900000000",
            INIT_3C => X"0000001700000000000000190000000000000014000000000000001e00000000",
            INIT_3D => X"00000009000000000000001b0000000000000024000000000000003000000000",
            INIT_3E => X"0000003400000000000000210000000000000011000000000000001300000000",
            INIT_3F => X"0000002200000000000000210000000000000026000000000000002600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000150000000000000016000000000000000b000000000000001700000000",
            INIT_41 => X"00000006000000000000000f0000000000000017000000000000001000000000",
            INIT_42 => X"000000030000000000000003000000000000000b000000000000000b00000000",
            INIT_43 => X"0000002500000000000000230000000000000027000000000000002a00000000",
            INIT_44 => X"00000000000000000000000b0000000000000002000000000000000400000000",
            INIT_45 => X"0000000c00000000000000180000000000000015000000000000000000000000",
            INIT_46 => X"0000001f0000000000000015000000000000000a000000000000000200000000",
            INIT_47 => X"000000000000000000000000000000000000001a000000000000003200000000",
            INIT_48 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"00000000000000000000002f0000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_4B => X"0000000300000000000000110000000000000000000000000000003800000000",
            INIT_4C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_4D => X"0000002000000000000000000000000000000016000000000000000000000000",
            INIT_4E => X"0000004600000000000000000000000000000006000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000001a000000000000002c00000000",
            INIT_52 => X"0000000000000000000000480000000000000004000000000000000000000000",
            INIT_53 => X"0000003300000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000002500000000000000130000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000002f0000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000027000000000000002c00000000",
            INIT_57 => X"0000000000000000000000360000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_59 => X"0000000000000000000000180000000000000004000000000000003a00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_5B => X"0000000000000000000000000000000000000030000000000000000000000000",
            INIT_5C => X"0000000f00000000000000000000000000000001000000000000002300000000",
            INIT_5D => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000013000000000000002200000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_62 => X"0000001400000000000000000000000000000000000000000000000900000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_64 => X"0000000800000000000000000000000000000004000000000000000500000000",
            INIT_65 => X"000000000000000000000000000000000000000e000000000000000500000000",
            INIT_66 => X"00000000000000000000000e0000000000000009000000000000000000000000",
            INIT_67 => X"000000180000000000000000000000000000000d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"000000020000000000000000000000000000001d000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_6E => X"0000000d00000000000000110000000000000000000000000000001200000000",
            INIT_6F => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000001d00000000000000190000000000000002000000000000000900000000",
            INIT_72 => X"0000001900000000000000000000000000000012000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_74 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000000e0000000000000006000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_7C => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_7D => X"0000000000000000000000140000000000000037000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "samplegold_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000004c000000000000001100000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000005000000000000000d000000000000000e000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000004000000000000000900000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000007000000000000000e0000000000000010000000000000000000000000",
            INIT_1D => X"000000000000000000000000000000000000000c000000000000000900000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000001100000000000000090000000000000002000000000000000000000000",
            INIT_21 => X"0000000000000000000000040000000000000006000000000000000b00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000500000000000000020000000000000001000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000b00000000000000090000000000000003000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_2C => X"0000000e000000000000000a0000000000000007000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000010000000000000009000000000000000e000000000000000000000000",
            INIT_30 => X"000000000000000000000007000000000000000a000000000000000000000000",
            INIT_31 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000400000000000000060000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000004000000000000000b00000000",
            INIT_35 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000070000000000000003000000000000000a000000000000000200000000",
            INIT_38 => X"0000007e00000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000620000000000000068000000000000005e000000000000005300000000",
            INIT_3A => X"0000009d00000000000000570000000000000074000000000000001000000000",
            INIT_3B => X"000000e5000000000000006400000000000000a0000000000000008d00000000",
            INIT_3C => X"0000008600000000000000a40000000000000063000000000000004200000000",
            INIT_3D => X"00000029000000000000005c000000000000007c000000000000009000000000",
            INIT_3E => X"000000880000000000000092000000000000004d000000000000004d00000000",
            INIT_3F => X"0000006f00000000000000ee000000000000006e000000000000009b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000800000000000000073000000000000009e00000000000000b400000000",
            INIT_41 => X"0000006c000000000000001c000000000000004a000000000000008100000000",
            INIT_42 => X"0000005b00000000000000960000000000000076000000000000009500000000",
            INIT_43 => X"000000ca00000000000000c10000000000000121000000000000009300000000",
            INIT_44 => X"0000007900000000000000ad000000000000005c000000000000007400000000",
            INIT_45 => X"0000005d00000000000000b90000000000000088000000000000003000000000",
            INIT_46 => X"000000bf00000000000000960000000000000077000000000000004a00000000",
            INIT_47 => X"0000008c00000000000000f800000000000000e6000000000000011800000000",
            INIT_48 => X"0000005d000000000000008600000000000000eb000000000000009700000000",
            INIT_49 => X"000000b2000000000000003100000000000000bd00000000000000cf00000000",
            INIT_4A => X"0000010c00000000000000bf00000000000000db00000000000000a500000000",
            INIT_4B => X"0000008c000000000000009500000000000000d900000000000000f100000000",
            INIT_4C => X"000000c500000000000000ae00000000000000c700000000000000ea00000000",
            INIT_4D => X"000000e400000000000000ef00000000000000d200000000000000b200000000",
            INIT_4E => X"000000de000000000000011600000000000000b200000000000000d800000000",
            INIT_4F => X"000000d10000000000000095000000000000009300000000000000d300000000",
            INIT_50 => X"000000c600000000000000d500000000000000f0000000000000010700000000",
            INIT_51 => X"000000d600000000000000d300000000000000d100000000000000e500000000",
            INIT_52 => X"000000cc00000000000000e200000000000000fa00000000000000f800000000",
            INIT_53 => X"000000f600000000000000ce0000000000000098000000000000009e00000000",
            INIT_54 => X"000000ed00000000000000ce00000000000000d800000000000000f600000000",
            INIT_55 => X"000000f400000000000000f200000000000000f100000000000000f700000000",
            INIT_56 => X"000000a300000000000000ba00000000000000e5000000000000012000000000",
            INIT_57 => X"000000e900000000000000d200000000000000d700000000000000d100000000",
            INIT_58 => X"00000114000000000000010300000000000000f100000000000000f600000000",
            INIT_59 => X"000000ff000000000000010900000000000000fe000000000000010c00000000",
            INIT_5A => X"000000c900000000000000d8000000000000009600000000000000d200000000",
            INIT_5B => X"000000c900000000000000c2000000000000009c00000000000000a700000000",
            INIT_5C => X"00000131000000000000011e000000000000011900000000000000fd00000000",
            INIT_5D => X"0000009100000000000000e50000000000000109000000000000010000000000",
            INIT_5E => X"000000ae000000000000008400000000000000db000000000000007e00000000",
            INIT_5F => X"000000d900000000000000c300000000000000bb000000000000009600000000",
            INIT_60 => X"000000ff00000000000001190000000000000132000000000000014200000000",
            INIT_61 => X"000000e200000000000000a800000000000000e200000000000000fa00000000",
            INIT_62 => X"000000ba0000000000000104000000000000011b00000000000000b500000000",
            INIT_63 => X"0000012c000000000000010900000000000000bc00000000000000d600000000",
            INIT_64 => X"0000010700000000000001070000000000000115000000000000012700000000",
            INIT_65 => X"000000df00000000000000d900000000000000be00000000000000e700000000",
            INIT_66 => X"000000e0000000000000011a000000000000014100000000000000ee00000000",
            INIT_67 => X"000000c4000000000000010d000000000000010600000000000000c600000000",
            INIT_68 => X"000000e400000000000001080000000000000121000000000000010f00000000",
            INIT_69 => X"0000007400000000000000ac00000000000000ce000000000000008600000000",
            INIT_6A => X"000000e80000000000000132000000000000012500000000000000b800000000",
            INIT_6B => X"0000010b00000000000000ba00000000000000ba00000000000000d500000000",
            INIT_6C => X"0000005a00000000000000bf0000000000000109000000000000010b00000000",
            INIT_6D => X"0000005e000000000000004900000000000000ab000000000000009e00000000",
            INIT_6E => X"000001170000000000000144000000000000013700000000000000d500000000",
            INIT_6F => X"000000e800000000000000d000000000000000d700000000000000f400000000",
            INIT_70 => X"000000cc0000000000000096000000000000009b00000000000000be00000000",
            INIT_71 => X"0000000000000000000000030000000000000003000000000000001700000000",
            INIT_72 => X"00000004000000000000000f0000000000000000000000000000001000000000",
            INIT_73 => X"000000000000000000000029000000000000001c000000000000002200000000",
            INIT_74 => X"00000010000000000000000c0000000000000003000000000000004f00000000",
            INIT_75 => X"0000000e00000000000000050000000000000010000000000000000f00000000",
            INIT_76 => X"0000001e0000000000000000000000000000000b000000000000000000000000",
            INIT_77 => X"0000004c00000000000000000000000000000027000000000000000f00000000",
            INIT_78 => X"0000001d0000000000000029000000000000001a000000000000000200000000",
            INIT_79 => X"000000000000000000000006000000000000000e000000000000000e00000000",
            INIT_7A => X"0000001d0000000000000006000000000000001a000000000000000300000000",
            INIT_7B => X"0000001800000000000000540000000000000000000000000000001d00000000",
            INIT_7C => X"0000001d00000000000000000000000000000017000000000000003200000000",
            INIT_7D => X"0000002e00000000000000120000000000000000000000000000000e00000000",
            INIT_7E => X"0000001900000000000000100000000000000004000000000000000900000000",
            INIT_7F => X"0000004700000000000000280000000000000056000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "samplegold_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000023000000000000002f000000000000000d000000000000001000000000",
            INIT_01 => X"0000000000000000000000270000000000000023000000000000000500000000",
            INIT_02 => X"0000001e000000000000003b000000000000001c000000000000001b00000000",
            INIT_03 => X"000000190000000000000046000000000000002b000000000000004400000000",
            INIT_04 => X"000000180000000000000010000000000000002f000000000000001300000000",
            INIT_05 => X"0000002f000000000000001f0000000000000040000000000000002e00000000",
            INIT_06 => X"00000046000000000000001a000000000000003b000000000000002f00000000",
            INIT_07 => X"0000000b00000000000000170000000000000046000000000000002900000000",
            INIT_08 => X"000000420000000000000047000000000000003a000000000000001f00000000",
            INIT_09 => X"00000046000000000000004b0000000000000039000000000000004100000000",
            INIT_0A => X"0000002400000000000000480000000000000034000000000000003e00000000",
            INIT_0B => X"000000180000000000000011000000000000001c000000000000003b00000000",
            INIT_0C => X"00000044000000000000003b0000000000000044000000000000004000000000",
            INIT_0D => X"00000043000000000000003e0000000000000049000000000000005b00000000",
            INIT_0E => X"0000002a0000000000000036000000000000004a000000000000004f00000000",
            INIT_0F => X"0000002b00000000000000270000000000000016000000000000001600000000",
            INIT_10 => X"0000005100000000000000440000000000000047000000000000003e00000000",
            INIT_11 => X"0000004000000000000000630000000000000058000000000000004e00000000",
            INIT_12 => X"00000025000000000000001e0000000000000033000000000000006c00000000",
            INIT_13 => X"0000002900000000000000260000000000000020000000000000002600000000",
            INIT_14 => X"0000005b000000000000004c000000000000003f000000000000004e00000000",
            INIT_15 => X"0000004a0000000000000058000000000000004f000000000000005c00000000",
            INIT_16 => X"00000020000000000000002f000000000000000f000000000000002000000000",
            INIT_17 => X"0000001900000000000000170000000000000010000000000000002100000000",
            INIT_18 => X"00000061000000000000005b0000000000000057000000000000004300000000",
            INIT_19 => X"0000001a000000000000004a0000000000000058000000000000004e00000000",
            INIT_1A => X"00000038000000000000002e0000000000000018000000000000002300000000",
            INIT_1B => X"000000400000000000000021000000000000002f000000000000001200000000",
            INIT_1C => X"0000004e00000000000000590000000000000056000000000000006800000000",
            INIT_1D => X"0000002700000000000000280000000000000058000000000000005f00000000",
            INIT_1E => X"00000040000000000000005d0000000000000057000000000000003a00000000",
            INIT_1F => X"0000006c00000000000000460000000000000035000000000000002700000000",
            INIT_20 => X"00000055000000000000005d0000000000000054000000000000004500000000",
            INIT_21 => X"0000003100000000000000280000000000000016000000000000005a00000000",
            INIT_22 => X"0000004a00000000000000570000000000000049000000000000001f00000000",
            INIT_23 => X"000000190000000000000033000000000000003d000000000000002b00000000",
            INIT_24 => X"0000004b00000000000000610000000000000058000000000000005600000000",
            INIT_25 => X"0000000a000000000000003a0000000000000004000000000000001700000000",
            INIT_26 => X"0000004000000000000000610000000000000045000000000000001700000000",
            INIT_27 => X"000000510000000000000047000000000000002f000000000000003f00000000",
            INIT_28 => X"00000007000000000000001e0000000000000041000000000000005a00000000",
            INIT_29 => X"0000000000000000000000140000000000000004000000000000002400000000",
            INIT_2A => X"000000030000000000000000000000000000003b000000000000000000000000",
            INIT_2B => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"000000000000000000000000000000000000006e000000000000000000000000",
            INIT_2D => X"000000000000000000000009000000000000000b000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000004000000000",
            INIT_2F => X"0000000000000000000000270000000000000000000000000000000400000000",
            INIT_30 => X"0000000b000000000000000d0000000000000000000000000000006200000000",
            INIT_31 => X"0000003400000000000000050000000000000005000000000000000000000000",
            INIT_32 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_33 => X"0000003200000000000000000000000000000000000000000000002500000000",
            INIT_34 => X"0000000000000000000000220000000000000012000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000001b000000000000001600000000",
            INIT_36 => X"0000002300000000000000000000000000000029000000000000001700000000",
            INIT_37 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_38 => X"0000003a00000000000000000000000000000020000000000000004900000000",
            INIT_39 => X"0000004f00000000000000000000000000000000000000000000001700000000",
            INIT_3A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000007d0000000000000000000000000000000b000000000000000000000000",
            INIT_3C => X"0000004400000000000000000000000000000000000000000000003800000000",
            INIT_3D => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000130000000000000000000000000000000800000000",
            INIT_3F => X"0000002c00000000000000830000000000000000000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000018000000000000000d0000000000000000000000000000000000000000",
            INIT_41 => X"0000000c00000000000000000000000000000008000000000000000000000000",
            INIT_42 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"00000000000000000000001c0000000000000067000000000000000000000000",
            INIT_44 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000002f0000000000000000000000000000000800000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000005a00000000",
            INIT_48 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_49 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000003f00000000000000120000000000000027000000000000000000000000",
            INIT_4B => X"0000000000000000000000160000000000000008000000000000000000000000",
            INIT_4C => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_4D => X"0000000f0000000000000003000000000000000d000000000000000000000000",
            INIT_4E => X"000000390000000000000000000000000000000a000000000000002f00000000",
            INIT_4F => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_50 => X"0000000700000000000000040000000000000000000000000000000900000000",
            INIT_51 => X"0000001c000000000000000b0000000000000002000000000000001200000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000000b0000000000000000000000000000003600000000",
            INIT_54 => X"0000002000000000000000040000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000210000000000000009000000000000000000000000",
            INIT_56 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000000000000000000001a000000000000001e00000000",
            INIT_58 => X"0000000000000000000000040000000000000000000000000000001d00000000",
            INIT_59 => X"0000000000000000000000000000000000000025000000000000002300000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_5B => X"0000001500000000000000000000000000000003000000000000002b00000000",
            INIT_5C => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000003700000000000000000000000000000000000000000000004900000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_5F => X"0000000b00000000000000000000000000000012000000000000001c00000000",
            INIT_60 => X"0000002a000000000000000f0000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_66 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6B => X"0000000000000000000000160000000000000001000000000000000000000000",
            INIT_6C => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000c00000000000000110000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "samplegold_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000001c0000000000000000000000000000000200000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001100000000000000020000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_11 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000002800000000000000210000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_16 => X"0000000300000000000000160000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_1B => X"00000000000000000000000c0000000000000000000000000000002f00000000",
            INIT_1C => X"0000000000000000000000390000000000000000000000000000000600000000",
            INIT_1D => X"0000000000000000000000000000000000000004000000000000001e00000000",
            INIT_1E => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000018000000000000000200000000",
            INIT_20 => X"0000001500000000000000000000000000000045000000000000000000000000",
            INIT_21 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_22 => X"0000000100000000000000270000000000000000000000000000000000000000",
            INIT_23 => X"0000002100000000000000000000000000000010000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_25 => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000011000000000000000100000000",
            INIT_27 => X"0000001800000000000000150000000000000000000000000000002a00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000003200000000000000000000000000000000000000000000003f00000000",
            INIT_2A => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_2B => X"00000000000000000000000a0000000000000000000000000000000600000000",
            INIT_2C => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_30 => X"0000000c000000000000001d0000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000800000000000000040000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_35 => X"0000000200000000000000180000000000000000000000000000000000000000",
            INIT_36 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000200000000000000000000000000000001000000000000000000000000",
            INIT_38 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000b00000000000000010000000000000012000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000005000000000000000a00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000000000000000000001f0000000000000000000000000000001c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002e00000000000000000000000000000000000000000000001100000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_44 => X"00000000000000000000000c000000000000000a000000000000000000000000",
            INIT_45 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_48 => X"0000002900000000000000000000000000000000000000000000000d00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000d00000000000000000000000000000000000000000000001200000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000004900000000",
            INIT_4C => X"0000000400000000000000090000000000000000000000000000000000000000",
            INIT_4D => X"0000002b00000000000000000000000000000000000000000000000600000000",
            INIT_4E => X"0000002600000000000000000000000000000000000000000000001200000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_50 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_51 => X"0000002800000000000000000000000000000000000000000000000200000000",
            INIT_52 => X"0000000000000000000000070000000000000009000000000000000a00000000",
            INIT_53 => X"0000000200000000000000050000000000000004000000000000000000000000",
            INIT_54 => X"0000000400000000000000050000000000000000000000000000000600000000",
            INIT_55 => X"0000000400000000000000040000000000000000000000000000001400000000",
            INIT_56 => X"0000000200000000000000000000000000000003000000000000000d00000000",
            INIT_57 => X"0000000600000000000000040000000000000000000000000000000100000000",
            INIT_58 => X"0000001400000000000000050000000000000004000000000000000600000000",
            INIT_59 => X"0000000000000000000000020000000000000009000000000000000e00000000",
            INIT_5A => X"0000000500000000000000010000000000000000000000000000000000000000",
            INIT_5B => X"0000000200000000000000000000000000000008000000000000000b00000000",
            INIT_5C => X"0000000600000000000000150000000000000007000000000000000000000000",
            INIT_5D => X"0000000b00000000000000020000000000000000000000000000000c00000000",
            INIT_5E => X"00000005000000000000000c0000000000000007000000000000000800000000",
            INIT_5F => X"00000013000000000000000c0000000000000002000000000000000000000000",
            INIT_60 => X"000000090000000000000009000000000000000d000000000000000600000000",
            INIT_61 => X"0000000c000000000000000a0000000000000000000000000000000400000000",
            INIT_62 => X"0000000a0000000000000009000000000000000e000000000000000c00000000",
            INIT_63 => X"000000030000000000000011000000000000000a000000000000000c00000000",
            INIT_64 => X"0000000800000000000000060000000000000005000000000000000e00000000",
            INIT_65 => X"0000000d000000000000000d0000000000000001000000000000000000000000",
            INIT_66 => X"00000015000000000000001a0000000000000025000000000000001200000000",
            INIT_67 => X"0000000b00000000000000120000000000000012000000000000001300000000",
            INIT_68 => X"00000003000000000000000c000000000000000e000000000000000200000000",
            INIT_69 => X"0000001f0000000000000020000000000000000f000000000000000000000000",
            INIT_6A => X"0000001e00000000000000200000000000000021000000000000002800000000",
            INIT_6B => X"0000000500000000000000120000000000000022000000000000002400000000",
            INIT_6C => X"0000000400000000000000000000000000000003000000000000000b00000000",
            INIT_6D => X"0000001a0000000000000020000000000000001b000000000000000700000000",
            INIT_6E => X"00000025000000000000002a0000000000000028000000000000002800000000",
            INIT_6F => X"00000001000000000000000d0000000000000026000000000000001e00000000",
            INIT_70 => X"0000000000000000000000010000000000000008000000000000000900000000",
            INIT_71 => X"0000002400000000000000230000000000000022000000000000000b00000000",
            INIT_72 => X"0000001f00000000000000260000000000000020000000000000002400000000",
            INIT_73 => X"0000000900000000000000070000000000000010000000000000001f00000000",
            INIT_74 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_75 => X"000000260000000000000022000000000000001c000000000000000f00000000",
            INIT_76 => X"0000001900000000000000210000000000000022000000000000002300000000",
            INIT_77 => X"0000000a00000000000000050000000000000001000000000000000c00000000",
            INIT_78 => X"0000000400000000000000070000000000000002000000000000000a00000000",
            INIT_79 => X"0000002200000000000000210000000000000021000000000000001500000000",
            INIT_7A => X"0000000d00000000000000220000000000000023000000000000002000000000",
            INIT_7B => X"0000001d00000000000000270000000000000011000000000000000a00000000",
            INIT_7C => X"0000001600000000000000070000000000000005000000000000000900000000",
            INIT_7D => X"0000002400000000000000220000000000000020000000000000002400000000",
            INIT_7E => X"0000000000000000000000100000000000000023000000000000002800000000",
            INIT_7F => X"0000001a000000000000001e0000000000000005000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "samplegold_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001b0000000000000011000000000000000b000000000000000c00000000",
            INIT_01 => X"0000002500000000000000250000000000000022000000000000000f00000000",
            INIT_02 => X"0000000a00000000000000000000000000000008000000000000002300000000",
            INIT_03 => X"0000001b00000000000000190000000000000000000000000000000000000000",
            INIT_04 => X"00000011000000000000000f0000000000000009000000000000000d00000000",
            INIT_05 => X"0000001200000000000000240000000000000022000000000000001d00000000",
            INIT_06 => X"00000006000000000000000b0000000000000000000000000000000800000000",
            INIT_07 => X"00000019000000000000001b0000000000000000000000000000000400000000",
            INIT_08 => X"0000001500000000000000130000000000000009000000000000001400000000",
            INIT_09 => X"0000000b0000000000000015000000000000000f000000000000001400000000",
            INIT_0A => X"0000000000000000000000050000000000000000000000000000000e00000000",
            INIT_0B => X"0000000000000000000000060000000000000007000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000001000000000000000900000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000001a000000000000001b00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000021000000000000000c000000000000000b000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "samplegold_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_01 => X"0000003300000000000000210000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_03 => X"00000031000000000000002d0000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000030000000000000006000000000000000f000000000000000000000000",
            INIT_06 => X"00000000000000000000000a0000000000000025000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000001b000000000000002000000000",
            INIT_08 => X"0000000000000000000000260000000000000011000000000000000000000000",
            INIT_09 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000c00000000000000000000000000000018000000000000000000000000",
            INIT_0B => X"0000001500000000000000370000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000000000000000000001c0000000000000046000000000000000000000000",
            INIT_0F => X"0000000000000000000000060000000000000010000000000000000d00000000",
            INIT_10 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_12 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000600000000000000000000000000000000000000000000000300000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_17 => X"00000000000000000000000a000000000000002a000000000000000c00000000",
            INIT_18 => X"0000001400000000000000000000000000000000000000000000001500000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_1F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000300000000000000000000000000000000000000000000001300000000",
            INIT_21 => X"0000000000000000000000000000000000000005000000000000000200000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000009000000000000000e0000000000000002000000000000000000000000",
            INIT_24 => X"00000003000000000000003d0000000000000060000000000000004000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000110000000000000015000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_30 => X"0000001300000000000000240000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000a0000000000000035000000000000003f000000000000000000000000",
            INIT_33 => X"00000023000000000000002a0000000000000017000000000000001d00000000",
            INIT_34 => X"0000002500000000000000200000000000000033000000000000000c00000000",
            INIT_35 => X"0000003500000000000000150000000000000028000000000000002900000000",
            INIT_36 => X"0000001e000000000000001d0000000000000032000000000000000600000000",
            INIT_37 => X"00000007000000000000001f0000000000000022000000000000001900000000",
            INIT_38 => X"00000021000000000000002b0000000000000022000000000000003000000000",
            INIT_39 => X"0000000a000000000000003d0000000000000019000000000000002600000000",
            INIT_3A => X"0000001d0000000000000011000000000000001d000000000000002e00000000",
            INIT_3B => X"0000003500000000000000090000000000000016000000000000001b00000000",
            INIT_3C => X"00000011000000000000002a0000000000000020000000000000003000000000",
            INIT_3D => X"00000023000000000000000f000000000000003e000000000000002d00000000",
            INIT_3E => X"00000013000000000000003d000000000000001a000000000000001800000000",
            INIT_3F => X"00000026000000000000003f000000000000001e000000000000001300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004200000000000000110000000000000032000000000000001a00000000",
            INIT_41 => X"00000006000000000000001c0000000000000019000000000000003600000000",
            INIT_42 => X"00000013000000000000000c000000000000003e000000000000001300000000",
            INIT_43 => X"0000002d0000000000000013000000000000002b000000000000002e00000000",
            INIT_44 => X"00000037000000000000002b0000000000000031000000000000003400000000",
            INIT_45 => X"0000000600000000000000000000000000000018000000000000001f00000000",
            INIT_46 => X"00000037000000000000000b000000000000001c000000000000003b00000000",
            INIT_47 => X"0000001e000000000000002a0000000000000005000000000000002100000000",
            INIT_48 => X"0000001a0000000000000032000000000000001c000000000000002800000000",
            INIT_49 => X"00000034000000000000000b0000000000000000000000000000001f00000000",
            INIT_4A => X"0000001900000000000000120000000000000014000000000000002800000000",
            INIT_4B => X"000000120000000000000013000000000000001f000000000000001500000000",
            INIT_4C => X"000000260000000000000015000000000000001c000000000000001400000000",
            INIT_4D => X"0000001e000000000000002e0000000000000012000000000000000000000000",
            INIT_4E => X"0000001f000000000000000d0000000000000014000000000000001700000000",
            INIT_4F => X"0000001000000000000000180000000000000014000000000000000f00000000",
            INIT_50 => X"00000000000000000000001e0000000000000000000000000000001800000000",
            INIT_51 => X"0000001e00000000000000190000000000000022000000000000001f00000000",
            INIT_52 => X"0000000f00000000000000180000000000000000000000000000001e00000000",
            INIT_53 => X"00000010000000000000000b0000000000000012000000000000001300000000",
            INIT_54 => X"00000016000000000000000a000000000000000f000000000000000200000000",
            INIT_55 => X"0000001f00000000000000210000000000000011000000000000001800000000",
            INIT_56 => X"0000000a000000000000000e0000000000000009000000000000002000000000",
            INIT_57 => X"00000008000000000000000b000000000000000c000000000000000a00000000",
            INIT_58 => X"00000028000000000000000a0000000000000029000000000000001700000000",
            INIT_59 => X"0000001400000000000000200000000000000031000000000000001600000000",
            INIT_5A => X"000000040000000000000006000000000000000b000000000000002800000000",
            INIT_5B => X"0000001d000000000000000d000000000000000e000000000000000e00000000",
            INIT_5C => X"0000001b000000000000002d000000000000001f000000000000002400000000",
            INIT_5D => X"0000001c0000000000000025000000000000001a000000000000003100000000",
            INIT_5E => X"0000001300000000000000000000000000000009000000000000000e00000000",
            INIT_5F => X"000000260000000000000020000000000000000f000000000000000b00000000",
            INIT_60 => X"0000002100000000000000210000000000000030000000000000001d00000000",
            INIT_61 => X"00000005000000000000001b0000000000000026000000000000002400000000",
            INIT_62 => X"000000070000000000000011000000000000000a000000000000001600000000",
            INIT_63 => X"0000001600000000000000230000000000000027000000000000000b00000000",
            INIT_64 => X"00000023000000000000002b000000000000003f000000000000002f00000000",
            INIT_65 => X"00000027000000000000001e000000000000002d000000000000002f00000000",
            INIT_66 => X"000000040000000000000002000000000000000b000000000000001100000000",
            INIT_67 => X"0000002500000000000000110000000000000039000000000000002500000000",
            INIT_68 => X"00000027000000000000002a0000000000000040000000000000004600000000",
            INIT_69 => X"0000001400000000000000180000000000000030000000000000002f00000000",
            INIT_6A => X"0000003800000000000000120000000000000012000000000000000f00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_6C => X"000000040000000000000000000000000000001b000000000000000900000000",
            INIT_6D => X"0000000e00000000000000020000000000000008000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_6F => X"0000000c000000000000000a0000000000000000000000000000000200000000",
            INIT_70 => X"0000000000000000000000080000000000000000000000000000001200000000",
            INIT_71 => X"00000000000000000000000e0000000000000000000000000000000100000000",
            INIT_72 => X"0000001a000000000000000d0000000000000000000000000000000000000000",
            INIT_73 => X"0000000800000000000000120000000000000004000000000000000200000000",
            INIT_74 => X"00000009000000000000000f0000000000000000000000000000000000000000",
            INIT_75 => X"0000000800000000000000000000000000000000000000000000001b00000000",
            INIT_76 => X"00000000000000000000000e0000000000000005000000000000000400000000",
            INIT_77 => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_78 => X"000000000000000000000000000000000000000a000000000000000e00000000",
            INIT_79 => X"0000000500000000000000120000000000000000000000000000000000000000",
            INIT_7A => X"000000120000000000000000000000000000000b000000000000003300000000",
            INIT_7B => X"0000000d00000000000000000000000000000000000000000000000700000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000003200000000000000120000000000000007000000000000000000000000",
            INIT_7E => X"00000000000000000000000d0000000000000005000000000000001000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "samplegold_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000220000000000000014000000000000000a00000000",
            INIT_02 => X"00000000000000000000000d0000000000000008000000000000000100000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000100000000000000070000000000000013000000000000000900000000",
            INIT_06 => X"0000000000000000000000000000000000000011000000000000000100000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000001600000000000000000000000000000000000000000000002400000000",
            INIT_0A => X"000000000000000000000000000000000000000a000000000000001100000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"00000005000000000000000c0000000000000004000000000000000000000000",
            INIT_0D => X"00000006000000000000000f0000000000000016000000000000000f00000000",
            INIT_0E => X"0000000000000000000000000000000000000007000000000000001400000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000002300000000000000000000000000000000000000000000000200000000",
            INIT_11 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_15 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000040000000000000022000000000000000e00000000",
            INIT_19 => X"0000000b00000000000000030000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_1B => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000000000000000000000000000e000000000000001200000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001700000000000000000000000000000000000000000000001300000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000012000000000000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000002000000000000000a000000000000000000000000",
            INIT_3C => X"000000000000000000000003000000000000000b000000000000000100000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000001000000000000000b000000000000000f000000000000000300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000800000000000000020000000000000006000000000000000900000000",
            INIT_44 => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_47 => X"0000000400000000000000000000000000000002000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_4B => X"0000000300000000000000050000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_4F => X"0000000100000000000000090000000000000001000000000000000000000000",
            INIT_50 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"000000000000000000000018000000000000000b000000000000000000000000",
            INIT_53 => X"0000000000000000000000030000000000000000000000000000000400000000",
            INIT_54 => X"0000000a00000000000000100000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000900000000000000090000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_58 => X"00000002000000000000000d0000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000130000000000000009000000000000000000000000",
            INIT_5B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000004000000000000000a0000000000000004000000000000002100000000",
            INIT_5D => X"0000000d00000000000000200000000000000009000000000000001500000000",
            INIT_5E => X"00000000000000000000002b0000000000000008000000000000001b00000000",
            INIT_5F => X"0000002f0000000000000013000000000000001b000000000000000900000000",
            INIT_60 => X"0000000900000000000000170000000000000009000000000000000b00000000",
            INIT_61 => X"00000018000000000000000d0000000000000022000000000000000700000000",
            INIT_62 => X"0000001700000000000000040000000000000021000000000000000500000000",
            INIT_63 => X"000000100000000000000019000000000000000b000000000000000200000000",
            INIT_64 => X"000000180000000000000012000000000000001f000000000000001300000000",
            INIT_65 => X"000000030000000000000013000000000000000f000000000000001000000000",
            INIT_66 => X"0000000c00000000000000120000000000000004000000000000002800000000",
            INIT_67 => X"0000000b00000000000000140000000000000001000000000000000800000000",
            INIT_68 => X"0000001b0000000000000011000000000000000f000000000000003400000000",
            INIT_69 => X"0000002a00000000000000030000000000000020000000000000001000000000",
            INIT_6A => X"0000001a00000000000000000000000000000015000000000000000300000000",
            INIT_6B => X"00000022000000000000001c0000000000000003000000000000000000000000",
            INIT_6C => X"0000000c000000000000002e000000000000000d000000000000001d00000000",
            INIT_6D => X"00000010000000000000003a0000000000000013000000000000001d00000000",
            INIT_6E => X"0000000000000000000000200000000000000000000000000000000900000000",
            INIT_6F => X"000000230000000000000011000000000000001b000000000000000d00000000",
            INIT_70 => X"0000002500000000000000250000000000000010000000000000003900000000",
            INIT_71 => X"0000000a00000000000000130000000000000039000000000000002400000000",
            INIT_72 => X"0000001f00000000000000010000000000000025000000000000000000000000",
            INIT_73 => X"0000002d000000000000001d000000000000002e000000000000001a00000000",
            INIT_74 => X"0000002600000000000000220000000000000028000000000000001700000000",
            INIT_75 => X"0000001300000000000000150000000000000028000000000000002600000000",
            INIT_76 => X"0000000e0000000000000019000000000000000a000000000000001c00000000",
            INIT_77 => X"0000002c00000000000000170000000000000037000000000000001000000000",
            INIT_78 => X"0000001e00000000000000220000000000000021000000000000001f00000000",
            INIT_79 => X"0000001f00000000000000160000000000000012000000000000001a00000000",
            INIT_7A => X"000000150000000000000015000000000000001d000000000000001600000000",
            INIT_7B => X"0000001600000000000000200000000000000022000000000000001a00000000",
            INIT_7C => X"0000001a000000000000001c000000000000002f000000000000001b00000000",
            INIT_7D => X"0000001600000000000000130000000000000015000000000000001900000000",
            INIT_7E => X"000000200000000000000003000000000000000c000000000000001900000000",
            INIT_7F => X"0000000c00000000000000260000000000000015000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "samplegold_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000e0000000000000006000000000000001a000000000000002900000000",
            INIT_01 => X"0000001c000000000000001c0000000000000008000000000000002100000000",
            INIT_02 => X"00000017000000000000000c000000000000001d000000000000000500000000",
            INIT_03 => X"00000017000000000000001b0000000000000012000000000000001200000000",
            INIT_04 => X"000000060000000000000020000000000000001d000000000000001e00000000",
            INIT_05 => X"0000001d00000000000000270000000000000011000000000000002f00000000",
            INIT_06 => X"00000019000000000000000e0000000000000015000000000000001300000000",
            INIT_07 => X"00000020000000000000000a0000000000000023000000000000001600000000",
            INIT_08 => X"0000000c000000000000001c000000000000001e000000000000002600000000",
            INIT_09 => X"000000190000000000000033000000000000002f000000000000001f00000000",
            INIT_0A => X"0000001e000000000000000e000000000000000f000000000000001f00000000",
            INIT_0B => X"00000018000000000000001e0000000000000016000000000000001b00000000",
            INIT_0C => X"0000001c00000000000000020000000000000018000000000000003400000000",
            INIT_0D => X"00000021000000000000002e0000000000000030000000000000001700000000",
            INIT_0E => X"0000000f00000000000000200000000000000014000000000000001b00000000",
            INIT_0F => X"0000001d000000000000000d0000000000000023000000000000001e00000000",
            INIT_10 => X"0000001e00000000000000050000000000000007000000000000001300000000",
            INIT_11 => X"00000029000000000000002f000000000000002d000000000000001a00000000",
            INIT_12 => X"0000000f000000000000000b000000000000002d000000000000001600000000",
            INIT_13 => X"0000002100000000000000070000000000000025000000000000001600000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_17 => X"0000000d00000000000000070000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000110000000000000000000000000000000700000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000100000000000000030000000000000000000000000000000000000000",
            INIT_1F => X"000000020000000000000004000000000000000c000000000000000300000000",
            INIT_20 => X"0000000000000000000000010000000000000003000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000200000000000000030000000000000004000000000000001300000000",
            INIT_24 => X"0000000000000000000000030000000000000002000000000000000000000000",
            INIT_25 => X"0000000c00000000000000060000000000000000000000000000000600000000",
            INIT_26 => X"0000000000000000000000050000000000000003000000000000000000000000",
            INIT_27 => X"0000000500000000000000040000000000000000000000000000000b00000000",
            INIT_28 => X"00000018000000000000001a000000000000001f000000000000000000000000",
            INIT_29 => X"0000000000000000000000040000000000000011000000000000000000000000",
            INIT_2A => X"0000000e00000000000000000000000000000001000000000000000100000000",
            INIT_2B => X"0000001c00000000000000000000000000000013000000000000001500000000",
            INIT_2C => X"000000080000000000000000000000000000000b000000000000001e00000000",
            INIT_2D => X"0000000000000000000000000000000000000007000000000000001600000000",
            INIT_2E => X"0000001b00000000000000000000000000000009000000000000000100000000",
            INIT_2F => X"0000001100000000000000120000000000000014000000000000000f00000000",
            INIT_30 => X"0000001a000000000000001f0000000000000022000000000000001800000000",
            INIT_31 => X"0000000200000000000000000000000000000000000000000000000e00000000",
            INIT_32 => X"0000001f0000000000000014000000000000000c000000000000000200000000",
            INIT_33 => X"0000002200000000000000230000000000000018000000000000002900000000",
            INIT_34 => X"0000000200000000000000260000000000000030000000000000002900000000",
            INIT_35 => X"0000000c00000000000000190000000000000003000000000000000000000000",
            INIT_36 => X"0000000000000000000000350000000000000022000000000000000400000000",
            INIT_37 => X"000000100000000000000000000000000000001a000000000000002600000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_39 => X"0000001100000000000000110000000000000020000000000000000000000000",
            INIT_3A => X"0000000d00000000000000060000000000000013000000000000002b00000000",
            INIT_3B => X"0000000900000000000000110000000000000014000000000000001000000000",
            INIT_3C => X"0000000700000000000000000000000000000000000000000000000500000000",
            INIT_3D => X"000000110000000000000014000000000000000c000000000000002300000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000f00000000000000110000000000000000000000000000000000000000",
            INIT_41 => X"0000000a0000000000000017000000000000000b000000000000000c00000000",
            INIT_42 => X"0000000000000000000000000000000000000014000000000000000600000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000001100000000000000020000000000000000000000000000000000000000",
            INIT_45 => X"0000001000000000000000180000000000000014000000000000000b00000000",
            INIT_46 => X"00000000000000000000000f0000000000000005000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_48 => X"0000000c00000000000000000000000000000003000000000000000000000000",
            INIT_49 => X"0000000700000000000000080000000000000004000000000000000a00000000",
            INIT_4A => X"00000003000000000000000d0000000000000009000000000000000b00000000",
            INIT_4B => X"0000000400000000000000050000000000000000000000000000000100000000",
            INIT_4C => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000100000000000000000000000000000000000000000000000500000000",
            INIT_4F => X"000000000000000000000014000000000000000b000000000000000000000000",
            INIT_50 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_52 => X"00000004000000000000000b0000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000040000000000000000000000000000000600000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_56 => X"0000000300000000000000000000000000000021000000000000000000000000",
            INIT_57 => X"0000000400000000000000000000000000000002000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000070000000000000000000000000000000300000000",
            INIT_5C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5D => X"00000000000000000000000a0000000000000000000000000000000100000000",
            INIT_5E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_5F => X"0000000000000000000000120000000000000000000000000000003d00000000",
            INIT_60 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_62 => X"0000005300000000000000060000000000000000000000000000000e00000000",
            INIT_63 => X"0000001100000000000000000000000000000000000000000000000d00000000",
            INIT_64 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000e00000000000000000000000000000000000000000000001000000000",
            INIT_66 => X"0000004100000000000000000000000000000001000000000000000700000000",
            INIT_67 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_69 => X"0000001700000000000000130000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000025000000000000002f000000000000000000000000",
            INIT_6E => X"000000000000000000000000000000000000003f000000000000000000000000",
            INIT_6F => X"0000001a00000000000000000000000000000000000000000000003000000000",
            INIT_70 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_71 => X"000000000000000000000000000000000000003f000000000000002600000000",
            INIT_72 => X"0000001500000000000000000000000000000000000000000000001f00000000",
            INIT_73 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_74 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000600000000000000000000000000000000000000000000003f00000000",
            INIT_76 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_78 => X"00000016000000000000001a000000000000000b000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_7A => X"0000000900000000000000000000000000000000000000000000000900000000",
            INIT_7B => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_7C => X"000000140000000000000003000000000000001e000000000000001600000000",
            INIT_7D => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_7E => X"0000000000000000000000160000000000000008000000000000000000000000",
            INIT_7F => X"0000001800000000000000080000000000000000000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "samplegold_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000200000000000000000000000000000016000000000000000900000000",
            INIT_01 => X"00000001000000000000000e0000000000000000000000000000001400000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_03 => X"00000000000000000000000a000000000000000b000000000000000000000000",
            INIT_04 => X"0000002500000000000000310000000000000012000000000000000000000000",
            INIT_05 => X"0000004800000000000000480000000000000041000000000000003f00000000",
            INIT_06 => X"0000001500000000000000240000000000000036000000000000004400000000",
            INIT_07 => X"0000001500000000000000190000000000000018000000000000001900000000",
            INIT_08 => X"00000047000000000000003e0000000000000033000000000000001400000000",
            INIT_09 => X"00000051000000000000004e0000000000000049000000000000004400000000",
            INIT_0A => X"000000190000000000000019000000000000003f000000000000004b00000000",
            INIT_0B => X"0000001c000000000000001f000000000000001d000000000000001b00000000",
            INIT_0C => X"0000004a0000000000000043000000000000003b000000000000002b00000000",
            INIT_0D => X"0000005300000000000000540000000000000052000000000000004a00000000",
            INIT_0E => X"00000021000000000000001a0000000000000028000000000000004c00000000",
            INIT_0F => X"0000002d00000000000000200000000000000026000000000000002600000000",
            INIT_10 => X"0000004c00000000000000460000000000000044000000000000002d00000000",
            INIT_11 => X"00000047000000000000004d0000000000000053000000000000005700000000",
            INIT_12 => X"000000270000000000000035000000000000003f000000000000004900000000",
            INIT_13 => X"00000032000000000000001e0000000000000025000000000000002700000000",
            INIT_14 => X"0000004d0000000000000051000000000000004b000000000000004100000000",
            INIT_15 => X"0000004700000000000000370000000000000036000000000000003a00000000",
            INIT_16 => X"000000210000000000000023000000000000002b000000000000003f00000000",
            INIT_17 => X"0000003d00000000000000310000000000000029000000000000002300000000",
            INIT_18 => X"0000000900000000000000330000000000000044000000000000004100000000",
            INIT_19 => X"00000029000000000000002a000000000000002b000000000000001300000000",
            INIT_1A => X"0000002300000000000000210000000000000012000000000000002000000000",
            INIT_1B => X"00000030000000000000002a0000000000000032000000000000000b00000000",
            INIT_1C => X"0000001300000000000000240000000000000020000000000000002d00000000",
            INIT_1D => X"0000000a0000000000000014000000000000000f000000000000000500000000",
            INIT_1E => X"00000021000000000000001e000000000000001f000000000000000700000000",
            INIT_1F => X"0000001f00000000000000240000000000000027000000000000001e00000000",
            INIT_20 => X"0000000b000000000000001f000000000000002e000000000000001e00000000",
            INIT_21 => X"000000040000000000000005000000000000000e000000000000000c00000000",
            INIT_22 => X"0000001b00000000000000310000000000000011000000000000001300000000",
            INIT_23 => X"0000002f0000000000000025000000000000001f000000000000001e00000000",
            INIT_24 => X"00000022000000000000002c0000000000000037000000000000002d00000000",
            INIT_25 => X"0000001900000000000000070000000000000010000000000000001f00000000",
            INIT_26 => X"0000000f00000000000000230000000000000036000000000000000f00000000",
            INIT_27 => X"0000002c000000000000001d000000000000000c000000000000001b00000000",
            INIT_28 => X"0000000700000000000000140000000000000025000000000000001f00000000",
            INIT_29 => X"0000000100000000000000150000000000000006000000000000000400000000",
            INIT_2A => X"0000001700000000000000160000000000000026000000000000003300000000",
            INIT_2B => X"0000003b00000000000000280000000000000019000000000000000c00000000",
            INIT_2C => X"0000000d00000000000000090000000000000013000000000000002d00000000",
            INIT_2D => X"0000003500000000000000080000000000000013000000000000001000000000",
            INIT_2E => X"00000014000000000000001d0000000000000018000000000000002c00000000",
            INIT_2F => X"0000000a00000000000000170000000000000014000000000000000e00000000",
            INIT_30 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"000000340000000000000038000000000000001c000000000000001a00000000",
            INIT_32 => X"0000002d0000000000000028000000000000001e000000000000002800000000",
            INIT_33 => X"000000000000000000000006000000000000001f000000000000003000000000",
            INIT_34 => X"0000001800000000000000010000000000000000000000000000000000000000",
            INIT_35 => X"0000002c00000000000000320000000000000032000000000000001f00000000",
            INIT_36 => X"0000002c000000000000002b000000000000001f000000000000002a00000000",
            INIT_37 => X"0000001400000000000000110000000000000021000000000000003300000000",
            INIT_38 => X"0000001100000000000000180000000000000012000000000000001100000000",
            INIT_39 => X"0000002c0000000000000034000000000000002a000000000000003500000000",
            INIT_3A => X"000000350000000000000039000000000000002e000000000000002700000000",
            INIT_3B => X"0000003200000000000000310000000000000032000000000000003300000000",
            INIT_3C => X"000000c90000000000000025000000000000002c000000000000002e00000000",
            INIT_3D => X"000000c200000000000000be00000000000000c400000000000000bc00000000",
            INIT_3E => X"00000099000000000000009d00000000000000a800000000000000b900000000",
            INIT_3F => X"000000620000000000000071000000000000006a000000000000006100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ed00000000000000ea000000000000007f000000000000007c00000000",
            INIT_41 => X"000000ca00000000000000d200000000000000d100000000000000c300000000",
            INIT_42 => X"0000005f00000000000000a400000000000000b300000000000000c200000000",
            INIT_43 => X"0000009600000000000000890000000000000074000000000000005900000000",
            INIT_44 => X"000000da00000000000000cf0000000000000101000000000000007600000000",
            INIT_45 => X"000000d600000000000000e300000000000000e200000000000000dd00000000",
            INIT_46 => X"0000008d00000000000000aa00000000000000c000000000000000b700000000",
            INIT_47 => X"0000008d00000000000000840000000000000089000000000000009400000000",
            INIT_48 => X"000000e100000000000000e200000000000000e700000000000000db00000000",
            INIT_49 => X"000000ca00000000000000e200000000000000e900000000000000f300000000",
            INIT_4A => X"000000a800000000000000c100000000000000d000000000000000c500000000",
            INIT_4B => X"000000cb000000000000008d0000000000000074000000000000007800000000",
            INIT_4C => X"000000ea00000000000000e900000000000000ea00000000000000d700000000",
            INIT_4D => X"000000d000000000000000d500000000000000d700000000000000eb00000000",
            INIT_4E => X"0000006900000000000000c600000000000000c800000000000000b200000000",
            INIT_4F => X"000000f5000000000000003f000000000000008c000000000000008600000000",
            INIT_50 => X"000000db00000000000000ee00000000000000fc00000000000000e600000000",
            INIT_51 => X"000000aa00000000000000bf00000000000000e6000000000000012600000000",
            INIT_52 => X"000000710000000000000059000000000000008700000000000000c800000000",
            INIT_53 => X"0000012100000000000000ce0000000000000079000000000000007e00000000",
            INIT_54 => X"000000fd000000000000012800000000000000da000000000000010700000000",
            INIT_55 => X"000000d200000000000000e400000000000000cb00000000000000de00000000",
            INIT_56 => X"0000007a0000000000000067000000000000004d000000000000006e00000000",
            INIT_57 => X"000000f5000000000000011b00000000000000a800000000000000ab00000000",
            INIT_58 => X"0000011700000000000001180000000000000131000000000000010c00000000",
            INIT_59 => X"0000007a00000000000000f60000000000000120000000000000012800000000",
            INIT_5A => X"000000b70000000000000099000000000000008a000000000000004600000000",
            INIT_5B => X"0000010600000000000000f8000000000000011700000000000000c600000000",
            INIT_5C => X"000000e300000000000000e4000000000000012300000000000000f000000000",
            INIT_5D => X"0000002e000000000000003400000000000000a600000000000000e200000000",
            INIT_5E => X"000000bc00000000000000c800000000000000c000000000000000a200000000",
            INIT_5F => X"000000f800000000000000710000000000000109000000000000012400000000",
            INIT_60 => X"0000006300000000000000eb00000000000000c700000000000000ee00000000",
            INIT_61 => X"000000a800000000000000420000000000000051000000000000003e00000000",
            INIT_62 => X"0000011200000000000000c600000000000000df000000000000010000000000",
            INIT_63 => X"00000063000000000000005b000000000000004800000000000000c500000000",
            INIT_64 => X"0000003500000000000000430000000000000081000000000000009000000000",
            INIT_65 => X"0000010d00000000000000a30000000000000056000000000000003500000000",
            INIT_66 => X"000000c900000000000000d600000000000000d300000000000000c800000000",
            INIT_67 => X"0000008f000000000000008a000000000000007200000000000000aa00000000",
            INIT_68 => X"000000120000000000000011000000000000000f000000000000002d00000000",
            INIT_69 => X"000000c000000000000000b70000000000000085000000000000002a00000000",
            INIT_6A => X"000000d400000000000000d000000000000000da00000000000000d300000000",
            INIT_6B => X"0000006900000000000000a2000000000000009600000000000000b900000000",
            INIT_6C => X"00000044000000000000001c000000000000002b000000000000004100000000",
            INIT_6D => X"000000ac00000000000000cc0000000000000084000000000000004600000000",
            INIT_6E => X"0000009c00000000000000bd00000000000000b700000000000000e100000000",
            INIT_6F => X"00000098000000000000009200000000000000c700000000000000ba00000000",
            INIT_70 => X"0000008600000000000000880000000000000087000000000000007d00000000",
            INIT_71 => X"000000c900000000000000cf00000000000000ae000000000000009500000000",
            INIT_72 => X"000000c500000000000000d400000000000000c400000000000000c200000000",
            INIT_73 => X"000000a5000000000000009900000000000000b300000000000000b400000000",
            INIT_74 => X"0000008b00000000000000b200000000000000bf00000000000000b600000000",
            INIT_75 => X"0000006b00000000000000680000000000000048000000000000005c00000000",
            INIT_76 => X"0000004b00000000000000670000000000000068000000000000006d00000000",
            INIT_77 => X"0000002f0000000000000034000000000000002d000000000000005000000000",
            INIT_78 => X"0000006e000000000000003b0000000000000035000000000000002d00000000",
            INIT_79 => X"00000075000000000000006e0000000000000064000000000000007700000000",
            INIT_7A => X"0000005f00000000000000670000000000000071000000000000007500000000",
            INIT_7B => X"000000410000000000000040000000000000002f000000000000002c00000000",
            INIT_7C => X"0000006c0000000000000071000000000000003b000000000000004500000000",
            INIT_7D => X"0000007d00000000000000770000000000000077000000000000006b00000000",
            INIT_7E => X"00000042000000000000006e0000000000000073000000000000007b00000000",
            INIT_7F => X"0000004a00000000000000480000000000000043000000000000003d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "samplegold_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000730000000000000067000000000000005c000000000000004000000000",
            INIT_01 => X"000000830000000000000082000000000000007e000000000000007600000000",
            INIT_02 => X"0000005c0000000000000071000000000000006f000000000000007300000000",
            INIT_03 => X"00000047000000000000003f0000000000000043000000000000005a00000000",
            INIT_04 => X"0000007100000000000000730000000000000068000000000000005500000000",
            INIT_05 => X"000000610000000000000069000000000000007c000000000000008400000000",
            INIT_06 => X"00000066000000000000006a000000000000006d000000000000006500000000",
            INIT_07 => X"0000002900000000000000450000000000000045000000000000003b00000000",
            INIT_08 => X"0000007800000000000000770000000000000075000000000000005e00000000",
            INIT_09 => X"0000005e0000000000000074000000000000005e000000000000005c00000000",
            INIT_0A => X"000000300000000000000048000000000000005e000000000000004e00000000",
            INIT_0B => X"0000005f00000000000000280000000000000040000000000000003c00000000",
            INIT_0C => X"0000006700000000000000590000000000000071000000000000007800000000",
            INIT_0D => X"0000004300000000000000400000000000000047000000000000006e00000000",
            INIT_0E => X"000000350000000000000021000000000000002e000000000000005100000000",
            INIT_0F => X"0000007600000000000000480000000000000045000000000000003e00000000",
            INIT_10 => X"0000006b000000000000007a000000000000005b000000000000006700000000",
            INIT_11 => X"0000006100000000000000600000000000000065000000000000006700000000",
            INIT_12 => X"0000003e00000000000000370000000000000018000000000000003100000000",
            INIT_13 => X"00000061000000000000006e0000000000000043000000000000006000000000",
            INIT_14 => X"00000072000000000000008c0000000000000061000000000000006c00000000",
            INIT_15 => X"000000230000000000000063000000000000006f000000000000007200000000",
            INIT_16 => X"00000061000000000000004e000000000000003e000000000000000e00000000",
            INIT_17 => X"000000540000000000000070000000000000006a000000000000004d00000000",
            INIT_18 => X"0000005b000000000000005f0000000000000079000000000000005600000000",
            INIT_19 => X"000000190000000000000021000000000000001d000000000000003200000000",
            INIT_1A => X"00000051000000000000006c000000000000005c000000000000003900000000",
            INIT_1B => X"0000003e00000000000000040000000000000063000000000000006a00000000",
            INIT_1C => X"000000200000000000000069000000000000005c000000000000004c00000000",
            INIT_1D => X"0000003a00000000000000200000000000000029000000000000002200000000",
            INIT_1E => X"00000059000000000000005a0000000000000067000000000000007200000000",
            INIT_1F => X"00000033000000000000002c000000000000003d000000000000005200000000",
            INIT_20 => X"00000007000000000000000d0000000000000018000000000000003d00000000",
            INIT_21 => X"0000005f0000000000000038000000000000001e000000000000000700000000",
            INIT_22 => X"0000006c00000000000000540000000000000064000000000000006000000000",
            INIT_23 => X"0000004b00000000000000500000000000000051000000000000006500000000",
            INIT_24 => X"0000000000000000000000020000000000000008000000000000002000000000",
            INIT_25 => X"00000069000000000000003f0000000000000020000000000000001600000000",
            INIT_26 => X"0000006500000000000000440000000000000072000000000000005800000000",
            INIT_27 => X"0000004500000000000000650000000000000058000000000000004800000000",
            INIT_28 => X"0000003100000000000000300000000000000031000000000000003b00000000",
            INIT_29 => X"0000005b000000000000005e0000000000000046000000000000003300000000",
            INIT_2A => X"000000630000000000000050000000000000005a000000000000006700000000",
            INIT_2B => X"00000055000000000000005a0000000000000067000000000000006900000000",
            INIT_2C => X"00000058000000000000005a000000000000005a000000000000005600000000",
            INIT_2D => X"0000000700000000000000000000000000000039000000000000004100000000",
            INIT_2E => X"0000001300000000000000080000000000000010000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000030000000000000000000000000",
            INIT_30 => X"0000002100000000000000000000000000000004000000000000000c00000000",
            INIT_31 => X"0000000700000000000000060000000000000016000000000000000500000000",
            INIT_32 => X"000000030000000000000016000000000000000b000000000000000200000000",
            INIT_33 => X"0000000000000000000000000000000000000018000000000000003100000000",
            INIT_34 => X"000000200000000000000008000000000000000f000000000000000000000000",
            INIT_35 => X"0000000100000000000000000000000000000002000000000000000000000000",
            INIT_36 => X"0000000f00000000000000000000000000000017000000000000000a00000000",
            INIT_37 => X"0000000000000000000000170000000000000000000000000000003600000000",
            INIT_38 => X"0000000000000000000000290000000000000003000000000000000200000000",
            INIT_39 => X"0000000800000000000000090000000000000000000000000000000300000000",
            INIT_3A => X"0000000a00000000000000000000000000000011000000000000001200000000",
            INIT_3B => X"000000000000000000000006000000000000002d000000000000001200000000",
            INIT_3C => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000900000000000000080000000000000003000000000000000300000000",
            INIT_3E => X"000000040000000000000000000000000000001b000000000000000400000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000004800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000040000000000000000000000000000000d000000000000000000000000",
            INIT_41 => X"00000003000000000000001f0000000000000000000000000000000900000000",
            INIT_42 => X"0000004100000000000000120000000000000000000000000000002300000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000000000000000000010000000000000000d000000000000000000000000",
            INIT_45 => X"000000000000000000000029000000000000001f000000000000000000000000",
            INIT_46 => X"00000000000000000000002b0000000000000037000000000000000000000000",
            INIT_47 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_48 => X"0000001300000000000000000000000000000000000000000000001400000000",
            INIT_49 => X"0000000b00000000000000060000000000000000000000000000000e00000000",
            INIT_4A => X"000000000000000000000000000000000000002f000000000000004c00000000",
            INIT_4B => X"0000000a0000000000000000000000000000001a000000000000002900000000",
            INIT_4C => X"0000003100000000000000000000000000000000000000000000002300000000",
            INIT_4D => X"00000047000000000000000d0000000000000000000000000000000400000000",
            INIT_4E => X"0000006500000000000000000000000000000000000000000000002000000000",
            INIT_4F => X"0000007f00000000000000030000000000000000000000000000002000000000",
            INIT_50 => X"0000000000000000000000450000000000000000000000000000000000000000",
            INIT_51 => X"000000110000000000000011000000000000001e000000000000004200000000",
            INIT_52 => X"0000001f00000000000000800000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000007a000000000000000d000000000000000000000000",
            INIT_54 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000001000000000000001800000000",
            INIT_56 => X"0000000000000000000000140000000000000064000000000000000000000000",
            INIT_57 => X"0000000a00000000000000260000000000000030000000000000000000000000",
            INIT_58 => X"00000006000000000000001d0000000000000027000000000000000200000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_5A => X"0000000b00000000000000030000000000000000000000000000000000000000",
            INIT_5B => X"000000000000000000000010000000000000002e000000000000000000000000",
            INIT_5C => X"0000001600000000000000150000000000000028000000000000002e00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000230000000000000000000000000000001200000000",
            INIT_5F => X"0000002700000000000000000000000000000000000000000000001e00000000",
            INIT_60 => X"0000000000000000000000140000000000000015000000000000000f00000000",
            INIT_61 => X"00000007000000000000000d0000000000000000000000000000001500000000",
            INIT_62 => X"0000001200000000000000000000000000000016000000000000000000000000",
            INIT_63 => X"0000000d00000000000000070000000000000009000000000000000400000000",
            INIT_64 => X"0000001000000000000000000000000000000000000000000000000e00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "samplegold_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000001a000000000000002100000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_09 => X"0000000400000000000000100000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001400000000000000220000000000000044000000000000000000000000",
            INIT_0D => X"00000007000000000000000f0000000000000000000000000000002800000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001100000000000000090000000000000008000000000000001d00000000",
            INIT_12 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_17 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000000b0000000000000000000000000000000200000000",
            INIT_1F => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_20 => X"000000090000000000000000000000000000000a000000000000000500000000",
            INIT_21 => X"0000000000000000000000010000000000000000000000000000000f00000000",
            INIT_22 => X"0000000200000000000000040000000000000001000000000000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_24 => X"0000000000000000000000100000000000000008000000000000001400000000",
            INIT_25 => X"0000000000000000000000100000000000000000000000000000000600000000",
            INIT_26 => X"0000000000000000000000000000000000000006000000000000000500000000",
            INIT_27 => X"0000000800000000000000000000000000000002000000000000000a00000000",
            INIT_28 => X"00000008000000000000000c0000000000000008000000000000000000000000",
            INIT_29 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000200000000000000000000000000000001000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000004000000000000000c00000000",
            INIT_2C => X"00000000000000000000000a0000000000000012000000000000000400000000",
            INIT_2D => X"0000000300000000000000030000000000000002000000000000000c00000000",
            INIT_2E => X"00000000000000000000000b0000000000000004000000000000000200000000",
            INIT_2F => X"000000150000000000000000000000000000000e000000000000001b00000000",
            INIT_30 => X"000000000000000000000060000000000000000b000000000000000800000000",
            INIT_31 => X"0000002900000000000000000000000000000000000000000000000e00000000",
            INIT_32 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000900000000000000140000000000000000000000000000000000000000",
            INIT_34 => X"00000000000000000000002c0000000000000037000000000000001000000000",
            INIT_35 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_37 => X"00000008000000000000000a000000000000000c000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000047000000000000000000000000",
            INIT_39 => X"0000001100000000000000000000000000000000000000000000001b00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000018000000000000001900000000",
            INIT_3C => X"0000001d00000000000000000000000000000000000000000000003a00000000",
            INIT_3D => X"0000000c00000000000000080000000000000000000000000000001700000000",
            INIT_3E => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000003e00000000000000000000000000000000000000000000002e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000012000000000000004d0000000000000000000000000000000200000000",
            INIT_41 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_42 => X"0000004800000000000000270000000000000000000000000000000100000000",
            INIT_43 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_44 => X"00000010000000000000000d0000000000000011000000000000000000000000",
            INIT_45 => X"0000000700000000000000000000000000000000000000000000002500000000",
            INIT_46 => X"0000000000000000000000470000000000000017000000000000001500000000",
            INIT_47 => X"00000000000000000000000e000000000000000e000000000000000000000000",
            INIT_48 => X"0000000000000000000000020000000000000005000000000000000000000000",
            INIT_49 => X"0000001100000000000000020000000000000004000000000000000000000000",
            INIT_4A => X"0000000e000000000000001a0000000000000015000000000000002b00000000",
            INIT_4B => X"0000000000000000000000170000000000000000000000000000000900000000",
            INIT_4C => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_4D => X"0000000e00000000000000090000000000000000000000000000000000000000",
            INIT_4E => X"0000002400000000000000000000000000000018000000000000000e00000000",
            INIT_4F => X"0000000c0000000000000000000000000000000c000000000000000000000000",
            INIT_50 => X"0000000000000000000000060000000000000000000000000000001500000000",
            INIT_51 => X"0000000400000000000000000000000000000007000000000000000000000000",
            INIT_52 => X"00000000000000000000000d000000000000000d000000000000000000000000",
            INIT_53 => X"0000000400000000000000000000000000000000000000000000000b00000000",
            INIT_54 => X"0000000e00000000000000060000000000000000000000000000000400000000",
            INIT_55 => X"0000001200000000000000000000000000000000000000000000000e00000000",
            INIT_56 => X"00000042000000000000003d0000000000000040000000000000003d00000000",
            INIT_57 => X"0000003800000000000000420000000000000042000000000000004200000000",
            INIT_58 => X"000000240000000000000022000000000000001f000000000000003000000000",
            INIT_59 => X"0000003b00000000000000270000000000000027000000000000002300000000",
            INIT_5A => X"000000460000000000000043000000000000003d000000000000003c00000000",
            INIT_5B => X"0000003e0000000000000047000000000000004a000000000000004800000000",
            INIT_5C => X"0000002d0000000000000028000000000000001d000000000000002400000000",
            INIT_5D => X"0000003300000000000000350000000000000029000000000000002e00000000",
            INIT_5E => X"0000004600000000000000450000000000000042000000000000003f00000000",
            INIT_5F => X"0000003e00000000000000470000000000000046000000000000004800000000",
            INIT_60 => X"0000002d000000000000002e0000000000000035000000000000003900000000",
            INIT_61 => X"0000003d0000000000000035000000000000002d000000000000002d00000000",
            INIT_62 => X"0000004a00000000000000480000000000000046000000000000004200000000",
            INIT_63 => X"000000400000000000000043000000000000003f000000000000004300000000",
            INIT_64 => X"0000002c000000000000002b0000000000000029000000000000003500000000",
            INIT_65 => X"00000040000000000000003f0000000000000037000000000000002900000000",
            INIT_66 => X"0000003900000000000000340000000000000040000000000000004500000000",
            INIT_67 => X"0000002f000000000000003b0000000000000039000000000000003800000000",
            INIT_68 => X"0000001600000000000000290000000000000029000000000000002300000000",
            INIT_69 => X"0000003a000000000000003e000000000000003d000000000000003500000000",
            INIT_6A => X"000000250000000000000029000000000000002d000000000000003000000000",
            INIT_6B => X"0000001b000000000000001e000000000000002e000000000000002b00000000",
            INIT_6C => X"0000002a00000000000000240000000000000027000000000000002400000000",
            INIT_6D => X"0000003300000000000000340000000000000034000000000000003800000000",
            INIT_6E => X"0000002b000000000000002e0000000000000031000000000000002f00000000",
            INIT_6F => X"000000220000000000000019000000000000001c000000000000002800000000",
            INIT_70 => X"0000003600000000000000290000000000000030000000000000002500000000",
            INIT_71 => X"00000041000000000000003b000000000000002f000000000000003000000000",
            INIT_72 => X"00000030000000000000002c000000000000002e000000000000003500000000",
            INIT_73 => X"0000002900000000000000270000000000000016000000000000001d00000000",
            INIT_74 => X"0000002e00000000000000350000000000000030000000000000003d00000000",
            INIT_75 => X"0000002a000000000000003a0000000000000025000000000000002300000000",
            INIT_76 => X"0000001000000000000000160000000000000021000000000000002800000000",
            INIT_77 => X"0000003a00000000000000280000000000000022000000000000001400000000",
            INIT_78 => X"000000110000000000000028000000000000002d000000000000002c00000000",
            INIT_79 => X"00000039000000000000003e0000000000000032000000000000002600000000",
            INIT_7A => X"0000001d0000000000000022000000000000001a000000000000001900000000",
            INIT_7B => X"0000002f000000000000003f000000000000002a000000000000002200000000",
            INIT_7C => X"0000000600000000000000110000000000000025000000000000002800000000",
            INIT_7D => X"0000001500000000000000210000000000000020000000000000001300000000",
            INIT_7E => X"0000001f00000000000000230000000000000017000000000000000d00000000",
            INIT_7F => X"0000002900000000000000390000000000000039000000000000002900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "samplegold_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000038000000000000003a000000000000003c000000000000003b00000000",
            INIT_01 => X"000000060000000000000008000000000000000e000000000000002600000000",
            INIT_02 => X"0000002300000000000000200000000000000010000000000000000300000000",
            INIT_03 => X"0000002b0000000000000033000000000000003c000000000000003d00000000",
            INIT_04 => X"0000003c0000000000000034000000000000002e000000000000003800000000",
            INIT_05 => X"000000130000000000000018000000000000001d000000000000002c00000000",
            INIT_06 => X"00000036000000000000001d0000000000000016000000000000001600000000",
            INIT_07 => X"0000002c000000000000002e000000000000003c000000000000002f00000000",
            INIT_08 => X"00000036000000000000003d0000000000000037000000000000003000000000",
            INIT_09 => X"0000003600000000000000380000000000000035000000000000003600000000",
            INIT_0A => X"0000003f000000000000003a000000000000002c000000000000003300000000",
            INIT_0B => X"00000040000000000000003b000000000000003f000000000000003e00000000",
            INIT_0C => X"0000003700000000000000370000000000000039000000000000003c00000000",
            INIT_0D => X"00000038000000000000003c000000000000003b000000000000003a00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000011000000000000000d0000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000001000000000000000500000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000017000000000000000e0000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000013000000000000001f00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000200000000000000019000000000000000b000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000007000000000000001d00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000002b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "samplegold_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000b00000000000000050000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000d0000000000000000000000000000000100000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000002900000000000000360000000000000004000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000100000000000000060000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000a00000000000000000000000000000000000000000000000800000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_17 => X"0000000000000000000000230000000000000049000000000000003500000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000060000000000000002000000000000000000000000",
            INIT_1B => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_1C => X"000000080000000000000009000000000000001c000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000007000000000000001a000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000017000000000000001500000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_28 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"00000000000000000000002c000000000000003b000000000000001f00000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"000000300000000000000029000000000000000a000000000000000000000000",
            INIT_2E => X"000000000000000000000025000000000000002b000000000000003000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000001d00000000000000170000000000000000000000000000000000000000",
            INIT_32 => X"0000001c00000000000000340000000000000034000000000000002a00000000",
            INIT_33 => X"00000000000000000000000c0000000000000002000000000000000000000000",
            INIT_34 => X"0000000000000000000000060000000000000016000000000000000e00000000",
            INIT_35 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000c00000000000000040000000000000007000000000000000100000000",
            INIT_37 => X"00000019000000000000001a0000000000000024000000000000000c00000000",
            INIT_38 => X"0000001b0000000000000016000000000000001c000000000000001a00000000",
            INIT_39 => X"0000001300000000000000140000000000000015000000000000000c00000000",
            INIT_3A => X"0000001300000000000000060000000000000016000000000000001500000000",
            INIT_3B => X"0000001e000000000000001e0000000000000018000000000000001700000000",
            INIT_3C => X"00000013000000000000001c0000000000000018000000000000001b00000000",
            INIT_3D => X"0000001300000000000000100000000000000019000000000000001200000000",
            INIT_3E => X"0000002000000000000000100000000000000010000000000000000e00000000",
            INIT_3F => X"0000001c000000000000001d000000000000001c000000000000001c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c0000000000000017000000000000001f000000000000001800000000",
            INIT_41 => X"000000110000000000000012000000000000000e000000000000001e00000000",
            INIT_42 => X"0000001a0000000000000022000000000000000a000000000000001100000000",
            INIT_43 => X"00000014000000000000001a0000000000000019000000000000001e00000000",
            INIT_44 => X"000000180000000000000016000000000000001b000000000000001700000000",
            INIT_45 => X"0000001100000000000000160000000000000014000000000000000a00000000",
            INIT_46 => X"0000001f000000000000001a000000000000001b000000000000001600000000",
            INIT_47 => X"000000150000000000000013000000000000001c000000000000001c00000000",
            INIT_48 => X"000000010000000000000012000000000000001b000000000000000f00000000",
            INIT_49 => X"0000002c00000000000000130000000000000013000000000000001700000000",
            INIT_4A => X"0000001b0000000000000018000000000000001f000000000000001b00000000",
            INIT_4B => X"0000000800000000000000090000000000000007000000000000002200000000",
            INIT_4C => X"0000001d0000000000000002000000000000000c000000000000001d00000000",
            INIT_4D => X"0000001a00000000000000330000000000000016000000000000001400000000",
            INIT_4E => X"00000017000000000000001b0000000000000012000000000000001200000000",
            INIT_4F => X"00000015000000000000001e000000000000000c000000000000000900000000",
            INIT_50 => X"00000019000000000000001a0000000000000004000000000000000000000000",
            INIT_51 => X"0000000b000000000000002d000000000000000f000000000000001500000000",
            INIT_52 => X"0000000e000000000000000c000000000000001d000000000000001400000000",
            INIT_53 => X"00000000000000000000000e000000000000000c000000000000001200000000",
            INIT_54 => X"000000070000000000000020000000000000001c000000000000000000000000",
            INIT_55 => X"00000003000000000000000b0000000000000028000000000000000600000000",
            INIT_56 => X"0000001000000000000000000000000000000017000000000000001d00000000",
            INIT_57 => X"0000000b00000000000000000000000000000006000000000000000c00000000",
            INIT_58 => X"0000000900000000000000000000000000000025000000000000002400000000",
            INIT_59 => X"0000002f0000000000000000000000000000000a000000000000002600000000",
            INIT_5A => X"00000002000000000000001d0000000000000000000000000000001300000000",
            INIT_5B => X"00000023000000000000000f000000000000000e000000000000000b00000000",
            INIT_5C => X"0000001a00000000000000030000000000000000000000000000002f00000000",
            INIT_5D => X"0000001700000000000000230000000000000000000000000000000a00000000",
            INIT_5E => X"0000000a0000000000000000000000000000001b000000000000000d00000000",
            INIT_5F => X"0000002e000000000000001a0000000000000016000000000000001100000000",
            INIT_60 => X"00000015000000000000000e0000000000000006000000000000000000000000",
            INIT_61 => X"00000013000000000000000e000000000000000f000000000000000300000000",
            INIT_62 => X"000000140000000000000014000000000000000e000000000000000f00000000",
            INIT_63 => X"000000150000000000000019000000000000001f000000000000001e00000000",
            INIT_64 => X"00000019000000000000000d000000000000000f000000000000000b00000000",
            INIT_65 => X"000000030000000000000010000000000000000d000000000000000000000000",
            INIT_66 => X"0000001e00000000000000130000000000000013000000000000000a00000000",
            INIT_67 => X"00000008000000000000001e0000000000000016000000000000002200000000",
            INIT_68 => X"0000000700000000000000110000000000000001000000000000001100000000",
            INIT_69 => X"0000000d00000000000000020000000000000017000000000000001400000000",
            INIT_6A => X"000000120000000000000018000000000000000f000000000000000a00000000",
            INIT_6B => X"00000012000000000000000d0000000000000013000000000000001600000000",
            INIT_6C => X"00000010000000000000000b000000000000000d000000000000000600000000",
            INIT_6D => X"0000000b000000000000000e000000000000000b000000000000000e00000000",
            INIT_6E => X"0000000d000000000000000c0000000000000014000000000000001200000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "samplegold_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000f00000000000000050000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000002300000000000000100000000000000000000000000000000000000000",
            INIT_28 => X"000000380000000000000032000000000000003a000000000000003100000000",
            INIT_29 => X"0000001f0000000000000015000000000000002d000000000000003500000000",
            INIT_2A => X"0000002400000000000000190000000000000019000000000000002000000000",
            INIT_2B => X"000000320000000000000028000000000000002a000000000000001600000000",
            INIT_2C => X"0000003900000000000000380000000000000038000000000000003200000000",
            INIT_2D => X"000000250000000000000018000000000000001f000000000000003e00000000",
            INIT_2E => X"0000002000000000000000220000000000000029000000000000002900000000",
            INIT_2F => X"000000380000000000000031000000000000002a000000000000001a00000000",
            INIT_30 => X"000000430000000000000039000000000000003a000000000000003600000000",
            INIT_31 => X"0000002100000000000000220000000000000010000000000000003300000000",
            INIT_32 => X"000000130000000000000025000000000000002c000000000000002d00000000",
            INIT_33 => X"0000003800000000000000380000000000000032000000000000002600000000",
            INIT_34 => X"00000041000000000000003b000000000000003e000000000000004000000000",
            INIT_35 => X"000000280000000000000021000000000000002a000000000000003700000000",
            INIT_36 => X"0000002a00000000000000260000000000000028000000000000002b00000000",
            INIT_37 => X"0000003000000000000000390000000000000030000000000000003000000000",
            INIT_38 => X"00000044000000000000002b0000000000000024000000000000002a00000000",
            INIT_39 => X"0000002800000000000000290000000000000016000000000000003500000000",
            INIT_3A => X"000000290000000000000019000000000000003e000000000000002800000000",
            INIT_3B => X"00000007000000000000001a000000000000002f000000000000002c00000000",
            INIT_3C => X"00000024000000000000002a000000000000001f000000000000002600000000",
            INIT_3D => X"0000002900000000000000250000000000000025000000000000000f00000000",
            INIT_3E => X"0000001e000000000000001c0000000000000031000000000000003400000000",
            INIT_3F => X"000000000000000000000015000000000000001a000000000000001e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000000000090000000000000008000000000000000400000000",
            INIT_41 => X"000000190000000000000025000000000000001f000000000000001a00000000",
            INIT_42 => X"00000019000000000000001d000000000000001b000000000000003800000000",
            INIT_43 => X"0000000900000000000000140000000000000020000000000000001300000000",
            INIT_44 => X"0000001a000000000000000a0000000000000000000000000000000600000000",
            INIT_45 => X"0000002b000000000000002a0000000000000012000000000000001700000000",
            INIT_46 => X"0000002100000000000000210000000000000018000000000000001500000000",
            INIT_47 => X"00000029000000000000002b000000000000002f000000000000002500000000",
            INIT_48 => X"0000001c00000000000000240000000000000010000000000000001700000000",
            INIT_49 => X"0000000f00000000000000300000000000000029000000000000000000000000",
            INIT_4A => X"0000001e00000000000000270000000000000038000000000000000000000000",
            INIT_4B => X"0000001100000000000000190000000000000014000000000000002f00000000",
            INIT_4C => X"00000000000000000000001e0000000000000028000000000000001100000000",
            INIT_4D => X"0000000000000000000000130000000000000032000000000000002d00000000",
            INIT_4E => X"0000003d00000000000000340000000000000029000000000000001600000000",
            INIT_4F => X"0000001e00000000000000190000000000000016000000000000002700000000",
            INIT_50 => X"0000003200000000000000000000000000000032000000000000002300000000",
            INIT_51 => X"000000110000000000000009000000000000001b000000000000002c00000000",
            INIT_52 => X"0000001000000000000000130000000000000021000000000000001c00000000",
            INIT_53 => X"0000002600000000000000170000000000000008000000000000000f00000000",
            INIT_54 => X"0000002b000000000000003b0000000000000017000000000000003500000000",
            INIT_55 => X"000000290000000000000022000000000000002d000000000000002300000000",
            INIT_56 => X"0000000000000000000000060000000000000018000000000000003000000000",
            INIT_57 => X"0000001e000000000000001c0000000000000003000000000000000000000000",
            INIT_58 => X"0000002a000000000000003e0000000000000031000000000000002500000000",
            INIT_59 => X"0000003600000000000000250000000000000024000000000000002d00000000",
            INIT_5A => X"00000016000000000000001b0000000000000021000000000000002a00000000",
            INIT_5B => X"0000001900000000000000200000000000000013000000000000001800000000",
            INIT_5C => X"0000002f00000000000000300000000000000033000000000000002d00000000",
            INIT_5D => X"000000360000000000000036000000000000002e000000000000002300000000",
            INIT_5E => X"000000310000000000000033000000000000002f000000000000003100000000",
            INIT_5F => X"00000045000000000000002a0000000000000026000000000000002a00000000",
            INIT_60 => X"0000003000000000000000300000000000000032000000000000003400000000",
            INIT_61 => X"0000002500000000000000330000000000000038000000000000003200000000",
            INIT_62 => X"0000002000000000000000190000000000000019000000000000001e00000000",
            INIT_63 => X"0000002f000000000000003a0000000000000022000000000000001e00000000",
            INIT_64 => X"0000003c00000000000000340000000000000032000000000000004000000000",
            INIT_65 => X"00000024000000000000002d0000000000000035000000000000003b00000000",
            INIT_66 => X"0000001a000000000000001c0000000000000023000000000000001700000000",
            INIT_67 => X"0000003900000000000000280000000000000026000000000000002600000000",
            INIT_68 => X"00000037000000000000003f0000000000000036000000000000003b00000000",
            INIT_69 => X"0000002a0000000000000032000000000000003f000000000000004000000000",
            INIT_6A => X"000000210000000000000023000000000000001a000000000000002a00000000",
            INIT_6B => X"0000003b00000000000000360000000000000027000000000000003b00000000",
            INIT_6C => X"0000003b000000000000003b0000000000000042000000000000003b00000000",
            INIT_6D => X"0000002c00000000000000370000000000000038000000000000003500000000",
            INIT_6E => X"0000003100000000000000200000000000000020000000000000001a00000000",
            INIT_6F => X"0000003f00000000000000370000000000000035000000000000002f00000000",
            INIT_70 => X"0000002d00000000000000240000000000000027000000000000003100000000",
            INIT_71 => X"0000001c000000000000001e0000000000000039000000000000002e00000000",
            INIT_72 => X"00000028000000000000003a000000000000001b000000000000001d00000000",
            INIT_73 => X"0000003400000000000000380000000000000035000000000000003000000000",
            INIT_74 => X"0000001a000000000000001c000000000000001f000000000000001800000000",
            INIT_75 => X"0000001e00000000000000140000000000000020000000000000001f00000000",
            INIT_76 => X"0000002600000000000000340000000000000016000000000000001b00000000",
            INIT_77 => X"000000390000000000000021000000000000003f000000000000002400000000",
            INIT_78 => X"0000001e000000000000001a0000000000000018000000000000001700000000",
            INIT_79 => X"00000016000000000000001b0000000000000017000000000000001d00000000",
            INIT_7A => X"0000003300000000000000270000000000000025000000000000001b00000000",
            INIT_7B => X"0000001d000000000000003d0000000000000034000000000000002800000000",
            INIT_7C => X"0000001a000000000000001b000000000000001b000000000000002200000000",
            INIT_7D => X"0000002c00000000000000200000000000000016000000000000001e00000000",
            INIT_7E => X"0000000000000000000000370000000000000027000000000000001e00000000",
            INIT_7F => X"0000001b000000000000001b000000000000002b000000000000003600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "samplegold_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f00000000000000120000000000000011000000000000001b00000000",
            INIT_01 => X"00000028000000000000001e0000000000000016000000000000001300000000",
            INIT_02 => X"0000001c0000000000000013000000000000000e000000000000001900000000",
            INIT_03 => X"00000020000000000000001a000000000000001a000000000000002c00000000",
            INIT_04 => X"00000017000000000000001b000000000000000e000000000000001e00000000",
            INIT_05 => X"00000010000000000000002c0000000000000023000000000000000000000000",
            INIT_06 => X"0000001400000000000000110000000000000002000000000000001b00000000",
            INIT_07 => X"0000000b00000000000000160000000000000025000000000000000600000000",
            INIT_08 => X"00000003000000000000001f000000000000001b000000000000001100000000",
            INIT_09 => X"000000350000000000000021000000000000001d000000000000003100000000",
            INIT_0A => X"0000000400000000000000250000000000000031000000000000002f00000000",
            INIT_0B => X"0000000100000000000000030000000000000011000000000000001400000000",
            INIT_0C => X"0000003000000000000000130000000000000024000000000000001800000000",
            INIT_0D => X"0000003d000000000000002f0000000000000028000000000000002300000000",
            INIT_0E => X"00000021000000000000002d0000000000000020000000000000001300000000",
            INIT_0F => X"0000000d00000000000000100000000000000011000000000000001500000000",
            INIT_10 => X"0000002d00000000000000180000000000000007000000000000001e00000000",
            INIT_11 => X"0000001f0000000000000025000000000000002b000000000000002a00000000",
            INIT_12 => X"00000029000000000000002b0000000000000027000000000000001f00000000",
            INIT_13 => X"0000002600000000000000290000000000000024000000000000002c00000000",
            INIT_14 => X"0000002e00000000000000210000000000000028000000000000001300000000",
            INIT_15 => X"000000270000000000000021000000000000002e000000000000002f00000000",
            INIT_16 => X"00000028000000000000002c0000000000000025000000000000002700000000",
            INIT_17 => X"000000300000000000000023000000000000002c000000000000002800000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000004100000000000000180000000000000000000000000000000000000000",
            INIT_2D => X"00000000000000000000002c0000000000000028000000000000004200000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000001000000000000001e0000000000000031000000000000003f00000000",
            INIT_31 => X"0000000000000000000000040000000000000045000000000000003200000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000140000000000000009000000000000000c000000000000000000000000",
            INIT_34 => X"0000005a000000000000001b0000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000002b000000000000005f00000000",
            INIT_36 => X"0000000d00000000000000080000000000000000000000000000000000000000",
            INIT_37 => X"000000320000000000000000000000000000000d000000000000002400000000",
            INIT_38 => X"0000003600000000000000790000000000000067000000000000006900000000",
            INIT_39 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_3A => X"0000001700000000000000150000000000000033000000000000000000000000",
            INIT_3B => X"0000005a0000000000000051000000000000001d000000000000000200000000",
            INIT_3C => X"0000002900000000000000380000000000000055000000000000007500000000",
            INIT_3D => X"0000004700000000000000000000000000000050000000000000004200000000",
            INIT_3E => X"000000000000000000000005000000000000001e000000000000004500000000",
            INIT_3F => X"0000004700000000000000790000000000000052000000000000001100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005600000000000000680000000000000039000000000000003500000000",
            INIT_41 => X"0000001c000000000000001f0000000000000006000000000000004500000000",
            INIT_42 => X"0000002c00000000000000110000000000000000000000000000001600000000",
            INIT_43 => X"00000000000000000000000e0000000000000052000000000000005700000000",
            INIT_44 => X"0000000000000000000000420000000000000040000000000000001b00000000",
            INIT_45 => X"00000014000000000000001f0000000000000014000000000000000000000000",
            INIT_46 => X"0000005600000000000000360000000000000012000000000000000000000000",
            INIT_47 => X"0000001500000000000000100000000000000002000000000000004700000000",
            INIT_48 => X"000000000000000000000000000000000000002d000000000000002b00000000",
            INIT_49 => X"0000004400000000000000350000000000000032000000000000001300000000",
            INIT_4A => X"00000042000000000000006a0000000000000066000000000000005c00000000",
            INIT_4B => X"0000000d000000000000000b000000000000001f000000000000001f00000000",
            INIT_4C => X"0000000b00000000000000000000000000000000000000000000000300000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000008000000000000002600000000",
            INIT_50 => X"000000060000000000000005000000000000001d000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000100000000000000030000000000000000000000000000000800000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000110000000000000000000000000000000300000000",
            INIT_57 => X"0000000000000000000000040000000000000029000000000000000000000000",
            INIT_58 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000800000000000000070000000000000008000000000000000500000000",
            INIT_5A => X"0000000100000000000000000000000000000009000000000000001400000000",
            INIT_5B => X"0000000c00000000000000050000000000000000000000000000002200000000",
            INIT_5C => X"0000000e000000000000000d0000000000000009000000000000000b00000000",
            INIT_5D => X"0000000f000000000000000e000000000000000f000000000000000c00000000",
            INIT_5E => X"00000003000000000000000e000000000000000f000000000000000000000000",
            INIT_5F => X"0000000b000000000000000d000000000000000e000000000000000000000000",
            INIT_60 => X"0000000a00000000000000100000000000000011000000000000000800000000",
            INIT_61 => X"0000000000000000000000030000000000000021000000000000000c00000000",
            INIT_62 => X"0000000400000000000000000000000000000000000000000000002500000000",
            INIT_63 => X"00000006000000000000000b000000000000000b000000000000000e00000000",
            INIT_64 => X"0000000500000000000000370000000000000030000000000000001700000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000c00000000000000040000000000000000000000000000001d00000000",
            INIT_67 => X"0000001c00000000000000140000000000000001000000000000000a00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000500000000000000000000000000000039000000000000006100000000",
            INIT_6A => X"00000008000000000000000b0000000000000000000000000000000400000000",
            INIT_6B => X"000000110000000000000000000000000000000b000000000000002200000000",
            INIT_6C => X"0000006a00000000000000730000000000000029000000000000000000000000",
            INIT_6D => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"00000000000000000000001a0000000000000008000000000000003300000000",
            INIT_6F => X"0000005400000000000000040000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_71 => X"00000023000000000000004e000000000000002c000000000000000000000000",
            INIT_72 => X"0000000e00000000000000000000000000000057000000000000002800000000",
            INIT_73 => X"000000040000000000000060000000000000001d000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000004300000000000000000000000000000000000000000000001e00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"000000000000000000000000000000000000007b000000000000002e00000000",
            INIT_78 => X"0000000000000000000000340000000000000001000000000000000000000000",
            INIT_79 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_7A => X"0000002f00000000000000180000000000000000000000000000000000000000",
            INIT_7B => X"0000000100000000000000000000000000000000000000000000005100000000",
            INIT_7C => X"0000000000000000000000000000000000000047000000000000000000000000",
            INIT_7D => X"000000060000000000000008000000000000000b000000000000000000000000",
            INIT_7E => X"00000040000000000000002a000000000000004a000000000000000000000000",
            INIT_7F => X"0000000000000000000000250000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "samplegold_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b0000000000000000000000000000000e000000000000000700000000",
            INIT_01 => X"0000000000000000000000000000000000000009000000000000000a00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_04 => X"00000008000000000000000a0000000000000000000000000000000000000000",
            INIT_05 => X"0000000c00000000000000030000000000000009000000000000000000000000",
            INIT_06 => X"0000000000000000000000010000000000000007000000000000000a00000000",
            INIT_07 => X"0000000400000000000000000000000000000000000000000000002300000000",
            INIT_08 => X"000000d000000000000000bf0000000000000010000000000000000600000000",
            INIT_09 => X"000000c700000000000000da00000000000000e200000000000000dc00000000",
            INIT_0A => X"0000007b000000000000009b00000000000000b200000000000000bd00000000",
            INIT_0B => X"0000001e000000000000001a0000000000000057000000000000007600000000",
            INIT_0C => X"000000bb00000000000000c200000000000000d3000000000000004800000000",
            INIT_0D => X"00000092000000000000009800000000000000aa00000000000000b900000000",
            INIT_0E => X"0000005e0000000000000071000000000000007e000000000000008b00000000",
            INIT_0F => X"0000005300000000000000170000000000000008000000000000003500000000",
            INIT_10 => X"00000088000000000000008e0000000000000091000000000000009100000000",
            INIT_11 => X"0000007600000000000000770000000000000078000000000000008100000000",
            INIT_12 => X"000000000000000000000028000000000000006c000000000000006f00000000",
            INIT_13 => X"0000006e00000000000000570000000000000033000000000000001300000000",
            INIT_14 => X"00000073000000000000006f000000000000006f000000000000006e00000000",
            INIT_15 => X"0000006e00000000000000720000000000000073000000000000007500000000",
            INIT_16 => X"0000003a00000000000000000000000000000009000000000000005c00000000",
            INIT_17 => X"0000006f00000000000000640000000000000062000000000000005b00000000",
            INIT_18 => X"0000006900000000000000710000000000000070000000000000007100000000",
            INIT_19 => X"000000320000000000000052000000000000005d000000000000005c00000000",
            INIT_1A => X"0000005e00000000000000420000000000000000000000000000000000000000",
            INIT_1B => X"00000070000000000000006f000000000000006d000000000000005c00000000",
            INIT_1C => X"0000000000000000000000410000000000000064000000000000007000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000051000000000000002f0000000000000002000000000000000000000000",
            INIT_1F => X"00000062000000000000006d0000000000000070000000000000007100000000",
            INIT_20 => X"0000000000000000000000000000000000000007000000000000003600000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000006f000000000000002a0000000000000000000000000000000000000000",
            INIT_23 => X"000000060000000000000025000000000000004d000000000000006f00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000058000000000000006d0000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000130000000000000060000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000bd00000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000b300000000000000ba00000000000000bb00000000000000bc00000000",
            INIT_42 => X"0000007e000000000000008b0000000000000094000000000000009c00000000",
            INIT_43 => X"0000005800000000000000560000000000000068000000000000007f00000000",
            INIT_44 => X"000000a900000000000000a80000000000000049000000000000002000000000",
            INIT_45 => X"00000072000000000000007c000000000000008800000000000000a300000000",
            INIT_46 => X"0000005c0000000000000062000000000000006a000000000000007000000000",
            INIT_47 => X"00000029000000000000002d0000000000000069000000000000005600000000",
            INIT_48 => X"00000066000000000000007c000000000000008a000000000000005200000000",
            INIT_49 => X"000000630000000000000060000000000000005d000000000000006300000000",
            INIT_4A => X"0000007d00000000000000600000000000000062000000000000006200000000",
            INIT_4B => X"0000006900000000000000580000000000000046000000000000006100000000",
            INIT_4C => X"0000005d000000000000005d0000000000000054000000000000004f00000000",
            INIT_4D => X"0000007a000000000000006c0000000000000067000000000000005f00000000",
            INIT_4E => X"0000001c000000000000007a000000000000007c000000000000007900000000",
            INIT_4F => X"0000005500000000000000530000000000000067000000000000006100000000",
            INIT_50 => X"000000630000000000000062000000000000005f000000000000005a00000000",
            INIT_51 => X"0000009a000000000000008f000000000000008b000000000000007500000000",
            INIT_52 => X"000000610000000000000050000000000000007500000000000000c300000000",
            INIT_53 => X"0000005f000000000000005b000000000000004d000000000000005300000000",
            INIT_54 => X"00000078000000000000005e000000000000005f000000000000006100000000",
            INIT_55 => X"0000010a0000000000000125000000000000010a00000000000000cd00000000",
            INIT_56 => X"0000006e000000000000001c00000000000000e6000000000000010900000000",
            INIT_57 => X"0000006500000000000000650000000000000060000000000000004b00000000",
            INIT_58 => X"000000b000000000000000b20000000000000077000000000000005400000000",
            INIT_59 => X"0000015400000000000000260000000000000039000000000000006400000000",
            INIT_5A => X"000000360000000000000033000000000000004f000000000000014b00000000",
            INIT_5B => X"0000008b00000000000000550000000000000066000000000000006400000000",
            INIT_5C => X"000000560000000000000084000000000000005d000000000000008300000000",
            INIT_5D => X"0000017e000000000000019b000000000000013d000000000000009b00000000",
            INIT_5E => X"000000640000000000000056000000000000001b000000000000007200000000",
            INIT_5F => X"0000008a00000000000000600000000000000082000000000000005a00000000",
            INIT_60 => X"000001b00000000000000148000000000000003c000000000000003900000000",
            INIT_61 => X"0000005000000000000000dd00000000000001b900000000000001a200000000",
            INIT_62 => X"000000a7000000000000004f000000000000010b000000000000008400000000",
            INIT_63 => X"0000000d0000000000000048000000000000004b00000000000000fe00000000",
            INIT_64 => X"00000186000000000000016d0000000000000163000000000000005c00000000",
            INIT_65 => X"0000012f00000000000001240000000000000136000000000000012400000000",
            INIT_66 => X"000000cb00000000000000fe000000000000004f000000000000012300000000",
            INIT_67 => X"00000085000000000000000a000000000000000c000000000000006100000000",
            INIT_68 => X"000000650000000000000088000000000000017d000000000000015a00000000",
            INIT_69 => X"000000ad00000000000001160000000000000153000000000000009d00000000",
            INIT_6A => X"0000006c00000000000000a00000000000000056000000000000005100000000",
            INIT_6B => X"0000017500000000000000bb0000000000000068000000000000000700000000",
            INIT_6C => X"00000048000000000000003a0000000000000039000000000000014c00000000",
            INIT_6D => X"0000002f000000000000000e00000000000000e400000000000000d200000000",
            INIT_6E => X"0000004f000000000000006d000000000000009f000000000000005b00000000",
            INIT_6F => X"00000127000000000000015e000000000000012100000000000000ce00000000",
            INIT_70 => X"0000007d000000000000003e0000000000000080000000000000004700000000",
            INIT_71 => X"0000005500000000000000380000000000000009000000000000007400000000",
            INIT_72 => X"0000009b00000000000000710000000000000058000000000000008900000000",
            INIT_73 => X"00000049000000000000007d00000000000000b500000000000000ad00000000",
            INIT_74 => X"00000000000000000000001c0000000000000035000000000000007700000000",
            INIT_75 => X"0000002f000000000000004a0000000000000049000000000000000000000000",
            INIT_76 => X"00000021000000000000001d0000000000000019000000000000003700000000",
            INIT_77 => X"00000053000000000000001f000000000000000e000000000000001a00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_79 => X"000000d900000000000000d900000000000000ca00000000000000be00000000",
            INIT_7A => X"000000ab00000000000000b800000000000000bd00000000000000d200000000",
            INIT_7B => X"000000610000000000000072000000000000008b000000000000009000000000",
            INIT_7C => X"000000c8000000000000004f000000000000002b000000000000003900000000",
            INIT_7D => X"000000a600000000000000b100000000000000b900000000000000be00000000",
            INIT_7E => X"0000007b00000000000000880000000000000091000000000000009500000000",
            INIT_7F => X"0000001900000000000000470000000000000059000000000000007100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "samplegold_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009300000000000000990000000000000058000000000000001c00000000",
            INIT_01 => X"00000076000000000000007d0000000000000086000000000000008f00000000",
            INIT_02 => X"0000006900000000000000710000000000000075000000000000007800000000",
            INIT_03 => X"00000046000000000000001c000000000000002b000000000000005000000000",
            INIT_04 => X"0000006e000000000000006d000000000000006a000000000000006400000000",
            INIT_05 => X"0000007100000000000000750000000000000070000000000000007000000000",
            INIT_06 => X"0000003600000000000000630000000000000073000000000000007600000000",
            INIT_07 => X"000000660000000000000065000000000000004d000000000000000500000000",
            INIT_08 => X"000000730000000000000071000000000000006e000000000000006500000000",
            INIT_09 => X"00000067000000000000006f0000000000000079000000000000007200000000",
            INIT_0A => X"000000110000000000000018000000000000004c000000000000004d00000000",
            INIT_0B => X"0000006c000000000000005d0000000000000061000000000000005200000000",
            INIT_0C => X"0000006000000000000000720000000000000072000000000000007000000000",
            INIT_0D => X"0000005f00000000000000590000000000000055000000000000004800000000",
            INIT_0E => X"00000023000000000000001d000000000000001f000000000000005b00000000",
            INIT_0F => X"0000007200000000000000700000000000000053000000000000004400000000",
            INIT_10 => X"0000003600000000000000560000000000000060000000000000007300000000",
            INIT_11 => X"00000000000000000000001d0000000000000024000000000000003a00000000",
            INIT_12 => X"0000002e0000000000000000000000000000004f000000000000003400000000",
            INIT_13 => X"0000005600000000000000720000000000000071000000000000003a00000000",
            INIT_14 => X"000000110000000000000018000000000000002d000000000000004000000000",
            INIT_15 => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000090000000000000000000000000000001a000000000000008200000000",
            INIT_17 => X"00000022000000000000002e0000000000000055000000000000007100000000",
            INIT_18 => X"0000002c00000000000000000000000000000000000000000000002000000000",
            INIT_19 => X"0000004900000000000000580000000000000050000000000000004900000000",
            INIT_1A => X"0000005700000000000000220000000000000000000000000000000600000000",
            INIT_1B => X"0000000c00000000000000000000000000000026000000000000003600000000",
            INIT_1C => X"0000003b00000000000000370000000000000000000000000000000000000000",
            INIT_1D => X"00000014000000000000002f0000000000000055000000000000006600000000",
            INIT_1E => X"0000004700000000000000420000000000000047000000000000002900000000",
            INIT_1F => X"0000000000000000000000000000000000000005000000000000003700000000",
            INIT_20 => X"0000002100000000000000600000000000000030000000000000000000000000",
            INIT_21 => X"00000045000000000000003e000000000000002c000000000000000200000000",
            INIT_22 => X"0000001c00000000000000000000000000000039000000000000003900000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_24 => X"0000000500000000000000000000000000000060000000000000003300000000",
            INIT_25 => X"0000000900000000000000380000000000000024000000000000000000000000",
            INIT_26 => X"00000000000000000000000d0000000000000004000000000000002600000000",
            INIT_27 => X"0000003200000000000000040000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000070000000000000000000000000000005100000000",
            INIT_29 => X"0000002000000000000000020000000000000026000000000000001a00000000",
            INIT_2A => X"0000000a000000000000000f000000000000001c000000000000001300000000",
            INIT_2B => X"000000460000000000000040000000000000003c000000000000003200000000",
            INIT_2C => X"00000000000000000000000a0000000000000018000000000000000000000000",
            INIT_2D => X"0000000300000000000000270000000000000000000000000000000400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000001000000000000001400000000",
            INIT_31 => X"0000000600000000000000140000000000000007000000000000000000000000",
            INIT_32 => X"0000000800000000000000150000000000000019000000000000001100000000",
            INIT_33 => X"00000014000000000000001f0000000000000006000000000000001c00000000",
            INIT_34 => X"0000000d00000000000000000000000000000019000000000000000b00000000",
            INIT_35 => X"0000001200000000000000150000000000000016000000000000000900000000",
            INIT_36 => X"0000001200000000000000070000000000000011000000000000001000000000",
            INIT_37 => X"0000001b00000000000000000000000000000011000000000000000c00000000",
            INIT_38 => X"00000008000000000000000f0000000000000000000000000000002b00000000",
            INIT_39 => X"000000090000000000000010000000000000000d000000000000001300000000",
            INIT_3A => X"0000000a000000000000000c000000000000000a000000000000000c00000000",
            INIT_3B => X"0000000a00000000000000200000000000000000000000000000000300000000",
            INIT_3C => X"0000000800000000000000080000000000000015000000000000000000000000",
            INIT_3D => X"0000000a0000000000000006000000000000000f000000000000000b00000000",
            INIT_3E => X"000000000000000000000007000000000000000b000000000000000700000000",
            INIT_3F => X"0000001000000000000000040000000000000000000000000000004100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000a0000000000000004000000000000001200000000",
            INIT_41 => X"0000000000000000000000010000000000000001000000000000000e00000000",
            INIT_42 => X"0000003e00000000000000270000000000000000000000000000000000000000",
            INIT_43 => X"0000000a000000000000000a0000000000000003000000000000000000000000",
            INIT_44 => X"0000000d000000000000000e000000000000000b000000000000000800000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000008700000000000000000000000000000001000000000000000000000000",
            INIT_47 => X"00000009000000000000000b0000000000000015000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000014000000000000000d00000000",
            INIT_49 => X"00000009000000000000002b000000000000001b000000000000000000000000",
            INIT_4A => X"0000001600000000000000c00000000000000000000000000000000000000000",
            INIT_4B => X"0000000f000000000000000a0000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_4E => X"0000000000000000000000550000000000000085000000000000000000000000",
            INIT_4F => X"0000000e0000000000000000000000000000000c000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_51 => X"0000003300000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"000000000000000000000000000000000000000000000000000000a500000000",
            INIT_53 => X"00000000000000000000008c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_55 => X"0000003a00000000000000000000000000000018000000000000000000000000",
            INIT_56 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_57 => X"000000200000000000000016000000000000006a000000000000000000000000",
            INIT_58 => X"0000004800000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000002000000000000000000000000000000000000000000000005c00000000",
            INIT_5A => X"000000090000000000000000000000000000005d000000000000002a00000000",
            INIT_5B => X"0000000000000000000000000000000000000044000000000000000000000000",
            INIT_5C => X"0000000000000000000000b50000000000000000000000000000000000000000",
            INIT_5D => X"0000006e00000000000000000000000000000000000000000000001900000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_60 => X"00000033000000000000000000000000000000b2000000000000000000000000",
            INIT_61 => X"00000000000000000000006f0000000000000000000000000000000000000000",
            INIT_62 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000002b000000000000001e0000000000000000000000000000005600000000",
            INIT_65 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_66 => X"0000000000000000000000140000000000000007000000000000001100000000",
            INIT_67 => X"0000000b00000000000000080000000000000004000000000000000000000000",
            INIT_68 => X"00000002000000000000002b000000000000000e000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000f00000000000000000000000000000001000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000160000000000000009000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000026000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "samplegold_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000005000000000000000310000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000028000000000000004000000000",
            INIT_03 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"000000160000000000000000000000000000002c000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_0A => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000010000000000000000d000000000000000600000000",
            INIT_0D => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_11 => X"00000052000000000000002d0000000000000048000000000000000000000000",
            INIT_12 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_13 => X"0000000200000000000000000000000000000000000000000000000d00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000800000000000000020000000000000011000000000000000000000000",
            INIT_16 => X"000000020000000000000008000000000000001b000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001a00000000000000150000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000030000000000000000000000000000000600000000",
            INIT_1B => X"0000004900000000000000410000000000000010000000000000001000000000",
            INIT_1C => X"0000001a0000000000000000000000000000004b000000000000004e00000000",
            INIT_1D => X"00000001000000000000002e000000000000001b000000000000001400000000",
            INIT_1E => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000001300000000000000000000000000000014000000000000000800000000",
            INIT_21 => X"0000000f00000000000000010000000000000003000000000000000400000000",
            INIT_22 => X"000000160000000000000019000000000000001a000000000000000f00000000",
            INIT_23 => X"000000170000000000000011000000000000001d000000000000001800000000",
            INIT_24 => X"000000000000000000000011000000000000000a000000000000001200000000",
            INIT_25 => X"0000001700000000000000230000000000000004000000000000001600000000",
            INIT_26 => X"00000019000000000000001c000000000000001c000000000000000d00000000",
            INIT_27 => X"0000001200000000000000140000000000000015000000000000001a00000000",
            INIT_28 => X"0000001800000000000000000000000000000000000000000000002400000000",
            INIT_29 => X"000000190000000000000013000000000000001a000000000000000700000000",
            INIT_2A => X"0000001400000000000000160000000000000018000000000000001700000000",
            INIT_2B => X"0000002b00000000000000170000000000000012000000000000001300000000",
            INIT_2C => X"00000003000000000000000e0000000000000000000000000000000000000000",
            INIT_2D => X"0000001300000000000000150000000000000017000000000000001600000000",
            INIT_2E => X"00000015000000000000001b0000000000000017000000000000001500000000",
            INIT_2F => X"0000001000000000000000000000000000000013000000000000001100000000",
            INIT_30 => X"00000014000000000000000b000000000000000b000000000000000500000000",
            INIT_31 => X"0000001c00000000000000150000000000000016000000000000001600000000",
            INIT_32 => X"00000027000000000000001e000000000000001d000000000000001f00000000",
            INIT_33 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001600000000000000160000000000000010000000000000000c00000000",
            INIT_35 => X"0000003d00000000000000280000000000000014000000000000001400000000",
            INIT_36 => X"0000000000000000000000040000000000000004000000000000002a00000000",
            INIT_37 => X"0000000000000000000000280000000000000000000000000000001e00000000",
            INIT_38 => X"0000001000000000000000140000000000000017000000000000000c00000000",
            INIT_39 => X"000000000000000000000009000000000000002f000000000000002400000000",
            INIT_3A => X"0000002a000000000000006a0000000000000008000000000000000000000000",
            INIT_3B => X"0000000800000000000000150000000000000000000000000000000000000000",
            INIT_3C => X"0000000c00000000000000340000000000000015000000000000001600000000",
            INIT_3D => X"0000002000000000000000000000000000000015000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000020000000000000002200000000",
            INIT_3F => X"00000015000000000000002c0000000000000013000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000170000000000000000000000000000003000000000",
            INIT_41 => X"00000000000000000000003f0000000000000046000000000000001400000000",
            INIT_42 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000006a00000000000000340000000000000009000000000000002800000000",
            INIT_44 => X"000000220000000000000000000000000000000d000000000000000000000000",
            INIT_45 => X"000000000000000000000000000000000000000c000000000000006c00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_47 => X"00000000000000000000000a0000000000000056000000000000000000000000",
            INIT_48 => X"0000005500000000000000370000000000000000000000000000000000000000",
            INIT_49 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_4B => X"00000000000000000000000a0000000000000012000000000000002c00000000",
            INIT_4C => X"00000000000000000000005a000000000000002a000000000000001a00000000",
            INIT_4D => X"0000003e0000000000000000000000000000000b000000000000000000000000",
            INIT_4E => X"0000002400000000000000020000000000000000000000000000002000000000",
            INIT_4F => X"0000003800000000000000000000000000000016000000000000001800000000",
            INIT_50 => X"000000000000000000000000000000000000001e000000000000000800000000",
            INIT_51 => X"0000003800000000000000000000000000000000000000000000002500000000",
            INIT_52 => X"000000170000000000000013000000000000000e000000000000000000000000",
            INIT_53 => X"0000000a00000000000000120000000000000000000000000000000000000000",
            INIT_54 => X"0000003000000000000000000000000000000001000000000000000a00000000",
            INIT_55 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_56 => X"000000030000000000000006000000000000000f000000000000000c00000000",
            INIT_57 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_58 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_59 => X"0000000f00000000000000050000000000000004000000000000000000000000",
            INIT_5A => X"00000089000000000000008a000000000000008e000000000000009500000000",
            INIT_5B => X"0000006b00000000000000710000000000000076000000000000008000000000",
            INIT_5C => X"0000003f000000000000004d000000000000004d000000000000005d00000000",
            INIT_5D => X"0000007d000000000000003d0000000000000015000000000000001c00000000",
            INIT_5E => X"00000066000000000000006d0000000000000072000000000000007600000000",
            INIT_5F => X"000000520000000000000058000000000000005c000000000000005e00000000",
            INIT_60 => X"0000001800000000000000320000000000000044000000000000005100000000",
            INIT_61 => X"0000005200000000000000550000000000000047000000000000002600000000",
            INIT_62 => X"0000005500000000000000550000000000000058000000000000005600000000",
            INIT_63 => X"0000004f00000000000000540000000000000056000000000000005600000000",
            INIT_64 => X"0000003c00000000000000240000000000000012000000000000002f00000000",
            INIT_65 => X"000000540000000000000052000000000000004a000000000000004800000000",
            INIT_66 => X"0000005b00000000000000590000000000000056000000000000005500000000",
            INIT_67 => X"0000001c00000000000000450000000000000055000000000000005800000000",
            INIT_68 => X"00000049000000000000004a000000000000003d000000000000000e00000000",
            INIT_69 => X"0000005700000000000000570000000000000056000000000000004f00000000",
            INIT_6A => X"0000004700000000000000470000000000000054000000000000005500000000",
            INIT_6B => X"00000014000000000000001a0000000000000038000000000000003e00000000",
            INIT_6C => X"0000005600000000000000450000000000000042000000000000003300000000",
            INIT_6D => X"0000004800000000000000540000000000000055000000000000005600000000",
            INIT_6E => X"000000110000000000000024000000000000002f000000000000003900000000",
            INIT_6F => X"0000000400000000000000170000000000000010000000000000000500000000",
            INIT_70 => X"000000570000000000000056000000000000003c000000000000002a00000000",
            INIT_71 => X"0000000e00000000000000370000000000000045000000000000005300000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000030000000000000007000000000000001b000000000000000600000000",
            INIT_74 => X"0000004200000000000000530000000000000055000000000000002000000000",
            INIT_75 => X"0000000b000000000000000f0000000000000012000000000000002c00000000",
            INIT_76 => X"00000006000000000000001c000000000000001d000000000000000600000000",
            INIT_77 => X"0000001200000000000000050000000000000010000000000000001400000000",
            INIT_78 => X"00000000000000000000001b0000000000000041000000000000005400000000",
            INIT_79 => X"0000001000000000000000000000000000000000000000000000000100000000",
            INIT_7A => X"00000014000000000000000a0000000000000003000000000000000800000000",
            INIT_7B => X"000000440000000000000012000000000000001c000000000000001500000000",
            INIT_7C => X"0000000300000000000000000000000000000014000000000000003200000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001100000000000000130000000000000000000000000000000400000000",
            INIT_7F => X"000000020000000000000037000000000000000a000000000000000600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "samplegold_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_01 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000000000003000000000000002f000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_05 => X"000000050000000000000000000000000000000a000000000000000300000000",
            INIT_06 => X"0000000900000000000000040000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000003000000000000002200000000",
            INIT_08 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_09 => X"00000000000000000000000a0000000000000000000000000000000c00000000",
            INIT_0A => X"0000002400000000000000070000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_0E => X"0000000c00000000000000200000000000000003000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_10 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_11 => X"0000000300000000000000030000000000000001000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000200000000000000000000000000000005000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000011000000000000001400000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000006000000000000000100000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000002000000000000000f000000000000000000000000",
            INIT_2F => X"0000001e000000000000000f0000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000006000000000000000c000000000000000000000000",
            INIT_34 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000017000000000000001400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"00000020000000000000000f0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000250000000000000014000000000000000000000000",
            INIT_3D => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_3F => X"000000000000000000000003000000000000000b000000000000001800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000000d000000000000001200000000",
            INIT_41 => X"0000001200000000000000090000000000000000000000000000000000000000",
            INIT_42 => X"0000001c00000000000000030000000000000000000000000000001600000000",
            INIT_43 => X"0000000000000000000000000000000000000003000000000000001000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000b0000000000000028000000000000001e000000000000000e00000000",
            INIT_47 => X"0000002b00000000000000280000000000000018000000000000001200000000",
            INIT_48 => X"0000002700000000000000260000000000000026000000000000002900000000",
            INIT_49 => X"0000002e00000000000000210000000000000008000000000000000e00000000",
            INIT_4A => X"0000000000000000000000000000000000000026000000000000002d00000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "samplegold_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000400000000000000000000000000000006000000000000000900000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000100000000000000030000000000000000000000000000000000000000",
            INIT_0D => X"00000000000000000000000e000000000000001a000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000014000000000000000b0000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000009000000000000001000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000004500000000000000090000000000000000000000000000000600000000",
            INIT_14 => X"000000000000000000000019000000000000004c000000000000006e00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000009000000000000004e00000000",
            INIT_18 => X"000000050000000000000000000000000000003b000000000000005700000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_1B => X"0000000400000000000000070000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000000000000000000000000001b000000000000005f00000000",
            INIT_1D => X"00000026000000000000001c0000000000000000000000000000000000000000",
            INIT_1E => X"00000092000000000000000a0000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000004000000000000009500000000000000f000000000",
            INIT_20 => X"00000000000000000000005a0000000000000014000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_22 => X"000000000000000000000025000000000000000a000000000000000000000000",
            INIT_23 => X"0000004400000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000007800000000000000130000000000000024000000000000008700000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000b000000000000005b000000000000005e000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000002900000000000000370000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000800000000000000010000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000006000000000000001f00000000",
            INIT_2E => X"00000000000000000000000d0000000000000005000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000005b00000000000000310000000000000000000000000000000000000000",
            INIT_31 => X"0000000e00000000000000000000000000000025000000000000007200000000",
            INIT_32 => X"0000000000000000000000000000000000000036000000000000001200000000",
            INIT_33 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000002c00000000000000100000000000000006000000000000000000000000",
            INIT_38 => X"0000002000000000000000290000000000000026000000000000004400000000",
            INIT_39 => X"0000000000000000000000000000000000000010000000000000001500000000",
            INIT_3A => X"0000000c00000000000000090000000000000008000000000000000000000000",
            INIT_3B => X"0000002a000000000000002c0000000000000027000000000000002900000000",
            INIT_3C => X"0000001c00000000000000230000000000000020000000000000002300000000",
            INIT_3D => X"0000001900000000000000170000000000000019000000000000001c00000000",
            INIT_3E => X"0000002500000000000000120000000000000014000000000000000900000000",
            INIT_3F => X"000000160000000000000018000000000000001c000000000000001b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001600000000000000170000000000000019000000000000001500000000",
            INIT_41 => X"0000000800000000000000070000000000000022000000000000001600000000",
            INIT_42 => X"0000001100000000000000150000000000000014000000000000001e00000000",
            INIT_43 => X"0000001200000000000000140000000000000010000000000000001100000000",
            INIT_44 => X"0000001a00000000000000170000000000000017000000000000001400000000",
            INIT_45 => X"0000001f000000000000000f0000000000000003000000000000001200000000",
            INIT_46 => X"0000001200000000000000110000000000000012000000000000001000000000",
            INIT_47 => X"0000001700000000000000130000000000000013000000000000001100000000",
            INIT_48 => X"0000000200000000000000160000000000000017000000000000001700000000",
            INIT_49 => X"0000001200000000000000150000000000000012000000000000001600000000",
            INIT_4A => X"0000000f000000000000000f0000000000000010000000000000001200000000",
            INIT_4B => X"0000001b00000000000000180000000000000012000000000000001300000000",
            INIT_4C => X"000000160000000000000000000000000000000a000000000000002300000000",
            INIT_4D => X"0000001100000000000000140000000000000010000000000000001400000000",
            INIT_4E => X"000000190000000000000010000000000000000f000000000000000e00000000",
            INIT_4F => X"000000000000000000000000000000000000000f000000000000001f00000000",
            INIT_50 => X"0000001d00000000000000000000000000000006000000000000000000000000",
            INIT_51 => X"0000000d000000000000000f000000000000000f000000000000000b00000000",
            INIT_52 => X"0000000d000000000000000e0000000000000016000000000000000c00000000",
            INIT_53 => X"0000002c000000000000000b0000000000000000000000000000000000000000",
            INIT_54 => X"0000001900000000000000060000000000000000000000000000001a00000000",
            INIT_55 => X"00000019000000000000000c000000000000000e000000000000000f00000000",
            INIT_56 => X"0000000b000000000000000e0000000000000006000000000000000a00000000",
            INIT_57 => X"00000000000000000000001a0000000000000029000000000000002100000000",
            INIT_58 => X"00000021000000000000001b0000000000000000000000000000000000000000",
            INIT_59 => X"0000000800000000000000090000000000000018000000000000000b00000000",
            INIT_5A => X"0000001a000000000000001f0000000000000019000000000000000100000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"000000190000000000000011000000000000000d000000000000001a00000000",
            INIT_5D => X"00000000000000000000000d0000000000000000000000000000001e00000000",
            INIT_5E => X"0000000000000000000000050000000000000027000000000000001700000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000a00000000000000140000000000000000000000000000000000000000",
            INIT_61 => X"0000002500000000000000060000000000000002000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_63 => X"000000000000000000000000000000000000001c000000000000001100000000",
            INIT_64 => X"0000000c00000000000000000000000000000012000000000000000000000000",
            INIT_65 => X"0000001b000000000000001e000000000000001a000000000000000000000000",
            INIT_66 => X"0000000700000000000000100000000000000000000000000000000000000000",
            INIT_67 => X"0000000800000000000000000000000000000000000000000000002500000000",
            INIT_68 => X"000000000000000000000013000000000000000d000000000000001000000000",
            INIT_69 => X"0000000000000000000000170000000000000010000000000000002400000000",
            INIT_6A => X"000000080000000000000000000000000000001b000000000000000000000000",
            INIT_6B => X"0000000f00000000000000190000000000000000000000000000001b00000000",
            INIT_6C => X"0000000d00000000000000000000000000000007000000000000000a00000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001e00000000000000000000000000000000000000000000001c00000000",
            INIT_6F => X"0000000d000000000000000e000000000000001a000000000000000600000000",
            INIT_70 => X"000000120000000000000012000000000000000a000000000000001200000000",
            INIT_71 => X"0000001f00000000000000120000000000000010000000000000001100000000",
            INIT_72 => X"0000001900000000000000170000000000000005000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "samplegold_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000001b0000000000000006000000000000003a000000000000003200000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000f0000000000000029000000000000002e000000000000001300000000",
            INIT_0C => X"0000000900000000000000250000000000000027000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_10 => X"00000000000000000000000d0000000000000063000000000000003700000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000012000000000000002e000000000000000900000000",
            INIT_13 => X"0000004c00000000000000350000000000000040000000000000001900000000",
            INIT_14 => X"0000001800000000000000000000000000000000000000000000000c00000000",
            INIT_15 => X"0000001100000000000000270000000000000000000000000000000000000000",
            INIT_16 => X"0000003c00000000000000000000000000000000000000000000001700000000",
            INIT_17 => X"0000001000000000000000400000000000000064000000000000003500000000",
            INIT_18 => X"000000000000000000000038000000000000002d000000000000001500000000",
            INIT_19 => X"0000000300000000000000200000000000000038000000000000004b00000000",
            INIT_1A => X"0000006900000000000000390000000000000000000000000000000000000000",
            INIT_1B => X"0000004f000000000000002a000000000000002c000000000000003200000000",
            INIT_1C => X"0000000100000000000000000000000000000045000000000000004700000000",
            INIT_1D => X"0000001700000000000000000000000000000020000000000000002a00000000",
            INIT_1E => X"00000008000000000000005b0000000000000038000000000000000a00000000",
            INIT_1F => X"0000004b000000000000002a0000000000000013000000000000000700000000",
            INIT_20 => X"0000002c000000000000000d0000000000000000000000000000000000000000",
            INIT_21 => X"0000002000000000000000050000000000000000000000000000000e00000000",
            INIT_22 => X"0000000d00000000000000030000000000000042000000000000003200000000",
            INIT_23 => X"00000000000000000000002d000000000000002f000000000000000c00000000",
            INIT_24 => X"00000030000000000000003c0000000000000004000000000000000000000000",
            INIT_25 => X"000000610000000000000060000000000000005b000000000000004900000000",
            INIT_26 => X"0000001100000000000000230000000000000016000000000000004200000000",
            INIT_27 => X"0000000000000000000000000000000000000003000000000000001e00000000",
            INIT_28 => X"0000000600000000000000020000000000000000000000000000000000000000",
            INIT_29 => X"0000000100000000000000050000000000000005000000000000000500000000",
            INIT_2A => X"0000000000000000000000060000000000000025000000000000000d00000000",
            INIT_2B => X"000000a1000000000000009a0000000000000000000000000000000000000000",
            INIT_2C => X"0000009e00000000000000a700000000000000b100000000000000af00000000",
            INIT_2D => X"000000650000000000000082000000000000008c000000000000009a00000000",
            INIT_2E => X"0000003c00000000000000210000000000000042000000000000005d00000000",
            INIT_2F => X"0000009b000000000000009800000000000000a4000000000000004900000000",
            INIT_30 => X"0000008300000000000000860000000000000091000000000000009c00000000",
            INIT_31 => X"0000004e00000000000000650000000000000070000000000000007800000000",
            INIT_32 => X"000000500000000000000037000000000000000b000000000000003100000000",
            INIT_33 => X"0000007d00000000000000830000000000000080000000000000008600000000",
            INIT_34 => X"0000006c00000000000000710000000000000072000000000000007700000000",
            INIT_35 => X"0000000e0000000000000030000000000000005d000000000000006500000000",
            INIT_36 => X"0000006b00000000000000530000000000000046000000000000001d00000000",
            INIT_37 => X"0000006f000000000000006c000000000000006e000000000000006e00000000",
            INIT_38 => X"0000005f00000000000000610000000000000066000000000000006c00000000",
            INIT_39 => X"0000004700000000000000210000000000000006000000000000004e00000000",
            INIT_3A => X"0000007000000000000000680000000000000059000000000000005600000000",
            INIT_3B => X"00000064000000000000006e000000000000006e000000000000007100000000",
            INIT_3C => X"00000002000000000000002b0000000000000049000000000000005800000000",
            INIT_3D => X"0000005800000000000000410000000000000018000000000000000000000000",
            INIT_3E => X"0000006e0000000000000070000000000000006d000000000000005900000000",
            INIT_3F => X"00000018000000000000002e000000000000005e000000000000006b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000010000000000000020000000000000001a00000000",
            INIT_41 => X"0000005300000000000000310000000000000025000000000000000000000000",
            INIT_42 => X"0000005c0000000000000068000000000000006f000000000000007000000000",
            INIT_43 => X"0000000000000000000000000000000000000023000000000000004200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_45 => X"00000070000000000000003c000000000000001d000000000000000000000000",
            INIT_46 => X"0000000000000000000000230000000000000047000000000000006900000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000004e000000000000006e0000000000000000000000000000000000000000",
            INIT_4A => X"0000000100000000000000000000000000000004000000000000001900000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000150000000000000056000000000000000000000000",
            INIT_4E => X"0000000400000000000000040000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000000a000000000000005100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000c00000000000000050000000000000000000000000000000000000000",
            INIT_54 => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_58 => X"00000000000000000000002e0000000000000009000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000080000000000000026000000000000001300000000",
            INIT_5D => X"0000000c00000000000000090000000000000007000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_5F => X"0000000600000000000000000000000000000001000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000010000000000000004000000000000000000000000",
            INIT_63 => X"0000006c00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000064000000000000006c0000000000000066000000000000006700000000",
            INIT_65 => X"0000004600000000000000520000000000000055000000000000005a00000000",
            INIT_66 => X"000000000000000000000030000000000000003d000000000000003000000000",
            INIT_67 => X"0000005c000000000000005d000000000000002e000000000000001d00000000",
            INIT_68 => X"000000410000000000000046000000000000004d000000000000005200000000",
            INIT_69 => X"0000003b000000000000003b000000000000003e000000000000003f00000000",
            INIT_6A => X"0000001e00000000000000190000000000000022000000000000002700000000",
            INIT_6B => X"0000003e00000000000000380000000000000039000000000000002c00000000",
            INIT_6C => X"000000380000000000000038000000000000003a000000000000003800000000",
            INIT_6D => X"00000003000000000000003d000000000000003a000000000000003b00000000",
            INIT_6E => X"0000002b00000000000000250000000000000023000000000000001200000000",
            INIT_6F => X"0000003900000000000000370000000000000038000000000000003300000000",
            INIT_70 => X"0000003800000000000000340000000000000039000000000000003b00000000",
            INIT_71 => X"0000002300000000000000000000000000000031000000000000003c00000000",
            INIT_72 => X"000000320000000000000032000000000000002f000000000000003700000000",
            INIT_73 => X"0000003800000000000000380000000000000038000000000000003800000000",
            INIT_74 => X"0000002200000000000000280000000000000024000000000000003100000000",
            INIT_75 => X"00000014000000000000001b0000000000000011000000000000000d00000000",
            INIT_76 => X"000000370000000000000035000000000000002d000000000000002f00000000",
            INIT_77 => X"0000001e000000000000002c0000000000000035000000000000003600000000",
            INIT_78 => X"0000000300000000000000010000000000000012000000000000001500000000",
            INIT_79 => X"000000090000000000000017000000000000001b000000000000000000000000",
            INIT_7A => X"0000003000000000000000380000000000000038000000000000002a00000000",
            INIT_7B => X"0000000000000000000000000000000000000018000000000000002d00000000",
            INIT_7C => X"0000000000000000000000210000000000000000000000000000000400000000",
            INIT_7D => X"000000170000000000000000000000000000001a000000000000000000000000",
            INIT_7E => X"0000000f00000000000000270000000000000034000000000000003900000000",
            INIT_7F => X"0000000000000000000000000000000000000016000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "samplegold_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000005000000000000001300000000",
            INIT_01 => X"000000340000000000000000000000000000000f000000000000000b00000000",
            INIT_02 => X"0000000000000000000000080000000000000007000000000000002700000000",
            INIT_03 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_04 => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000360000000000000000000000000000001f00000000",
            INIT_06 => X"0000000e00000000000000120000000000000000000000000000000100000000",
            INIT_07 => X"0000000100000000000000000000000000000000000000000000001800000000",
            INIT_08 => X"0000000000000000000000000000000000000001000000000000000600000000",
            INIT_09 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_0A => X"0000001200000000000000000000000000000013000000000000000000000000",
            INIT_0B => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000300000000000000000000000000000012000000000000001400000000",
            INIT_0E => X"0000000000000000000000030000000000000000000000000000000600000000",
            INIT_0F => X"0000000900000000000000060000000000000000000000000000000000000000",
            INIT_10 => X"00000017000000000000001e0000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_14 => X"0000000500000000000000140000000000000007000000000000001000000000",
            INIT_15 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000120000000000000000000000000000000d000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000f000000000000000200000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_1B => X"0000000700000000000000050000000000000005000000000000000d00000000",
            INIT_1C => X"0000001c00000000000000140000000000000015000000000000001500000000",
            INIT_1D => X"00000011000000000000000e0000000000000007000000000000001200000000",
            INIT_1E => X"00000008000000000000000a000000000000000b000000000000000d00000000",
            INIT_1F => X"0000001500000000000000000000000000000000000000000000000300000000",
            INIT_20 => X"00000005000000000000000d0000000000000013000000000000001300000000",
            INIT_21 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_23 => X"0000001200000000000000140000000000000001000000000000000000000000",
            INIT_24 => X"000000000000000000000000000000000000000f000000000000001200000000",
            INIT_25 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000012000000000000000c000000000000000a000000000000000700000000",
            INIT_27 => X"00000005000000000000000c000000000000000d000000000000000f00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000002000000000000000b000000000000000c000000000000000b00000000",
            INIT_2B => X"00000003000000000000001b0000000000000005000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000002900000000000000000000000000000004000000000000000400000000",
            INIT_2F => X"0000000000000000000000000000000000000028000000000000003200000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000003300000000000000340000000000000009000000000000000900000000",
            INIT_33 => X"000000000000000000000000000000000000001f000000000000002400000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000002c00000000000000250000000000000027000000000000001300000000",
            INIT_37 => X"0000000000000000000000000000000000000010000000000000001300000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001b00000000000000180000000000000024000000000000002400000000",
            INIT_3B => X"000000000000000000000000000000000000001f000000000000001e00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000002600000000000000100000000000000000000000000000000000000000",
            INIT_3E => X"00000020000000000000005a0000000000000061000000000000004400000000",
            INIT_3F => X"0000000000000000000000000000000000000002000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000006800000000000000600000000000000000000000000000000000000000",
            INIT_42 => X"0000000a0000000000000015000000000000001f000000000000006100000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000030000000000000005d000000000000007a000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"00000016000000000000001e000000000000002b000000000000002b00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000a00000000000000180000000000000017000000000000001100000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000001200000000000000160000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000900000000000000010000000000000000000000000000000000000000",
            INIT_5B => X"000000000000000000000003000000000000000d000000000000000e00000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000020000000000000001d000000000000000000000000",
            INIT_64 => X"00000000000000000000000b0000000000000004000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000200000000000000010000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_68 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_6B => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_6E => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000001000000000000000100000000000000006000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000f000000000000002700000000",
            INIT_77 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000100000000000000010000000000000000000000000000000900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "samplegold_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000130000000000000007000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_09 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0B => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000f000000000000000f0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000002e0000000000000024000000000000001c000000000000000c00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000034000000000000002e0000000000000026000000000000001f00000000",
            INIT_1A => X"0000000000000000000000090000000000000003000000000000001a00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000f000000000000000e0000000000000000000000000000000000000000",
            INIT_1D => X"0000003500000000000000350000000000000021000000000000001000000000",
            INIT_1E => X"00000008000000000000000b000000000000001f000000000000002c00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_20 => X"0000001100000000000000080000000000000008000000000000000000000000",
            INIT_21 => X"00000038000000000000002f0000000000000027000000000000001e00000000",
            INIT_22 => X"0000000f00000000000000170000000000000020000000000000002c00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000002000000000000000150000000000000009000000000000000000000000",
            INIT_25 => X"0000002c000000000000002d000000000000001c000000000000001b00000000",
            INIT_26 => X"0000000000000000000000050000000000000016000000000000002700000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000170000000000000021000000000000000f000000000000000000000000",
            INIT_29 => X"00000023000000000000002e0000000000000024000000000000001200000000",
            INIT_2A => X"0000000000000000000000000000000000000004000000000000001100000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000001100000000000000180000000000000019000000000000000800000000",
            INIT_2D => X"00000014000000000000001f0000000000000026000000000000001c00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_2F => X"0000000900000000000000040000000000000000000000000000000000000000",
            INIT_30 => X"00000017000000000000000f0000000000000017000000000000001d00000000",
            INIT_31 => X"0000001e00000000000000200000000000000021000000000000002100000000",
            INIT_32 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000019000000000000001d000000000000001c000000000000000f00000000",
            INIT_34 => X"00000025000000000000001c0000000000000019000000000000001a00000000",
            INIT_35 => X"000000000000000000000018000000000000001c000000000000002400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000001600000000000000040000000000000015000000000000001700000000",
            INIT_38 => X"0000002600000000000000190000000000000010000000000000001c00000000",
            INIT_39 => X"0000000000000000000000000000000000000020000000000000002100000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000c00000000000000070000000000000012000000000000000a00000000",
            INIT_3C => X"0000002a00000000000000290000000000000012000000000000000200000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_3E => X"0000000c00000000000000100000000000000016000000000000000c00000000",
            INIT_3F => X"0000000c00000000000000130000000000000014000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000026000000000000002e0000000000000024000000000000001200000000",
            INIT_41 => X"0000001e000000000000001c000000000000000f000000000000000000000000",
            INIT_42 => X"0000002500000000000000180000000000000017000000000000001f00000000",
            INIT_43 => X"0000001c0000000000000019000000000000001f000000000000002500000000",
            INIT_44 => X"00000097000000000000002a000000000000002d000000000000002600000000",
            INIT_45 => X"00000097000000000000009d000000000000008e000000000000009200000000",
            INIT_46 => X"00000078000000000000007e0000000000000094000000000000009600000000",
            INIT_47 => X"0000003e0000000000000050000000000000005f000000000000006d00000000",
            INIT_48 => X"0000008f00000000000000930000000000000034000000000000003500000000",
            INIT_49 => X"00000084000000000000008e0000000000000076000000000000008b00000000",
            INIT_4A => X"00000067000000000000006d0000000000000081000000000000008c00000000",
            INIT_4B => X"0000006b0000000000000061000000000000005e000000000000006100000000",
            INIT_4C => X"0000008300000000000000860000000000000088000000000000006d00000000",
            INIT_4D => X"0000006e0000000000000064000000000000006b000000000000005e00000000",
            INIT_4E => X"0000009d000000000000009a0000000000000073000000000000006e00000000",
            INIT_4F => X"0000007a000000000000008d0000000000000094000000000000009f00000000",
            INIT_50 => X"0000005000000000000000780000000000000081000000000000007e00000000",
            INIT_51 => X"000000780000000000000064000000000000005f000000000000005400000000",
            INIT_52 => X"000000a4000000000000009f000000000000008a000000000000008600000000",
            INIT_53 => X"000000aa00000000000000730000000000000085000000000000008900000000",
            INIT_54 => X"0000005b000000000000007300000000000000fe00000000000000d200000000",
            INIT_55 => X"0000007f0000000000000094000000000000009d000000000000006e00000000",
            INIT_56 => X"0000009700000000000000930000000000000084000000000000007f00000000",
            INIT_57 => X"0000012000000000000001120000000000000096000000000000009c00000000",
            INIT_58 => X"0000007e0000000000000067000000000000007f000000000000011800000000",
            INIT_59 => X"000000870000000000000086000000000000009200000000000000ad00000000",
            INIT_5A => X"000000b10000000000000096000000000000007e000000000000008400000000",
            INIT_5B => X"000000fe0000000000000109000000000000010a00000000000000ad00000000",
            INIT_5C => X"000000a50000000000000085000000000000007100000000000000ca00000000",
            INIT_5D => X"0000008600000000000000960000000000000094000000000000008d00000000",
            INIT_5E => X"0000009900000000000000990000000000000097000000000000007500000000",
            INIT_5F => X"000000e40000000000000118000000000000010100000000000000f300000000",
            INIT_60 => X"0000008f00000000000000ab000000000000007900000000000000db00000000",
            INIT_61 => X"0000007a000000000000008d00000000000000b000000000000000a700000000",
            INIT_62 => X"00000110000000000000007f000000000000007e000000000000007f00000000",
            INIT_63 => X"0000012500000000000001400000000000000148000000000000012800000000",
            INIT_64 => X"000000a100000000000000b500000000000000b8000000000000010800000000",
            INIT_65 => X"000000770000000000000086000000000000009600000000000000ac00000000",
            INIT_66 => X"000001b5000000000000017a000000000000008a000000000000008b00000000",
            INIT_67 => X"0000011a000000000000011b000000000000018c00000000000001c200000000",
            INIT_68 => X"000000a9000000000000009f00000000000000bc00000000000000ba00000000",
            INIT_69 => X"00000077000000000000007c000000000000009700000000000000a800000000",
            INIT_6A => X"0000016200000000000001d500000000000001d4000000000000004c00000000",
            INIT_6B => X"0000009700000000000000ac00000000000000bd00000000000000dd00000000",
            INIT_6C => X"000000a600000000000000a800000000000000a0000000000000008d00000000",
            INIT_6D => X"0000006a0000000000000075000000000000007a000000000000008e00000000",
            INIT_6E => X"000000d600000000000000e60000000000000137000000000000018b00000000",
            INIT_6F => X"0000008d0000000000000072000000000000005d000000000000009f00000000",
            INIT_70 => X"000000a50000000000000098000000000000007a000000000000006400000000",
            INIT_71 => X"000000c900000000000000860000000000000078000000000000008300000000",
            INIT_72 => X"000000ac00000000000000b200000000000000b200000000000000c300000000",
            INIT_73 => X"00000071000000000000007f0000000000000089000000000000009200000000",
            INIT_74 => X"0000009000000000000000ae00000000000000c3000000000000008600000000",
            INIT_75 => X"000000a10000000000000096000000000000007a000000000000007600000000",
            INIT_76 => X"000000790000000000000073000000000000009900000000000000ad00000000",
            INIT_77 => X"0000008300000000000000770000000000000084000000000000007800000000",
            INIT_78 => X"0000006a000000000000008d0000000000000097000000000000009300000000",
            INIT_79 => X"00000065000000000000007d0000000000000098000000000000007000000000",
            INIT_7A => X"00000084000000000000007e0000000000000055000000000000005a00000000",
            INIT_7B => X"00000065000000000000005d000000000000005f000000000000007100000000",
            INIT_7C => X"0000005a0000000000000056000000000000006d000000000000007600000000",
            INIT_7D => X"0000002200000000000000150000000000000017000000000000001800000000",
            INIT_7E => X"0000001c00000000000000230000000000000029000000000000002a00000000",
            INIT_7F => X"0000000c000000000000000f0000000000000014000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "samplegold_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001600000000000000000000000000000000000000000000000600000000",
            INIT_01 => X"000000340000000000000017000000000000001a000000000000001800000000",
            INIT_02 => X"0000001900000000000000260000000000000037000000000000003500000000",
            INIT_03 => X"0000000b000000000000000d000000000000000e000000000000001300000000",
            INIT_04 => X"0000001800000000000000170000000000000011000000000000000c00000000",
            INIT_05 => X"000000300000000000000031000000000000001a000000000000002300000000",
            INIT_06 => X"0000002000000000000000230000000000000039000000000000003800000000",
            INIT_07 => X"0000002600000000000000260000000000000029000000000000002300000000",
            INIT_08 => X"0000001300000000000000110000000000000015000000000000002500000000",
            INIT_09 => X"0000003200000000000000280000000000000027000000000000001800000000",
            INIT_0A => X"00000037000000000000003c000000000000003b000000000000004200000000",
            INIT_0B => X"0000002500000000000000260000000000000026000000000000003400000000",
            INIT_0C => X"0000002000000000000000410000000000000019000000000000000f00000000",
            INIT_0D => X"000000400000000000000035000000000000002a000000000000002600000000",
            INIT_0E => X"0000003e00000000000000430000000000000040000000000000004700000000",
            INIT_0F => X"0000003300000000000000350000000000000036000000000000002d00000000",
            INIT_10 => X"0000001c000000000000001f0000000000000053000000000000003f00000000",
            INIT_11 => X"0000003e0000000000000043000000000000003d000000000000002300000000",
            INIT_12 => X"0000003c00000000000000380000000000000046000000000000004500000000",
            INIT_13 => X"0000003d000000000000003c0000000000000043000000000000004600000000",
            INIT_14 => X"0000003300000000000000320000000000000024000000000000003f00000000",
            INIT_15 => X"000000400000000000000039000000000000003b000000000000004600000000",
            INIT_16 => X"00000041000000000000003e0000000000000037000000000000004700000000",
            INIT_17 => X"0000004700000000000000350000000000000031000000000000003a00000000",
            INIT_18 => X"0000003c00000000000000160000000000000026000000000000004800000000",
            INIT_19 => X"000000430000000000000041000000000000003c000000000000003f00000000",
            INIT_1A => X"0000002b0000000000000027000000000000003a000000000000003a00000000",
            INIT_1B => X"0000003d000000000000003c0000000000000031000000000000003300000000",
            INIT_1C => X"00000044000000000000004b000000000000004c000000000000005300000000",
            INIT_1D => X"0000003e000000000000003f000000000000003f000000000000003900000000",
            INIT_1E => X"00000040000000000000003e0000000000000033000000000000003000000000",
            INIT_1F => X"0000005800000000000000830000000000000073000000000000005200000000",
            INIT_20 => X"00000037000000000000004e0000000000000043000000000000006f00000000",
            INIT_21 => X"0000002f00000000000000420000000000000042000000000000003a00000000",
            INIT_22 => X"0000007a00000000000000670000000000000032000000000000003100000000",
            INIT_23 => X"00000058000000000000004d000000000000005e000000000000005a00000000",
            INIT_24 => X"00000040000000000000003f0000000000000044000000000000004100000000",
            INIT_25 => X"0000003300000000000000320000000000000040000000000000004300000000",
            INIT_26 => X"00000050000000000000005e000000000000006f000000000000003200000000",
            INIT_27 => X"00000026000000000000002b0000000000000030000000000000003900000000",
            INIT_28 => X"0000003700000000000000320000000000000032000000000000002200000000",
            INIT_29 => X"0000003e000000000000003b000000000000003b000000000000003c00000000",
            INIT_2A => X"00000032000000000000002d000000000000002c000000000000003d00000000",
            INIT_2B => X"00000035000000000000002f0000000000000026000000000000003c00000000",
            INIT_2C => X"0000004400000000000000390000000000000025000000000000002900000000",
            INIT_2D => X"000000260000000000000045000000000000003c000000000000004100000000",
            INIT_2E => X"00000035000000000000003d000000000000003a000000000000002c00000000",
            INIT_2F => X"00000031000000000000003c0000000000000026000000000000003900000000",
            INIT_30 => X"00000043000000000000003a0000000000000040000000000000002d00000000",
            INIT_31 => X"000000360000000000000034000000000000003d000000000000003e00000000",
            INIT_32 => X"0000003c000000000000002e0000000000000035000000000000003700000000",
            INIT_33 => X"000000330000000000000037000000000000003d000000000000003b00000000",
            INIT_34 => X"0000003a000000000000003e000000000000003a000000000000002d00000000",
            INIT_35 => X"0000000000000000000000040000000000000000000000000000003c00000000",
            INIT_36 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000900000000000000050000000000000008000000000000000700000000",
            INIT_38 => X"0000000a00000000000000000000000000000009000000000000000c00000000",
            INIT_39 => X"0000000300000000000000000000000000000008000000000000000000000000",
            INIT_3A => X"0000000700000000000000070000000000000000000000000000000100000000",
            INIT_3B => X"0000000400000000000000040000000000000002000000000000000900000000",
            INIT_3C => X"0000000000000000000000080000000000000000000000000000000100000000",
            INIT_3D => X"000000050000000000000000000000000000000e000000000000000200000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000500000000000000040000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000000e000000000000000800000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000d00000000000000050000000000000011000000000000000000000000",
            INIT_44 => X"0000002e00000000000000000000000000000000000000000000000900000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_47 => X"00000006000000000000000b0000000000000000000000000000000000000000",
            INIT_48 => X"0000002400000000000000450000000000000000000000000000000000000000",
            INIT_49 => X"0000000d00000000000000050000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000000d0000000000000003000000000000000000000000",
            INIT_4C => X"0000000000000000000000590000000000000011000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000007000000000000000700000000",
            INIT_4F => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_50 => X"000000000000000000000045000000000000000b000000000000000600000000",
            INIT_51 => X"0000000e00000000000000000000000000000000000000000000001000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_54 => X"000000000000000000000032000000000000000e000000000000002500000000",
            INIT_55 => X"0000000700000000000000070000000000000000000000000000000f00000000",
            INIT_56 => X"0000001400000000000000000000000000000000000000000000000800000000",
            INIT_57 => X"0000004f00000000000000010000000000000000000000000000000000000000",
            INIT_58 => X"0000002000000000000000000000000000000032000000000000000000000000",
            INIT_59 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_5A => X"00000000000000000000000b000000000000001b000000000000000000000000",
            INIT_5B => X"0000000000000000000000130000000000000069000000000000001600000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_5D => X"0000000300000000000000100000000000000005000000000000000000000000",
            INIT_5E => X"0000002000000000000000150000000000000013000000000000000500000000",
            INIT_5F => X"00000000000000000000002d0000000000000013000000000000002800000000",
            INIT_60 => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_61 => X"000000000000000000000010000000000000000c000000000000000000000000",
            INIT_62 => X"000000040000000000000000000000000000000c000000000000002900000000",
            INIT_63 => X"000000000000000000000012000000000000001c000000000000000100000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_65 => X"0000000000000000000000000000000000000017000000000000000800000000",
            INIT_66 => X"0000000f00000000000000060000000000000000000000000000000100000000",
            INIT_67 => X"0000000300000000000000020000000000000004000000000000000600000000",
            INIT_68 => X"0000000800000000000000000000000000000000000000000000000200000000",
            INIT_69 => X"0000000900000000000000000000000000000005000000000000000c00000000",
            INIT_6A => X"00000000000000000000000c000000000000000b000000000000000d00000000",
            INIT_6B => X"0000000a0000000000000012000000000000000c000000000000000000000000",
            INIT_6C => X"0000001500000000000000010000000000000000000000000000000700000000",
            INIT_6D => X"0000000000000000000000000000000000000005000000000000000100000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000500000000000000050000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "samplegold_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000b00000000000000000000000000000015000000000000001000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000013000000000000002500000000",
            INIT_18 => X"0000001e00000000000000000000000000000000000000000000001300000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_1A => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_20 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000f0000000000000004000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000700000000000000010000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_26 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2F => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_34 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000200000000000000050000000000000004000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_3F => X"00000000000000000000000a0000000000000000000000000000000500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_43 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_45 => X"0000000200000000000000000000000000000008000000000000000000000000",
            INIT_46 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000004000000000000000b00000000",
            INIT_52 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_56 => X"000000000000000000000000000000000000000c000000000000000200000000",
            INIT_57 => X"0000000600000000000000010000000000000000000000000000000000000000",
            INIT_58 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_5B => X"00000000000000000000000c000000000000000f000000000000000000000000",
            INIT_5C => X"0000000300000000000000010000000000000000000000000000000000000000",
            INIT_5D => X"0000000700000000000000050000000000000000000000000000000000000000",
            INIT_5E => X"0000000a00000000000000050000000000000006000000000000000500000000",
            INIT_5F => X"0000000b000000000000000f000000000000000f000000000000000f00000000",
            INIT_60 => X"0000000600000000000000070000000000000008000000000000000800000000",
            INIT_61 => X"0000000500000000000000080000000000000006000000000000000600000000",
            INIT_62 => X"00000015000000000000000a0000000000000006000000000000000600000000",
            INIT_63 => X"0000000e00000000000000150000000000000017000000000000001300000000",
            INIT_64 => X"000000140000000000000012000000000000000e000000000000000b00000000",
            INIT_65 => X"0000000500000000000000040000000000000015000000000000001500000000",
            INIT_66 => X"000000170000000000000013000000000000000b000000000000000900000000",
            INIT_67 => X"00000019000000000000001b000000000000001b000000000000001900000000",
            INIT_68 => X"0000001100000000000000130000000000000017000000000000001600000000",
            INIT_69 => X"0000000e00000000000000060000000000000006000000000000001100000000",
            INIT_6A => X"0000001b00000000000000140000000000000010000000000000001500000000",
            INIT_6B => X"000000170000000000000018000000000000001e000000000000002200000000",
            INIT_6C => X"0000001900000000000000150000000000000014000000000000001600000000",
            INIT_6D => X"00000018000000000000001f0000000000000019000000000000001300000000",
            INIT_6E => X"00000020000000000000001b0000000000000013000000000000001200000000",
            INIT_6F => X"0000001b00000000000000200000000000000021000000000000002300000000",
            INIT_70 => X"0000001300000000000000260000000000000025000000000000001d00000000",
            INIT_71 => X"0000001200000000000000160000000000000012000000000000001100000000",
            INIT_72 => X"0000001d00000000000000180000000000000016000000000000001600000000",
            INIT_73 => X"0000001e00000000000000170000000000000022000000000000002200000000",
            INIT_74 => X"0000000c000000000000000a0000000000000022000000000000002600000000",
            INIT_75 => X"0000000e0000000000000014000000000000001b000000000000001100000000",
            INIT_76 => X"0000001d0000000000000019000000000000001a000000000000001900000000",
            INIT_77 => X"000000180000000000000018000000000000001a000000000000002000000000",
            INIT_78 => X"000000180000000000000013000000000000000d000000000000001400000000",
            INIT_79 => X"00000021000000000000001d0000000000000023000000000000001c00000000",
            INIT_7A => X"0000001e000000000000001a000000000000001a000000000000001f00000000",
            INIT_7B => X"0000001b00000000000000130000000000000014000000000000001b00000000",
            INIT_7C => X"00000026000000000000001f0000000000000014000000000000001200000000",
            INIT_7D => X"0000002400000000000000210000000000000026000000000000002100000000",
            INIT_7E => X"0000001b000000000000001c0000000000000015000000000000001500000000",
            INIT_7F => X"00000023000000000000001d0000000000000019000000000000001500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "samplegold_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000013000000000000001d000000000000001c000000000000002200000000",
            INIT_01 => X"000000160000000000000022000000000000001d000000000000001f00000000",
            INIT_02 => X"00000014000000000000001d000000000000001c000000000000001500000000",
            INIT_03 => X"0000001800000000000000150000000000000020000000000000001700000000",
            INIT_04 => X"00000011000000000000000d0000000000000007000000000000000b00000000",
            INIT_05 => X"00000018000000000000001a0000000000000016000000000000001200000000",
            INIT_06 => X"000000200000000000000018000000000000001a000000000000001a00000000",
            INIT_07 => X"0000000f00000000000000000000000000000000000000000000002800000000",
            INIT_08 => X"00000010000000000000000d0000000000000011000000000000001200000000",
            INIT_09 => X"00000019000000000000000f000000000000000d000000000000001500000000",
            INIT_0A => X"000000280000000000000023000000000000001f000000000000001b00000000",
            INIT_0B => X"00000015000000000000000a0000000000000005000000000000000700000000",
            INIT_0C => X"000000180000000000000013000000000000001d000000000000001f00000000",
            INIT_0D => X"0000001800000000000000170000000000000011000000000000001700000000",
            INIT_0E => X"0000000d00000000000000250000000000000026000000000000002100000000",
            INIT_0F => X"0000001800000000000000170000000000000017000000000000001500000000",
            INIT_10 => X"0000001c000000000000001c000000000000001e000000000000002000000000",
            INIT_11 => X"000000180000000000000011000000000000000d000000000000001000000000",
            INIT_12 => X"0000001600000000000000150000000000000025000000000000002400000000",
            INIT_13 => X"0000002400000000000000230000000000000022000000000000001b00000000",
            INIT_14 => X"0000002400000000000000280000000000000025000000000000002300000000",
            INIT_15 => X"000000260000000000000020000000000000001e000000000000001f00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000013000000000000000f000000000000000b000000000000000400000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000020000000000000004000000000000000300000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "samplegold_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000010000000000000000200000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000002700000000000000290000000000000023000000000000001200000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000d00000000000000190000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_12 => X"0000000900000000000000230000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000004300000000000000030000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000050000000000000029000000000000004c00000000",
            INIT_17 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000040000000000000010000000000000000e00000000",
            INIT_1A => X"00000007000000000000000f000000000000000d000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_22 => X"00000000000000000000000d0000000000000036000000000000004900000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000500000000000000040000000000000000000000000000000000000000",
            INIT_25 => X"00000014000000000000004b0000000000000059000000000000001d00000000",
            INIT_26 => X"0000000000000000000000000000000000000002000000000000001800000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002700000000000000560000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000800000000000000020000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_34 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000e00000000000000140000000000000010000000000000001100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001600000000000000160000000000000021000000000000001c00000000",
            INIT_41 => X"0000001200000000000000130000000000000013000000000000001300000000",
            INIT_42 => X"0000001100000000000000150000000000000017000000000000001400000000",
            INIT_43 => X"0000002400000000000000150000000000000015000000000000001000000000",
            INIT_44 => X"0000001a00000000000000280000000000000029000000000000002f00000000",
            INIT_45 => X"000000180000000000000019000000000000001a000000000000001900000000",
            INIT_46 => X"0000001300000000000000130000000000000012000000000000001600000000",
            INIT_47 => X"0000003b0000000000000030000000000000001e000000000000000d00000000",
            INIT_48 => X"0000001e000000000000002c000000000000003d000000000000004100000000",
            INIT_49 => X"0000000e00000000000000110000000000000016000000000000001700000000",
            INIT_4A => X"0000001000000000000000180000000000000016000000000000000e00000000",
            INIT_4B => X"000000430000000000000042000000000000003e000000000000002600000000",
            INIT_4C => X"00000025000000000000002e000000000000003a000000000000004300000000",
            INIT_4D => X"0000001500000000000000100000000000000012000000000000001d00000000",
            INIT_4E => X"0000001700000000000000060000000000000018000000000000001b00000000",
            INIT_4F => X"00000039000000000000003a0000000000000040000000000000003900000000",
            INIT_50 => X"0000003000000000000000400000000000000040000000000000004400000000",
            INIT_51 => X"0000000e00000000000000170000000000000014000000000000001e00000000",
            INIT_52 => X"0000003200000000000000100000000000000000000000000000000a00000000",
            INIT_53 => X"0000004200000000000000390000000000000035000000000000004500000000",
            INIT_54 => X"0000002800000000000000420000000000000044000000000000004200000000",
            INIT_55 => X"0000000700000000000000090000000000000011000000000000001600000000",
            INIT_56 => X"0000003300000000000000250000000000000000000000000000000800000000",
            INIT_57 => X"0000003900000000000000400000000000000040000000000000003000000000",
            INIT_58 => X"0000001c000000000000002c0000000000000046000000000000003f00000000",
            INIT_59 => X"00000008000000000000000e0000000000000010000000000000000c00000000",
            INIT_5A => X"0000002c000000000000002f000000000000000d000000000000000900000000",
            INIT_5B => X"0000003f0000000000000034000000000000003e000000000000003e00000000",
            INIT_5C => X"0000001400000000000000260000000000000039000000000000004400000000",
            INIT_5D => X"00000002000000000000000e0000000000000015000000000000001300000000",
            INIT_5E => X"000000310000000000000025000000000000000b000000000000001200000000",
            INIT_5F => X"00000041000000000000003d0000000000000037000000000000004000000000",
            INIT_60 => X"0000000a00000000000000110000000000000023000000000000004200000000",
            INIT_61 => X"0000002100000000000000000000000000000000000000000000000100000000",
            INIT_62 => X"00000040000000000000002b000000000000002f000000000000000e00000000",
            INIT_63 => X"0000003f000000000000003e000000000000003b000000000000003b00000000",
            INIT_64 => X"0000000000000000000000000000000000000014000000000000001d00000000",
            INIT_65 => X"0000002b00000000000000240000000000000019000000000000000000000000",
            INIT_66 => X"00000039000000000000003a000000000000002e000000000000003300000000",
            INIT_67 => X"000000200000000000000035000000000000003c000000000000003700000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_69 => X"00000037000000000000003c000000000000001e000000000000001400000000",
            INIT_6A => X"00000037000000000000003e000000000000003d000000000000002300000000",
            INIT_6B => X"0000000f00000000000000260000000000000028000000000000003600000000",
            INIT_6C => X"000000110000000000000010000000000000000e000000000000000500000000",
            INIT_6D => X"00000024000000000000002f000000000000001e000000000000001100000000",
            INIT_6E => X"0000003200000000000000300000000000000042000000000000003c00000000",
            INIT_6F => X"00000014000000000000001e0000000000000023000000000000002700000000",
            INIT_70 => X"0000001700000000000000130000000000000014000000000000001400000000",
            INIT_71 => X"0000002e00000000000000270000000000000026000000000000001c00000000",
            INIT_72 => X"0000002c00000000000000330000000000000031000000000000003200000000",
            INIT_73 => X"0000001400000000000000110000000000000020000000000000001f00000000",
            INIT_74 => X"00000020000000000000001e0000000000000019000000000000001900000000",
            INIT_75 => X"000000240000000000000020000000000000001c000000000000001c00000000",
            INIT_76 => X"0000001e00000000000000200000000000000027000000000000002b00000000",
            INIT_77 => X"00000007000000000000000c000000000000000c000000000000001b00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_79 => X"0000000600000000000000050000000000000006000000000000000400000000",
            INIT_7A => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_7B => X"000000000000000000000009000000000000000b000000000000000c00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000000f000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "samplegold_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000200000000000000050000000000000000000000000000000100000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000001d000000000000000f000000000000000800000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000008000000000000001200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000100000000000000070000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000026000000000000002f000000000000000c000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000000000000d0000000000000030000000000000003200000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000003c00000000000000540000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000007000000000000000900000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000600000000000000170000000000000014000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000700000000000000060000000000000001000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000b000000000000000f0000000000000003000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_3E => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000a000000000000000b0000000000000001000000000000000000000000",
            INIT_41 => X"0000000700000000000000030000000000000000000000000000000800000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"00000008000000000000000a0000000000000002000000000000000000000000",
            INIT_45 => X"0000000e00000000000000120000000000000011000000000000000800000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000000000000000000000e000000000000000900000000",
            INIT_48 => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000090000000000000010000000000000000a00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_4C => X"0000000100000000000000040000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000004000000000000000200000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_50 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000001e000000000000000b0000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000d00000000000000050000000000000000000000000000000500000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000018000000000000000f000000000000000600000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000400000000000000000000000000000000000000000000000400000000",
            INIT_5B => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000011000000000000001f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_5F => X"00000020000000000000000a0000000000000000000000000000000000000000",
            INIT_60 => X"0000000600000000000000000000000000000000000000000000001b00000000",
            INIT_61 => X"00000006000000000000000c0000000000000015000000000000001100000000",
            INIT_62 => X"00000001000000000000000d000000000000000d000000000000000d00000000",
            INIT_63 => X"000000250000000000000023000000000000000e000000000000000000000000",
            INIT_64 => X"0000001d00000000000000190000000000000015000000000000000b00000000",
            INIT_65 => X"0000001d00000000000000140000000000000019000000000000002500000000",
            INIT_66 => X"0000001900000000000000170000000000000018000000000000002000000000",
            INIT_67 => X"0000000a0000000000000028000000000000002a000000000000001b00000000",
            INIT_68 => X"00000016000000000000000d000000000000000a000000000000000b00000000",
            INIT_69 => X"0000000c000000000000000d0000000000000015000000000000001a00000000",
            INIT_6A => X"0000000b000000000000000b000000000000000b000000000000000b00000000",
            INIT_6B => X"00000009000000000000000a000000000000000c000000000000000a00000000",
            INIT_6C => X"00000028000000000000001c0000000000000023000000000000000600000000",
            INIT_6D => X"0000000e0000000000000015000000000000001f000000000000002500000000",
            INIT_6E => X"0000001100000000000000160000000000000015000000000000001300000000",
            INIT_6F => X"0000000c0000000000000008000000000000000a000000000000001100000000",
            INIT_70 => X"0000003200000000000000300000000000000027000000000000001a00000000",
            INIT_71 => X"000000170000000000000014000000000000002c000000000000003900000000",
            INIT_72 => X"00000010000000000000000d0000000000000015000000000000001400000000",
            INIT_73 => X"0000002a00000000000000070000000000000009000000000000000d00000000",
            INIT_74 => X"0000003e0000000000000037000000000000002b000000000000002d00000000",
            INIT_75 => X"0000001900000000000000210000000000000026000000000000003300000000",
            INIT_76 => X"0000001500000000000000190000000000000015000000000000001200000000",
            INIT_77 => X"0000003000000000000000350000000000000000000000000000001600000000",
            INIT_78 => X"0000003b000000000000003d000000000000002a000000000000002500000000",
            INIT_79 => X"0000001900000000000000280000000000000036000000000000003b00000000",
            INIT_7A => X"0000000e000000000000000e0000000000000022000000000000002300000000",
            INIT_7B => X"000000270000000000000022000000000000003c000000000000000000000000",
            INIT_7C => X"0000004000000000000000310000000000000036000000000000002e00000000",
            INIT_7D => X"0000001e00000000000000290000000000000032000000000000003a00000000",
            INIT_7E => X"0000000f000000000000000e000000000000000b000000000000001b00000000",
            INIT_7F => X"0000003100000000000000280000000000000023000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "samplegold_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003800000000000000340000000000000028000000000000003600000000",
            INIT_01 => X"0000001000000000000000120000000000000022000000000000003f00000000",
            INIT_02 => X"0000002c000000000000000f0000000000000013000000000000001000000000",
            INIT_03 => X"0000003a000000000000002b0000000000000030000000000000000e00000000",
            INIT_04 => X"00000038000000000000003a000000000000002f000000000000002b00000000",
            INIT_05 => X"00000012000000000000001f000000000000001b000000000000002100000000",
            INIT_06 => X"0000000d00000000000000350000000000000015000000000000001200000000",
            INIT_07 => X"0000002c000000000000003d000000000000001e000000000000000d00000000",
            INIT_08 => X"0000002e00000000000000370000000000000037000000000000002e00000000",
            INIT_09 => X"0000000f00000000000000190000000000000017000000000000002a00000000",
            INIT_0A => X"00000005000000000000001a0000000000000009000000000000001b00000000",
            INIT_0B => X"00000031000000000000002f000000000000003e000000000000002800000000",
            INIT_0C => X"000000210000000000000032000000000000003a000000000000003500000000",
            INIT_0D => X"0000002100000000000000040000000000000009000000000000001e00000000",
            INIT_0E => X"0000002700000000000000260000000000000029000000000000000f00000000",
            INIT_0F => X"0000002f00000000000000320000000000000031000000000000003800000000",
            INIT_10 => X"00000021000000000000001d0000000000000036000000000000003800000000",
            INIT_11 => X"0000001100000000000000270000000000000000000000000000000000000000",
            INIT_12 => X"0000001d00000000000000230000000000000032000000000000001e00000000",
            INIT_13 => X"0000002c000000000000002b0000000000000031000000000000002700000000",
            INIT_14 => X"00000016000000000000001e0000000000000024000000000000003700000000",
            INIT_15 => X"00000023000000000000001b0000000000000010000000000000000b00000000",
            INIT_16 => X"0000002d0000000000000023000000000000001d000000000000002600000000",
            INIT_17 => X"0000002d0000000000000030000000000000001d000000000000003300000000",
            INIT_18 => X"0000001a00000000000000160000000000000021000000000000002700000000",
            INIT_19 => X"0000001b0000000000000022000000000000001a000000000000001800000000",
            INIT_1A => X"000000280000000000000032000000000000002b000000000000002900000000",
            INIT_1B => X"0000002a0000000000000029000000000000002e000000000000002100000000",
            INIT_1C => X"0000002200000000000000190000000000000016000000000000002400000000",
            INIT_1D => X"00000025000000000000001b0000000000000027000000000000002400000000",
            INIT_1E => X"0000002c0000000000000027000000000000002c000000000000002a00000000",
            INIT_1F => X"0000001f0000000000000027000000000000002a000000000000002c00000000",
            INIT_20 => X"0000001900000000000000150000000000000000000000000000000000000000",
            INIT_21 => X"0000000c0000000000000012000000000000000e000000000000001800000000",
            INIT_22 => X"000000180000000000000003000000000000001b000000000000000f00000000",
            INIT_23 => X"0000000000000000000000190000000000000018000000000000001800000000",
            INIT_24 => X"00000027000000000000001b000000000000000e000000000000000400000000",
            INIT_25 => X"0000002e00000000000000250000000000000022000000000000002200000000",
            INIT_26 => X"00000026000000000000002c000000000000000a000000000000002500000000",
            INIT_27 => X"0000000600000000000000000000000000000022000000000000002300000000",
            INIT_28 => X"000000450000000000000038000000000000001c000000000000000000000000",
            INIT_29 => X"0000001700000000000000330000000000000029000000000000002c00000000",
            INIT_2A => X"0000002d00000000000000340000000000000032000000000000002700000000",
            INIT_2B => X"0000000100000000000000000000000000000000000000000000002b00000000",
            INIT_2C => X"00000025000000000000003a000000000000003d000000000000002d00000000",
            INIT_2D => X"0000004000000000000000210000000000000014000000000000002000000000",
            INIT_2E => X"0000003d00000000000000530000000000000049000000000000003000000000",
            INIT_2F => X"0000002a000000000000002d0000000000000021000000000000001700000000",
            INIT_30 => X"00000038000000000000003f0000000000000044000000000000002a00000000",
            INIT_31 => X"0000003b000000000000002f0000000000000029000000000000002000000000",
            INIT_32 => X"000000300000000000000030000000000000003e000000000000004b00000000",
            INIT_33 => X"0000003000000000000000270000000000000036000000000000003300000000",
            INIT_34 => X"0000002100000000000000250000000000000046000000000000004600000000",
            INIT_35 => X"0000004900000000000000360000000000000039000000000000002800000000",
            INIT_36 => X"0000002e000000000000002f0000000000000023000000000000003900000000",
            INIT_37 => X"0000002e0000000000000038000000000000002a000000000000003500000000",
            INIT_38 => X"0000003400000000000000320000000000000027000000000000003600000000",
            INIT_39 => X"0000003c0000000000000048000000000000003b000000000000003100000000",
            INIT_3A => X"0000003500000000000000310000000000000031000000000000002800000000",
            INIT_3B => X"0000003200000000000000480000000000000039000000000000001b00000000",
            INIT_3C => X"00000045000000000000002c0000000000000033000000000000004200000000",
            INIT_3D => X"0000003d0000000000000051000000000000004b000000000000003c00000000",
            INIT_3E => X"0000003100000000000000210000000000000027000000000000003500000000",
            INIT_3F => X"00000036000000000000003d000000000000003a000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002c00000000000000280000000000000034000000000000001c00000000",
            INIT_41 => X"0000002c0000000000000032000000000000003e000000000000002500000000",
            INIT_42 => X"0000004200000000000000420000000000000038000000000000002700000000",
            INIT_43 => X"000000310000000000000037000000000000004d000000000000005100000000",
            INIT_44 => X"00000019000000000000001b0000000000000031000000000000001f00000000",
            INIT_45 => X"0000003b00000000000000360000000000000033000000000000002300000000",
            INIT_46 => X"00000045000000000000003a000000000000003b000000000000003300000000",
            INIT_47 => X"0000003a000000000000003b0000000000000048000000000000003800000000",
            INIT_48 => X"00000029000000000000002d000000000000001a000000000000001d00000000",
            INIT_49 => X"000000310000000000000038000000000000003a000000000000002200000000",
            INIT_4A => X"00000032000000000000003d000000000000004b000000000000004700000000",
            INIT_4B => X"00000017000000000000002a000000000000003e000000000000003b00000000",
            INIT_4C => X"00000021000000000000002b000000000000002c000000000000002b00000000",
            INIT_4D => X"0000004a000000000000002f000000000000002c000000000000003800000000",
            INIT_4E => X"0000003c00000000000000330000000000000032000000000000004f00000000",
            INIT_4F => X"00000027000000000000001f0000000000000029000000000000003800000000",
            INIT_50 => X"0000003700000000000000220000000000000027000000000000002e00000000",
            INIT_51 => X"0000003400000000000000410000000000000023000000000000002900000000",
            INIT_52 => X"0000002900000000000000300000000000000036000000000000002d00000000",
            INIT_53 => X"000000200000000000000021000000000000001a000000000000001c00000000",
            INIT_54 => X"000000220000000000000033000000000000001e000000000000001900000000",
            INIT_55 => X"0000003a00000000000000420000000000000042000000000000001e00000000",
            INIT_56 => X"0000001200000000000000220000000000000024000000000000003200000000",
            INIT_57 => X"000000190000000000000018000000000000001c000000000000001b00000000",
            INIT_58 => X"00000008000000000000005e0000000000000000000000000000002300000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000004800000000000000000000000000000000000000000000000300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_5C => X"0000000300000000000000190000000000000034000000000000000200000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000620000000000000000000000000000000000000000",
            INIT_5F => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"00000011000000000000000d0000000000000047000000000000001000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000024000000000000000100000000",
            INIT_63 => X"0000005700000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000100000000000000000000000000000005200000000",
            INIT_65 => X"0000003400000000000000060000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_67 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_69 => X"0000000d000000000000001c0000000000000002000000000000000000000000",
            INIT_6A => X"0000000200000000000000000000000000000000000000000000001100000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_6D => X"000000160000000000000009000000000000001b000000000000000400000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000000f0000000000000000000000000000000700000000",
            INIT_71 => X"0000000000000000000000150000000000000010000000000000000400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_74 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_78 => X"0000000000000000000000000000000000000028000000000000000000000000",
            INIT_79 => X"0000000f0000000000000000000000000000001d000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_7E => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000008000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "samplegold_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_05 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_0B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_11 => X"0000001e000000000000000b0000000000000016000000000000002000000000",
            INIT_12 => X"0000000000000000000000090000000000000019000000000000001f00000000",
            INIT_13 => X"00000020000000000000001e0000000000000007000000000000000000000000",
            INIT_14 => X"0000001d00000000000000000000000000000000000000000000002400000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_16 => X"0000000000000000000000000000000000000002000000000000000300000000",
            INIT_17 => X"0000001b0000000000000016000000000000000e000000000000000000000000",
            INIT_18 => X"00000011000000000000000a0000000000000000000000000000000000000000",
            INIT_19 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000400000000000000030000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000700000000000000060000000000000007000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000500000000000000000000000000000000000000000000000a00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000100000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_41 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000040000000000000008000000000000000700000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_46 => X"0000000800000000000000010000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000006000000000000000700000000",
            INIT_48 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"00000104000000000000010f00000000000000f5000000000000002e00000000",
            INIT_4A => X"00000110000000000000010b000000000000011100000000000000fc00000000",
            INIT_4B => X"0000013d0000000000000139000000000000007f00000000000000d700000000",
            INIT_4C => X"0000002500000000000000170000000000000139000000000000013c00000000",
            INIT_4D => X"00000120000000000000012200000000000000f100000000000000c300000000",
            INIT_4E => X"000000f80000000000000143000000000000012a000000000000010f00000000",
            INIT_4F => X"00000154000000000000015f000000000000016600000000000000c400000000",
            INIT_50 => X"0000007c0000000000000022000000000000001c000000000000014f00000000",
            INIT_51 => X"000000e70000000000000151000000000000013200000000000000fa00000000",
            INIT_52 => X"0000013900000000000000d200000000000000fd00000000000000e700000000",
            INIT_53 => X"0000017000000000000001710000000000000175000000000000015d00000000",
            INIT_54 => X"0000013100000000000000fe000000000000004300000000000000a200000000",
            INIT_55 => X"000000f3000000000000011b0000000000000152000000000000011f00000000",
            INIT_56 => X"0000015a000000000000015900000000000000df00000000000000c200000000",
            INIT_57 => X"0000013a000000000000016800000000000001a300000000000001a500000000",
            INIT_58 => X"00000103000000000000012c0000000000000159000000000000012e00000000",
            INIT_59 => X"000000c800000000000001140000000000000151000000000000015200000000",
            INIT_5A => X"000001ac0000000000000183000000000000013800000000000000e200000000",
            INIT_5B => X"000001560000000000000160000000000000014b000000000000018b00000000",
            INIT_5C => X"00000152000000000000012d0000000000000128000000000000016500000000",
            INIT_5D => X"000000ef00000000000000ea00000000000000e4000000000000014200000000",
            INIT_5E => X"0000019800000000000001b90000000000000176000000000000013600000000",
            INIT_5F => X"0000015500000000000001530000000000000168000000000000014d00000000",
            INIT_60 => X"0000013700000000000001130000000000000135000000000000012200000000",
            INIT_61 => X"000001290000000000000114000000000000013100000000000000ee00000000",
            INIT_62 => X"0000018000000000000001b000000000000001b6000000000000017b00000000",
            INIT_63 => X"00000112000000000000013f0000000000000149000000000000016b00000000",
            INIT_64 => X"000001270000000000000129000000000000014d000000000000016500000000",
            INIT_65 => X"0000013c00000000000001430000000000000123000000000000010900000000",
            INIT_66 => X"00000173000000000000017a00000000000001bb000000000000017900000000",
            INIT_67 => X"000001610000000000000145000000000000012e000000000000012600000000",
            INIT_68 => X"000000eb000000000000013c000000000000015f000000000000017400000000",
            INIT_69 => X"000000fc00000000000001040000000000000127000000000000011600000000",
            INIT_6A => X"0000014800000000000001790000000000000149000000000000013f00000000",
            INIT_6B => X"000001700000000000000162000000000000015f000000000000015b00000000",
            INIT_6C => X"0000010700000000000001380000000000000159000000000000016400000000",
            INIT_6D => X"0000012100000000000000f600000000000000f5000000000000012f00000000",
            INIT_6E => X"00000146000000000000016b0000000000000181000000000000011c00000000",
            INIT_6F => X"00000134000000000000016b000000000000016f000000000000017200000000",
            INIT_70 => X"000000df0000000000000143000000000000015b000000000000015800000000",
            INIT_71 => X"000000f900000000000001140000000000000121000000000000010700000000",
            INIT_72 => X"000001820000000000000140000000000000016b000000000000017c00000000",
            INIT_73 => X"00000155000000000000014b0000000000000154000000000000018a00000000",
            INIT_74 => X"0000011600000000000000e40000000000000118000000000000015900000000",
            INIT_75 => X"0000017600000000000000f30000000000000119000000000000011d00000000",
            INIT_76 => X"0000017b0000000000000179000000000000013f000000000000015b00000000",
            INIT_77 => X"000001390000000000000149000000000000013b00000000000000f100000000",
            INIT_78 => X"0000010800000000000000fd00000000000000e900000000000000fa00000000",
            INIT_79 => X"00000149000000000000016f00000000000000f800000000000000f000000000",
            INIT_7A => X"000001210000000000000168000000000000016c000000000000012200000000",
            INIT_7B => X"000000cb00000000000000ff0000000000000118000000000000014400000000",
            INIT_7C => X"000000cc00000000000000df00000000000000e700000000000000e000000000",
            INIT_7D => X"00000110000000000000012c000000000000014000000000000000f600000000",
            INIT_7E => X"000001150000000000000156000000000000016c000000000000015000000000",
            INIT_7F => X"000000d500000000000000a800000000000000de00000000000000ea00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "samplegold_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ed00000000000000de00000000000000d900000000000000e100000000",
            INIT_01 => X"0000005d00000000000000680000000000000000000000000000000000000000",
            INIT_02 => X"0000006000000000000000660000000000000064000000000000005900000000",
            INIT_03 => X"0000006300000000000000190000000000000036000000000000005400000000",
            INIT_04 => X"0000000000000000000000760000000000000072000000000000007200000000",
            INIT_05 => X"000000440000000000000048000000000000005c000000000000000000000000",
            INIT_06 => X"000000620000000000000058000000000000005c000000000000004b00000000",
            INIT_07 => X"0000007000000000000000670000000000000017000000000000005300000000",
            INIT_08 => X"0000000000000000000000000000000000000077000000000000007400000000",
            INIT_09 => X"000000530000000000000046000000000000003f000000000000003000000000",
            INIT_0A => X"00000039000000000000005e0000000000000058000000000000004100000000",
            INIT_0B => X"0000006700000000000000670000000000000060000000000000003b00000000",
            INIT_0C => X"0000002e00000000000000000000000000000001000000000000006700000000",
            INIT_0D => X"000000360000000000000057000000000000003f000000000000005900000000",
            INIT_0E => X"0000005c00000000000000270000000000000033000000000000003800000000",
            INIT_0F => X"0000006200000000000000710000000000000065000000000000005000000000",
            INIT_10 => X"00000055000000000000005c0000000000000031000000000000005d00000000",
            INIT_11 => X"0000004b000000000000005e0000000000000052000000000000003200000000",
            INIT_12 => X"0000005500000000000000540000000000000029000000000000003400000000",
            INIT_13 => X"0000006300000000000000590000000000000075000000000000007200000000",
            INIT_14 => X"0000004200000000000000520000000000000069000000000000005800000000",
            INIT_15 => X"00000030000000000000003a0000000000000056000000000000005100000000",
            INIT_16 => X"00000073000000000000005e0000000000000047000000000000002600000000",
            INIT_17 => X"0000005c0000000000000066000000000000005d000000000000007600000000",
            INIT_18 => X"0000003d000000000000003f0000000000000059000000000000006c00000000",
            INIT_19 => X"0000003400000000000000450000000000000031000000000000005400000000",
            INIT_1A => X"0000007500000000000000720000000000000059000000000000004400000000",
            INIT_1B => X"0000006b000000000000005d000000000000006c000000000000005a00000000",
            INIT_1C => X"0000004e00000000000000440000000000000059000000000000005100000000",
            INIT_1D => X"000000550000000000000043000000000000004d000000000000003c00000000",
            INIT_1E => X"00000064000000000000007e000000000000006a000000000000007000000000",
            INIT_1F => X"000000460000000000000060000000000000004d000000000000006c00000000",
            INIT_20 => X"0000005800000000000000410000000000000049000000000000005700000000",
            INIT_21 => X"0000003f00000000000000610000000000000048000000000000003b00000000",
            INIT_22 => X"0000006b00000000000000600000000000000077000000000000004f00000000",
            INIT_23 => X"00000052000000000000005a0000000000000057000000000000004b00000000",
            INIT_24 => X"0000003e000000000000004c000000000000005b000000000000006400000000",
            INIT_25 => X"0000003e0000000000000057000000000000005f000000000000004f00000000",
            INIT_26 => X"0000005c0000000000000067000000000000004c000000000000005800000000",
            INIT_27 => X"0000005a000000000000005b0000000000000057000000000000005100000000",
            INIT_28 => X"0000006200000000000000690000000000000057000000000000004e00000000",
            INIT_29 => X"00000057000000000000004f000000000000004a000000000000004a00000000",
            INIT_2A => X"0000004700000000000000690000000000000065000000000000005300000000",
            INIT_2B => X"0000005100000000000000650000000000000068000000000000006100000000",
            INIT_2C => X"0000003e000000000000005e0000000000000061000000000000005700000000",
            INIT_2D => X"0000004700000000000000550000000000000055000000000000005000000000",
            INIT_2E => X"0000005a0000000000000048000000000000006c000000000000006700000000",
            INIT_2F => X"0000006100000000000000660000000000000045000000000000007000000000",
            INIT_30 => X"0000004c00000000000000460000000000000055000000000000006700000000",
            INIT_31 => X"000000690000000000000049000000000000004f000000000000005500000000",
            INIT_32 => X"0000006700000000000000590000000000000043000000000000006800000000",
            INIT_33 => X"0000005d000000000000005c0000000000000063000000000000004700000000",
            INIT_34 => X"0000004900000000000000450000000000000044000000000000004100000000",
            INIT_35 => X"000000620000000000000062000000000000004e000000000000003900000000",
            INIT_36 => X"00000066000000000000005d0000000000000050000000000000003f00000000",
            INIT_37 => X"0000003400000000000000500000000000000052000000000000006300000000",
            INIT_38 => X"00000041000000000000003f0000000000000047000000000000003f00000000",
            INIT_39 => X"0000000000000000000000000000000000000006000000000000004700000000",
            INIT_3A => X"0000000100000000000000000000000000000002000000000000000a00000000",
            INIT_3B => X"000000000000000000000045000000000000001d000000000000000000000000",
            INIT_3C => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_3E => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_3F => X"000000000000000000000000000000000000005e000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000300000000000000060000000000000002000000000000000400000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000800000000000000000000000000000002000000000000004a00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"00000000000000000000003f0000000000000001000000000000000000000000",
            INIT_45 => X"000000250000000000000000000000000000001f000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000001c000000000000002700000000",
            INIT_47 => X"0000001600000000000000010000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_49 => X"0000001b00000000000000000000000000000000000000000000003d00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_4B => X"0000000000000000000000360000000000000002000000000000000000000000",
            INIT_4C => X"0000002500000000000000080000000000000000000000000000000600000000",
            INIT_4D => X"0000001d00000000000000290000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000700000000000000000000000000000034000000000000000100000000",
            INIT_50 => X"0000000800000000000000000000000000000024000000000000000000000000",
            INIT_51 => X"0000001100000000000000000000000000000026000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000140000000000000018000000000000001500000000",
            INIT_54 => X"0000000100000000000000140000000000000000000000000000004800000000",
            INIT_55 => X"0000000000000000000000000000000000000010000000000000001000000000",
            INIT_56 => X"0000000e00000000000000000000000000000000000000000000000900000000",
            INIT_57 => X"0000000b0000000000000000000000000000002d000000000000000000000000",
            INIT_58 => X"0000001300000000000000000000000000000003000000000000000000000000",
            INIT_59 => X"0000000000000000000000140000000000000000000000000000003a00000000",
            INIT_5A => X"0000000000000000000000040000000000000000000000000000002300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_5C => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"00000000000000000000001a0000000000000000000000000000002600000000",
            INIT_5E => X"0000000400000000000000000000000000000006000000000000000000000000",
            INIT_5F => X"0000000000000000000000010000000000000000000000000000001f00000000",
            INIT_60 => X"0000001b00000000000000000000000000000000000000000000002b00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_62 => X"0000002a00000000000000000000000000000002000000000000001800000000",
            INIT_63 => X"00000016000000000000000d0000000000000000000000000000000000000000",
            INIT_64 => X"0000003d00000000000000110000000000000000000000000000000000000000",
            INIT_65 => X"0000001700000000000000000000000000000001000000000000000000000000",
            INIT_66 => X"0000000000000000000000190000000000000006000000000000001800000000",
            INIT_67 => X"0000000000000000000000000000000000000035000000000000000000000000",
            INIT_68 => X"00000000000000000000001f000000000000001c000000000000000300000000",
            INIT_69 => X"0000000800000000000000020000000000000000000000000000000400000000",
            INIT_6A => X"000000000000000000000000000000000000001b000000000000000f00000000",
            INIT_6B => X"00000008000000000000000f0000000000000000000000000000002c00000000",
            INIT_6C => X"000000020000000000000000000000000000000c000000000000001900000000",
            INIT_6D => X"0000000d00000000000000000000000000000000000000000000001800000000",
            INIT_6E => X"0000001000000000000000000000000000000000000000000000000d00000000",
            INIT_6F => X"0000002300000000000000000000000000000021000000000000001900000000",
            INIT_70 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "samplegold_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000017000000000000001a0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000001e000000000000005100000000",
            INIT_2B => X"0000000000000000000000080000000000000000000000000000000b00000000",
            INIT_2C => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_2D => X"0000003000000000000000040000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000040000000000000013000000000000003700000000",
            INIT_2F => X"0000000000000000000000000000000000000008000000000000000a00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_31 => X"0000005700000000000000120000000000000001000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000022000000000000000900000000",
            INIT_33 => X"0000001500000000000000180000000000000000000000000000001000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_35 => X"0000000000000000000000220000000000000028000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_37 => X"0000001e0000000000000000000000000000002e000000000000000400000000",
            INIT_38 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_39 => X"0000002f00000000000000000000000000000000000000000000000a00000000",
            INIT_3A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000150000000000000013000000000000001e00000000",
            INIT_3C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_3D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_3E => X"0000001600000000000000030000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000023000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000060000000000000000000000000000001700000000",
            INIT_42 => X"0000000a00000000000000070000000000000000000000000000001100000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_44 => X"0000004500000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000b00000000000000000000000000000000000000000000001400000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_48 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_49 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000090000000000000006000000000000000000000000",
            INIT_4F => X"0000001400000000000000000000000000000000000000000000000700000000",
            INIT_50 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_53 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_57 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000012000000000000000100000000",
            INIT_59 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_5B => X"0000000000000000000000000000000000000006000000000000001100000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000001300000000000000000000000000000000000000000000000800000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_60 => X"0000000000000000000000160000000000000000000000000000000200000000",
            INIT_61 => X"0000000200000000000000030000000000000000000000000000000200000000",
            INIT_62 => X"0000002700000000000000290000000000000008000000000000000500000000",
            INIT_63 => X"00000029000000000000002d0000000000000027000000000000002200000000",
            INIT_64 => X"0000002f0000000000000010000000000000001f000000000000002600000000",
            INIT_65 => X"0000000500000000000000370000000000000036000000000000003600000000",
            INIT_66 => X"0000001b000000000000001e000000000000001c000000000000000500000000",
            INIT_67 => X"000000260000000000000024000000000000001e000000000000001c00000000",
            INIT_68 => X"0000002c0000000000000026000000000000001b000000000000002500000000",
            INIT_69 => X"0000000500000000000000070000000000000032000000000000003000000000",
            INIT_6A => X"0000001a00000000000000170000000000000020000000000000001100000000",
            INIT_6B => X"0000001400000000000000110000000000000012000000000000001100000000",
            INIT_6C => X"00000020000000000000001d0000000000000016000000000000001900000000",
            INIT_6D => X"00000027000000000000001a0000000000000024000000000000002400000000",
            INIT_6E => X"00000021000000000000001b000000000000000f000000000000001d00000000",
            INIT_6F => X"0000001a00000000000000120000000000000015000000000000001b00000000",
            INIT_70 => X"0000001800000000000000210000000000000023000000000000001800000000",
            INIT_71 => X"0000001d00000000000000210000000000000023000000000000002800000000",
            INIT_72 => X"00000018000000000000001c0000000000000013000000000000001100000000",
            INIT_73 => X"000000180000000000000019000000000000000f000000000000001100000000",
            INIT_74 => X"0000002100000000000000190000000000000023000000000000002100000000",
            INIT_75 => X"000000180000000000000020000000000000001e000000000000001e00000000",
            INIT_76 => X"0000001500000000000000130000000000000015000000000000001500000000",
            INIT_77 => X"0000001d00000000000000140000000000000016000000000000001000000000",
            INIT_78 => X"000000200000000000000020000000000000001d000000000000002300000000",
            INIT_79 => X"0000000f0000000000000013000000000000001d000000000000002300000000",
            INIT_7A => X"0000001000000000000000190000000000000014000000000000001800000000",
            INIT_7B => X"00000022000000000000001e0000000000000019000000000000001700000000",
            INIT_7C => X"00000028000000000000001c000000000000001f000000000000002000000000",
            INIT_7D => X"000000140000000000000013000000000000001d000000000000001e00000000",
            INIT_7E => X"0000001a000000000000001b0000000000000016000000000000001a00000000",
            INIT_7F => X"0000001b000000000000001e0000000000000014000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60 : if BRAM_NAME = "samplegold_layersamples_instance60" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002200000000000000240000000000000014000000000000001e00000000",
            INIT_01 => X"0000001b0000000000000019000000000000001c000000000000001800000000",
            INIT_02 => X"000000200000000000000022000000000000001b000000000000001900000000",
            INIT_03 => X"0000001f00000000000000170000000000000013000000000000001100000000",
            INIT_04 => X"00000013000000000000001e000000000000001b000000000000001b00000000",
            INIT_05 => X"00000022000000000000001b0000000000000014000000000000001200000000",
            INIT_06 => X"0000002400000000000000210000000000000020000000000000001f00000000",
            INIT_07 => X"0000001a000000000000001b0000000000000017000000000000002500000000",
            INIT_08 => X"0000001b000000000000001e000000000000001e000000000000001400000000",
            INIT_09 => X"00000022000000000000001d0000000000000018000000000000001500000000",
            INIT_0A => X"0000001e000000000000001e0000000000000020000000000000001a00000000",
            INIT_0B => X"00000014000000000000001c000000000000001a000000000000001f00000000",
            INIT_0C => X"000000210000000000000020000000000000001e000000000000001a00000000",
            INIT_0D => X"0000001e00000000000000200000000000000020000000000000001f00000000",
            INIT_0E => X"0000001e0000000000000022000000000000001e000000000000001d00000000",
            INIT_0F => X"000000170000000000000013000000000000001d000000000000001c00000000",
            INIT_10 => X"0000001e00000000000000210000000000000019000000000000001b00000000",
            INIT_11 => X"0000001b000000000000001a000000000000001e000000000000001f00000000",
            INIT_12 => X"0000001e000000000000001e0000000000000018000000000000001a00000000",
            INIT_13 => X"0000001e0000000000000015000000000000000f000000000000001e00000000",
            INIT_14 => X"0000001e000000000000001d0000000000000024000000000000002c00000000",
            INIT_15 => X"0000001c000000000000001a000000000000001b000000000000001900000000",
            INIT_16 => X"0000001d0000000000000017000000000000001f000000000000001800000000",
            INIT_17 => X"0000001e0000000000000019000000000000000f000000000000000f00000000",
            INIT_18 => X"00000018000000000000001d000000000000001c000000000000001e00000000",
            INIT_19 => X"0000001e000000000000001d000000000000001c000000000000001900000000",
            INIT_1A => X"0000000000000000000000000000000000000022000000000000001900000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000005000000000000002100000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000005000000000000000d0000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61 : if BRAM_NAME = "samplegold_layersamples_instance61" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"00000005000000000000000d0000000000000000000000000000001800000000",
            INIT_0E => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_0F => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_10 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000003000000000000002000000000",
            INIT_12 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_13 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_14 => X"0000000f00000000000000010000000000000000000000000000000000000000",
            INIT_15 => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000046000000000000007c000000000000008c00000000",
            INIT_17 => X"00000016000000000000003f0000000000000012000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_19 => X"0000002600000000000000000000000000000000000000000000000300000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000300000000000000160000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_24 => X"0000001000000000000000030000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000003000000000000000f000000000000000000000000",
            INIT_2A => X"00000000000000000000000b000000000000001e000000000000002500000000",
            INIT_2B => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000030000000000000001d000000000000000000000000",
            INIT_2F => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000f000000000000001f0000000000000033000000000000001100000000",
            INIT_44 => X"0000001900000000000000150000000000000018000000000000001000000000",
            INIT_45 => X"0000001900000000000000280000000000000000000000000000000c00000000",
            INIT_46 => X"0000001100000000000000120000000000000014000000000000001200000000",
            INIT_47 => X"00000008000000000000000f000000000000002e000000000000002200000000",
            INIT_48 => X"000000070000000000000011000000000000000e000000000000000500000000",
            INIT_49 => X"0000000e00000000000000100000000000000034000000000000000000000000",
            INIT_4A => X"000000170000000000000011000000000000000e000000000000001000000000",
            INIT_4B => X"000000000000000000000008000000000000000f000000000000004300000000",
            INIT_4C => X"0000000c00000000000000050000000000000010000000000000000900000000",
            INIT_4D => X"0000000900000000000000080000000000000011000000000000001f00000000",
            INIT_4E => X"00000034000000000000002b000000000000000f000000000000000a00000000",
            INIT_4F => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_50 => X"0000000a0000000000000019000000000000000f000000000000000500000000",
            INIT_51 => X"0000001100000000000000000000000000000000000000000000001500000000",
            INIT_52 => X"000000000000000000000011000000000000001b000000000000000600000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_54 => X"0000001a00000000000000120000000000000011000000000000000b00000000",
            INIT_55 => X"0000000d000000000000001d0000000000000001000000000000000200000000",
            INIT_56 => X"0000000f0000000000000000000000000000000e000000000000001000000000",
            INIT_57 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"00000009000000000000001d0000000000000010000000000000000d00000000",
            INIT_59 => X"000000100000000000000011000000000000001c000000000000000400000000",
            INIT_5A => X"0000000600000000000000080000000000000010000000000000000200000000",
            INIT_5B => X"0000000d00000000000000010000000000000004000000000000000000000000",
            INIT_5C => X"00000007000000000000000b000000000000001c000000000000000c00000000",
            INIT_5D => X"00000000000000000000000e000000000000000d000000000000000f00000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_5F => X"000000040000000000000008000000000000000d000000000000000000000000",
            INIT_60 => X"0000000d00000000000000040000000000000015000000000000001400000000",
            INIT_61 => X"0000001100000000000000000000000000000014000000000000000900000000",
            INIT_62 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_63 => X"00000009000000000000000b0000000000000000000000000000001900000000",
            INIT_64 => X"0000000d0000000000000020000000000000000b000000000000002500000000",
            INIT_65 => X"0000000900000000000000030000000000000007000000000000000d00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000e00000000000000100000000000000006000000000000000c00000000",
            INIT_68 => X"00000002000000000000000f0000000000000019000000000000000d00000000",
            INIT_69 => X"0000000000000000000000010000000000000004000000000000001100000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_6B => X"00000003000000000000000a0000000000000012000000000000000d00000000",
            INIT_6C => X"0000001a0000000000000005000000000000000f000000000000000a00000000",
            INIT_6D => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001a00000000000000000000000000000000000000000000000200000000",
            INIT_6F => X"000000080000000000000001000000000000000b000000000000000900000000",
            INIT_70 => X"00000001000000000000001c0000000000000010000000000000000f00000000",
            INIT_71 => X"00000004000000000000000d0000000000000000000000000000000000000000",
            INIT_72 => X"0000000800000000000000160000000000000001000000000000000000000000",
            INIT_73 => X"0000000e000000000000000b000000000000000a000000000000000900000000",
            INIT_74 => X"0000000000000000000000070000000000000022000000000000001300000000",
            INIT_75 => X"0000000300000000000000080000000000000007000000000000000000000000",
            INIT_76 => X"00000006000000000000000b0000000000000016000000000000000b00000000",
            INIT_77 => X"00000019000000000000000f000000000000000d000000000000001700000000",
            INIT_78 => X"000000000000000000000000000000000000000e000000000000001b00000000",
            INIT_79 => X"000000140000000000000005000000000000000d000000000000000000000000",
            INIT_7A => X"00000012000000000000000b000000000000000f000000000000001100000000",
            INIT_7B => X"0000000000000000000000000000000000000004000000000000001000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62 : if BRAM_NAME = "samplegold_layersamples_instance62" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000800000000000000000000000000000000000000000000000200000000",
            INIT_04 => X"0000000d0000000000000005000000000000000c000000000000001c00000000",
            INIT_05 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000c00000000000000110000000000000002000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_09 => X"0000001c00000000000000090000000000000000000000000000001100000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0B => X"0000001200000000000000140000000000000002000000000000000000000000",
            INIT_0C => X"0000000200000000000000000000000000000002000000000000001600000000",
            INIT_0D => X"0000000000000000000000070000000000000008000000000000000100000000",
            INIT_0E => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_0F => X"00000000000000000000001b000000000000001a000000000000000700000000",
            INIT_10 => X"0000000000000000000000090000000000000000000000000000000200000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_12 => X"0000000a00000000000000000000000000000006000000000000000000000000",
            INIT_13 => X"0000001300000000000000000000000000000016000000000000000000000000",
            INIT_14 => X"0000000900000000000000000000000000000001000000000000000e00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_16 => X"00000019000000000000000f0000000000000000000000000000000000000000",
            INIT_17 => X"0000000300000000000000020000000000000012000000000000000f00000000",
            INIT_18 => X"0000001800000000000000080000000000000015000000000000001400000000",
            INIT_19 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_1A => X"0000000d000000000000000a0000000000000007000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_1C => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_1D => X"00000006000000000000000a0000000000000000000000000000000000000000",
            INIT_1E => X"000000080000000000000017000000000000001f000000000000001100000000",
            INIT_1F => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_20 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000200000000000000020000000000000004000000000000000a00000000",
            INIT_22 => X"0000000e000000000000000e000000000000000a000000000000001600000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_24 => X"0000000800000000000000050000000000000000000000000000000000000000",
            INIT_25 => X"0000000900000000000000140000000000000011000000000000000200000000",
            INIT_26 => X"00000000000000000000000c0000000000000001000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000023000000000000001400000000",
            INIT_2A => X"0000000000000000000000000000000000000009000000000000000500000000",
            INIT_2B => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_2C => X"0000001000000000000000000000000000000000000000000000000400000000",
            INIT_2D => X"0000000000000000000000060000000000000000000000000000000b00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000f00000000000000140000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000007000000000000000e00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000018000000000000000c0000000000000008000000000000001c00000000",
            INIT_35 => X"000000000000000000000000000000000000000d000000000000001200000000",
            INIT_36 => X"00000011000000000000000f0000000000000006000000000000001700000000",
            INIT_37 => X"00000026000000000000001f0000000000000000000000000000001300000000",
            INIT_38 => X"0000000c00000000000000000000000000000000000000000000000800000000",
            INIT_39 => X"0000000b00000000000000000000000000000000000000000000000400000000",
            INIT_3A => X"0000000b00000000000000060000000000000000000000000000000000000000",
            INIT_3B => X"000000040000000000000020000000000000000c000000000000000000000000",
            INIT_3C => X"0000001400000000000000030000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_58 => X"0000000a00000000000000000000000000000000000000000000000700000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000300000000",
            INIT_63 => X"0000000300000000000000050000000000000001000000000000000800000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000600000000000000050000000000000004000000000000000500000000",
            INIT_67 => X"0000000100000000000000090000000000000000000000000000000200000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000c00000000000000050000000000000000000000000000000000000000",
            INIT_6A => X"000000030000000000000004000000000000000d000000000000000300000000",
            INIT_6B => X"0000000100000000000000040000000000000007000000000000000000000000",
            INIT_6C => X"00000018000000000000001d0000000000000018000000000000002600000000",
            INIT_6D => X"0000001600000000000000250000000000000026000000000000002800000000",
            INIT_6E => X"0000002b000000000000001a0000000000000029000000000000001900000000",
            INIT_6F => X"0000001a0000000000000004000000000000002d000000000000002d00000000",
            INIT_70 => X"0000001e00000000000000060000000000000028000000000000000100000000",
            INIT_71 => X"000000210000000000000018000000000000001e000000000000001d00000000",
            INIT_72 => X"0000002a0000000000000023000000000000001c000000000000001500000000",
            INIT_73 => X"0000000000000000000000080000000000000007000000000000002a00000000",
            INIT_74 => X"00000012000000000000000a0000000000000002000000000000002700000000",
            INIT_75 => X"000000000000000000000020000000000000000a000000000000001000000000",
            INIT_76 => X"0000001d000000000000001a0000000000000019000000000000001b00000000",
            INIT_77 => X"000000220000000000000009000000000000002c000000000000000e00000000",
            INIT_78 => X"0000000900000000000000180000000000000010000000000000000000000000",
            INIT_79 => X"0000001d0000000000000002000000000000001c000000000000000d00000000",
            INIT_7A => X"0000002700000000000000210000000000000011000000000000001b00000000",
            INIT_7B => X"0000000000000000000000280000000000000016000000000000001d00000000",
            INIT_7C => X"0000000b000000000000000d000000000000000f000000000000000b00000000",
            INIT_7D => X"0000001c000000000000000c0000000000000013000000000000001700000000",
            INIT_7E => X"0000002100000000000000210000000000000024000000000000002500000000",
            INIT_7F => X"0000000e0000000000000007000000000000002f000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63 : if BRAM_NAME = "samplegold_layersamples_instance63" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000130000000000000000000000000000001c000000000000000400000000",
            INIT_01 => X"00000025000000000000001a000000000000000f000000000000001200000000",
            INIT_02 => X"0000002900000000000000280000000000000023000000000000002a00000000",
            INIT_03 => X"0000000400000000000000170000000000000005000000000000000900000000",
            INIT_04 => X"0000001b00000000000000060000000000000000000000000000002200000000",
            INIT_05 => X"00000032000000000000001e0000000000000020000000000000000f00000000",
            INIT_06 => X"00000002000000000000001e0000000000000023000000000000002700000000",
            INIT_07 => X"0000000a00000000000000130000000000000003000000000000001600000000",
            INIT_08 => X"0000002c0000000000000009000000000000002a000000000000000f00000000",
            INIT_09 => X"0000001c00000000000000300000000000000012000000000000001300000000",
            INIT_0A => X"00000014000000000000000f0000000000000014000000000000002100000000",
            INIT_0B => X"0000002a00000000000000000000000000000012000000000000000600000000",
            INIT_0C => X"0000001b000000000000001f0000000000000008000000000000002800000000",
            INIT_0D => X"0000002a00000000000000220000000000000029000000000000001a00000000",
            INIT_0E => X"0000000d00000000000000100000000000000013000000000000000a00000000",
            INIT_0F => X"0000001b00000000000000190000000000000014000000000000000e00000000",
            INIT_10 => X"0000001600000000000000260000000000000019000000000000000f00000000",
            INIT_11 => X"0000000f000000000000001f0000000000000021000000000000001700000000",
            INIT_12 => X"0000000c000000000000000e000000000000001b000000000000001800000000",
            INIT_13 => X"00000023000000000000000b0000000000000014000000000000001700000000",
            INIT_14 => X"0000001b000000000000001b000000000000000f000000000000001500000000",
            INIT_15 => X"000000120000000000000011000000000000001a000000000000002100000000",
            INIT_16 => X"0000001a00000000000000100000000000000028000000000000000f00000000",
            INIT_17 => X"00000018000000000000001a0000000000000020000000000000001200000000",
            INIT_18 => X"000000220000000000000017000000000000001d000000000000000c00000000",
            INIT_19 => X"00000000000000000000000a000000000000001c000000000000002400000000",
            INIT_1A => X"00000016000000000000001b000000000000000a000000000000003b00000000",
            INIT_1B => X"0000000e000000000000001d0000000000000012000000000000002000000000",
            INIT_1C => X"0000002600000000000000250000000000000015000000000000001800000000",
            INIT_1D => X"0000002700000000000000150000000000000008000000000000002700000000",
            INIT_1E => X"00000026000000000000001c0000000000000019000000000000001000000000",
            INIT_1F => X"000000180000000000000019000000000000001a000000000000001100000000",
            INIT_20 => X"00000033000000000000001e0000000000000027000000000000001800000000",
            INIT_21 => X"0000002200000000000000100000000000000017000000000000000000000000",
            INIT_22 => X"0000001700000000000000200000000000000014000000000000001500000000",
            INIT_23 => X"000000130000000000000017000000000000001b000000000000001500000000",
            INIT_24 => X"00000048000000000000004d0000000000000047000000000000004600000000",
            INIT_25 => X"0000003500000000000000300000000000000036000000000000003900000000",
            INIT_26 => X"0000004b00000000000000510000000000000050000000000000004900000000",
            INIT_27 => X"0000005a00000000000000360000000000000037000000000000004000000000",
            INIT_28 => X"00000052000000000000005d0000000000000059000000000000005800000000",
            INIT_29 => X"000000620000000000000063000000000000005b000000000000005800000000",
            INIT_2A => X"00000052000000000000004b0000000000000046000000000000005a00000000",
            INIT_2B => X"0000006100000000000000610000000000000038000000000000004b00000000",
            INIT_2C => X"00000047000000000000003a000000000000005c000000000000005d00000000",
            INIT_2D => X"0000004a0000000000000049000000000000004e000000000000004a00000000",
            INIT_2E => X"000000460000000000000053000000000000004a000000000000003200000000",
            INIT_2F => X"0000005c00000000000000650000000000000061000000000000002e00000000",
            INIT_30 => X"0000007a00000000000000610000000000000045000000000000005e00000000",
            INIT_31 => X"0000006200000000000000540000000000000067000000000000006e00000000",
            INIT_32 => X"0000003c00000000000000350000000000000048000000000000004600000000",
            INIT_33 => X"00000060000000000000006f0000000000000060000000000000006100000000",
            INIT_34 => X"00000069000000000000006c000000000000006f000000000000005000000000",
            INIT_35 => X"0000003f0000000000000066000000000000006f000000000000006a00000000",
            INIT_36 => X"0000005a00000000000000270000000000000048000000000000005400000000",
            INIT_37 => X"00000046000000000000005e0000000000000058000000000000006500000000",
            INIT_38 => X"000000660000000000000066000000000000005c000000000000005800000000",
            INIT_39 => X"0000004e00000000000000640000000000000066000000000000006400000000",
            INIT_3A => X"0000005e00000000000000560000000000000061000000000000006200000000",
            INIT_3B => X"00000059000000000000003c000000000000003f000000000000005000000000",
            INIT_3C => X"0000005b000000000000004a000000000000004f000000000000006400000000",
            INIT_3D => X"0000005e000000000000005b0000000000000048000000000000005100000000",
            INIT_3E => X"0000002600000000000000510000000000000059000000000000006400000000",
            INIT_3F => X"0000003b0000000000000050000000000000005e000000000000005300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003e0000000000000048000000000000004b000000000000004600000000",
            INIT_41 => X"0000004b0000000000000057000000000000004b000000000000004a00000000",
            INIT_42 => X"00000041000000000000003a000000000000003f000000000000004300000000",
            INIT_43 => X"0000002c0000000000000047000000000000003b000000000000003900000000",
            INIT_44 => X"00000000000000000000001d0000000000000007000000000000000000000000",
            INIT_45 => X"000000540000000000000052000000000000004e000000000000001a00000000",
            INIT_46 => X"00000033000000000000002e0000000000000030000000000000005000000000",
            INIT_47 => X"00000064000000000000003d000000000000003c000000000000003a00000000",
            INIT_48 => X"000000530000000000000055000000000000005e000000000000005300000000",
            INIT_49 => X"0000004600000000000000540000000000000040000000000000005100000000",
            INIT_4A => X"0000001e00000000000000230000000000000028000000000000002200000000",
            INIT_4B => X"0000004100000000000000340000000000000042000000000000002200000000",
            INIT_4C => X"0000003600000000000000380000000000000032000000000000003d00000000",
            INIT_4D => X"00000017000000000000005e0000000000000061000000000000004200000000",
            INIT_4E => X"0000003a00000000000000200000000000000024000000000000002100000000",
            INIT_4F => X"000000390000000000000043000000000000001d000000000000003300000000",
            INIT_50 => X"0000003500000000000000360000000000000051000000000000004b00000000",
            INIT_51 => X"000000410000000000000022000000000000003a000000000000006100000000",
            INIT_52 => X"0000000e000000000000000b0000000000000012000000000000002d00000000",
            INIT_53 => X"0000004a00000000000000450000000000000010000000000000000e00000000",
            INIT_54 => X"0000005800000000000000310000000000000011000000000000002900000000",
            INIT_55 => X"00000034000000000000003d0000000000000054000000000000006200000000",
            INIT_56 => X"0000001800000000000000060000000000000003000000000000002300000000",
            INIT_57 => X"000000180000000000000050000000000000004c000000000000004200000000",
            INIT_58 => X"0000005a0000000000000062000000000000003c000000000000001300000000",
            INIT_59 => X"0000002000000000000000300000000000000037000000000000004b00000000",
            INIT_5A => X"00000029000000000000001a0000000000000011000000000000000e00000000",
            INIT_5B => X"0000001500000000000000180000000000000038000000000000004100000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_5D => X"0000000800000000000000030000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000005000000000000001400000000",
            INIT_5F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000300000000000000010000000000000010000000000000001100000000",
            INIT_66 => X"0000000000000000000000000000000000000028000000000000000800000000",
            INIT_67 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_68 => X"0000000a000000000000003b0000000000000000000000000000000000000000",
            INIT_69 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001100000000000000000000000000000001000000000000003200000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_71 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_73 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000c00000000000000000000000000000000000000000000000200000000",
            INIT_75 => X"00000002000000000000000f0000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_79 => X"0000000d00000000000000060000000000000000000000000000000000000000",
            INIT_7A => X"0000001900000000000000000000000000000000000000000000003400000000",
            INIT_7B => X"00000000000000000000000f000000000000000e000000000000000000000000",
            INIT_7C => X"0000000000000000000000430000000000000036000000000000000000000000",
            INIT_7D => X"00000042000000000000000b0000000000000040000000000000002b00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000002700000000000000010000000000000000000000000000000e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64 : if BRAM_NAME = "samplegold_layersamples_instance64" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000000000000000000005d0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_03 => X"0000001700000000000000000000000000000023000000000000001300000000",
            INIT_04 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000054000000000000000c00000000",
            INIT_06 => X"0000000000000000000000000000000000000005000000000000001500000000",
            INIT_07 => X"0000000000000000000000460000000000000000000000000000000a00000000",
            INIT_08 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_09 => X"0000002300000000000000000000000000000000000000000000005d00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000060000000000000001e000000000000000700000000",
            INIT_0C => X"0000006500000000000000170000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0E => X"0000001300000000000000090000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000000000000000000000000000f000000000000001800000000",
            INIT_10 => X"00000000000000000000004e000000000000002b000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000b00000000000000070000000000000004000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000009000000000000000a00000000",
            INIT_14 => X"0000000000000000000000000000000000000061000000000000001c00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000019a00000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"00000138000000000000016a000000000000019a000000000000019900000000",
            INIT_4E => X"000001a200000000000001720000000000000154000000000000013f00000000",
            INIT_4F => X"00000192000000000000019700000000000001a500000000000001ab00000000",
            INIT_50 => X"000001c400000000000001c50000000000000168000000000000018300000000",
            INIT_51 => X"0000010a0000000000000113000000000000016500000000000001c500000000",
            INIT_52 => X"000001590000000000000145000000000000012e000000000000011200000000",
            INIT_53 => X"0000019500000000000001a2000000000000018c000000000000017000000000",
            INIT_54 => X"000001bc00000000000001c900000000000001ca000000000000016800000000",
            INIT_55 => X"000000ee00000000000000ee00000000000000af000000000000014e00000000",
            INIT_56 => X"0000011800000000000000f700000000000000ef00000000000000fa00000000",
            INIT_57 => X"00000144000000000000017000000000000001a6000000000000019a00000000",
            INIT_58 => X"0000015c000000000000019600000000000001cc00000000000001c800000000",
            INIT_59 => X"0000011b0000000000000163000000000000014000000000000000d100000000",
            INIT_5A => X"0000014f00000000000001510000000000000113000000000000011900000000",
            INIT_5B => X"000001c2000000000000014d000000000000017f000000000000018900000000",
            INIT_5C => X"000000d90000000000000103000000000000018f00000000000001c800000000",
            INIT_5D => X"000001140000000000000102000000000000010e000000000000010b00000000",
            INIT_5E => X"000001a100000000000001430000000000000136000000000000011b00000000",
            INIT_5F => X"000001c10000000000000195000000000000017200000000000001af00000000",
            INIT_60 => X"000000cc00000000000000930000000000000110000000000000014a00000000",
            INIT_61 => X"000000de00000000000000d800000000000000d600000000000000e300000000",
            INIT_62 => X"000001cb0000000000000167000000000000011600000000000000f900000000",
            INIT_63 => X"000001280000000000000179000000000000017700000000000001c900000000",
            INIT_64 => X"000000e200000000000000e600000000000000d100000000000000de00000000",
            INIT_65 => X"000000d300000000000000ec00000000000000bd00000000000000be00000000",
            INIT_66 => X"000001ad0000000000000161000000000000013100000000000000d600000000",
            INIT_67 => X"0000014000000000000000c3000000000000011e000000000000017100000000",
            INIT_68 => X"00000091000000000000008f00000000000000aa00000000000000bb00000000",
            INIT_69 => X"0000006d000000000000006f0000000000000066000000000000006f00000000",
            INIT_6A => X"0000016a000000000000014c00000000000000df000000000000008600000000",
            INIT_6B => X"0000008a00000000000000d400000000000000ee000000000000010900000000",
            INIT_6C => X"000000ab00000000000000cb00000000000000ce00000000000000c600000000",
            INIT_6D => X"000000d500000000000000ba00000000000000fa00000000000000c400000000",
            INIT_6E => X"00000119000000000000017e0000000000000130000000000000010800000000",
            INIT_6F => X"0000008e000000000000007d000000000000008300000000000000af00000000",
            INIT_70 => X"000000e200000000000001110000000000000093000000000000008800000000",
            INIT_71 => X"000000ce00000000000000f800000000000000e200000000000000f400000000",
            INIT_72 => X"0000009d000000000000011b000000000000017500000000000000c600000000",
            INIT_73 => X"00000081000000000000004b000000000000005a000000000000007c00000000",
            INIT_74 => X"000000a300000000000000c9000000000000006f00000000000000c300000000",
            INIT_75 => X"000000e000000000000000a300000000000000cd00000000000000ad00000000",
            INIT_76 => X"000000b30000000000000066000000000000010e000000000000016e00000000",
            INIT_77 => X"0000006200000000000000610000000000000048000000000000009200000000",
            INIT_78 => X"0000010300000000000000dd00000000000000c6000000000000006200000000",
            INIT_79 => X"00000143000000000000007f000000000000008a00000000000000a800000000",
            INIT_7A => X"0000009900000000000000e800000000000000cf000000000000010a00000000",
            INIT_7B => X"00000037000000000000002b0000000000000027000000000000005f00000000",
            INIT_7C => X"000000760000000000000136000000000000015200000000000000a400000000",
            INIT_7D => X"00000146000000000000013f00000000000000a0000000000000003f00000000",
            INIT_7E => X"0000007a000000000000009d00000000000000dd000000000000010300000000",
            INIT_7F => X"000000c4000000000000005d0000000000000037000000000000002f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65 : if BRAM_NAME = "samplegold_layersamples_instance65" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000470000000000000047000000000000011100000000000000e300000000",
            INIT_01 => X"0000010d0000000000000120000000000000013500000000000000a500000000",
            INIT_02 => X"000000510000000000000070000000000000008b00000000000000bb00000000",
            INIT_03 => X"000000a3000000000000007a000000000000005f000000000000005400000000",
            INIT_04 => X"000000a30000000000000048000000000000005f00000000000000b800000000",
            INIT_05 => X"00000059000000000000005f000000000000004f000000000000005a00000000",
            INIT_06 => X"0000003d000000000000003e0000000000000042000000000000004d00000000",
            INIT_07 => X"0000005f00000000000000610000000000000062000000000000004900000000",
            INIT_08 => X"00000060000000000000004c0000000000000053000000000000005a00000000",
            INIT_09 => X"000000330000000000000054000000000000006e000000000000005f00000000",
            INIT_0A => X"0000005800000000000000480000000000000034000000000000003500000000",
            INIT_0B => X"00000067000000000000005c000000000000005e000000000000005c00000000",
            INIT_0C => X"0000006300000000000000630000000000000059000000000000007000000000",
            INIT_0D => X"0000000000000000000000000000000000000036000000000000006a00000000",
            INIT_0E => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000006d000000000000006b000000000000005c000000000000003a00000000",
            INIT_10 => X"0000005500000000000000670000000000000063000000000000005300000000",
            INIT_11 => X"00000014000000000000001b0000000000000005000000000000004a00000000",
            INIT_12 => X"0000001d00000000000000070000000000000006000000000000000a00000000",
            INIT_13 => X"0000004900000000000000680000000000000060000000000000005900000000",
            INIT_14 => X"0000002d0000000000000055000000000000006b000000000000006300000000",
            INIT_15 => X"000000000000000000000018000000000000000a000000000000000000000000",
            INIT_16 => X"0000003400000000000000210000000000000003000000000000000c00000000",
            INIT_17 => X"0000006000000000000000440000000000000061000000000000005200000000",
            INIT_18 => X"00000000000000000000001b000000000000003b000000000000007300000000",
            INIT_19 => X"0000000200000000000000020000000000000001000000000000000000000000",
            INIT_1A => X"0000004d000000000000001a000000000000001b000000000000000100000000",
            INIT_1B => X"0000006800000000000000520000000000000063000000000000006300000000",
            INIT_1C => X"0000000000000000000000000000000000000027000000000000004500000000",
            INIT_1D => X"0000001400000000000000000000000000000000000000000000000b00000000",
            INIT_1E => X"00000059000000000000003d0000000000000013000000000000000c00000000",
            INIT_1F => X"0000002f000000000000004c0000000000000064000000000000005d00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_21 => X"0000000c00000000000000000000000000000008000000000000000b00000000",
            INIT_22 => X"0000004700000000000000100000000000000000000000000000000c00000000",
            INIT_23 => X"0000003400000000000000280000000000000037000000000000005800000000",
            INIT_24 => X"000000000000000000000004000000000000001e000000000000000100000000",
            INIT_25 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_26 => X"000000570000000000000020000000000000001a000000000000000000000000",
            INIT_27 => X"00000000000000000000000c0000000000000032000000000000003f00000000",
            INIT_28 => X"0000001d00000000000000130000000000000000000000000000000700000000",
            INIT_29 => X"00000035000000000000001f0000000000000026000000000000001c00000000",
            INIT_2A => X"0000004100000000000000540000000000000001000000000000001400000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000000000000b00000000",
            INIT_2C => X"0000000d0000000000000000000000000000000d000000000000000000000000",
            INIT_2D => X"0000000900000000000000180000000000000000000000000000000500000000",
            INIT_2E => X"00000016000000000000003f0000000000000045000000000000000000000000",
            INIT_2F => X"0000000900000000000000000000000000000007000000000000000700000000",
            INIT_30 => X"0000001900000000000000230000000000000003000000000000002200000000",
            INIT_31 => X"000000000000000000000011000000000000001a000000000000003700000000",
            INIT_32 => X"0000002900000000000000000000000000000025000000000000003000000000",
            INIT_33 => X"0000000000000000000000000000000000000004000000000000001000000000",
            INIT_34 => X"0000004100000000000000290000000000000011000000000000000000000000",
            INIT_35 => X"0000002d00000000000000000000000000000000000000000000000700000000",
            INIT_36 => X"0000000e000000000000002d0000000000000029000000000000003400000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_38 => X"00000006000000000000004e000000000000002a000000000000000a00000000",
            INIT_39 => X"0000002200000000000000250000000000000000000000000000000000000000",
            INIT_3A => X"0000000d000000000000000a0000000000000018000000000000002800000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000034000000000000000a00000000",
            INIT_3D => X"0000000b00000000000000000000000000000001000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_3F => X"0000000200000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001a0000000000000000000000000000001b000000000000000000000000",
            INIT_41 => X"0000005100000000000000190000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_45 => X"000000000000000000000090000000000000001d000000000000000000000000",
            INIT_46 => X"00000001000000000000000f0000000000000000000000000000000000000000",
            INIT_47 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000800000000000000000000000000000000000000000000002600000000",
            INIT_49 => X"0000000000000000000000000000000000000086000000000000000f00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_4B => X"00000024000000000000000e0000000000000000000000000000000000000000",
            INIT_4C => X"0000002a00000000000000130000000000000000000000000000000000000000",
            INIT_4D => X"0000001a00000000000000000000000000000000000000000000006000000000",
            INIT_4E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000100000000000000220000000000000000000000000000000000000000",
            INIT_50 => X"0000006800000000000000360000000000000020000000000000000000000000",
            INIT_51 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"00000000000000000000004a000000000000000b000000000000003100000000",
            INIT_55 => X"00000000000000000000000a0000000000000013000000000000000000000000",
            INIT_56 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_57 => X"0000004a00000000000000080000000000000000000000000000000000000000",
            INIT_58 => X"00000017000000000000000a0000000000000035000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000017000000000000000500000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_5B => X"0000000000000000000000590000000000000019000000000000000000000000",
            INIT_5C => X"0000000200000000000000000000000000000000000000000000005500000000",
            INIT_5D => X"0000002700000000000000000000000000000000000000000000002000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_5F => X"0000003f0000000000000000000000000000007b000000000000001e00000000",
            INIT_60 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_61 => X"00000000000000000000000c0000000000000000000000000000001500000000",
            INIT_62 => X"000000070000000000000000000000000000002e000000000000000000000000",
            INIT_63 => X"0000000b000000000000001c0000000000000006000000000000008900000000",
            INIT_64 => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_65 => X"0000002600000000000000000000000000000008000000000000001c00000000",
            INIT_66 => X"00000093000000000000000a0000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000040000000000000000a000000000000000000000000",
            INIT_68 => X"0000000a00000000000000000000000000000042000000000000000000000000",
            INIT_69 => X"00000000000000000000005e0000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_6B => X"0000000100000000000000290000000000000033000000000000000b00000000",
            INIT_6C => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000030000000000000005900000000",
            INIT_6E => X"0000000e00000000000000370000000000000017000000000000000000000000",
            INIT_6F => X"000000000000000000000001000000000000003f000000000000000a00000000",
            INIT_70 => X"0000006600000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000800000000000000000000000000000000000000000000002900000000",
            INIT_72 => X"000000040000000000000025000000000000002e000000000000000a00000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000001d00000000",
            INIT_74 => X"0000002800000000000000300000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000001300000000000000050000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000000f000000000000001b00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_7F => X"0000000000000000000000080000000000000008000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66 : if BRAM_NAME = "samplegold_layersamples_instance66" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_0A => X"0000000b00000000000000030000000000000001000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000012000000000000000600000000",
            INIT_10 => X"0000000000000000000000000000000000000007000000000000000700000000",
            INIT_11 => X"0000001400000000000000160000000000000027000000000000000c00000000",
            INIT_12 => X"00000013000000000000000c000000000000001d000000000000001900000000",
            INIT_13 => X"0000000000000000000000000000000000000004000000000000000e00000000",
            INIT_14 => X"000000000000000000000000000000000000002c000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000014000000000000000a0000000000000000000000000000000000000000",
            INIT_19 => X"0000001f00000000000000280000000000000000000000000000002700000000",
            INIT_1A => X"0000000000000000000000150000000000000017000000000000002000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000016000000000000000300000000",
            INIT_1D => X"00000000000000000000000f0000000000000006000000000000001a00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_1F => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_20 => X"00000000000000000000002c0000000000000023000000000000000000000000",
            INIT_21 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000018000000000000001700000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_25 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000000e000000000000000400000000",
            INIT_2A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000001000000000000000130000000000000004000000000000000a00000000",
            INIT_34 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_36 => X"0000000000000000000000030000000000000026000000000000000000000000",
            INIT_37 => X"00000037000000000000000a0000000000000000000000000000000000000000",
            INIT_38 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000000000000000000000d000000000000004000000000",
            INIT_3B => X"0000002a00000000000000000000000000000003000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000200000000000000010000000000000000000000000000000800000000",
            INIT_3F => X"0000000900000000000000210000000000000000000000000000000700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_41 => X"0000000d000000000000001c0000000000000000000000000000000000000000",
            INIT_42 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000310000000000000013000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_47 => X"0000000e000000000000001b0000000000000021000000000000001e00000000",
            INIT_48 => X"0000000000000000000000390000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_4A => X"0000000800000000000000000000000000000005000000000000000000000000",
            INIT_4B => X"00000000000000000000004d0000000000000021000000000000003100000000",
            INIT_4C => X"0000002b00000000000000000000000000000023000000000000000000000000",
            INIT_4D => X"0000000700000000000000000000000000000007000000000000000300000000",
            INIT_4E => X"0000001300000000000000000000000000000000000000000000000c00000000",
            INIT_4F => X"0000000000000000000000000000000000000046000000000000000000000000",
            INIT_50 => X"0000000000000000000000190000000000000000000000000000001800000000",
            INIT_51 => X"0000000b00000000000000000000000000000033000000000000000c00000000",
            INIT_52 => X"0000000000000000000000090000000000000005000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_54 => X"0000002100000000000000180000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000000000000000000003c000000000000000000000000",
            INIT_56 => X"0000003b00000000000000240000000000000000000000000000002200000000",
            INIT_57 => X"00000006000000000000002c0000000000000000000000000000000000000000",
            INIT_58 => X"00000000000000000000001d0000000000000001000000000000000000000000",
            INIT_59 => X"0000000000000000000000040000000000000008000000000000004000000000",
            INIT_5A => X"00000000000000000000006f0000000000000008000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000019000000000000000c0000000000000003000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000006600000000",
            INIT_5E => X"000000000000000000000000000000000000005d000000000000002200000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"00000022000000000000001a000000000000000e000000000000000300000000",
            INIT_61 => X"0000002d00000000000000000000000000000000000000000000001d00000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000005100000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000014000000000000000e0000000000000009000000000000000500000000",
            INIT_65 => X"0000006600000000000000240000000000000000000000000000000000000000",
            INIT_66 => X"0000001700000000000000190000000000000016000000000000001900000000",
            INIT_67 => X"0000001f000000000000001d0000000000000019000000000000001000000000",
            INIT_68 => X"0000001600000000000000180000000000000018000000000000001800000000",
            INIT_69 => X"00000017000000000000001a000000000000001e000000000000001e00000000",
            INIT_6A => X"00000000000000000000000e0000000000000018000000000000001600000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"000000170000000000000014000000000000000e000000000000000100000000",
            INIT_6D => X"0000001300000000000000140000000000000017000000000000001c00000000",
            INIT_6E => X"0000000000000000000000000000000000000008000000000000001500000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000019000000000000001b0000000000000019000000000000000000000000",
            INIT_71 => X"0000000f00000000000000130000000000000014000000000000000e00000000",
            INIT_72 => X"0000000000000000000000030000000000000000000000000000000b00000000",
            INIT_73 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000001800000000000000230000000000000017000000000000000400000000",
            INIT_75 => X"0000000000000000000000070000000000000015000000000000001400000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000120000000000000020000000000000001b000000000000001300000000",
            INIT_79 => X"00000000000000000000000a000000000000000f000000000000001500000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001300000000000000130000000000000014000000000000001400000000",
            INIT_7D => X"0000000000000000000000000000000000000009000000000000000c00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67 : if BRAM_NAME = "samplegold_layersamples_instance67" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b000000000000000f000000000000001c000000000000000c00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000c0000000000000019000000000000001d00000000",
            INIT_05 => X"0000000b00000000000000020000000000000008000000000000000000000000",
            INIT_06 => X"0000001a000000000000001c0000000000000018000000000000001800000000",
            INIT_07 => X"000000160000000000000001000000000000000b000000000000001000000000",
            INIT_08 => X"0000000000000000000000060000000000000000000000000000001200000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000001500000000000000130000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000001000000000000000700000000",
            INIT_0D => X"0000000100000000000000000000000000000005000000000000000000000000",
            INIT_0E => X"0000000200000000000000050000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000080000000000000005000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000009000000000000000b00000000",
            INIT_11 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_13 => X"00000002000000000000000b0000000000000011000000000000000100000000",
            INIT_14 => X"0000000000000000000000010000000000000007000000000000000400000000",
            INIT_15 => X"000000160000000000000019000000000000000e000000000000000000000000",
            INIT_16 => X"0000000100000000000000000000000000000000000000000000000500000000",
            INIT_17 => X"0000000000000000000000000000000000000006000000000000000200000000",
            INIT_18 => X"0000000300000000000000030000000000000004000000000000000700000000",
            INIT_19 => X"0000000200000000000000050000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000300000000000000000000000000000000000000000000000200000000",
            INIT_1C => X"0000000000000000000000000000000000000001000000000000000200000000",
            INIT_1D => X"0000000000000000000000050000000000000004000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000006000000000000000c0000000000000012000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000002000000000000001400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000001100000000000000050000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000010000000000000006000000000000000300000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000001200000000000000140000000000000001000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000001f000000000000001d0000000000000004000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000012000000000000001b00000000",
            INIT_4E => X"00000000000000000000000f000000000000000e000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000001c00000000000000200000000000000011000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_52 => X"000000000000000000000000000000000000000e000000000000001400000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000d00000000000000140000000000000017000000000000000900000000",
            INIT_55 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68 : if BRAM_NAME = "samplegold_layersamples_instance68" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000003000000000000000900000000",
            INIT_10 => X"0000000900000000000000360000000000000021000000000000001000000000",
            INIT_11 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000000a000000000000000d00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000040000000000000003a0000000000000014000000000000000c00000000",
            INIT_18 => X"000000000000000000000000000000000000001d000000000000004300000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000024000000000000000e00000000",
            INIT_1D => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000055000000000000001e00000000",
            INIT_22 => X"000000000000000000000000000000000000000d000000000000000600000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000039000000000000001300000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2E => X"000000a500000000000000500000000000000009000000000000000000000000",
            INIT_2F => X"0000007900000000000000ae000000000000009a000000000000009e00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_31 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001000000000000000130000000000000000000000000000000000000000",
            INIT_35 => X"0000003500000000000000000000000000000000000000000000000100000000",
            INIT_36 => X"00000003000000000000000c0000000000000000000000000000000900000000",
            INIT_37 => X"0000000000000000000000190000000000000000000000000000002a00000000",
            INIT_38 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_3A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000001b0000000000000000000000000000004b000000000000006900000000",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000001b00000000",
            INIT_3E => X"0000000000000000000000260000000000000037000000000000003400000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001300000000000000000000000000000000000000000000000100000000",
            INIT_41 => X"0000000000000000000000020000000000000011000000000000001400000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000001400000000000000050000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000005000000000000001100000000",
            INIT_46 => X"0000000b00000000000000000000000000000012000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_48 => X"0000000500000000000000030000000000000000000000000000000000000000",
            INIT_49 => X"0000000300000000000000000000000000000000000000000000000600000000",
            INIT_4A => X"000000000000000000000005000000000000000b000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000050000000000000008000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000009000000000000000c00000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000f00000000000000000000000000000000000000000000000900000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000f00000000000000000000000000000004000000000000000000000000",
            INIT_65 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000140000000000000000000000000000000100000000",
            INIT_69 => X"000000040000000000000000000000000000000a000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_6D => X"0000000400000000000000000000000000000000000000000000000100000000",
            INIT_6E => X"00000000000000000000000b0000000000000000000000000000000100000000",
            INIT_6F => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_70 => X"0000000d00000000000000000000000000000000000000000000000b00000000",
            INIT_71 => X"0000000500000000000000040000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_73 => X"0000001100000000000000070000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000b00000000000000090000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000001a000000000000000b00000000",
            INIT_77 => X"000000000000000000000014000000000000000b000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000008000000000000000b000000000000000c000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_7B => X"000000000000000000000000000000000000000a000000000000000f00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000030000000000000005000000000000000500000000",
            INIT_7E => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000017000000000000000e0000000000000010000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69 : if BRAM_NAME = "samplegold_layersamples_instance69" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000000000080000000000000011000000000000001800000000",
            INIT_01 => X"00000017000000000000001a0000000000000017000000000000000400000000",
            INIT_02 => X"0000000100000000000000050000000000000006000000000000001100000000",
            INIT_03 => X"0000003d0000000000000028000000000000001d000000000000001e00000000",
            INIT_04 => X"000000520000000000000048000000000000004b000000000000004900000000",
            INIT_05 => X"000000130000000000000016000000000000002e000000000000004c00000000",
            INIT_06 => X"0000002400000000000000000000000000000012000000000000001800000000",
            INIT_07 => X"000000320000000000000038000000000000002c000000000000002400000000",
            INIT_08 => X"00000044000000000000003e0000000000000039000000000000003a00000000",
            INIT_09 => X"0000001b0000000000000016000000000000000a000000000000003a00000000",
            INIT_0A => X"0000002b00000000000000240000000000000001000000000000001200000000",
            INIT_0B => X"0000004700000000000000390000000000000050000000000000002200000000",
            INIT_0C => X"0000004700000000000000550000000000000060000000000000006000000000",
            INIT_0D => X"0000000900000000000000100000000000000016000000000000004800000000",
            INIT_0E => X"0000004d00000000000000290000000000000023000000000000000d00000000",
            INIT_0F => X"0000005b000000000000005a000000000000004c000000000000004e00000000",
            INIT_10 => X"000000540000000000000057000000000000005a000000000000005e00000000",
            INIT_11 => X"0000000000000000000000130000000000000019000000000000002000000000",
            INIT_12 => X"00000053000000000000001c0000000000000035000000000000001c00000000",
            INIT_13 => X"0000005a0000000000000052000000000000004a000000000000004000000000",
            INIT_14 => X"0000003d0000000000000054000000000000004f000000000000005b00000000",
            INIT_15 => X"0000001d00000000000000240000000000000025000000000000001500000000",
            INIT_16 => X"0000003a00000000000000190000000000000021000000000000003100000000",
            INIT_17 => X"00000046000000000000004b000000000000005e000000000000005200000000",
            INIT_18 => X"0000004400000000000000390000000000000044000000000000005c00000000",
            INIT_19 => X"0000002c00000000000000250000000000000024000000000000003300000000",
            INIT_1A => X"0000003c000000000000004d0000000000000037000000000000000000000000",
            INIT_1B => X"0000003e0000000000000044000000000000003d000000000000003500000000",
            INIT_1C => X"0000003b000000000000003e0000000000000042000000000000003700000000",
            INIT_1D => X"0000001500000000000000190000000000000014000000000000001e00000000",
            INIT_1E => X"0000002c000000000000002a0000000000000027000000000000003400000000",
            INIT_1F => X"0000000b00000000000000000000000000000000000000000000001c00000000",
            INIT_20 => X"00000029000000000000003a0000000000000004000000000000000000000000",
            INIT_21 => X"0000001100000000000000290000000000000031000000000000001f00000000",
            INIT_22 => X"000000240000000000000036000000000000002e000000000000003400000000",
            INIT_23 => X"00000044000000000000004c0000000000000040000000000000005200000000",
            INIT_24 => X"000000200000000000000012000000000000003b000000000000004900000000",
            INIT_25 => X"0000001c000000000000001c0000000000000017000000000000002700000000",
            INIT_26 => X"0000001d0000000000000038000000000000000f000000000000001900000000",
            INIT_27 => X"0000002f00000000000000120000000000000028000000000000002b00000000",
            INIT_28 => X"00000042000000000000003a000000000000001b000000000000001900000000",
            INIT_29 => X"0000001a000000000000001e0000000000000012000000000000001200000000",
            INIT_2A => X"0000002a000000000000001a0000000000000028000000000000003100000000",
            INIT_2B => X"0000003d000000000000002e0000000000000041000000000000002a00000000",
            INIT_2C => X"000000160000000000000015000000000000003c000000000000000400000000",
            INIT_2D => X"0000000f0000000000000014000000000000001f000000000000003800000000",
            INIT_2E => X"0000002700000000000000000000000000000007000000000000000f00000000",
            INIT_2F => X"00000012000000000000000b0000000000000022000000000000003e00000000",
            INIT_30 => X"0000003b00000000000000380000000000000046000000000000003800000000",
            INIT_31 => X"000000070000000000000005000000000000001c000000000000002a00000000",
            INIT_32 => X"0000004c0000000000000033000000000000003e000000000000001000000000",
            INIT_33 => X"00000048000000000000001c000000000000000f000000000000000e00000000",
            INIT_34 => X"000000290000000000000032000000000000003c000000000000004000000000",
            INIT_35 => X"00000015000000000000000f000000000000000c000000000000001a00000000",
            INIT_36 => X"0000001200000000000000350000000000000031000000000000002100000000",
            INIT_37 => X"000000000000000000000000000000000000000f000000000000001000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_5C => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000150000000000000000000000000000000c000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000b000000000000001e0000000000000006000000000000001200000000",
            INIT_71 => X"0000000700000000000000150000000000000017000000000000001000000000",
            INIT_72 => X"0000001c00000000000000150000000000000015000000000000001100000000",
            INIT_73 => X"0000000e000000000000000e0000000000000022000000000000001e00000000",
            INIT_74 => X"0000000000000000000000000000000000000016000000000000000400000000",
            INIT_75 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000002100000000000000120000000000000009000000000000001600000000",
            INIT_77 => X"00000009000000000000000a000000000000000b000000000000001d00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_79 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000002200000000000000190000000000000011000000000000000300000000",
            INIT_7B => X"0000000000000000000000150000000000000001000000000000000c00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000b000000000000001a0000000000000018000000000000001300000000",
            INIT_7F => X"0000000000000000000000000000000000000008000000000000000300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70 : if BRAM_NAME = "samplegold_layersamples_instance70" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000800000000000000030000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000000b000000000000001e000000000000000a00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000b00000000000000070000000000000000000000000000000000000000",
            INIT_06 => X"0000000c00000000000000080000000000000001000000000000000a00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000160000000000000014000000000000000100000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000180000000000000000000000000000002500000000",
            INIT_0F => X"0000000400000000000000000000000000000000000000000000000400000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_11 => X"0000001700000000000000070000000000000000000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000210000000000000005000000000000000c00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001700000000000000000000000000000012000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_1A => X"0000000200000000000000000000000000000000000000000000000500000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000001e0000000000000000000000000000001300000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_1E => X"0000000800000000000000000000000000000000000000000000000300000000",
            INIT_1F => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000001000000000000000100000000",
            INIT_23 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70;

MEM_EMPTY_36Kb : if BRAM_NAME(1 to 7) = "default" generate
    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
        BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
        DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
        DO_REG => 0,                     -- Optional output register (0 or 1)
        INIT => X"000000000000000000",   -- Initial values on output port
        INIT_FILE => "NONE",
        WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        SRVAL => X"000000000000000000",  -- Set/Reset value for port output
        WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    )
    port map (
        DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
        ADDR => bram_addr,  -- Input address, width defined by read/write port depth
        CLK => CLK,    -- 1-bit input clock
        DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
        EN => EN,      -- 1-bit input RAM enable
        REGCE => '1', -- 1-bit input output register enable
        RST => RST,    -- 1-bit input reset
        WE => bram_wr_en       -- Input write enable, width defined by write port depth
    );
-- End of BRAM_SINGLE_MACRO_inst instantiation
end generate;


end a1;