library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    27622, 8918, -10166, -5123, -19765, -7146, -31934, -8966, 32049, 4956,

    -- weights
    -- filter=0 channel=0
    -9, 3, -17, 6, -3, -11, -14, 6, -20, -12, -5, -2, -3, 5, 0, -4, -13, -15, 0, -17, -6, -21, 3, 8, 2, 6, -2, -14, -2, -5, 2, -11, -9, 1, -11, -1, -3, 0, -16, -20, 1, -15, -17, -11, 0, -12, -15, -1, -21, -10, 3, -22, -13, 4, -7, -9, 0, -5, -13, 14, -14, 2, -21, -13, -6, -13, 8, 7, -4, -13, 11, -12, -10, -8, 0, -21, -25, -23, -19, -26, -8, -23, -6, 10, 4, 2, -6, 3, -3, -4, -4, 1, -14, -23, -9, -17, -5, -9, -16, -15, 6, -20, 4, -18, 0, -14, -4, 1, -12, -3, 2, 7, -22, 9, 9, -21, -13, -18, -19, -5, -15, -9, -26, -7, -15, -13, -25, -16, -7, -6, 0, 8, -4, -3, 3, -9, -16, -19, -11, -10, -15, 1, 4, -12, -15, 8, -13, 3, 7, 11, -7, -19, -11, -10, -15, -3, -17, -17, -10, -10, -6, 5, 2, 2, 8, -12, -10, -7, -22, -14, 4, -1, -3, 8, -14, 8, -19, -5, -10, -8, 12, -26, -3, -21, -16, -24, -15, -20, -13, 6, 5, -10, -1, -2, -17, 4, -20, -2, -1, 0, -1, -19, -8, 1, -21, 2, -4, 7, 12, 7, 8, -21, -5, -13, -7, -6, -19, -7, -9, -10, 1, 3, -10, -6, 1,
    -- filter=0 channel=1
    2, 26, -6, 12, -6, 9, 11, 14, 8, 5, 0, -13, 14, -1, -4, 4, 15, -3, -1, -7, 13, 2, 14, 1, 3, -5, 4, 15, 0, -12, 24, 0, 15, 12, 20, 0, -4, -15, -21, -20, -16, 4, 6, -12, -13, 10, 26, 7, 13, -2, -10, -17, -21, 8, -19, -10, -13, 3, 9, -17, 23, 19, 9, -7, 12, -2, -15, -15, -14, -20, -21, 2, -10, 8, 15, 21, 16, 9, -4, 11, -20, -14, -8, -12, 3, -11, 2, 11, -5, 4, 24, 2, 5, -18, -1, 3, -27, -8, -25, -14, 0, 2, 0, 0, -12, -5, 23, 3, -13, 5, -12, -23, -21, -19, -17, -17, 3, -16, -16, -8, 12, -5, 13, -8, 1, -26, -28, -23, -23, -5, -12, 6, -22, 2, -7, 18, -6, 3, 5, -6, -17, -9, -21, -7, -7, -20, -16, -5, -3, -10, 9, 20, -7, -12, 5, -12, -2, -15, 2, -6, -4, 1, -20, -4, -10, 26, 14, 9, -6, 6, -19, 6, -15, -17, 5, -10, 0, -4, -15, 13, -2, 18, 3, 5, 19, 13, -2, -11, 4, 8, -15, 1, -12, -12, -6, 6, 15, 17, 23, 1, 18, -1, -19, -22, -12, 7, 6, 13, -6, -2, -5, 17, 2, 13, 5, -1, 0, 10, 0, 10, 12, 11, -15, 9, -3,
    -- filter=0 channel=2
    18, 16, -4, 16, 18, 0, -5, -1, 9, 7, -14, 5, 0, 4, -9, -7, 16, 23, 23, -9, -5, 15, 6, -4, 14, 6, 2, 6, -6, 16, 19, 11, 20, 1, 7, 18, 19, 15, 10, -11, -11, 17, -12, 17, -10, 15, 14, 0, 7, -11, -9, -13, 4, -11, -10, 4, 0, -10, 5, 7, 5, -1, 9, 6, 1, -9, 10, 7, -5, 6, -9, -2, -5, -1, 13, 18, 20, -3, 15, 3, -6, -16, 7, 7, 8, -4, -18, 6, 11, -11, 16, 2, -2, 18, -1, 12, 14, -20, 10, 1, 8, -7, -1, 1, -8, -3, -6, 8, -2, 15, -9, 4, -14, 10, 5, 6, -16, 4, -14, -4, 10, 21, 3, 1, 10, -2, 11, 6, 0, -9, -3, 7, 9, 13, 0, 0, 7, 20, -13, 15, -6, -3, 6, -16, -13, -4, 2, -9, -10, -12, 14, 15, -1, 13, 2, -2, -14, -6, -9, -12, -11, 9, 0, 5, -13, 12, 12, 15, -4, 3, 2, -5, 3, 5, 0, 11, -6, 14, 7, 15, 9, 24, 24, 22, 0, -10, -3, 11, -5, 5, 13, -13, 9, 14, 6, -9, 15, 11, 23, 7, 15, -9, 6, 6, 20, -2, -4, -3, 4, 11, 9, 22, -2, -6, 17, 18, 3, 9, 14, 8, 13, -10, 9, -10, 5,
    -- filter=0 channel=3
    0, 0, 9, -4, 15, 17, 9, 9, 2, 0, -13, 6, -4, -15, 9, 16, -6, 18, -5, 3, 19, 11, 0, -6, 3, -14, 2, 6, 0, -6, 19, 5, 18, -9, -8, -12, 7, -1, -9, -6, 5, 7, -13, 10, 1, -8, -2, 8, 15, 6, 18, 6, 11, -12, 13, 4, 10, -9, -12, -12, 10, 2, 23, 0, -6, 6, 17, -9, 9, -17, 0, -17, 10, -10, 3, 11, 0, -9, 13, 15, 17, 18, -15, 10, 12, -7, -6, 0, -22, 8, -3, -4, -1, -2, 2, -5, -11, -2, 6, -16, -8, -11, -19, -4, 1, 11, 4, 18, -5, -1, -10, 17, 4, -17, 3, 3, -2, -15, 3, -22, 13, 6, -10, 15, 11, -9, -3, -9, -6, 12, -6, 5, -17, -11, -10, -3, 6, 0, 8, -8, 21, 0, 14, -14, -8, -17, -16, 0, 8, -15, 0, 22, 14, 21, 16, -10, 17, 1, 16, 11, 1, -3, -3, 7, -3, 19, 0, 5, -10, -3, 1, -3, -11, -13, 14, -15, -4, 9, -8, -20, 6, 19, 8, -1, 7, -8, -6, 10, -4, 15, -9, 3, 3, 1, 7, -2, 12, -9, -7, 2, 16, -12, -12, 2, 8, -16, 8, 4, -22, -21, 1, 11, 0, 14, -14, -8, -7, 14, 5, -2, -5, -13, 10, -13, -3,
    -- filter=0 channel=4
    0, 13, 0, -5, 1, 11, 10, 10, -17, -16, 10, 3, 3, 7, -13, -5, -9, 3, -4, 7, 16, 13, 7, 11, 14, -7, 10, -1, -1, 14, 11, 15, 14, 14, 17, 17, 15, 1, 5, -4, 10, -7, 1, 13, 10, -11, -4, 3, 15, -2, 18, 12, -3, -10, 20, -9, 2, 4, 7, 12, 4, -8, -10, -2, 6, -4, -10, 13, -3, 2, -7, 11, 11, 13, 21, 12, -1, 9, -6, 10, -6, 8, 4, -3, 9, -12, -12, -10, 0, -10, -7, 2, -10, 18, 9, 13, -13, -8, 12, -6, -9, 0, -2, 4, 0, -12, 6, 17, 18, -2, -4, 11, 3, -6, -9, -10, 0, 0, 6, 14, -13, -5, 1, 4, 15, -8, -7, 16, -1, 8, 5, 3, 6, 7, -9, -12, 9, -2, 0, -6, -9, 9, -11, -14, 6, 15, 13, 2, -1, 23, -8, -13, 4, -10, 1, -10, 19, 2, 5, -4, -4, 5, 21, 5, -7, 12, -1, 14, -1, -8, 11, 1, 19, 14, 7, -9, 0, 17, 5, -5, -13, 10, -9, -9, 7, -10, 8, 9, 0, 9, 0, 0, -8, -8, 19, -5, 6, 16, 7, 2, 14, 7, -7, 9, 4, 2, -8, 8, 21, -4, 10, -4, -2, 4, 16, -8, -9, -5, -5, 12, 9, -14, 13, 9, 16,
    -- filter=0 channel=5
    10, 14, 18, 22, 8, 5, -5, 18, 0, 2, 9, 17, -13, 14, 14, 4, 8, 0, 4, 11, -5, 16, -3, 14, -4, -7, 8, 14, -12, -5, 0, 19, 11, -1, -3, -4, -9, 14, -11, 1, -4, 17, -1, -2, 2, 15, 1, -1, 11, 2, 2, 7, 3, 8, -5, -5, -10, -13, -13, 7, 1, 23, 10, -6, 14, -11, 0, 0, -15, -3, -12, -8, 12, -5, -9, -8, -5, -3, 16, 3, 13, 6, -12, -5, 13, -6, -2, 11, 6, 0, -5, -3, 17, -2, 8, 20, 14, -11, 12, -12, -9, 8, 0, 11, -1, -8, 9, -1, 3, 19, -12, -13, -11, -20, -15, 10, -2, -10, -15, 2, 22, 14, 7, 7, -9, 7, 11, 1, 2, -19, -7, -1, 4, 3, -16, 0, 0, 23, 16, 3, 8, -10, -16, 12, 14, -2, -1, 1, -12, 0, 20, 0, 2, 13, -7, -8, -13, 5, -5, -14, -6, -3, -11, 10, -5, -9, 11, -4, 6, -8, 21, 0, 12, -4, -3, -13, -4, 7, -2, 11, 2, 6, 10, 3, 21, 5, 20, -5, -11, -9, -10, -10, 8, 8, -12, 1, 24, 16, -3, 5, 9, 23, -6, 1, -12, -14, -8, 8, 5, -4, 0, 0, 17, 16, 22, -2, -3, 16, 17, -8, 0, 0, 4, -17, 0,
    -- filter=0 channel=6
    -8, 20, -10, -7, -2, -1, -24, -20, -26, -10, -20, 3, -19, -21, -21, 18, 23, 22, 0, 5, 5, -22, -4, -8, -22, -14, -21, -15, -4, -24, -4, 2, 24, 22, 8, 9, 16, 4, -12, -1, 6, -23, -7, -20, -25, -8, 6, 0, 4, 20, 5, 24, 20, 1, 4, -13, -4, 5, -7, -14, 15, 17, 32, 13, 21, 36, 33, 22, 7, 23, 14, 10, 6, -2, -10, 18, 14, 10, 17, 27, 42, 39, 31, 23, 3, 11, 9, 9, -17, -11, -5, 4, 17, 28, 29, 40, 27, 31, 11, 22, 14, 9, 14, -16, 6, 5, 28, 8, 40, 44, 31, 39, 38, 17, 37, 19, 14, 2, 6, 0, -1, 5, 34, 14, 47, 42, 43, 47, 22, 24, 3, 12, -16, -4, -8, 2, 21, 18, 30, 43, 47, 43, 34, 36, 23, -2, -6, -4, -7, -14, 2, -2, 27, 18, 28, 28, 42, 34, 8, 27, 18, -12, 9, 5, -6, 9, 4, 18, 0, 16, 13, 24, 0, 11, -12, 0, 13, -21, 4, -12, 5, 15, 22, 15, -3, 16, 4, 6, -6, -8, -3, -2, 0, -11, -7, 8, -4, 6, 3, 20, 0, 12, 0, -3, -11, 5, -15, -9, -4, -26, 17, 12, -9, 4, -13, -6, -15, -4, -19, 0, -9, -12, -15, -16, -6,
    -- filter=0 channel=7
    -13, 0, -25, -18, -16, 3, 0, 18, 21, 4, 3, 30, 5, 19, 10, -11, -29, -27, -26, 0, 2, 13, 3, 30, 18, 11, 23, 37, 11, 12, -14, -22, -13, -25, 4, -13, 18, 24, 19, 19, 12, 13, 27, 12, 29, -22, -23, -10, -28, -6, -19, 16, 1, 16, 11, 23, 15, 29, 38, 34, -7, -19, -4, -11, -21, -4, 2, 15, 2, -7, 7, 27, 33, 11, 12, -27, -9, -25, -19, 1, -12, 1, 6, 9, 12, 10, 18, 28, 9, 10, -17, -18, -8, -26, -11, -4, -12, -5, -15, 5, 25, 19, 20, 35, 22, -28, -31, -32, -7, -24, -24, 3, -14, -12, -7, 31, 21, 21, 38, 38, -28, -11, -19, -4, 3, -8, -4, -14, -10, 3, 6, 11, 36, 11, 37, -21, -24, -21, -15, -9, 0, -11, 0, -15, 16, 16, 23, 35, 32, 18, -5, -11, -36, -31, -4, 0, 7, -20, 7, -8, 25, 29, 34, 36, 28, -9, -28, -34, -4, -18, -13, -9, 14, 3, 23, 22, 34, 13, 28, 20, -6, -28, -15, -12, 6, 5, 9, 12, -4, 10, 25, 30, 39, 42, 7, -15, -32, -29, -8, 0, 9, 0, 1, 13, 19, 7, 15, 26, 30, 6, -33, -9, -24, -16, 2, -8, 2, 22, 14, 33, 17, 19, 28, 12, 27,
    -- filter=0 channel=8
    -15, -15, -5, -21, -22, -9, -17, 4, -13, -10, -17, 12, 5, -13, -14, 6, 0, -12, 2, -18, 0, -3, -25, -23, -18, -21, -16, -21, 0, 3, 13, -2, -2, -3, 3, -8, -11, 4, 0, 7, -11, -11, 0, -19, 0, -10, 5, -15, -19, -4, -20, 3, 0, -2, 7, 8, -14, -4, 1, 9, -16, -2, -18, -12, -23, -9, -2, 1, -14, -8, -9, 10, 11, -14, 1, 2, -6, -3, -7, -12, -8, -4, 10, -18, -6, -2, -16, -16, 6, 4, 4, 0, -26, -12, -2, -10, -8, -19, -19, -8, -11, -12, 10, -7, 2, 1, -24, -22, -5, -5, -5, -1, 10, 0, 1, 1, -12, -5, 10, -2, -5, -21, -25, -6, -8, -1, 0, 0, 1, -13, 10, 6, 5, -2, -21, 11, -11, -4, -17, -20, -22, -24, 11, -6, 13, -6, -17, 3, -15, 0, 0, -11, -5, -20, -12, -4, -7, -7, -6, 1, -15, -11, -9, -9, 10, 0, 1, -6, -21, -8, 2, -5, 4, 2, 1, -8, -7, -14, -20, 2, 7, -10, -4, 5, 2, -10, -1, -4, -7, 9, -19, 0, 2, -6, 8, 13, -22, -3, -9, -11, 1, -10, -25, -13, 0, -16, -19, -15, 1, -9, -4, 5, -3, 0, -5, -16, -13, 0, -20, -15, 6, -11, -15, -11, 6,
    -- filter=0 channel=9
    12, -10, -18, -11, -15, -13, 3, 3, 3, 3, 21, 5, -9, 0, -10, 2, -1, -2, -14, -1, 3, -11, 6, 0, 11, 15, 18, 2, 14, -1, 9, -22, -14, -17, -5, -16, -16, -11, -10, -2, -13, 0, 10, -12, 17, -5, -18, -23, -16, -15, 4, -2, -7, 10, 0, 2, 0, 10, -11, 5, 10, 1, -11, 5, 7, -19, 11, 0, 9, 4, -6, -5, 0, -9, -12, 8, 2, -2, 4, -16, -1, 2, 2, 0, 17, -1, -16, 10, -5, -12, -16, -19, -5, -18, -18, -16, -6, 3, 14, 2, 7, -1, 3, 2, -1, 2, -14, -16, 8, 1, 6, 2, -15, 12, 10, 4, -2, -11, -11, -3, -18, -2, 4, -9, -10, -16, -5, 0, 12, 5, -4, 7, 11, -4, -11, 7, -21, 8, 0, -23, -3, 0, -6, 5, 6, 14, 12, 11, -11, 10, 7, -4, -21, 7, 2, -22, -8, 15, -2, -12, -6, -15, 12, -4, -15, 5, -5, 4, -8, -15, -17, 10, 9, -3, -15, 3, 4, 13, -17, 9, 8, -9, -21, -12, -10, -20, 0, 0, 10, 13, -8, -15, 0, 10, -4, -2, -16, -8, -7, -18, 0, 1, -5, -10, 2, 8, -4, 6, -9, -13, -14, 5, -2, -15, 8, -13, -10, -3, 5, -1, -1, 0, -10, -9, 15,

    others => 0);
end iwght_package;
