library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    2234, 6329, 1451, -57756, -288, -5744, 9721, -565, -12213, 26697, 27066, -4754, 8085, 4736, -2394, -6962, -20683, -10580, 36140, 14609, 10691, 13620, -4596, 18860, -3134, -518, 1603, -13151, 4587, -16439, -1333, 15775, 3953, -1920, -509, 11282, 17640, -27361, -17249, -5160, -10529, -29829, -5452, 1396, 3559, -11769, -1087, 1150, -1551, 18144, -100, 32913, 4435, -75, -2904, -8590, -267, -12498, 34788, -37673, -22803, -16482, -32601, 708,

    -- weights
    -- filter=0 channel=0
    0, 33, 28, -37, 54, 38, 6, 0, 26,
    -- filter=0 channel=1
    37, 80, 42, 42, 77, 78, 6, 43, 90,
    -- filter=0 channel=2
    -79, -57, -24, -37, -69, -2, -93, -58, -60,
    -- filter=1 channel=0
    67, 86, 10, 73, 102, 73, 24, 38, 22,
    -- filter=1 channel=1
    -30, -92, -103, -89, -55, -93, -121, -78, -136,
    -- filter=1 channel=2
    67, 70, 52, 31, 47, 34, 63, 45, -17,
    -- filter=2 channel=0
    21, 36, 42, 75, 122, 28, 67, 122, 85,
    -- filter=2 channel=1
    -147, -101, -65, -41, -107, -78, -105, -77, -10,
    -- filter=2 channel=2
    20, 48, 55, 35, 31, 99, 68, 83, 61,
    -- filter=3 channel=0
    -46, -9, 67, -21, 38, 99, 5, 68, 63,
    -- filter=3 channel=1
    -58, 34, -8, 1, -11, -56, -23, 23, -66,
    -- filter=3 channel=2
    40, 17, 70, -12, 87, 40, 27, 39, 59,
    -- filter=4 channel=0
    -13, -45, 18, -33, -4, -29, -38, 13, 5,
    -- filter=4 channel=1
    71, 14, 69, 49, 104, 52, 82, 70, 24,
    -- filter=4 channel=2
    -62, -9, -11, 20, -57, -22, 17, -27, -51,
    -- filter=5 channel=0
    68, -58, -57, 35, 22, 1, 50, -51, -60,
    -- filter=5 channel=1
    42, -20, -44, 65, -40, -53, 41, 7, -13,
    -- filter=5 channel=2
    14, 40, -24, 19, 31, -61, 88, 22, 22,
    -- filter=6 channel=0
    3, 55, 39, 6, -14, 0, -8, 10, 61,
    -- filter=6 channel=1
    -26, -17, 20, 35, -19, -15, -3, 9, 39,
    -- filter=6 channel=2
    -61, -20, 2, -35, 14, 31, 26, 9, -2,
    -- filter=7 channel=0
    64, -15, -37, 1, 12, -28, 89, -51, -34,
    -- filter=7 channel=1
    39, -41, -37, 72, -30, -11, 62, -16, -44,
    -- filter=7 channel=2
    30, -36, 4, -9, 31, -8, 34, -32, -18,
    -- filter=8 channel=0
    -14, 9, 4, -28, 26, 39, 4, -21, 31,
    -- filter=8 channel=1
    62, 46, 74, 105, 108, 58, 101, 138, 60,
    -- filter=8 channel=2
    -49, -17, -74, 35, 7, 6, 36, 8, -50,
    -- filter=9 channel=0
    -170, -198, -127, -172, -151, -168, -170, -147, -162,
    -- filter=9 channel=1
    51, 17, -12, -13, -4, 61, 26, 24, 27,
    -- filter=9 channel=2
    142, 179, 174, 171, 202, 215, 114, 169, 124,
    -- filter=10 channel=0
    55, 39, 53, 21, 61, 22, 65, -6, 0,
    -- filter=10 channel=1
    41, -30, 24, 17, 15, 17, -34, 4, 14,
    -- filter=10 channel=2
    -60, -69, -2, -100, -70, -6, -74, -76, -22,
    -- filter=11 channel=0
    -18, 59, 27, 42, 78, -6, 37, 6, -21,
    -- filter=11 channel=1
    -29, 39, 30, 56, 53, -18, 42, 38, -49,
    -- filter=11 channel=2
    40, 20, -38, 49, 3, -24, -51, -52, 4,
    -- filter=12 channel=0
    -29, -24, 1, -31, -23, 0, -25, 0, -34,
    -- filter=12 channel=1
    39, 12, -10, -33, 23, -8, -41, 19, -43,
    -- filter=12 channel=2
    16, 24, -21, -8, 46, 19, -31, -45, -11,
    -- filter=13 channel=0
    -41, 15, 5, -30, -15, 33, -99, -79, -27,
    -- filter=13 channel=1
    -4, 21, 94, 73, 35, 86, -11, 66, 59,
    -- filter=13 channel=2
    30, 53, 14, 19, 35, -3, -48, -5, -14,
    -- filter=14 channel=0
    72, -38, -19, 67, 5, -73, 62, -51, -62,
    -- filter=14 channel=1
    1, 10, -21, 47, 12, -19, 35, 37, -15,
    -- filter=14 channel=2
    62, -40, -48, 22, -8, -11, -12, 0, -24,
    -- filter=15 channel=0
    -22, -57, -4, -29, 20, 17, -73, 51, 44,
    -- filter=15 channel=1
    33, 45, 40, -1, 127, 110, 50, 108, 109,
    -- filter=15 channel=2
    -33, 7, -21, -48, 51, 5, -40, 48, 46,
    -- filter=16 channel=0
    -36, 1, 59, 17, 63, 30, 28, 24, 56,
    -- filter=16 channel=1
    15, -4, -2, -20, 26, 32, -16, 53, 20,
    -- filter=16 channel=2
    70, 27, 59, 88, 110, 70, 80, 22, 69,
    -- filter=17 channel=0
    -10, -20, 0, 59, 62, 7, 18, -11, -44,
    -- filter=17 channel=1
    43, 33, -24, 108, 78, 69, 93, 106, -15,
    -- filter=17 channel=2
    12, -36, -61, -4, 49, 4, -29, 10, -39,
    -- filter=18 channel=0
    -101, -93, -64, -7, -79, -6, -32, -87, -53,
    -- filter=18 channel=1
    9, 81, 77, 29, 101, 107, 103, 120, 91,
    -- filter=18 channel=2
    -31, 13, -41, -6, -28, -48, -54, -51, -61,
    -- filter=19 channel=0
    30, 11, -65, 94, 58, -67, 40, 21, -42,
    -- filter=19 channel=1
    -61, -16, -82, -7, -74, -111, -15, -91, -130,
    -- filter=19 channel=2
    76, 85, 33, 66, 77, 30, 75, 83, 62,
    -- filter=20 channel=0
    -94, -9, 5, -62, -69, -13, -60, -31, 4,
    -- filter=20 channel=1
    -49, -50, 91, -32, 29, 73, -28, -21, 0,
    -- filter=20 channel=2
    -44, 12, 96, -44, 20, 91, 3, 53, 52,
    -- filter=21 channel=0
    20, -30, -29, -31, -49, -22, -6, 2, 12,
    -- filter=21 channel=1
    -11, -9, -49, 42, 5, -37, -44, 40, -33,
    -- filter=21 channel=2
    -3, -50, 30, -17, 38, -1, 32, -19, 27,
    -- filter=22 channel=0
    -13, -31, 7, 4, 41, -8, -25, -34, -6,
    -- filter=22 channel=1
    1, 46, 5, -12, 12, -28, -7, -7, 48,
    -- filter=22 channel=2
    26, -18, 16, 27, 36, 14, 22, -30, -48,
    -- filter=23 channel=0
    43, 15, 32, 88, 92, 58, 37, 76, 53,
    -- filter=23 channel=1
    30, -20, 37, 44, -4, 15, -12, 8, -44,
    -- filter=23 channel=2
    -58, -45, -63, -99, -14, -66, -82, -56, -98,
    -- filter=24 channel=0
    -13, 0, 30, 49, -24, -22, 32, -22, -62,
    -- filter=24 channel=1
    79, 111, 55, 39, 65, -13, 53, 75, 11,
    -- filter=24 channel=2
    38, -33, 5, -5, -23, -51, 23, -5, -49,
    -- filter=25 channel=0
    79, 63, 95, 74, 143, 122, 99, 73, 154,
    -- filter=25 channel=1
    -173, -133, -144, -138, -62, -90, -161, -105, -139,
    -- filter=25 channel=2
    38, 21, 28, 16, 72, 108, 60, 71, 100,
    -- filter=26 channel=0
    -45, 52, 104, -43, -1, 100, -19, -4, 0,
    -- filter=26 channel=1
    -87, 37, -12, -118, 36, -5, -76, -37, 51,
    -- filter=26 channel=2
    -21, -24, 69, -69, 26, 40, -45, -6, 91,
    -- filter=27 channel=0
    79, 87, 25, 102, 151, 105, 42, 69, 118,
    -- filter=27 channel=1
    -67, -71, -64, 19, 38, -16, -26, 13, -25,
    -- filter=27 channel=2
    -49, -9, -13, 15, 28, 0, -11, 0, 4,
    -- filter=28 channel=0
    -53, 14, -84, 28, -8, -31, -36, -39, -18,
    -- filter=28 channel=1
    -8, 12, -29, 81, 55, 4, 46, 45, 25,
    -- filter=28 channel=2
    73, -1, -32, 82, 104, 8, 46, 100, 31,
    -- filter=29 channel=0
    -97, 21, -35, -25, 53, 42, -81, -11, 73,
    -- filter=29 channel=1
    -9, 1, 65, 14, 95, 53, 38, 59, 53,
    -- filter=29 channel=2
    -7, 74, 99, 67, 143, 117, 33, 61, 91,
    -- filter=30 channel=0
    124, 60, -120, 173, 60, -136, 125, 6, -120,
    -- filter=30 channel=1
    62, 10, -162, 120, -22, -209, 107, -48, -126,
    -- filter=30 channel=2
    47, 57, -88, 120, 56, -149, 74, 47, -103,
    -- filter=31 channel=0
    10, 35, 8, -41, 6, 20, -9, -9, -4,
    -- filter=31 channel=1
    -48, -6, 3, -21, 37, 16, 3, -42, 32,
    -- filter=31 channel=2
    -30, -13, -29, 31, -30, -43, -25, -20, -48,
    -- filter=32 channel=0
    130, 112, 19, 127, 65, 55, 66, 81, 45,
    -- filter=32 channel=1
    -58, -27, -56, -33, -92, -86, -37, -54, -70,
    -- filter=32 channel=2
    -15, -23, 17, -42, -56, 14, -1, -67, -11,
    -- filter=33 channel=0
    7, 48, -42, 14, -47, 40, -13, -34, 33,
    -- filter=33 channel=1
    6, -48, -2, -9, -28, -48, 6, 46, -13,
    -- filter=33 channel=2
    4, 15, 4, -5, -30, -19, -40, 37, -31,
    -- filter=34 channel=0
    -53, 0, 7, 1, 51, -9, -58, 65, -23,
    -- filter=34 channel=1
    -16, 19, 34, -62, 65, 8, -16, -17, 13,
    -- filter=34 channel=2
    -38, 39, -6, -28, 29, -34, -9, 16, 23,
    -- filter=35 channel=0
    102, 140, 44, 81, 153, 124, 100, 158, 121,
    -- filter=35 channel=1
    -82, -85, -15, -69, -6, -33, -91, 12, -33,
    -- filter=35 channel=2
    -108, -6, -84, -83, -92, -8, -48, -19, -84,
    -- filter=36 channel=0
    35, 20, -29, -33, -17, 48, 42, 41, -45,
    -- filter=36 channel=1
    -9, -39, -3, 19, 19, 41, -41, -34, -48,
    -- filter=36 channel=2
    -21, -12, -22, -21, -28, -22, -1, -32, -6,
    -- filter=37 channel=0
    -11, 17, -44, 21, -1, 39, -59, -28, -13,
    -- filter=37 channel=1
    -9, 49, -66, -24, 13, 0, -26, 0, -68,
    -- filter=37 channel=2
    67, 104, 31, 88, 124, 21, 52, 71, 34,
    -- filter=38 channel=0
    29, 113, 48, 28, 118, 79, 30, 80, 64,
    -- filter=38 channel=1
    -15, 67, 3, -5, -15, 33, -65, 9, 24,
    -- filter=38 channel=2
    -31, 64, 7, 18, -18, 14, 24, 5, -54,
    -- filter=39 channel=0
    -24, 42, -39, -22, -15, -17, -15, -8, 7,
    -- filter=39 channel=1
    -10, -4, -47, 31, 18, 4, 49, 9, 11,
    -- filter=39 channel=2
    -24, -21, -8, -46, -29, 24, 40, 24, 19,
    -- filter=40 channel=0
    8, 15, 3, 70, 58, 21, 42, -21, -3,
    -- filter=40 channel=1
    -65, -36, 8, 35, -30, 19, 6, 42, -18,
    -- filter=40 channel=2
    -4, -37, -14, -48, -21, 3, -15, 44, 19,
    -- filter=41 channel=0
    0, -14, 54, 36, 119, 57, 10, 106, 7,
    -- filter=41 channel=1
    -13, -6, -9, 40, 121, 90, -9, 103, 75,
    -- filter=41 channel=2
    -76, -27, -16, 10, 42, 40, 17, 37, 47,
    -- filter=42 channel=0
    -30, 1, 32, 22, -17, -48, -21, 38, -38,
    -- filter=42 channel=1
    -24, -2, -6, -7, -11, -25, 27, -31, -44,
    -- filter=42 channel=2
    -49, 42, -4, 8, 12, -49, -25, -41, 40,
    -- filter=43 channel=0
    113, 171, 87, -18, 59, -5, -20, -90, -95,
    -- filter=43 channel=1
    79, 43, 92, -45, -56, -21, -110, -168, -141,
    -- filter=43 channel=2
    69, 102, 138, 26, 23, 59, -113, -119, -95,
    -- filter=44 channel=0
    64, -11, 71, 110, 41, 54, 97, 52, 38,
    -- filter=44 channel=1
    -35, -90, -91, 47, -93, -120, 32, -91, -97,
    -- filter=44 channel=2
    59, 3, -51, 13, -58, 10, 43, 16, 7,
    -- filter=45 channel=0
    0, 48, -41, 23, 8, -11, -21, -42, -43,
    -- filter=45 channel=1
    3, -43, -41, -23, 30, -14, 12, -35, 22,
    -- filter=45 channel=2
    6, 0, -25, 2, 47, 38, -28, -34, 1,
    -- filter=46 channel=0
    -75, -28, 59, -66, -5, 52, -27, 35, 27,
    -- filter=46 channel=1
    -57, -6, 72, -27, 0, 54, -65, -13, 81,
    -- filter=46 channel=2
    -63, 37, 16, -72, 46, 38, -63, -12, 66,
    -- filter=47 channel=0
    -35, 45, 7, -24, 39, -41, 31, -2, -24,
    -- filter=47 channel=1
    -38, -7, 3, -35, 33, 33, -22, -18, -45,
    -- filter=47 channel=2
    -42, 21, -5, -46, -33, -4, 32, 10, -6,
    -- filter=48 channel=0
    -17, 16, 15, -58, -50, 47, -74, -12, 55,
    -- filter=48 channel=1
    -47, -4, -12, 2, 22, 38, -21, 2, 60,
    -- filter=48 channel=2
    49, 53, 4, -7, 20, 45, 5, 76, 44,
    -- filter=49 channel=0
    0, -42, -39, 32, 74, 11, 39, 78, 70,
    -- filter=49 channel=1
    -35, 3, -10, 34, 71, 81, 60, 76, 70,
    -- filter=49 channel=2
    -33, -70, -124, -73, -24, -63, -65, -67, -21,
    -- filter=50 channel=0
    54, 39, -67, 123, -41, -63, 111, -38, -44,
    -- filter=50 channel=1
    103, 14, -66, 32, -13, -64, 36, -88, -96,
    -- filter=50 channel=2
    78, 51, 29, 80, -10, -69, 19, -79, -50,
    -- filter=51 channel=0
    41, 13, -41, -12, 12, 8, -1, -17, -12,
    -- filter=51 channel=1
    87, 70, 64, 57, 35, 97, 22, 107, 88,
    -- filter=51 channel=2
    -89, -74, -51, -54, -117, -84, -87, -100, -91,
    -- filter=52 channel=0
    35, -2, -35, -35, -1, 45, -8, 9, -46,
    -- filter=52 channel=1
    32, -4, -2, -33, 38, 25, -20, -15, 4,
    -- filter=52 channel=2
    -22, 1, -11, -44, 8, -39, -31, 26, -48,
    -- filter=53 channel=0
    156, 28, -54, 162, -24, -35, 96, 22, 17,
    -- filter=53 channel=1
    89, -78, -141, 76, -60, -140, -32, -61, -35,
    -- filter=53 channel=2
    127, 16, -88, 31, 25, -110, 76, -55, -46,
    -- filter=54 channel=0
    -119, -61, -137, -100, -107, -158, -119, -116, -120,
    -- filter=54 channel=1
    0, -28, -13, 46, 58, 9, 16, 54, -15,
    -- filter=54 channel=2
    109, 82, 41, 141, 195, 126, 137, 192, 89,
    -- filter=55 channel=0
    -32, 26, -23, -6, -20, -3, -43, -10, 20,
    -- filter=55 channel=1
    -47, 37, 17, 43, 45, -42, -20, 0, 19,
    -- filter=55 channel=2
    -1, 15, -12, 11, 13, -7, 17, -40, -29,
    -- filter=56 channel=0
    -40, -45, 64, 21, -47, 43, 3, -21, -9,
    -- filter=56 channel=1
    36, -16, 14, 31, -3, 6, -16, 27, -31,
    -- filter=56 channel=2
    43, -55, 7, 23, -26, -27, 39, -12, -14,
    -- filter=57 channel=0
    41, 25, -30, -36, 3, 21, -43, -29, -3,
    -- filter=57 channel=1
    -9, 36, 27, -45, -22, -23, -25, -36, -7,
    -- filter=57 channel=2
    0, 37, 2, -41, -45, -34, -32, 24, 41,
    -- filter=58 channel=0
    0, -38, -10, 0, -5, -24, -25, 0, 5,
    -- filter=58 channel=1
    -14, -14, 18, -4, -11, -30, -21, -41, 27,
    -- filter=58 channel=2
    -27, 21, -27, -7, 7, 55, -49, -17, 49,
    -- filter=59 channel=0
    -4, 86, 90, 29, 40, 114, -5, 76, 102,
    -- filter=59 channel=1
    -21, -57, -24, -53, 9, 24, -9, 9, 34,
    -- filter=59 channel=2
    -1, 30, 50, 38, 14, 91, -1, 83, 18,
    -- filter=60 channel=0
    -24, -4, 52, -23, 39, 64, -87, 44, 34,
    -- filter=60 channel=1
    72, 141, 106, 95, 188, 145, 9, 166, 126,
    -- filter=60 channel=2
    -53, -39, -31, 26, 68, -30, -59, -15, -75,
    -- filter=61 channel=0
    38, 68, 27, 15, 52, 6, 19, -25, -4,
    -- filter=61 channel=1
    121, 121, 68, 93, 89, 35, 110, 122, 52,
    -- filter=61 channel=2
    -44, -63, -72, -29, 31, -29, -43, -43, -117,
    -- filter=62 channel=0
    -3, 42, -21, 5, 70, 74, 11, 36, 43,
    -- filter=62 channel=1
    -1, 28, -45, 43, -26, -57, 29, -10, -32,
    -- filter=62 channel=2
    52, 6, 31, 68, 73, -19, 79, 65, -33,
    -- filter=63 channel=0
    -8, -25, -3, 10, -41, 37, 3, -7, -33,
    -- filter=63 channel=1
    -41, -43, -3, -24, -17, -29, -38, -47, -6,
    -- filter=63 channel=2
    -9, 10, -40, 8, 31, 33, -34, 25, 23,

    others => 0);
end iwght_package;
